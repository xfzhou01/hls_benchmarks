// Processed by function `construct_kairos` in `verilog_tricks.py`.
// Machine A:
// Processed by function `add_clk_enable_signal` in `verilog_tricks.py`.
// Processed by function `remove_reset_signal` in `verilog_tricks.py`.
module top_A (
  ap_clk,
  ap_start,
  ap_done,
  ap_idle,
  ap_ready,
  op_0,
  op_1,
  op_4,
  op_6,
  op_8,
  op_11,
  op_15,
  op_28,
  op_28_ap_vld,
clk_enable
);
input clk_enable;


input ap_clk;
wire ap_rst;
assign ap_rst = op_28_ap_vld;
input ap_start;
input [1:0] op_0;
input [15:0] op_1;
input [31:0] op_11;
input [15:0] op_15;
input [7:0] op_4;
input [31:0] op_6;
input [7:0] op_8;
output ap_done;
output ap_idle;
output ap_ready;
output [31:0] op_28;
output op_28_ap_vld;


reg Range1_all_ones_1_reg_1647;
reg Range1_all_ones_reg_1706;
reg Range1_all_zeros_1_reg_1654;
reg Range1_all_zeros_reg_1713;
reg Range2_all_ones_1_reg_1642;
reg Range2_all_ones_reg_1701;
reg [8:0] \add_17ns_17ns_17_2_1_U10.top_add_17ns_17ns_17_2_1_Adder_5_U.ain_s1 ;
reg [8:0] \add_17ns_17ns_17_2_1_U10.top_add_17ns_17ns_17_2_1_Adder_5_U.bin_s1 ;
reg \add_17ns_17ns_17_2_1_U10.top_add_17ns_17ns_17_2_1_Adder_5_U.carry_s1 ;
reg [7:0] \add_17ns_17ns_17_2_1_U10.top_add_17ns_17ns_17_2_1_Adder_5_U.sum_s1 ;
reg [9:0] \add_19s_19ns_19_2_1_U12.top_add_19s_19ns_19_2_1_Adder_7_U.ain_s1 ;
reg [9:0] \add_19s_19ns_19_2_1_U12.top_add_19s_19ns_19_2_1_Adder_7_U.bin_s1 ;
reg \add_19s_19ns_19_2_1_U12.top_add_19s_19ns_19_2_1_Adder_7_U.carry_s1 ;
reg [8:0] \add_19s_19ns_19_2_1_U12.top_add_19s_19ns_19_2_1_Adder_7_U.sum_s1 ;
reg [12:0] \add_25s_25s_25_2_1_U11.top_add_25s_25s_25_2_1_Adder_6_U.ain_s1 ;
reg [12:0] \add_25s_25s_25_2_1_U11.top_add_25s_25s_25_2_1_Adder_6_U.bin_s1 ;
reg \add_25s_25s_25_2_1_U11.top_add_25s_25s_25_2_1_Adder_6_U.carry_s1 ;
reg [11:0] \add_25s_25s_25_2_1_U11.top_add_25s_25s_25_2_1_Adder_6_U.sum_s1 ;
reg \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_2_U.ain_s1 ;
reg \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_2_U.bin_s1 ;
reg \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_2_U.carry_s1 ;
reg \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_2_U.sum_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.ain_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.bin_s1 ;
reg \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.carry_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.sum_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.ain_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.bin_s1 ;
reg \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.carry_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.sum_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.ain_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.bin_s1 ;
reg \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.carry_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.sum_s1 ;
reg [15:0] \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_14_U.ain_s1 ;
reg [15:0] \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_14_U.bin_s1 ;
reg \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_14_U.carry_s1 ;
reg [15:0] \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_14_U.sum_s1 ;
reg [16:0] \add_33ns_33s_33_2_1_U6.top_add_33ns_33s_33_2_1_Adder_3_U.ain_s1 ;
reg [16:0] \add_33ns_33s_33_2_1_U6.top_add_33ns_33s_33_2_1_Adder_3_U.bin_s1 ;
reg \add_33ns_33s_33_2_1_U6.top_add_33ns_33s_33_2_1_Adder_3_U.carry_s1 ;
reg [15:0] \add_33ns_33s_33_2_1_U6.top_add_33ns_33s_33_2_1_Adder_3_U.sum_s1 ;
reg [17:0] \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.ain_s1 ;
reg [17:0] \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.bin_s1 ;
reg \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.carry_s1 ;
reg [16:0] \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.sum_s1 ;
reg [1:0] \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_8_U.ain_s1 ;
reg [1:0] \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_8_U.bin_s1 ;
reg \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_8_U.carry_s1 ;
reg \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_8_U.sum_s1 ;
reg [22:0] \add_46s_46s_46_2_1_U18.top_add_46s_46s_46_2_1_Adder_12_U.ain_s1 ;
reg [22:0] \add_46s_46s_46_2_1_U18.top_add_46s_46s_46_2_1_Adder_12_U.bin_s1 ;
reg \add_46s_46s_46_2_1_U18.top_add_46s_46s_46_2_1_Adder_12_U.carry_s1 ;
reg [22:0] \add_46s_46s_46_2_1_U18.top_add_46s_46s_46_2_1_Adder_12_U.sum_s1 ;
reg [1:0] \add_4ns_4ns_4_2_1_U7.top_add_4ns_4ns_4_2_1_Adder_4_U.ain_s1 ;
reg [1:0] \add_4ns_4ns_4_2_1_U7.top_add_4ns_4ns_4_2_1_Adder_4_U.bin_s1 ;
reg \add_4ns_4ns_4_2_1_U7.top_add_4ns_4ns_4_2_1_Adder_4_U.carry_s1 ;
reg [1:0] \add_4ns_4ns_4_2_1_U7.top_add_4ns_4ns_4_2_1_Adder_4_U.sum_s1 ;
reg [1:0] \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_4_U.ain_s1 ;
reg [1:0] \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_4_U.bin_s1 ;
reg \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_4_U.carry_s1 ;
reg [1:0] \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_4_U.sum_s1 ;
reg [1:0] \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.ain_s1 ;
reg [1:0] \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.bin_s1 ;
reg \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.carry_s1 ;
reg [1:0] \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.sum_s1 ;
reg [2:0] \add_5s_5s_5_2_1_U16.top_add_5s_5s_5_2_1_Adder_10_U.ain_s1 ;
reg [2:0] \add_5s_5s_5_2_1_U16.top_add_5s_5s_5_2_1_Adder_10_U.bin_s1 ;
reg \add_5s_5s_5_2_1_U16.top_add_5s_5s_5_2_1_Adder_10_U.carry_s1 ;
reg [1:0] \add_5s_5s_5_2_1_U16.top_add_5s_5s_5_2_1_Adder_10_U.sum_s1 ;
reg [2:0] \add_6ns_6ns_6_2_1_U19.top_add_6ns_6ns_6_2_1_Adder_13_U.ain_s1 ;
reg [2:0] \add_6ns_6ns_6_2_1_U19.top_add_6ns_6ns_6_2_1_Adder_13_U.bin_s1 ;
reg \add_6ns_6ns_6_2_1_U19.top_add_6ns_6ns_6_2_1_Adder_13_U.carry_s1 ;
reg [2:0] \add_6ns_6ns_6_2_1_U19.top_add_6ns_6ns_6_2_1_Adder_13_U.sum_s1 ;
reg [31:0] add_ln691_1_reg_2060;
reg [31:0] add_ln691_2_reg_2124;
reg [18:0] add_ln691_reg_1967;
reg [2:0] add_ln69_1_reg_2028;
reg [4:0] add_ln69_2_reg_2055;
reg [31:0] add_ln69_reg_2144;
reg and_ln406_reg_1696;
reg and_ln408_reg_1718;
reg and_ln785_1_reg_1924;
reg and_ln785_5_reg_1935;
reg and_ln786_1_reg_1900;
reg and_ln786_reg_1880;
reg [30:0] ap_CS_fsm = 31'h00000001;
reg carry_1_reg_1839;
reg carry_3_reg_1846;
reg deleted_zeros_1_reg_1888;
reg deleted_zeros_reg_1868;
reg icmp_ln1496_reg_1504;
reg icmp_ln851_1_reg_1723;
reg icmp_ln851_2_reg_2114;
reg icmp_ln851_3_reg_1686;
reg icmp_ln851_4_reg_1863;
reg icmp_ln851_5_reg_2023;
reg icmp_ln851_6_reg_2080;
reg icmp_ln851_reg_1590;
reg icmp_ln874_reg_1824;
reg lhs_V_4_reg_1585;
reg [3:0] \mul_4ns_4s_8_7_1_U14.top_mul_4ns_4s_8_7_1_Mul_DSP_2_U.a_reg0 ;
reg [3:0] \mul_4ns_4s_8_7_1_U14.top_mul_4ns_4s_8_7_1_Mul_DSP_2_U.b_reg0 ;
reg [7:0] \mul_4ns_4s_8_7_1_U14.top_mul_4ns_4s_8_7_1_Mul_DSP_2_U.buff0 ;
reg [7:0] \mul_4ns_4s_8_7_1_U14.top_mul_4ns_4s_8_7_1_Mul_DSP_2_U.buff1 ;
reg [7:0] \mul_4ns_4s_8_7_1_U14.top_mul_4ns_4s_8_7_1_Mul_DSP_2_U.buff2 ;
reg [7:0] \mul_4ns_4s_8_7_1_U14.top_mul_4ns_4s_8_7_1_Mul_DSP_2_U.buff3 ;
reg [7:0] \mul_4ns_4s_8_7_1_U14.top_mul_4ns_4s_8_7_1_Mul_DSP_2_U.buff4 ;
reg [7:0] \mul_8ns_8s_16_7_1_U2.top_mul_8ns_8s_16_7_1_Mul_DSP_1_U.a_reg0 ;
reg [7:0] \mul_8ns_8s_16_7_1_U2.top_mul_8ns_8s_16_7_1_Mul_DSP_1_U.b_reg0 ;
reg [15:0] \mul_8ns_8s_16_7_1_U2.top_mul_8ns_8s_16_7_1_Mul_DSP_1_U.buff0 ;
reg [15:0] \mul_8ns_8s_16_7_1_U2.top_mul_8ns_8s_16_7_1_Mul_DSP_1_U.buff1 ;
reg [15:0] \mul_8ns_8s_16_7_1_U2.top_mul_8ns_8s_16_7_1_Mul_DSP_1_U.buff2 ;
reg [15:0] \mul_8ns_8s_16_7_1_U2.top_mul_8ns_8s_16_7_1_Mul_DSP_1_U.buff3 ;
reg [15:0] \mul_8ns_8s_16_7_1_U2.top_mul_8ns_8s_16_7_1_Mul_DSP_1_U.buff4 ;
reg [7:0] \mul_8s_3ns_11_7_1_U1.top_mul_8s_3ns_11_7_1_Mul_DSP_0_U.a_reg0 ;
reg [2:0] \mul_8s_3ns_11_7_1_U1.top_mul_8s_3ns_11_7_1_Mul_DSP_0_U.b_reg0 ;
reg [10:0] \mul_8s_3ns_11_7_1_U1.top_mul_8s_3ns_11_7_1_Mul_DSP_0_U.buff0 ;
reg [10:0] \mul_8s_3ns_11_7_1_U1.top_mul_8s_3ns_11_7_1_Mul_DSP_0_U.buff1 ;
reg [10:0] \mul_8s_3ns_11_7_1_U1.top_mul_8s_3ns_11_7_1_Mul_DSP_0_U.buff2 ;
reg [10:0] \mul_8s_3ns_11_7_1_U1.top_mul_8s_3ns_11_7_1_Mul_DSP_0_U.buff3 ;
reg [10:0] \mul_8s_3ns_11_7_1_U1.top_mul_8s_3ns_11_7_1_Mul_DSP_0_U.buff4 ;
reg [3:0] op_14_V_reg_1972;
reg [3:0] op_16_V_reg_2003;
reg [3:0] op_9_V_reg_1977;
reg or_ln340_1_reg_1929;
reg or_ln340_reg_1918;
reg [9:0] p_Result_1_reg_1631;
reg p_Result_21_reg_1602;
reg p_Result_23_reg_1615;
reg p_Result_24_reg_1769;
reg p_Result_25_reg_1620;
reg p_Result_26_reg_1536;
reg p_Result_27_reg_1637;
reg p_Result_28_reg_1553;
reg p_Result_29_reg_1785;
reg p_Result_30_reg_1558;
reg [8:0] p_Result_s_22_reg_1626;
reg [3:0] p_Val2_2_reg_1610;
reg [3:0] p_Val2_3_reg_1760;
reg [3:0] p_Val2_6_reg_1543;
reg [3:0] p_Val2_7_reg_1776;
reg r_1_reg_1548;
reg [15:0] r_V_3_reg_1595;
reg [10:0] r_V_4_reg_1526;
reg [7:0] r_V_reg_2085;
reg [16:0] ret_V_12_reg_1733;
reg [16:0] ret_V_13_reg_1797;
reg [32:0] ret_V_18_reg_1509;
reg [1:0] ret_V_19_reg_1740;
reg [6:0] ret_V_21_reg_1659;
reg [3:0] ret_V_22_reg_1792;
reg [5:0] ret_V_23_reg_2129;
reg [32:0] ret_V_24_reg_1728;
reg [24:0] ret_V_25_reg_1908;
reg [34:0] ret_V_26_reg_2033;
reg [45:0] ret_V_27_reg_2102;
reg [31:0] ret_V_28_reg_2134;
reg [31:0] ret_V_34_cast_reg_2038;
reg [31:0] ret_V_36_cast_reg_2107;
reg [12:0] ret_V_3_reg_1802;
reg [3:0] ret_V_6_cast_reg_1664;
reg [3:0] ret_V_6_reg_1755;
reg [5:0] ret_V_7_reg_2090;
reg [5:0] ret_V_9_reg_2119;
reg [1:0] ret_V_cast_reg_1514;
reg [1:0] ret_V_reg_1691;
reg sel_tmp11_reg_1952;
reg sel_tmp25_reg_1962;
reg [3:0] select_ln340_1_reg_1957;
reg [3:0] select_ln340_reg_1947;
reg [31:0] select_ln353_1_reg_2065;
reg [18:0] select_ln353_reg_1983;
reg [16:0] select_ln850_5_reg_1829;
reg [18:0] sext_ln850_reg_1940;
reg signbit_reg_1488;
reg [16:0] \sub_33s_33s_33_2_1_U3.top_sub_33s_33s_33_2_1_Adder_0_U.ain_s1 ;
reg [16:0] \sub_33s_33s_33_2_1_U3.top_sub_33s_33s_33_2_1_Adder_0_U.bin_s1 ;
reg \sub_33s_33s_33_2_1_U3.top_sub_33s_33s_33_2_1_Adder_0_U.carry_s1 ;
reg [15:0] \sub_33s_33s_33_2_1_U3.top_sub_33s_33s_33_2_1_Adder_0_U.sum_s1 ;
reg [3:0] \sub_7ns_7ns_7_2_1_U4.top_sub_7ns_7ns_7_2_1_Adder_1_U.ain_s1 ;
reg [3:0] \sub_7ns_7ns_7_2_1_U4.top_sub_7ns_7ns_7_2_1_Adder_1_U.bin_s1 ;
reg \sub_7ns_7ns_7_2_1_U4.top_sub_7ns_7ns_7_2_1_Adder_1_U.carry_s1 ;
reg [2:0] \sub_7ns_7ns_7_2_1_U4.top_sub_7ns_7ns_7_2_1_Adder_1_U.sum_s1 ;
reg [3:0] tmp_1_reg_1564;
reg [4:0] tmp_2_reg_1569;
reg [17:0] tmp_3_reg_1913;
reg [1:0] trunc_ln1115_reg_1531;
reg [3:0] trunc_ln728_reg_1478;
reg [2:0] trunc_ln851_1_reg_1671;
reg [1:0] trunc_ln851_2_reg_2097;
reg [3:0] trunc_ln851_4_reg_1834;
reg [1:0] trunc_ln851_5_reg_1988;
reg [6:0] trunc_ln851_reg_1521;
reg xor_ln416_1_reg_1813;
reg xor_ln416_reg_1807;
reg xor_ln785_1_reg_1874;
reg xor_ln785_3_reg_1894;
reg [3:0] _700_;
wire _000_;
wire _001_;
wire _002_;
wire _003_;
wire _004_;
wire _005_;
wire [31:0] _006_;
wire [31:0] _007_;
wire [18:0] _008_;
wire [2:0] _009_;
wire [4:0] _010_;
wire [31:0] _011_;
wire _012_;
wire _013_;
wire _014_;
wire _015_;
wire _016_;
wire _017_;
wire [30:0] _018_;
wire _019_;
wire _020_;
wire _021_;
wire _022_;
wire _023_;
wire _024_;
wire _025_;
wire _026_;
wire _027_;
wire _028_;
wire _029_;
wire _030_;
wire _031_;
wire _032_;
wire [3:0] _033_;
wire [3:0] _034_;
wire [3:0] _035_;
wire _036_;
wire _037_;
wire [9:0] _038_;
wire _039_;
wire _040_;
wire _041_;
wire _042_;
wire _043_;
wire _044_;
wire _045_;
wire _046_;
wire _047_;
wire [8:0] _048_;
wire [3:0] _049_;
wire [3:0] _050_;
wire [3:0] _051_;
wire [3:0] _052_;
wire _053_;
wire [15:0] _054_;
wire [10:0] _055_;
wire [7:0] _056_;
wire [16:0] _057_;
wire [16:0] _058_;
wire [32:0] _059_;
wire [1:0] _060_;
wire [6:0] _061_;
wire [3:0] _062_;
wire [5:0] _063_;
wire [32:0] _064_;
wire [24:0] _065_;
wire [34:0] _066_;
wire [45:0] _067_;
wire [31:0] _068_;
wire [31:0] _069_;
wire [31:0] _070_;
wire [12:0] _071_;
wire [3:0] _072_;
wire [3:0] _073_;
wire [5:0] _074_;
wire [5:0] _075_;
wire [1:0] _076_;
wire [1:0] _077_;
wire _078_;
wire _079_;
wire [3:0] _080_;
wire [3:0] _081_;
wire [31:0] _082_;
wire [18:0] _083_;
wire [16:0] _084_;
wire [18:0] _085_;
wire _086_;
wire [3:0] _087_;
wire [4:0] _088_;
wire [17:0] _089_;
wire [1:0] _090_;
wire [3:0] _091_;
wire [2:0] _092_;
wire [1:0] _093_;
wire [3:0] _094_;
wire [1:0] _095_;
wire [6:0] _096_;
wire _097_;
wire _098_;
wire _099_;
wire _100_;
wire [3:0] _101_;
wire [1:0] _102_;
wire _103_;
wire _104_;
wire _105_;
wire _106_;
wire _107_;
wire _108_;
wire _109_;
wire _110_;
wire _111_;
wire _112_;
wire _113_;
wire _114_;
wire _115_;
wire _116_;
wire _117_;
wire _118_;
wire _119_;
wire _120_;
wire _121_;
wire _122_;
wire _123_;
wire _124_;
wire [8:0] _125_;
wire [8:0] _126_;
wire _127_;
wire [7:0] _128_;
wire [8:0] _129_;
wire [9:0] _130_;
wire [9:0] _131_;
wire [9:0] _132_;
wire _133_;
wire [8:0] _134_;
wire [9:0] _135_;
wire [10:0] _136_;
wire [12:0] _137_;
wire [12:0] _138_;
wire _139_;
wire [11:0] _140_;
wire [12:0] _141_;
wire [13:0] _142_;
wire _143_;
wire _144_;
wire _145_;
wire _146_;
wire [1:0] _147_;
wire [1:0] _148_;
wire [15:0] _149_;
wire [15:0] _150_;
wire _151_;
wire [15:0] _152_;
wire [16:0] _153_;
wire [16:0] _154_;
wire [15:0] _155_;
wire [15:0] _156_;
wire _157_;
wire [15:0] _158_;
wire [16:0] _159_;
wire [16:0] _160_;
wire [15:0] _161_;
wire [15:0] _162_;
wire _163_;
wire [15:0] _164_;
wire [16:0] _165_;
wire [16:0] _166_;
wire [15:0] _167_;
wire [15:0] _168_;
wire _169_;
wire [15:0] _170_;
wire [16:0] _171_;
wire [16:0] _172_;
wire [16:0] _173_;
wire [16:0] _174_;
wire _175_;
wire [15:0] _176_;
wire [16:0] _177_;
wire [17:0] _178_;
wire [17:0] _179_;
wire [17:0] _180_;
wire _181_;
wire [16:0] _182_;
wire [17:0] _183_;
wire [18:0] _184_;
wire [1:0] _185_;
wire [1:0] _186_;
wire _187_;
wire _188_;
wire [1:0] _189_;
wire [2:0] _190_;
wire [22:0] _191_;
wire [22:0] _192_;
wire _193_;
wire [22:0] _194_;
wire [23:0] _195_;
wire [23:0] _196_;
wire [1:0] _197_;
wire [1:0] _198_;
wire _199_;
wire [1:0] _200_;
wire [2:0] _201_;
wire [2:0] _202_;
wire [1:0] _203_;
wire [1:0] _204_;
wire _205_;
wire [1:0] _206_;
wire [2:0] _207_;
wire [2:0] _208_;
wire [1:0] _209_;
wire [1:0] _210_;
wire _211_;
wire [1:0] _212_;
wire [2:0] _213_;
wire [2:0] _214_;
wire [2:0] _215_;
wire [2:0] _216_;
wire _217_;
wire [1:0] _218_;
wire [2:0] _219_;
wire [3:0] _220_;
wire [2:0] _221_;
wire [2:0] _222_;
wire _223_;
wire [2:0] _224_;
wire [3:0] _225_;
wire [3:0] _226_;
wire [3:0] _227_;
wire [3:0] _228_;
wire [7:0] _229_;
wire [7:0] _230_;
wire [7:0] _231_;
wire [7:0] _232_;
wire [7:0] _233_;
wire [7:0] _234_;
wire [7:0] _235_;
wire [15:0] _236_;
wire [15:0] _237_;
wire [15:0] _238_;
wire [15:0] _239_;
wire [15:0] _240_;
wire [7:0] _241_;
wire [2:0] _242_;
wire [10:0] _243_;
wire [10:0] _244_;
wire [10:0] _245_;
wire [10:0] _246_;
wire [10:0] _247_;
wire [16:0] _248_;
wire [16:0] _249_;
wire _250_;
wire [15:0] _251_;
wire [16:0] _252_;
wire [17:0] _253_;
wire [3:0] _254_;
wire [3:0] _255_;
wire _256_;
wire [2:0] _257_;
wire [3:0] _258_;
wire [4:0] _259_;
wire _260_;
wire _261_;
wire _262_;
wire _263_;
wire _264_;
wire _265_;
wire _266_;
wire _267_;
wire _268_;
wire _269_;
wire _270_;
wire _271_;
wire _272_;
wire _273_;
wire _274_;
wire _275_;
wire _276_;
wire _277_;
wire _278_;
wire _279_;
wire _280_;
wire _281_;
wire _282_;
wire _283_;
wire _284_;
wire _285_;
wire _286_;
wire _287_;
wire _288_;
wire _289_;
wire _290_;
wire _291_;
wire _292_;
wire _293_;
wire _294_;
wire _295_;
wire _296_;
wire _297_;
wire Range1_all_ones_1_fu_515_p2;
wire Range1_all_ones_fu_596_p2;
wire Range1_all_zeros_1_fu_520_p2;
wire Range1_all_zeros_fu_601_p2;
wire Range2_all_ones_1_fu_510_p2;
wire Range2_all_ones_fu_591_p2;
wire \add_17ns_17ns_17_2_1_U10.ce ;
wire \add_17ns_17ns_17_2_1_U10.clk ;
wire [16:0] \add_17ns_17ns_17_2_1_U10.din0 ;
wire [16:0] \add_17ns_17ns_17_2_1_U10.din1 ;
wire [16:0] \add_17ns_17ns_17_2_1_U10.dout ;
wire \add_17ns_17ns_17_2_1_U10.reset ;
wire [16:0] \add_17ns_17ns_17_2_1_U10.top_add_17ns_17ns_17_2_1_Adder_5_U.a ;
wire [16:0] \add_17ns_17ns_17_2_1_U10.top_add_17ns_17ns_17_2_1_Adder_5_U.ain_s0 ;
wire [16:0] \add_17ns_17ns_17_2_1_U10.top_add_17ns_17ns_17_2_1_Adder_5_U.b ;
wire [16:0] \add_17ns_17ns_17_2_1_U10.top_add_17ns_17ns_17_2_1_Adder_5_U.bin_s0 ;
wire \add_17ns_17ns_17_2_1_U10.top_add_17ns_17ns_17_2_1_Adder_5_U.ce ;
wire \add_17ns_17ns_17_2_1_U10.top_add_17ns_17ns_17_2_1_Adder_5_U.clk ;
wire \add_17ns_17ns_17_2_1_U10.top_add_17ns_17ns_17_2_1_Adder_5_U.facout_s1 ;
wire \add_17ns_17ns_17_2_1_U10.top_add_17ns_17ns_17_2_1_Adder_5_U.facout_s2 ;
wire [7:0] \add_17ns_17ns_17_2_1_U10.top_add_17ns_17ns_17_2_1_Adder_5_U.fas_s1 ;
wire [8:0] \add_17ns_17ns_17_2_1_U10.top_add_17ns_17ns_17_2_1_Adder_5_U.fas_s2 ;
wire \add_17ns_17ns_17_2_1_U10.top_add_17ns_17ns_17_2_1_Adder_5_U.reset ;
wire [16:0] \add_17ns_17ns_17_2_1_U10.top_add_17ns_17ns_17_2_1_Adder_5_U.s ;
wire [7:0] \add_17ns_17ns_17_2_1_U10.top_add_17ns_17ns_17_2_1_Adder_5_U.u1.a ;
wire [7:0] \add_17ns_17ns_17_2_1_U10.top_add_17ns_17ns_17_2_1_Adder_5_U.u1.b ;
wire \add_17ns_17ns_17_2_1_U10.top_add_17ns_17ns_17_2_1_Adder_5_U.u1.cin ;
wire \add_17ns_17ns_17_2_1_U10.top_add_17ns_17ns_17_2_1_Adder_5_U.u1.cout ;
wire [7:0] \add_17ns_17ns_17_2_1_U10.top_add_17ns_17ns_17_2_1_Adder_5_U.u1.s ;
wire [8:0] \add_17ns_17ns_17_2_1_U10.top_add_17ns_17ns_17_2_1_Adder_5_U.u2.a ;
wire [8:0] \add_17ns_17ns_17_2_1_U10.top_add_17ns_17ns_17_2_1_Adder_5_U.u2.b ;
wire \add_17ns_17ns_17_2_1_U10.top_add_17ns_17ns_17_2_1_Adder_5_U.u2.cin ;
wire \add_17ns_17ns_17_2_1_U10.top_add_17ns_17ns_17_2_1_Adder_5_U.u2.cout ;
wire [8:0] \add_17ns_17ns_17_2_1_U10.top_add_17ns_17ns_17_2_1_Adder_5_U.u2.s ;
wire \add_19s_19ns_19_2_1_U12.ce ;
wire \add_19s_19ns_19_2_1_U12.clk ;
wire [18:0] \add_19s_19ns_19_2_1_U12.din0 ;
wire [18:0] \add_19s_19ns_19_2_1_U12.din1 ;
wire [18:0] \add_19s_19ns_19_2_1_U12.dout ;
wire \add_19s_19ns_19_2_1_U12.reset ;
wire [18:0] \add_19s_19ns_19_2_1_U12.top_add_19s_19ns_19_2_1_Adder_7_U.a ;
wire [18:0] \add_19s_19ns_19_2_1_U12.top_add_19s_19ns_19_2_1_Adder_7_U.ain_s0 ;
wire [18:0] \add_19s_19ns_19_2_1_U12.top_add_19s_19ns_19_2_1_Adder_7_U.b ;
wire [18:0] \add_19s_19ns_19_2_1_U12.top_add_19s_19ns_19_2_1_Adder_7_U.bin_s0 ;
wire \add_19s_19ns_19_2_1_U12.top_add_19s_19ns_19_2_1_Adder_7_U.ce ;
wire \add_19s_19ns_19_2_1_U12.top_add_19s_19ns_19_2_1_Adder_7_U.clk ;
wire \add_19s_19ns_19_2_1_U12.top_add_19s_19ns_19_2_1_Adder_7_U.facout_s1 ;
wire \add_19s_19ns_19_2_1_U12.top_add_19s_19ns_19_2_1_Adder_7_U.facout_s2 ;
wire [8:0] \add_19s_19ns_19_2_1_U12.top_add_19s_19ns_19_2_1_Adder_7_U.fas_s1 ;
wire [9:0] \add_19s_19ns_19_2_1_U12.top_add_19s_19ns_19_2_1_Adder_7_U.fas_s2 ;
wire \add_19s_19ns_19_2_1_U12.top_add_19s_19ns_19_2_1_Adder_7_U.reset ;
wire [18:0] \add_19s_19ns_19_2_1_U12.top_add_19s_19ns_19_2_1_Adder_7_U.s ;
wire [8:0] \add_19s_19ns_19_2_1_U12.top_add_19s_19ns_19_2_1_Adder_7_U.u1.a ;
wire [8:0] \add_19s_19ns_19_2_1_U12.top_add_19s_19ns_19_2_1_Adder_7_U.u1.b ;
wire \add_19s_19ns_19_2_1_U12.top_add_19s_19ns_19_2_1_Adder_7_U.u1.cin ;
wire \add_19s_19ns_19_2_1_U12.top_add_19s_19ns_19_2_1_Adder_7_U.u1.cout ;
wire [8:0] \add_19s_19ns_19_2_1_U12.top_add_19s_19ns_19_2_1_Adder_7_U.u1.s ;
wire [9:0] \add_19s_19ns_19_2_1_U12.top_add_19s_19ns_19_2_1_Adder_7_U.u2.a ;
wire [9:0] \add_19s_19ns_19_2_1_U12.top_add_19s_19ns_19_2_1_Adder_7_U.u2.b ;
wire \add_19s_19ns_19_2_1_U12.top_add_19s_19ns_19_2_1_Adder_7_U.u2.cin ;
wire \add_19s_19ns_19_2_1_U12.top_add_19s_19ns_19_2_1_Adder_7_U.u2.cout ;
wire [9:0] \add_19s_19ns_19_2_1_U12.top_add_19s_19ns_19_2_1_Adder_7_U.u2.s ;
wire \add_25s_25s_25_2_1_U11.ce ;
wire \add_25s_25s_25_2_1_U11.clk ;
wire [24:0] \add_25s_25s_25_2_1_U11.din0 ;
wire [24:0] \add_25s_25s_25_2_1_U11.din1 ;
wire [24:0] \add_25s_25s_25_2_1_U11.dout ;
wire \add_25s_25s_25_2_1_U11.reset ;
wire [24:0] \add_25s_25s_25_2_1_U11.top_add_25s_25s_25_2_1_Adder_6_U.a ;
wire [24:0] \add_25s_25s_25_2_1_U11.top_add_25s_25s_25_2_1_Adder_6_U.ain_s0 ;
wire [24:0] \add_25s_25s_25_2_1_U11.top_add_25s_25s_25_2_1_Adder_6_U.b ;
wire [24:0] \add_25s_25s_25_2_1_U11.top_add_25s_25s_25_2_1_Adder_6_U.bin_s0 ;
wire \add_25s_25s_25_2_1_U11.top_add_25s_25s_25_2_1_Adder_6_U.ce ;
wire \add_25s_25s_25_2_1_U11.top_add_25s_25s_25_2_1_Adder_6_U.clk ;
wire \add_25s_25s_25_2_1_U11.top_add_25s_25s_25_2_1_Adder_6_U.facout_s1 ;
wire \add_25s_25s_25_2_1_U11.top_add_25s_25s_25_2_1_Adder_6_U.facout_s2 ;
wire [11:0] \add_25s_25s_25_2_1_U11.top_add_25s_25s_25_2_1_Adder_6_U.fas_s1 ;
wire [12:0] \add_25s_25s_25_2_1_U11.top_add_25s_25s_25_2_1_Adder_6_U.fas_s2 ;
wire \add_25s_25s_25_2_1_U11.top_add_25s_25s_25_2_1_Adder_6_U.reset ;
wire [24:0] \add_25s_25s_25_2_1_U11.top_add_25s_25s_25_2_1_Adder_6_U.s ;
wire [11:0] \add_25s_25s_25_2_1_U11.top_add_25s_25s_25_2_1_Adder_6_U.u1.a ;
wire [11:0] \add_25s_25s_25_2_1_U11.top_add_25s_25s_25_2_1_Adder_6_U.u1.b ;
wire \add_25s_25s_25_2_1_U11.top_add_25s_25s_25_2_1_Adder_6_U.u1.cin ;
wire \add_25s_25s_25_2_1_U11.top_add_25s_25s_25_2_1_Adder_6_U.u1.cout ;
wire [11:0] \add_25s_25s_25_2_1_U11.top_add_25s_25s_25_2_1_Adder_6_U.u1.s ;
wire [12:0] \add_25s_25s_25_2_1_U11.top_add_25s_25s_25_2_1_Adder_6_U.u2.a ;
wire [12:0] \add_25s_25s_25_2_1_U11.top_add_25s_25s_25_2_1_Adder_6_U.u2.b ;
wire \add_25s_25s_25_2_1_U11.top_add_25s_25s_25_2_1_Adder_6_U.u2.cin ;
wire \add_25s_25s_25_2_1_U11.top_add_25s_25s_25_2_1_Adder_6_U.u2.cout ;
wire [12:0] \add_25s_25s_25_2_1_U11.top_add_25s_25s_25_2_1_Adder_6_U.u2.s ;
wire \add_2ns_2ns_2_2_1_U5.ce ;
wire \add_2ns_2ns_2_2_1_U5.clk ;
wire [1:0] \add_2ns_2ns_2_2_1_U5.din0 ;
wire [1:0] \add_2ns_2ns_2_2_1_U5.din1 ;
wire [1:0] \add_2ns_2ns_2_2_1_U5.dout ;
wire \add_2ns_2ns_2_2_1_U5.reset ;
wire [1:0] \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_2_U.a ;
wire [1:0] \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_2_U.ain_s0 ;
wire [1:0] \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_2_U.b ;
wire [1:0] \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_2_U.bin_s0 ;
wire \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_2_U.ce ;
wire \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_2_U.clk ;
wire \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_2_U.facout_s1 ;
wire \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_2_U.facout_s2 ;
wire \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_2_U.fas_s1 ;
wire \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_2_U.fas_s2 ;
wire \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_2_U.reset ;
wire [1:0] \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_2_U.s ;
wire \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_2_U.u1.a ;
wire \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_2_U.u1.b ;
wire \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_2_U.u1.cin ;
wire \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_2_U.u1.cout ;
wire \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_2_U.u1.s ;
wire \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_2_U.u2.a ;
wire \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_2_U.u2.b ;
wire \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_2_U.u2.cin ;
wire \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_2_U.u2.cout ;
wire \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_2_U.u2.s ;
wire \add_32ns_32ns_32_2_1_U17.ce ;
wire \add_32ns_32ns_32_2_1_U17.clk ;
wire [31:0] \add_32ns_32ns_32_2_1_U17.din0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U17.din1 ;
wire [31:0] \add_32ns_32ns_32_2_1_U17.dout ;
wire \add_32ns_32ns_32_2_1_U17.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.a ;
wire [31:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.ain_s0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.b ;
wire [31:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.bin_s0 ;
wire \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.ce ;
wire \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.clk ;
wire \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.facout_s1 ;
wire \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.facout_s2 ;
wire [15:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.fas_s1 ;
wire [15:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.fas_s2 ;
wire \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.b ;
wire \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.cin ;
wire \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.b ;
wire \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.cin ;
wire \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.s ;
wire \add_32ns_32ns_32_2_1_U20.ce ;
wire \add_32ns_32ns_32_2_1_U20.clk ;
wire [31:0] \add_32ns_32ns_32_2_1_U20.din0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U20.din1 ;
wire [31:0] \add_32ns_32ns_32_2_1_U20.dout ;
wire \add_32ns_32ns_32_2_1_U20.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.a ;
wire [31:0] \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.ain_s0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.b ;
wire [31:0] \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.bin_s0 ;
wire \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.ce ;
wire \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.clk ;
wire \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.facout_s1 ;
wire \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.facout_s2 ;
wire [15:0] \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.fas_s1 ;
wire [15:0] \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.fas_s2 ;
wire \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.b ;
wire \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.cin ;
wire \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.b ;
wire \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.cin ;
wire \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.s ;
wire \add_32ns_32ns_32_2_1_U21.ce ;
wire \add_32ns_32ns_32_2_1_U21.clk ;
wire [31:0] \add_32ns_32ns_32_2_1_U21.din0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U21.din1 ;
wire [31:0] \add_32ns_32ns_32_2_1_U21.dout ;
wire \add_32ns_32ns_32_2_1_U21.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.a ;
wire [31:0] \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.ain_s0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.b ;
wire [31:0] \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.bin_s0 ;
wire \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.ce ;
wire \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.clk ;
wire \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.facout_s1 ;
wire \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.facout_s2 ;
wire [15:0] \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.fas_s1 ;
wire [15:0] \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.fas_s2 ;
wire \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.b ;
wire \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.cin ;
wire \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.b ;
wire \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.cin ;
wire \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.s ;
wire \add_32s_32ns_32_2_1_U22.ce ;
wire \add_32s_32ns_32_2_1_U22.clk ;
wire [31:0] \add_32s_32ns_32_2_1_U22.din0 ;
wire [31:0] \add_32s_32ns_32_2_1_U22.din1 ;
wire [31:0] \add_32s_32ns_32_2_1_U22.dout ;
wire \add_32s_32ns_32_2_1_U22.reset ;
wire [31:0] \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_14_U.a ;
wire [31:0] \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_14_U.ain_s0 ;
wire [31:0] \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_14_U.b ;
wire [31:0] \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_14_U.bin_s0 ;
wire \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_14_U.ce ;
wire \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_14_U.clk ;
wire \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_14_U.facout_s1 ;
wire \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_14_U.facout_s2 ;
wire [15:0] \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_14_U.fas_s1 ;
wire [15:0] \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_14_U.fas_s2 ;
wire \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_14_U.reset ;
wire [31:0] \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_14_U.s ;
wire [15:0] \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_14_U.u1.a ;
wire [15:0] \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_14_U.u1.b ;
wire \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_14_U.u1.cin ;
wire \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_14_U.u1.cout ;
wire [15:0] \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_14_U.u1.s ;
wire [15:0] \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_14_U.u2.a ;
wire [15:0] \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_14_U.u2.b ;
wire \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_14_U.u2.cin ;
wire \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_14_U.u2.cout ;
wire [15:0] \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_14_U.u2.s ;
wire \add_33ns_33s_33_2_1_U6.ce ;
wire \add_33ns_33s_33_2_1_U6.clk ;
wire [32:0] \add_33ns_33s_33_2_1_U6.din0 ;
wire [32:0] \add_33ns_33s_33_2_1_U6.din1 ;
wire [32:0] \add_33ns_33s_33_2_1_U6.dout ;
wire \add_33ns_33s_33_2_1_U6.reset ;
wire [32:0] \add_33ns_33s_33_2_1_U6.top_add_33ns_33s_33_2_1_Adder_3_U.a ;
wire [32:0] \add_33ns_33s_33_2_1_U6.top_add_33ns_33s_33_2_1_Adder_3_U.ain_s0 ;
wire [32:0] \add_33ns_33s_33_2_1_U6.top_add_33ns_33s_33_2_1_Adder_3_U.b ;
wire [32:0] \add_33ns_33s_33_2_1_U6.top_add_33ns_33s_33_2_1_Adder_3_U.bin_s0 ;
wire \add_33ns_33s_33_2_1_U6.top_add_33ns_33s_33_2_1_Adder_3_U.ce ;
wire \add_33ns_33s_33_2_1_U6.top_add_33ns_33s_33_2_1_Adder_3_U.clk ;
wire \add_33ns_33s_33_2_1_U6.top_add_33ns_33s_33_2_1_Adder_3_U.facout_s1 ;
wire \add_33ns_33s_33_2_1_U6.top_add_33ns_33s_33_2_1_Adder_3_U.facout_s2 ;
wire [15:0] \add_33ns_33s_33_2_1_U6.top_add_33ns_33s_33_2_1_Adder_3_U.fas_s1 ;
wire [16:0] \add_33ns_33s_33_2_1_U6.top_add_33ns_33s_33_2_1_Adder_3_U.fas_s2 ;
wire \add_33ns_33s_33_2_1_U6.top_add_33ns_33s_33_2_1_Adder_3_U.reset ;
wire [32:0] \add_33ns_33s_33_2_1_U6.top_add_33ns_33s_33_2_1_Adder_3_U.s ;
wire [15:0] \add_33ns_33s_33_2_1_U6.top_add_33ns_33s_33_2_1_Adder_3_U.u1.a ;
wire [15:0] \add_33ns_33s_33_2_1_U6.top_add_33ns_33s_33_2_1_Adder_3_U.u1.b ;
wire \add_33ns_33s_33_2_1_U6.top_add_33ns_33s_33_2_1_Adder_3_U.u1.cin ;
wire \add_33ns_33s_33_2_1_U6.top_add_33ns_33s_33_2_1_Adder_3_U.u1.cout ;
wire [15:0] \add_33ns_33s_33_2_1_U6.top_add_33ns_33s_33_2_1_Adder_3_U.u1.s ;
wire [16:0] \add_33ns_33s_33_2_1_U6.top_add_33ns_33s_33_2_1_Adder_3_U.u2.a ;
wire [16:0] \add_33ns_33s_33_2_1_U6.top_add_33ns_33s_33_2_1_Adder_3_U.u2.b ;
wire \add_33ns_33s_33_2_1_U6.top_add_33ns_33s_33_2_1_Adder_3_U.u2.cin ;
wire \add_33ns_33s_33_2_1_U6.top_add_33ns_33s_33_2_1_Adder_3_U.u2.cout ;
wire [16:0] \add_33ns_33s_33_2_1_U6.top_add_33ns_33s_33_2_1_Adder_3_U.u2.s ;
wire \add_35s_35s_35_2_1_U15.ce ;
wire \add_35s_35s_35_2_1_U15.clk ;
wire [34:0] \add_35s_35s_35_2_1_U15.din0 ;
wire [34:0] \add_35s_35s_35_2_1_U15.din1 ;
wire [34:0] \add_35s_35s_35_2_1_U15.dout ;
wire \add_35s_35s_35_2_1_U15.reset ;
wire [34:0] \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.a ;
wire [34:0] \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.ain_s0 ;
wire [34:0] \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.b ;
wire [34:0] \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.bin_s0 ;
wire \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.ce ;
wire \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.clk ;
wire \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.facout_s1 ;
wire \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.facout_s2 ;
wire [16:0] \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.fas_s1 ;
wire [17:0] \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.fas_s2 ;
wire \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.reset ;
wire [34:0] \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.s ;
wire [16:0] \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.u1.a ;
wire [16:0] \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.u1.b ;
wire \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.u1.cin ;
wire \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.u1.cout ;
wire [16:0] \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.u1.s ;
wire [17:0] \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.u2.a ;
wire [17:0] \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.u2.b ;
wire \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.u2.cin ;
wire \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.u2.cout ;
wire [17:0] \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.u2.s ;
wire \add_3s_3ns_3_2_1_U13.ce ;
wire \add_3s_3ns_3_2_1_U13.clk ;
wire [2:0] \add_3s_3ns_3_2_1_U13.din0 ;
wire [2:0] \add_3s_3ns_3_2_1_U13.din1 ;
wire [2:0] \add_3s_3ns_3_2_1_U13.dout ;
wire \add_3s_3ns_3_2_1_U13.reset ;
wire [2:0] \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_8_U.a ;
wire [2:0] \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_8_U.ain_s0 ;
wire [2:0] \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_8_U.b ;
wire [2:0] \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_8_U.bin_s0 ;
wire \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_8_U.ce ;
wire \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_8_U.clk ;
wire \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_8_U.facout_s1 ;
wire \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_8_U.facout_s2 ;
wire \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_8_U.fas_s1 ;
wire [1:0] \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_8_U.fas_s2 ;
wire \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_8_U.reset ;
wire [2:0] \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_8_U.s ;
wire \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_8_U.u1.a ;
wire \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_8_U.u1.b ;
wire \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_8_U.u1.cin ;
wire \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_8_U.u1.cout ;
wire \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_8_U.u1.s ;
wire [1:0] \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_8_U.u2.a ;
wire [1:0] \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_8_U.u2.b ;
wire \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_8_U.u2.cin ;
wire \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_8_U.u2.cout ;
wire [1:0] \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_8_U.u2.s ;
wire \add_46s_46s_46_2_1_U18.ce ;
wire \add_46s_46s_46_2_1_U18.clk ;
wire [45:0] \add_46s_46s_46_2_1_U18.din0 ;
wire [45:0] \add_46s_46s_46_2_1_U18.din1 ;
wire [45:0] \add_46s_46s_46_2_1_U18.dout ;
wire \add_46s_46s_46_2_1_U18.reset ;
wire [45:0] \add_46s_46s_46_2_1_U18.top_add_46s_46s_46_2_1_Adder_12_U.a ;
wire [45:0] \add_46s_46s_46_2_1_U18.top_add_46s_46s_46_2_1_Adder_12_U.ain_s0 ;
wire [45:0] \add_46s_46s_46_2_1_U18.top_add_46s_46s_46_2_1_Adder_12_U.b ;
wire [45:0] \add_46s_46s_46_2_1_U18.top_add_46s_46s_46_2_1_Adder_12_U.bin_s0 ;
wire \add_46s_46s_46_2_1_U18.top_add_46s_46s_46_2_1_Adder_12_U.ce ;
wire \add_46s_46s_46_2_1_U18.top_add_46s_46s_46_2_1_Adder_12_U.clk ;
wire \add_46s_46s_46_2_1_U18.top_add_46s_46s_46_2_1_Adder_12_U.facout_s1 ;
wire \add_46s_46s_46_2_1_U18.top_add_46s_46s_46_2_1_Adder_12_U.facout_s2 ;
wire [22:0] \add_46s_46s_46_2_1_U18.top_add_46s_46s_46_2_1_Adder_12_U.fas_s1 ;
wire [22:0] \add_46s_46s_46_2_1_U18.top_add_46s_46s_46_2_1_Adder_12_U.fas_s2 ;
wire \add_46s_46s_46_2_1_U18.top_add_46s_46s_46_2_1_Adder_12_U.reset ;
wire [45:0] \add_46s_46s_46_2_1_U18.top_add_46s_46s_46_2_1_Adder_12_U.s ;
wire [22:0] \add_46s_46s_46_2_1_U18.top_add_46s_46s_46_2_1_Adder_12_U.u1.a ;
wire [22:0] \add_46s_46s_46_2_1_U18.top_add_46s_46s_46_2_1_Adder_12_U.u1.b ;
wire \add_46s_46s_46_2_1_U18.top_add_46s_46s_46_2_1_Adder_12_U.u1.cin ;
wire \add_46s_46s_46_2_1_U18.top_add_46s_46s_46_2_1_Adder_12_U.u1.cout ;
wire [22:0] \add_46s_46s_46_2_1_U18.top_add_46s_46s_46_2_1_Adder_12_U.u1.s ;
wire [22:0] \add_46s_46s_46_2_1_U18.top_add_46s_46s_46_2_1_Adder_12_U.u2.a ;
wire [22:0] \add_46s_46s_46_2_1_U18.top_add_46s_46s_46_2_1_Adder_12_U.u2.b ;
wire \add_46s_46s_46_2_1_U18.top_add_46s_46s_46_2_1_Adder_12_U.u2.cin ;
wire \add_46s_46s_46_2_1_U18.top_add_46s_46s_46_2_1_Adder_12_U.u2.cout ;
wire [22:0] \add_46s_46s_46_2_1_U18.top_add_46s_46s_46_2_1_Adder_12_U.u2.s ;
wire \add_4ns_4ns_4_2_1_U7.ce ;
wire \add_4ns_4ns_4_2_1_U7.clk ;
wire [3:0] \add_4ns_4ns_4_2_1_U7.din0 ;
wire [3:0] \add_4ns_4ns_4_2_1_U7.din1 ;
wire [3:0] \add_4ns_4ns_4_2_1_U7.dout ;
wire \add_4ns_4ns_4_2_1_U7.reset ;
wire [3:0] \add_4ns_4ns_4_2_1_U7.top_add_4ns_4ns_4_2_1_Adder_4_U.a ;
wire [3:0] \add_4ns_4ns_4_2_1_U7.top_add_4ns_4ns_4_2_1_Adder_4_U.ain_s0 ;
wire [3:0] \add_4ns_4ns_4_2_1_U7.top_add_4ns_4ns_4_2_1_Adder_4_U.b ;
wire [3:0] \add_4ns_4ns_4_2_1_U7.top_add_4ns_4ns_4_2_1_Adder_4_U.bin_s0 ;
wire \add_4ns_4ns_4_2_1_U7.top_add_4ns_4ns_4_2_1_Adder_4_U.ce ;
wire \add_4ns_4ns_4_2_1_U7.top_add_4ns_4ns_4_2_1_Adder_4_U.clk ;
wire \add_4ns_4ns_4_2_1_U7.top_add_4ns_4ns_4_2_1_Adder_4_U.facout_s1 ;
wire \add_4ns_4ns_4_2_1_U7.top_add_4ns_4ns_4_2_1_Adder_4_U.facout_s2 ;
wire [1:0] \add_4ns_4ns_4_2_1_U7.top_add_4ns_4ns_4_2_1_Adder_4_U.fas_s1 ;
wire [1:0] \add_4ns_4ns_4_2_1_U7.top_add_4ns_4ns_4_2_1_Adder_4_U.fas_s2 ;
wire \add_4ns_4ns_4_2_1_U7.top_add_4ns_4ns_4_2_1_Adder_4_U.reset ;
wire [3:0] \add_4ns_4ns_4_2_1_U7.top_add_4ns_4ns_4_2_1_Adder_4_U.s ;
wire [1:0] \add_4ns_4ns_4_2_1_U7.top_add_4ns_4ns_4_2_1_Adder_4_U.u1.a ;
wire [1:0] \add_4ns_4ns_4_2_1_U7.top_add_4ns_4ns_4_2_1_Adder_4_U.u1.b ;
wire \add_4ns_4ns_4_2_1_U7.top_add_4ns_4ns_4_2_1_Adder_4_U.u1.cin ;
wire \add_4ns_4ns_4_2_1_U7.top_add_4ns_4ns_4_2_1_Adder_4_U.u1.cout ;
wire [1:0] \add_4ns_4ns_4_2_1_U7.top_add_4ns_4ns_4_2_1_Adder_4_U.u1.s ;
wire [1:0] \add_4ns_4ns_4_2_1_U7.top_add_4ns_4ns_4_2_1_Adder_4_U.u2.a ;
wire [1:0] \add_4ns_4ns_4_2_1_U7.top_add_4ns_4ns_4_2_1_Adder_4_U.u2.b ;
wire \add_4ns_4ns_4_2_1_U7.top_add_4ns_4ns_4_2_1_Adder_4_U.u2.cin ;
wire \add_4ns_4ns_4_2_1_U7.top_add_4ns_4ns_4_2_1_Adder_4_U.u2.cout ;
wire [1:0] \add_4ns_4ns_4_2_1_U7.top_add_4ns_4ns_4_2_1_Adder_4_U.u2.s ;
wire \add_4ns_4ns_4_2_1_U8.ce ;
wire \add_4ns_4ns_4_2_1_U8.clk ;
wire [3:0] \add_4ns_4ns_4_2_1_U8.din0 ;
wire [3:0] \add_4ns_4ns_4_2_1_U8.din1 ;
wire [3:0] \add_4ns_4ns_4_2_1_U8.dout ;
wire \add_4ns_4ns_4_2_1_U8.reset ;
wire [3:0] \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_4_U.a ;
wire [3:0] \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_4_U.ain_s0 ;
wire [3:0] \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_4_U.b ;
wire [3:0] \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_4_U.bin_s0 ;
wire \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_4_U.ce ;
wire \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_4_U.clk ;
wire \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_4_U.facout_s1 ;
wire \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_4_U.facout_s2 ;
wire [1:0] \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_4_U.fas_s1 ;
wire [1:0] \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_4_U.fas_s2 ;
wire \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_4_U.reset ;
wire [3:0] \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_4_U.s ;
wire [1:0] \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_4_U.u1.a ;
wire [1:0] \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_4_U.u1.b ;
wire \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_4_U.u1.cin ;
wire \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_4_U.u1.cout ;
wire [1:0] \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_4_U.u1.s ;
wire [1:0] \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_4_U.u2.a ;
wire [1:0] \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_4_U.u2.b ;
wire \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_4_U.u2.cin ;
wire \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_4_U.u2.cout ;
wire [1:0] \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_4_U.u2.s ;
wire \add_4ns_4ns_4_2_1_U9.ce ;
wire \add_4ns_4ns_4_2_1_U9.clk ;
wire [3:0] \add_4ns_4ns_4_2_1_U9.din0 ;
wire [3:0] \add_4ns_4ns_4_2_1_U9.din1 ;
wire [3:0] \add_4ns_4ns_4_2_1_U9.dout ;
wire \add_4ns_4ns_4_2_1_U9.reset ;
wire [3:0] \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.a ;
wire [3:0] \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.ain_s0 ;
wire [3:0] \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.b ;
wire [3:0] \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.bin_s0 ;
wire \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.ce ;
wire \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.clk ;
wire \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.facout_s1 ;
wire \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.facout_s2 ;
wire [1:0] \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.fas_s1 ;
wire [1:0] \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.fas_s2 ;
wire \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.reset ;
wire [3:0] \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.s ;
wire [1:0] \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.u1.a ;
wire [1:0] \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.u1.b ;
wire \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.u1.cin ;
wire \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.u1.cout ;
wire [1:0] \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.u1.s ;
wire [1:0] \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.u2.a ;
wire [1:0] \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.u2.b ;
wire \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.u2.cin ;
wire \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.u2.cout ;
wire [1:0] \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.u2.s ;
wire \add_5s_5s_5_2_1_U16.ce ;
wire \add_5s_5s_5_2_1_U16.clk ;
wire [4:0] \add_5s_5s_5_2_1_U16.din0 ;
wire [4:0] \add_5s_5s_5_2_1_U16.din1 ;
wire [4:0] \add_5s_5s_5_2_1_U16.dout ;
wire \add_5s_5s_5_2_1_U16.reset ;
wire [4:0] \add_5s_5s_5_2_1_U16.top_add_5s_5s_5_2_1_Adder_10_U.a ;
wire [4:0] \add_5s_5s_5_2_1_U16.top_add_5s_5s_5_2_1_Adder_10_U.ain_s0 ;
wire [4:0] \add_5s_5s_5_2_1_U16.top_add_5s_5s_5_2_1_Adder_10_U.b ;
wire [4:0] \add_5s_5s_5_2_1_U16.top_add_5s_5s_5_2_1_Adder_10_U.bin_s0 ;
wire \add_5s_5s_5_2_1_U16.top_add_5s_5s_5_2_1_Adder_10_U.ce ;
wire \add_5s_5s_5_2_1_U16.top_add_5s_5s_5_2_1_Adder_10_U.clk ;
wire \add_5s_5s_5_2_1_U16.top_add_5s_5s_5_2_1_Adder_10_U.facout_s1 ;
wire \add_5s_5s_5_2_1_U16.top_add_5s_5s_5_2_1_Adder_10_U.facout_s2 ;
wire [1:0] \add_5s_5s_5_2_1_U16.top_add_5s_5s_5_2_1_Adder_10_U.fas_s1 ;
wire [2:0] \add_5s_5s_5_2_1_U16.top_add_5s_5s_5_2_1_Adder_10_U.fas_s2 ;
wire \add_5s_5s_5_2_1_U16.top_add_5s_5s_5_2_1_Adder_10_U.reset ;
wire [4:0] \add_5s_5s_5_2_1_U16.top_add_5s_5s_5_2_1_Adder_10_U.s ;
wire [1:0] \add_5s_5s_5_2_1_U16.top_add_5s_5s_5_2_1_Adder_10_U.u1.a ;
wire [1:0] \add_5s_5s_5_2_1_U16.top_add_5s_5s_5_2_1_Adder_10_U.u1.b ;
wire \add_5s_5s_5_2_1_U16.top_add_5s_5s_5_2_1_Adder_10_U.u1.cin ;
wire \add_5s_5s_5_2_1_U16.top_add_5s_5s_5_2_1_Adder_10_U.u1.cout ;
wire [1:0] \add_5s_5s_5_2_1_U16.top_add_5s_5s_5_2_1_Adder_10_U.u1.s ;
wire [2:0] \add_5s_5s_5_2_1_U16.top_add_5s_5s_5_2_1_Adder_10_U.u2.a ;
wire [2:0] \add_5s_5s_5_2_1_U16.top_add_5s_5s_5_2_1_Adder_10_U.u2.b ;
wire \add_5s_5s_5_2_1_U16.top_add_5s_5s_5_2_1_Adder_10_U.u2.cin ;
wire \add_5s_5s_5_2_1_U16.top_add_5s_5s_5_2_1_Adder_10_U.u2.cout ;
wire [2:0] \add_5s_5s_5_2_1_U16.top_add_5s_5s_5_2_1_Adder_10_U.u2.s ;
wire \add_6ns_6ns_6_2_1_U19.ce ;
wire \add_6ns_6ns_6_2_1_U19.clk ;
wire [5:0] \add_6ns_6ns_6_2_1_U19.din0 ;
wire [5:0] \add_6ns_6ns_6_2_1_U19.din1 ;
wire [5:0] \add_6ns_6ns_6_2_1_U19.dout ;
wire \add_6ns_6ns_6_2_1_U19.reset ;
wire [5:0] \add_6ns_6ns_6_2_1_U19.top_add_6ns_6ns_6_2_1_Adder_13_U.a ;
wire [5:0] \add_6ns_6ns_6_2_1_U19.top_add_6ns_6ns_6_2_1_Adder_13_U.ain_s0 ;
wire [5:0] \add_6ns_6ns_6_2_1_U19.top_add_6ns_6ns_6_2_1_Adder_13_U.b ;
wire [5:0] \add_6ns_6ns_6_2_1_U19.top_add_6ns_6ns_6_2_1_Adder_13_U.bin_s0 ;
wire \add_6ns_6ns_6_2_1_U19.top_add_6ns_6ns_6_2_1_Adder_13_U.ce ;
wire \add_6ns_6ns_6_2_1_U19.top_add_6ns_6ns_6_2_1_Adder_13_U.clk ;
wire \add_6ns_6ns_6_2_1_U19.top_add_6ns_6ns_6_2_1_Adder_13_U.facout_s1 ;
wire \add_6ns_6ns_6_2_1_U19.top_add_6ns_6ns_6_2_1_Adder_13_U.facout_s2 ;
wire [2:0] \add_6ns_6ns_6_2_1_U19.top_add_6ns_6ns_6_2_1_Adder_13_U.fas_s1 ;
wire [2:0] \add_6ns_6ns_6_2_1_U19.top_add_6ns_6ns_6_2_1_Adder_13_U.fas_s2 ;
wire \add_6ns_6ns_6_2_1_U19.top_add_6ns_6ns_6_2_1_Adder_13_U.reset ;
wire [5:0] \add_6ns_6ns_6_2_1_U19.top_add_6ns_6ns_6_2_1_Adder_13_U.s ;
wire [2:0] \add_6ns_6ns_6_2_1_U19.top_add_6ns_6ns_6_2_1_Adder_13_U.u1.a ;
wire [2:0] \add_6ns_6ns_6_2_1_U19.top_add_6ns_6ns_6_2_1_Adder_13_U.u1.b ;
wire \add_6ns_6ns_6_2_1_U19.top_add_6ns_6ns_6_2_1_Adder_13_U.u1.cin ;
wire \add_6ns_6ns_6_2_1_U19.top_add_6ns_6ns_6_2_1_Adder_13_U.u1.cout ;
wire [2:0] \add_6ns_6ns_6_2_1_U19.top_add_6ns_6ns_6_2_1_Adder_13_U.u1.s ;
wire [2:0] \add_6ns_6ns_6_2_1_U19.top_add_6ns_6ns_6_2_1_Adder_13_U.u2.a ;
wire [2:0] \add_6ns_6ns_6_2_1_U19.top_add_6ns_6ns_6_2_1_Adder_13_U.u2.b ;
wire \add_6ns_6ns_6_2_1_U19.top_add_6ns_6ns_6_2_1_Adder_13_U.u2.cin ;
wire \add_6ns_6ns_6_2_1_U19.top_add_6ns_6ns_6_2_1_Adder_13_U.u2.cout ;
wire [2:0] \add_6ns_6ns_6_2_1_U19.top_add_6ns_6ns_6_2_1_Adder_13_U.u2.s ;
wire and_ln340_1_fu_1133_p2;
wire and_ln340_fu_1056_p2;
wire and_ln406_fu_585_p2;
wire and_ln408_fu_606_p2;
wire and_ln780_1_fu_856_p2;
wire and_ln780_fu_825_p2;
wire and_ln781_1_fu_937_p2;
wire and_ln781_fu_887_p2;
wire and_ln785_1_fu_932_p2;
wire and_ln785_2_fu_1047_p2;
wire and_ln785_4_fu_973_p2;
wire and_ln785_5_fu_982_p2;
wire and_ln785_6_fu_1124_p2;
wire and_ln785_fu_923_p2;
wire and_ln786_1_fu_872_p2;
wire and_ln786_fu_841_p2;
wire ap_CS_fsm_state1;
wire ap_CS_fsm_state10;
wire ap_CS_fsm_state11;
wire ap_CS_fsm_state12;
wire ap_CS_fsm_state13;
wire ap_CS_fsm_state14;
wire ap_CS_fsm_state15;
wire ap_CS_fsm_state16;
wire ap_CS_fsm_state17;
wire ap_CS_fsm_state18;
wire ap_CS_fsm_state19;
wire ap_CS_fsm_state2;
wire ap_CS_fsm_state20;
wire ap_CS_fsm_state21;
wire ap_CS_fsm_state22;
wire ap_CS_fsm_state23;
wire ap_CS_fsm_state24;
wire ap_CS_fsm_state25;
wire ap_CS_fsm_state26;
wire ap_CS_fsm_state27;
wire ap_CS_fsm_state28;
wire ap_CS_fsm_state29;
wire ap_CS_fsm_state30;
wire ap_CS_fsm_state31;
wire ap_CS_fsm_state5;
wire ap_CS_fsm_state6;
wire ap_CS_fsm_state7;
wire ap_CS_fsm_state8;
wire ap_CS_fsm_state9;
wire [30:0] ap_NS_fsm;
wire ap_clk;
wire ap_done;
wire ap_idle;
wire ap_ready;
wire ap_rst;
wire ap_start;
wire carry_1_fu_773_p2;
wire carry_3_fu_777_p2;
wire deleted_ones_1_fu_861_p3;
wire deleted_ones_fu_830_p3;
wire deleted_zeros_1_fu_846_p3;
wire deleted_zeros_fu_815_p3;
wire [2:0] grp_fu_1201_p0;
wire [2:0] grp_fu_1201_p1;
wire [2:0] grp_fu_1201_p2;
wire [3:0] grp_fu_1236_p0;
wire [7:0] grp_fu_1236_p2;
wire [34:0] grp_fu_1255_p0;
wire [34:0] grp_fu_1255_p1;
wire [34:0] grp_fu_1255_p2;
wire [4:0] grp_fu_1282_p0;
wire [4:0] grp_fu_1282_p1;
wire [4:0] grp_fu_1282_p2;
wire [31:0] grp_fu_1288_p2;
wire [45:0] grp_fu_1327_p0;
wire [45:0] grp_fu_1327_p1;
wire [45:0] grp_fu_1327_p2;
wire [5:0] grp_fu_1372_p2;
wire [31:0] grp_fu_1377_p2;
wire [31:0] grp_fu_1427_p1;
wire [31:0] grp_fu_1427_p2;
wire [31:0] grp_fu_1435_p0;
wire [31:0] grp_fu_1435_p2;
wire [2:0] grp_fu_255_p1;
wire [10:0] grp_fu_255_p10;
wire [10:0] grp_fu_255_p2;
wire [7:0] grp_fu_268_p0;
wire [15:0] grp_fu_268_p00;
wire [15:0] grp_fu_268_p2;
wire [32:0] grp_fu_309_p0;
wire [32:0] grp_fu_309_p1;
wire [32:0] grp_fu_309_p2;
wire [6:0] grp_fu_430_p0;
wire [6:0] grp_fu_430_p1;
wire [6:0] grp_fu_430_p2;
wire [1:0] grp_fu_446_p2;
wire [32:0] grp_fu_554_p0;
wire [32:0] grp_fu_554_p1;
wire [32:0] grp_fu_554_p2;
wire [3:0] grp_fu_615_p2;
wire [3:0] grp_fu_652_p1;
wire [3:0] grp_fu_652_p2;
wire [3:0] grp_fu_660_p1;
wire [3:0] grp_fu_660_p2;
wire [16:0] grp_fu_665_p2;
wire [24:0] grp_fu_796_p0;
wire [24:0] grp_fu_796_p1;
wire [24:0] grp_fu_796_p2;
wire [18:0] grp_fu_990_p0;
wire [18:0] grp_fu_990_p2;
wire [31:0] icmp_ln1496_fu_326_p1;
wire icmp_ln1496_fu_326_p2;
wire icmp_ln851_1_fu_610_p2;
wire icmp_ln851_2_fu_1367_p2;
wire icmp_ln851_3_fu_564_p2;
wire icmp_ln851_4_fu_809_p2;
wire icmp_ln851_5_fu_1261_p2;
wire icmp_ln851_6_fu_1337_p2;
wire icmp_ln851_fu_441_p2;
wire icmp_ln874_fu_738_p2;
wire [5:0] lhs_V_2_fu_415_p3;
wire lhs_V_4_fu_436_p2;
wire [16:0] lhs_V_5_fu_539_p3;
wire [5:0] lhs_V_fu_1207_p3;
wire [21:0] lhs_fu_294_p3;
wire \mul_4ns_4s_8_7_1_U14.ce ;
wire \mul_4ns_4s_8_7_1_U14.clk ;
wire [3:0] \mul_4ns_4s_8_7_1_U14.din0 ;
wire [3:0] \mul_4ns_4s_8_7_1_U14.din1 ;
wire [7:0] \mul_4ns_4s_8_7_1_U14.dout ;
wire \mul_4ns_4s_8_7_1_U14.reset ;
wire [3:0] \mul_4ns_4s_8_7_1_U14.top_mul_4ns_4s_8_7_1_Mul_DSP_2_U.a ;
wire [3:0] \mul_4ns_4s_8_7_1_U14.top_mul_4ns_4s_8_7_1_Mul_DSP_2_U.b ;
wire \mul_4ns_4s_8_7_1_U14.top_mul_4ns_4s_8_7_1_Mul_DSP_2_U.ce ;
wire \mul_4ns_4s_8_7_1_U14.top_mul_4ns_4s_8_7_1_Mul_DSP_2_U.clk ;
wire [7:0] \mul_4ns_4s_8_7_1_U14.top_mul_4ns_4s_8_7_1_Mul_DSP_2_U.p ;
wire [7:0] \mul_4ns_4s_8_7_1_U14.top_mul_4ns_4s_8_7_1_Mul_DSP_2_U.tmp_product ;
wire \mul_8ns_8s_16_7_1_U2.ce ;
wire \mul_8ns_8s_16_7_1_U2.clk ;
wire [7:0] \mul_8ns_8s_16_7_1_U2.din0 ;
wire [7:0] \mul_8ns_8s_16_7_1_U2.din1 ;
wire [15:0] \mul_8ns_8s_16_7_1_U2.dout ;
wire \mul_8ns_8s_16_7_1_U2.reset ;
wire [7:0] \mul_8ns_8s_16_7_1_U2.top_mul_8ns_8s_16_7_1_Mul_DSP_1_U.a ;
wire [7:0] \mul_8ns_8s_16_7_1_U2.top_mul_8ns_8s_16_7_1_Mul_DSP_1_U.b ;
wire \mul_8ns_8s_16_7_1_U2.top_mul_8ns_8s_16_7_1_Mul_DSP_1_U.ce ;
wire \mul_8ns_8s_16_7_1_U2.top_mul_8ns_8s_16_7_1_Mul_DSP_1_U.clk ;
wire [15:0] \mul_8ns_8s_16_7_1_U2.top_mul_8ns_8s_16_7_1_Mul_DSP_1_U.p ;
wire [15:0] \mul_8ns_8s_16_7_1_U2.top_mul_8ns_8s_16_7_1_Mul_DSP_1_U.tmp_product ;
wire \mul_8s_3ns_11_7_1_U1.ce ;
wire \mul_8s_3ns_11_7_1_U1.clk ;
wire [7:0] \mul_8s_3ns_11_7_1_U1.din0 ;
wire [2:0] \mul_8s_3ns_11_7_1_U1.din1 ;
wire [10:0] \mul_8s_3ns_11_7_1_U1.dout ;
wire \mul_8s_3ns_11_7_1_U1.reset ;
wire [7:0] \mul_8s_3ns_11_7_1_U1.top_mul_8s_3ns_11_7_1_Mul_DSP_0_U.a ;
wire [2:0] \mul_8s_3ns_11_7_1_U1.top_mul_8s_3ns_11_7_1_Mul_DSP_0_U.b ;
wire \mul_8s_3ns_11_7_1_U1.top_mul_8s_3ns_11_7_1_Mul_DSP_0_U.ce ;
wire \mul_8s_3ns_11_7_1_U1.top_mul_8s_3ns_11_7_1_Mul_DSP_0_U.clk ;
wire [10:0] \mul_8s_3ns_11_7_1_U1.top_mul_8s_3ns_11_7_1_Mul_DSP_0_U.p ;
wire [10:0] \mul_8s_3ns_11_7_1_U1.top_mul_8s_3ns_11_7_1_Mul_DSP_0_U.tmp_product ;
wire neg_src_4_fu_947_p2;
wire neg_src_fu_897_p2;
wire [1:0] op_0;
wire [15:0] op_1;
wire [31:0] op_11;
wire [15:0] op_12_V_fu_766_p3;
wire [3:0] op_14_V_fu_1155_p3;
wire [15:0] op_15;
wire [31:0] op_28;
wire op_28_ap_vld;
wire [7:0] op_4;
wire [3:0] op_5_V_fu_408_p3;
wire [31:0] op_6;
wire [7:0] op_8;
wire [3:0] op_9_V_fu_1166_p3;
wire or_ln340_1_fu_967_p2;
wire or_ln340_2_fu_1036_p2;
wire or_ln340_3_fu_1061_p2;
wire or_ln340_4_fu_1113_p2;
wire or_ln340_5_fu_1138_p2;
wire or_ln340_fu_917_p2;
wire or_ln406_fu_580_p2;
wire or_ln785_1_fu_957_p2;
wire or_ln785_2_fu_927_p2;
wire or_ln785_3_fu_977_p2;
wire or_ln785_fu_907_p2;
wire overflow_1_fu_962_p2;
wire overflow_fu_912_p2;
wire [3:0] p_Result_14_fu_1104_p4;
wire p_Result_15_fu_686_p3;
wire p_Result_16_fu_1382_p3;
wire p_Result_17_fu_743_p3;
wire p_Result_18_fu_1172_p3;
wire p_Result_19_fu_1293_p3;
wire p_Result_20_fu_1401_p3;
wire p_Result_22_fu_570_p3;
wire p_Result_27_fu_505_p2;
wire [6:0] p_Result_5_fu_802_p3;
wire [3:0] p_Result_8_fu_1027_p4;
wire p_Result_s_fu_630_p3;
wire [2:0] p_Val2_4_fu_1022_p2;
wire [2:0] p_Val2_8_fu_1099_p2;
wire r_1_fu_368_p1;
wire r_fu_577_p1;
wire [1:0] ret_V_19_fu_642_p3;
wire [5:0] ret_V_20_fu_1217_p2;
wire [3:0] ret_V_22_fu_698_p3;
wire [5:0] ret_V_23_fu_1394_p3;
wire [31:0] ret_V_28_fu_1413_p3;
wire [12:0] ret_V_3_fu_719_p2;
wire [2:0] ret_fu_239_p3;
wire [23:0] rhs_3_fu_785_p3;
wire [44:0] rhs_4_fu_1316_p3;
wire [11:0] rhs_fu_708_p3;
wire sel_tmp11_fu_1067_p2;
wire sel_tmp25_fu_1144_p2;
wire [3:0] select_ln340_1_fu_1117_p3;
wire [3:0] select_ln340_fu_1040_p3;
wire [31:0] select_ln353_1_fu_1305_p3;
wire [18:0] select_ln353_fu_1184_p3;
wire [3:0] select_ln785_1_fu_1161_p3;
wire [3:0] select_ln785_fu_1150_p3;
wire [3:0] select_ln850_1_fu_693_p3;
wire [5:0] select_ln850_2_fu_1389_p3;
wire [16:0] select_ln850_4_fu_750_p3;
wire [16:0] select_ln850_5_fu_755_p3;
wire [31:0] select_ln850_6_fu_1408_p3;
wire [18:0] select_ln850_7_fu_1179_p3;
wire [31:0] select_ln850_8_fu_1300_p3;
wire [1:0] select_ln850_fu_637_p3;
wire [5:0] sext_ln1194_fu_1214_p1;
wire [15:0] sext_ln69_1_fu_1420_p1;
wire [7:0] sext_ln703_1_fu_705_p0;
wire [12:0] sext_ln703_1_fu_705_p1;
wire [31:0] sext_ln703_2_fu_550_p0;
wire [15:0] sext_ln703_4_fu_1312_p0;
wire [31:0] sext_ln703_fu_305_p0;
wire [18:0] sext_ln850_fu_987_p1;
wire [7:0] shl_ln_fu_315_p3;
wire signbit_fu_288_p2;
wire \sub_33s_33s_33_2_1_U3.ce ;
wire \sub_33s_33s_33_2_1_U3.clk ;
wire [32:0] \sub_33s_33s_33_2_1_U3.din0 ;
wire [32:0] \sub_33s_33s_33_2_1_U3.din1 ;
wire [32:0] \sub_33s_33s_33_2_1_U3.dout ;
wire \sub_33s_33s_33_2_1_U3.reset ;
wire [32:0] \sub_33s_33s_33_2_1_U3.top_sub_33s_33s_33_2_1_Adder_0_U.a ;
wire [32:0] \sub_33s_33s_33_2_1_U3.top_sub_33s_33s_33_2_1_Adder_0_U.ain_s0 ;
wire [32:0] \sub_33s_33s_33_2_1_U3.top_sub_33s_33s_33_2_1_Adder_0_U.b ;
wire [32:0] \sub_33s_33s_33_2_1_U3.top_sub_33s_33s_33_2_1_Adder_0_U.bin_s0 ;
wire \sub_33s_33s_33_2_1_U3.top_sub_33s_33s_33_2_1_Adder_0_U.ce ;
wire \sub_33s_33s_33_2_1_U3.top_sub_33s_33s_33_2_1_Adder_0_U.clk ;
wire \sub_33s_33s_33_2_1_U3.top_sub_33s_33s_33_2_1_Adder_0_U.facout_s1 ;
wire \sub_33s_33s_33_2_1_U3.top_sub_33s_33s_33_2_1_Adder_0_U.facout_s2 ;
wire [15:0] \sub_33s_33s_33_2_1_U3.top_sub_33s_33s_33_2_1_Adder_0_U.fas_s1 ;
wire [16:0] \sub_33s_33s_33_2_1_U3.top_sub_33s_33s_33_2_1_Adder_0_U.fas_s2 ;
wire \sub_33s_33s_33_2_1_U3.top_sub_33s_33s_33_2_1_Adder_0_U.reset ;
wire [32:0] \sub_33s_33s_33_2_1_U3.top_sub_33s_33s_33_2_1_Adder_0_U.s ;
wire [15:0] \sub_33s_33s_33_2_1_U3.top_sub_33s_33s_33_2_1_Adder_0_U.u1.a ;
wire [15:0] \sub_33s_33s_33_2_1_U3.top_sub_33s_33s_33_2_1_Adder_0_U.u1.b ;
wire \sub_33s_33s_33_2_1_U3.top_sub_33s_33s_33_2_1_Adder_0_U.u1.cin ;
wire \sub_33s_33s_33_2_1_U3.top_sub_33s_33s_33_2_1_Adder_0_U.u1.cout ;
wire [15:0] \sub_33s_33s_33_2_1_U3.top_sub_33s_33s_33_2_1_Adder_0_U.u1.s ;
wire [16:0] \sub_33s_33s_33_2_1_U3.top_sub_33s_33s_33_2_1_Adder_0_U.u2.a ;
wire [16:0] \sub_33s_33s_33_2_1_U3.top_sub_33s_33s_33_2_1_Adder_0_U.u2.b ;
wire \sub_33s_33s_33_2_1_U3.top_sub_33s_33s_33_2_1_Adder_0_U.u2.cin ;
wire \sub_33s_33s_33_2_1_U3.top_sub_33s_33s_33_2_1_Adder_0_U.u2.cout ;
wire [16:0] \sub_33s_33s_33_2_1_U3.top_sub_33s_33s_33_2_1_Adder_0_U.u2.s ;
wire \sub_7ns_7ns_7_2_1_U4.ce ;
wire \sub_7ns_7ns_7_2_1_U4.clk ;
wire [6:0] \sub_7ns_7ns_7_2_1_U4.din0 ;
wire [6:0] \sub_7ns_7ns_7_2_1_U4.din1 ;
wire [6:0] \sub_7ns_7ns_7_2_1_U4.dout ;
wire \sub_7ns_7ns_7_2_1_U4.reset ;
wire [6:0] \sub_7ns_7ns_7_2_1_U4.top_sub_7ns_7ns_7_2_1_Adder_1_U.a ;
wire [6:0] \sub_7ns_7ns_7_2_1_U4.top_sub_7ns_7ns_7_2_1_Adder_1_U.ain_s0 ;
wire [6:0] \sub_7ns_7ns_7_2_1_U4.top_sub_7ns_7ns_7_2_1_Adder_1_U.b ;
wire [6:0] \sub_7ns_7ns_7_2_1_U4.top_sub_7ns_7ns_7_2_1_Adder_1_U.bin_s0 ;
wire \sub_7ns_7ns_7_2_1_U4.top_sub_7ns_7ns_7_2_1_Adder_1_U.ce ;
wire \sub_7ns_7ns_7_2_1_U4.top_sub_7ns_7ns_7_2_1_Adder_1_U.clk ;
wire \sub_7ns_7ns_7_2_1_U4.top_sub_7ns_7ns_7_2_1_Adder_1_U.facout_s1 ;
wire \sub_7ns_7ns_7_2_1_U4.top_sub_7ns_7ns_7_2_1_Adder_1_U.facout_s2 ;
wire [2:0] \sub_7ns_7ns_7_2_1_U4.top_sub_7ns_7ns_7_2_1_Adder_1_U.fas_s1 ;
wire [3:0] \sub_7ns_7ns_7_2_1_U4.top_sub_7ns_7ns_7_2_1_Adder_1_U.fas_s2 ;
wire \sub_7ns_7ns_7_2_1_U4.top_sub_7ns_7ns_7_2_1_Adder_1_U.reset ;
wire [6:0] \sub_7ns_7ns_7_2_1_U4.top_sub_7ns_7ns_7_2_1_Adder_1_U.s ;
wire [2:0] \sub_7ns_7ns_7_2_1_U4.top_sub_7ns_7ns_7_2_1_Adder_1_U.u1.a ;
wire [2:0] \sub_7ns_7ns_7_2_1_U4.top_sub_7ns_7ns_7_2_1_Adder_1_U.u1.b ;
wire \sub_7ns_7ns_7_2_1_U4.top_sub_7ns_7ns_7_2_1_Adder_1_U.u1.cin ;
wire \sub_7ns_7ns_7_2_1_U4.top_sub_7ns_7ns_7_2_1_Adder_1_U.u1.cout ;
wire [2:0] \sub_7ns_7ns_7_2_1_U4.top_sub_7ns_7ns_7_2_1_Adder_1_U.u1.s ;
wire [3:0] \sub_7ns_7ns_7_2_1_U4.top_sub_7ns_7ns_7_2_1_Adder_1_U.u2.a ;
wire [3:0] \sub_7ns_7ns_7_2_1_U4.top_sub_7ns_7ns_7_2_1_Adder_1_U.u2.b ;
wire \sub_7ns_7ns_7_2_1_U4.top_sub_7ns_7ns_7_2_1_Adder_1_U.u2.cin ;
wire \sub_7ns_7ns_7_2_1_U4.top_sub_7ns_7ns_7_2_1_Adder_1_U.u2.cout ;
wire [3:0] \sub_7ns_7ns_7_2_1_U4.top_sub_7ns_7ns_7_2_1_Adder_1_U.u2.s ;
wire tmp_10_fu_1073_p3;
wire tmp_11_fu_1080_p3;
wire [14:0] tmp_13_fu_278_p4;
wire [20:0] tmp_18_fu_1244_p3;
wire tmp_4_fu_1003_p3;
wire tmp_fu_996_p3;
wire [1:0] trunc_ln1115_fu_346_p1;
wire [3:0] trunc_ln728_fu_274_p1;
wire [2:0] trunc_ln851_1_fu_535_p1;
wire [1:0] trunc_ln851_2_fu_1353_p1;
wire [31:0] trunc_ln851_3_fu_560_p0;
wire [15:0] trunc_ln851_3_fu_560_p1;
wire [3:0] trunc_ln851_4_fu_762_p1;
wire [1:0] trunc_ln851_5_fu_1191_p1;
wire [15:0] trunc_ln851_6_fu_1333_p0;
wire [12:0] trunc_ln851_6_fu_1333_p1;
wire [6:0] trunc_ln851_fu_342_p1;
wire xor_ln365_1_fu_1016_p2;
wire xor_ln365_2_fu_1087_p2;
wire xor_ln365_3_fu_1093_p2;
wire xor_ln365_fu_1010_p2;
wire xor_ln416_1_fu_730_p2;
wire xor_ln416_fu_725_p2;
wire xor_ln780_1_fu_851_p2;
wire xor_ln780_fu_820_p2;
wire xor_ln781_1_fu_941_p2;
wire xor_ln781_fu_891_p2;
wire xor_ln785_1_fu_836_p2;
wire xor_ln785_2_fu_952_p2;
wire xor_ln785_3_fu_867_p2;
wire xor_ln785_fu_902_p2;
wire xor_ln786_1_fu_1128_p2;
wire xor_ln786_fu_1051_p2;
wire [7:0] zext_ln1116_fu_735_p1;
wire [7:0] zext_ln1116_reg_1819;
wire [12:0] zext_ln1196_fu_715_p1;
wire [31:0] zext_ln1496_fu_322_p1;


assign _103_ = icmp_ln851_5_reg_2023 & ap_CS_fsm[20];
assign _104_ = icmp_ln851_6_reg_2080 & ap_CS_fsm[25];
assign _105_ = icmp_ln851_4_reg_1863 & ap_CS_fsm[15];
assign _106_ = ap_CS_fsm[10] & _111_;
assign _107_ = _112_ & ap_CS_fsm[15];
assign _108_ = _113_ & ap_CS_fsm[15];
assign _109_ = _114_ & ap_CS_fsm[0];
assign _110_ = ap_start & ap_CS_fsm[0];
assign and_ln340_1_fu_1133_p2 = xor_ln786_1_fu_1128_p2 & or_ln340_1_reg_1929;
assign and_ln340_fu_1056_p2 = xor_ln786_fu_1051_p2 & or_ln340_reg_1918;
assign and_ln406_fu_585_p2 = r_V_3_reg_1595[1] & or_ln406_fu_580_p2;
assign and_ln408_fu_606_p2 = r_1_reg_1548 & p_Result_27_reg_1637;
assign and_ln780_1_fu_856_p2 = xor_ln780_1_fu_851_p2 & Range2_all_ones_1_reg_1642;
assign and_ln780_fu_825_p2 = xor_ln780_fu_820_p2 & Range2_all_ones_reg_1701;
assign and_ln781_1_fu_937_p2 = carry_3_reg_1846 & Range1_all_ones_1_reg_1647;
assign and_ln781_fu_887_p2 = carry_1_reg_1839 & Range1_all_ones_reg_1706;
assign and_ln785_1_fu_932_p2 = or_ln785_2_fu_927_p2 & and_ln786_reg_1880;
assign and_ln785_2_fu_1047_p2 = xor_ln785_1_reg_1874 & and_ln786_reg_1880;
assign and_ln785_4_fu_973_p2 = xor_ln416_1_reg_1813 & deleted_zeros_1_reg_1888;
assign and_ln785_5_fu_982_p2 = or_ln785_3_fu_977_p2 & and_ln786_1_reg_1900;
assign and_ln785_6_fu_1124_p2 = xor_ln785_3_reg_1894 & and_ln786_1_reg_1900;
assign and_ln785_fu_923_p2 = xor_ln416_reg_1807 & deleted_zeros_reg_1868;
assign and_ln786_1_fu_872_p2 = p_Result_29_reg_1785 & deleted_ones_1_fu_861_p3;
assign and_ln786_fu_841_p2 = p_Result_24_reg_1769 & deleted_ones_fu_830_p3;
assign carry_1_fu_773_p2 = xor_ln416_reg_1807 & p_Result_23_reg_1615;
assign carry_3_fu_777_p2 = xor_ln416_1_reg_1813 & p_Result_28_reg_1553;
assign neg_src_4_fu_947_p2 = xor_ln781_1_fu_941_p2 & p_Result_26_reg_1536;
assign neg_src_fu_897_p2 = xor_ln781_fu_891_p2 & p_Result_21_reg_1602;
assign overflow_1_fu_962_p2 = xor_ln785_3_reg_1894 & or_ln785_1_fu_957_p2;
assign overflow_fu_912_p2 = xor_ln785_1_reg_1874 & or_ln785_fu_907_p2;
assign ret_V_20_fu_1217_p2 = { op_9_V_reg_1977[3], op_9_V_reg_1977[3], op_9_V_reg_1977 } & { trunc_ln728_reg_1478, 2'h0 };
assign sel_tmp11_fu_1067_p2 = xor_ln365_1_fu_1016_p2 & or_ln340_3_fu_1061_p2;
assign sel_tmp25_fu_1144_p2 = xor_ln365_3_fu_1093_p2 & or_ln340_5_fu_1138_p2;
assign xor_ln786_1_fu_1128_p2 = ~ and_ln786_1_reg_1900;
assign xor_ln786_fu_1051_p2 = ~ and_ln786_reg_1880;
assign xor_ln780_1_fu_851_p2 = ~ p_Result_30_reg_1558;
assign xor_ln780_fu_820_p2 = ~ p_Result_25_reg_1620;
assign lhs_V_4_fu_436_p2 = ~ icmp_ln1496_reg_1504;
assign xor_ln781_1_fu_941_p2 = ~ and_ln781_1_fu_937_p2;
assign xor_ln781_fu_891_p2 = ~ and_ln781_fu_887_p2;
assign xor_ln785_2_fu_952_p2 = ~ deleted_zeros_1_reg_1888;
assign xor_ln785_fu_902_p2 = ~ deleted_zeros_reg_1868;
assign xor_ln365_1_fu_1016_p2 = ~ xor_ln365_fu_1010_p2;
assign xor_ln365_3_fu_1093_p2 = ~ xor_ln365_2_fu_1087_p2;
assign xor_ln416_1_fu_730_p2 = ~ p_Result_29_reg_1785;
assign xor_ln416_fu_725_p2 = ~ p_Result_24_reg_1769;
assign xor_ln785_1_fu_836_p2 = ~ p_Result_21_reg_1602;
assign xor_ln785_3_fu_867_p2 = ~ p_Result_26_reg_1536;
assign p_Val2_4_fu_1022_p2 = ~ p_Val2_3_reg_1760[2:0];
assign p_Val2_8_fu_1099_p2 = ~ p_Val2_7_reg_1776[2:0];
assign _111_ = ~ icmp_ln851_3_reg_1686;
assign _112_ = ~ and_ln785_5_reg_1935;
assign _113_ = ~ and_ln785_1_reg_1924;
assign _114_ = ~ ap_start;
assign _115_ = tmp_2_reg_1569 == 5'h1f;
assign _116_ = p_Result_1_reg_1631 == 10'h3ff;
assign _117_ = ! tmp_2_reg_1569;
assign _118_ = ! p_Result_1_reg_1631;
assign _119_ = tmp_1_reg_1564 == 4'hf;
assign _120_ = p_Result_s_22_reg_1626 == 9'h1ff;
assign _121_ = ! trunc_ln851_1_reg_1671;
assign _122_ = ! trunc_ln851_2_reg_2097;
assign _123_ = ! op_11[15:0];
assign _124_ = ! trunc_ln851_reg_1521;
always @(posedge \add_17ns_17ns_17_2_1_U10.top_add_17ns_17ns_17_2_1_Adder_5_U.clk )
\add_17ns_17ns_17_2_1_U10.top_add_17ns_17ns_17_2_1_Adder_5_U.bin_s1  <= _126_;
always @(posedge \add_17ns_17ns_17_2_1_U10.top_add_17ns_17ns_17_2_1_Adder_5_U.clk )
\add_17ns_17ns_17_2_1_U10.top_add_17ns_17ns_17_2_1_Adder_5_U.ain_s1  <= _125_;
always @(posedge \add_17ns_17ns_17_2_1_U10.top_add_17ns_17ns_17_2_1_Adder_5_U.clk )
\add_17ns_17ns_17_2_1_U10.top_add_17ns_17ns_17_2_1_Adder_5_U.sum_s1  <= _128_;
always @(posedge \add_17ns_17ns_17_2_1_U10.top_add_17ns_17ns_17_2_1_Adder_5_U.clk )
\add_17ns_17ns_17_2_1_U10.top_add_17ns_17ns_17_2_1_Adder_5_U.carry_s1  <= _127_;
assign _126_ = \add_17ns_17ns_17_2_1_U10.top_add_17ns_17ns_17_2_1_Adder_5_U.ce  ? \add_17ns_17ns_17_2_1_U10.top_add_17ns_17ns_17_2_1_Adder_5_U.b [16:8] : \add_17ns_17ns_17_2_1_U10.top_add_17ns_17ns_17_2_1_Adder_5_U.bin_s1 ;
assign _125_ = \add_17ns_17ns_17_2_1_U10.top_add_17ns_17ns_17_2_1_Adder_5_U.ce  ? \add_17ns_17ns_17_2_1_U10.top_add_17ns_17ns_17_2_1_Adder_5_U.a [16:8] : \add_17ns_17ns_17_2_1_U10.top_add_17ns_17ns_17_2_1_Adder_5_U.ain_s1 ;
assign _127_ = \add_17ns_17ns_17_2_1_U10.top_add_17ns_17ns_17_2_1_Adder_5_U.ce  ? \add_17ns_17ns_17_2_1_U10.top_add_17ns_17ns_17_2_1_Adder_5_U.facout_s1  : \add_17ns_17ns_17_2_1_U10.top_add_17ns_17ns_17_2_1_Adder_5_U.carry_s1 ;
assign _128_ = \add_17ns_17ns_17_2_1_U10.top_add_17ns_17ns_17_2_1_Adder_5_U.ce  ? \add_17ns_17ns_17_2_1_U10.top_add_17ns_17ns_17_2_1_Adder_5_U.fas_s1  : \add_17ns_17ns_17_2_1_U10.top_add_17ns_17ns_17_2_1_Adder_5_U.sum_s1 ;
assign _129_ = \add_17ns_17ns_17_2_1_U10.top_add_17ns_17ns_17_2_1_Adder_5_U.u1.a  + \add_17ns_17ns_17_2_1_U10.top_add_17ns_17ns_17_2_1_Adder_5_U.u1.b ;
assign { \add_17ns_17ns_17_2_1_U10.top_add_17ns_17ns_17_2_1_Adder_5_U.u1.cout , \add_17ns_17ns_17_2_1_U10.top_add_17ns_17ns_17_2_1_Adder_5_U.u1.s  } = _129_ + \add_17ns_17ns_17_2_1_U10.top_add_17ns_17ns_17_2_1_Adder_5_U.u1.cin ;
assign _130_ = \add_17ns_17ns_17_2_1_U10.top_add_17ns_17ns_17_2_1_Adder_5_U.u2.a  + \add_17ns_17ns_17_2_1_U10.top_add_17ns_17ns_17_2_1_Adder_5_U.u2.b ;
assign { \add_17ns_17ns_17_2_1_U10.top_add_17ns_17ns_17_2_1_Adder_5_U.u2.cout , \add_17ns_17ns_17_2_1_U10.top_add_17ns_17ns_17_2_1_Adder_5_U.u2.s  } = _130_ + \add_17ns_17ns_17_2_1_U10.top_add_17ns_17ns_17_2_1_Adder_5_U.u2.cin ;
always @(posedge \add_19s_19ns_19_2_1_U12.top_add_19s_19ns_19_2_1_Adder_7_U.clk )
\add_19s_19ns_19_2_1_U12.top_add_19s_19ns_19_2_1_Adder_7_U.bin_s1  <= _132_;
always @(posedge \add_19s_19ns_19_2_1_U12.top_add_19s_19ns_19_2_1_Adder_7_U.clk )
\add_19s_19ns_19_2_1_U12.top_add_19s_19ns_19_2_1_Adder_7_U.ain_s1  <= _131_;
always @(posedge \add_19s_19ns_19_2_1_U12.top_add_19s_19ns_19_2_1_Adder_7_U.clk )
\add_19s_19ns_19_2_1_U12.top_add_19s_19ns_19_2_1_Adder_7_U.sum_s1  <= _134_;
always @(posedge \add_19s_19ns_19_2_1_U12.top_add_19s_19ns_19_2_1_Adder_7_U.clk )
\add_19s_19ns_19_2_1_U12.top_add_19s_19ns_19_2_1_Adder_7_U.carry_s1  <= _133_;
assign _132_ = \add_19s_19ns_19_2_1_U12.top_add_19s_19ns_19_2_1_Adder_7_U.ce  ? \add_19s_19ns_19_2_1_U12.top_add_19s_19ns_19_2_1_Adder_7_U.b [18:9] : \add_19s_19ns_19_2_1_U12.top_add_19s_19ns_19_2_1_Adder_7_U.bin_s1 ;
assign _131_ = \add_19s_19ns_19_2_1_U12.top_add_19s_19ns_19_2_1_Adder_7_U.ce  ? \add_19s_19ns_19_2_1_U12.top_add_19s_19ns_19_2_1_Adder_7_U.a [18:9] : \add_19s_19ns_19_2_1_U12.top_add_19s_19ns_19_2_1_Adder_7_U.ain_s1 ;
assign _133_ = \add_19s_19ns_19_2_1_U12.top_add_19s_19ns_19_2_1_Adder_7_U.ce  ? \add_19s_19ns_19_2_1_U12.top_add_19s_19ns_19_2_1_Adder_7_U.facout_s1  : \add_19s_19ns_19_2_1_U12.top_add_19s_19ns_19_2_1_Adder_7_U.carry_s1 ;
assign _134_ = \add_19s_19ns_19_2_1_U12.top_add_19s_19ns_19_2_1_Adder_7_U.ce  ? \add_19s_19ns_19_2_1_U12.top_add_19s_19ns_19_2_1_Adder_7_U.fas_s1  : \add_19s_19ns_19_2_1_U12.top_add_19s_19ns_19_2_1_Adder_7_U.sum_s1 ;
assign _135_ = \add_19s_19ns_19_2_1_U12.top_add_19s_19ns_19_2_1_Adder_7_U.u1.a  + \add_19s_19ns_19_2_1_U12.top_add_19s_19ns_19_2_1_Adder_7_U.u1.b ;
assign { \add_19s_19ns_19_2_1_U12.top_add_19s_19ns_19_2_1_Adder_7_U.u1.cout , \add_19s_19ns_19_2_1_U12.top_add_19s_19ns_19_2_1_Adder_7_U.u1.s  } = _135_ + \add_19s_19ns_19_2_1_U12.top_add_19s_19ns_19_2_1_Adder_7_U.u1.cin ;
assign _136_ = \add_19s_19ns_19_2_1_U12.top_add_19s_19ns_19_2_1_Adder_7_U.u2.a  + \add_19s_19ns_19_2_1_U12.top_add_19s_19ns_19_2_1_Adder_7_U.u2.b ;
assign { \add_19s_19ns_19_2_1_U12.top_add_19s_19ns_19_2_1_Adder_7_U.u2.cout , \add_19s_19ns_19_2_1_U12.top_add_19s_19ns_19_2_1_Adder_7_U.u2.s  } = _136_ + \add_19s_19ns_19_2_1_U12.top_add_19s_19ns_19_2_1_Adder_7_U.u2.cin ;
always @(posedge \add_25s_25s_25_2_1_U11.top_add_25s_25s_25_2_1_Adder_6_U.clk )
\add_25s_25s_25_2_1_U11.top_add_25s_25s_25_2_1_Adder_6_U.bin_s1  <= _138_;
always @(posedge \add_25s_25s_25_2_1_U11.top_add_25s_25s_25_2_1_Adder_6_U.clk )
\add_25s_25s_25_2_1_U11.top_add_25s_25s_25_2_1_Adder_6_U.ain_s1  <= _137_;
always @(posedge \add_25s_25s_25_2_1_U11.top_add_25s_25s_25_2_1_Adder_6_U.clk )
\add_25s_25s_25_2_1_U11.top_add_25s_25s_25_2_1_Adder_6_U.sum_s1  <= _140_;
always @(posedge \add_25s_25s_25_2_1_U11.top_add_25s_25s_25_2_1_Adder_6_U.clk )
\add_25s_25s_25_2_1_U11.top_add_25s_25s_25_2_1_Adder_6_U.carry_s1  <= _139_;
assign _138_ = \add_25s_25s_25_2_1_U11.top_add_25s_25s_25_2_1_Adder_6_U.ce  ? \add_25s_25s_25_2_1_U11.top_add_25s_25s_25_2_1_Adder_6_U.b [24:12] : \add_25s_25s_25_2_1_U11.top_add_25s_25s_25_2_1_Adder_6_U.bin_s1 ;
assign _137_ = \add_25s_25s_25_2_1_U11.top_add_25s_25s_25_2_1_Adder_6_U.ce  ? \add_25s_25s_25_2_1_U11.top_add_25s_25s_25_2_1_Adder_6_U.a [24:12] : \add_25s_25s_25_2_1_U11.top_add_25s_25s_25_2_1_Adder_6_U.ain_s1 ;
assign _139_ = \add_25s_25s_25_2_1_U11.top_add_25s_25s_25_2_1_Adder_6_U.ce  ? \add_25s_25s_25_2_1_U11.top_add_25s_25s_25_2_1_Adder_6_U.facout_s1  : \add_25s_25s_25_2_1_U11.top_add_25s_25s_25_2_1_Adder_6_U.carry_s1 ;
assign _140_ = \add_25s_25s_25_2_1_U11.top_add_25s_25s_25_2_1_Adder_6_U.ce  ? \add_25s_25s_25_2_1_U11.top_add_25s_25s_25_2_1_Adder_6_U.fas_s1  : \add_25s_25s_25_2_1_U11.top_add_25s_25s_25_2_1_Adder_6_U.sum_s1 ;
assign _141_ = \add_25s_25s_25_2_1_U11.top_add_25s_25s_25_2_1_Adder_6_U.u1.a  + \add_25s_25s_25_2_1_U11.top_add_25s_25s_25_2_1_Adder_6_U.u1.b ;
assign { \add_25s_25s_25_2_1_U11.top_add_25s_25s_25_2_1_Adder_6_U.u1.cout , \add_25s_25s_25_2_1_U11.top_add_25s_25s_25_2_1_Adder_6_U.u1.s  } = _141_ + \add_25s_25s_25_2_1_U11.top_add_25s_25s_25_2_1_Adder_6_U.u1.cin ;
assign _142_ = \add_25s_25s_25_2_1_U11.top_add_25s_25s_25_2_1_Adder_6_U.u2.a  + \add_25s_25s_25_2_1_U11.top_add_25s_25s_25_2_1_Adder_6_U.u2.b ;
assign { \add_25s_25s_25_2_1_U11.top_add_25s_25s_25_2_1_Adder_6_U.u2.cout , \add_25s_25s_25_2_1_U11.top_add_25s_25s_25_2_1_Adder_6_U.u2.s  } = _142_ + \add_25s_25s_25_2_1_U11.top_add_25s_25s_25_2_1_Adder_6_U.u2.cin ;
always @(posedge \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_2_U.clk )
\add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_2_U.bin_s1  <= _144_;
always @(posedge \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_2_U.clk )
\add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_2_U.ain_s1  <= _143_;
always @(posedge \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_2_U.clk )
\add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_2_U.sum_s1  <= _146_;
always @(posedge \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_2_U.clk )
\add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_2_U.carry_s1  <= _145_;
assign _144_ = \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_2_U.ce  ? \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_2_U.b [1] : \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_2_U.bin_s1 ;
assign _143_ = \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_2_U.ce  ? \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_2_U.a [1] : \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_2_U.ain_s1 ;
assign _145_ = \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_2_U.ce  ? \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_2_U.facout_s1  : \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_2_U.carry_s1 ;
assign _146_ = \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_2_U.ce  ? \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_2_U.fas_s1  : \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_2_U.sum_s1 ;
assign _147_ = \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_2_U.u1.a  + \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_2_U.u1.b ;
assign { \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_2_U.u1.cout , \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_2_U.u1.s  } = _147_ + \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_2_U.u1.cin ;
assign _148_ = \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_2_U.u2.a  + \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_2_U.u2.b ;
assign { \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_2_U.u2.cout , \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_2_U.u2.s  } = _148_ + \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_2_U.u2.cin ;
always @(posedge \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.clk )
\add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.bin_s1  <= _150_;
always @(posedge \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.clk )
\add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.ain_s1  <= _149_;
always @(posedge \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.clk )
\add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.sum_s1  <= _152_;
always @(posedge \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.clk )
\add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.carry_s1  <= _151_;
assign _150_ = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.ce  ? \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.b [31:16] : \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.bin_s1 ;
assign _149_ = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.ce  ? \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.a [31:16] : \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.ain_s1 ;
assign _151_ = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.ce  ? \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.facout_s1  : \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.carry_s1 ;
assign _152_ = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.ce  ? \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.fas_s1  : \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.sum_s1 ;
assign _153_ = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.a  + \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.b ;
assign { \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.cout , \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.s  } = _153_ + \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.cin ;
assign _154_ = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.a  + \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.b ;
assign { \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.cout , \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.s  } = _154_ + \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.cin ;
always @(posedge \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.clk )
\add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.bin_s1  <= _156_;
always @(posedge \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.clk )
\add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.ain_s1  <= _155_;
always @(posedge \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.clk )
\add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.sum_s1  <= _158_;
always @(posedge \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.clk )
\add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.carry_s1  <= _157_;
assign _156_ = \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.ce  ? \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.b [31:16] : \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.bin_s1 ;
assign _155_ = \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.ce  ? \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.a [31:16] : \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.ain_s1 ;
assign _157_ = \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.ce  ? \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.facout_s1  : \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.carry_s1 ;
assign _158_ = \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.ce  ? \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.fas_s1  : \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.sum_s1 ;
assign _159_ = \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.a  + \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.b ;
assign { \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.cout , \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.s  } = _159_ + \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.cin ;
assign _160_ = \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.a  + \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.b ;
assign { \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.cout , \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.s  } = _160_ + \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.cin ;
always @(posedge \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.clk )
\add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.bin_s1  <= _162_;
always @(posedge \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.clk )
\add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.ain_s1  <= _161_;
always @(posedge \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.clk )
\add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.sum_s1  <= _164_;
always @(posedge \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.clk )
\add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.carry_s1  <= _163_;
assign _162_ = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.ce  ? \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.b [31:16] : \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.bin_s1 ;
assign _161_ = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.ce  ? \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.a [31:16] : \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.ain_s1 ;
assign _163_ = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.ce  ? \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.facout_s1  : \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.carry_s1 ;
assign _164_ = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.ce  ? \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.fas_s1  : \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.sum_s1 ;
assign _165_ = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.a  + \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.b ;
assign { \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.cout , \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.s  } = _165_ + \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.cin ;
assign _166_ = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.a  + \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.b ;
assign { \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.cout , \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.s  } = _166_ + \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.cin ;
always @(posedge \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_14_U.clk )
\add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_14_U.bin_s1  <= _168_;
always @(posedge \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_14_U.clk )
\add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_14_U.ain_s1  <= _167_;
always @(posedge \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_14_U.clk )
\add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_14_U.sum_s1  <= _170_;
always @(posedge \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_14_U.clk )
\add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_14_U.carry_s1  <= _169_;
assign _168_ = \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_14_U.ce  ? \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_14_U.b [31:16] : \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_14_U.bin_s1 ;
assign _167_ = \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_14_U.ce  ? \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_14_U.a [31:16] : \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_14_U.ain_s1 ;
assign _169_ = \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_14_U.ce  ? \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_14_U.facout_s1  : \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_14_U.carry_s1 ;
assign _170_ = \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_14_U.ce  ? \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_14_U.fas_s1  : \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_14_U.sum_s1 ;
assign _171_ = \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_14_U.u1.a  + \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_14_U.u1.b ;
assign { \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_14_U.u1.cout , \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_14_U.u1.s  } = _171_ + \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_14_U.u1.cin ;
assign _172_ = \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_14_U.u2.a  + \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_14_U.u2.b ;
assign { \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_14_U.u2.cout , \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_14_U.u2.s  } = _172_ + \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_14_U.u2.cin ;
always @(posedge \add_33ns_33s_33_2_1_U6.top_add_33ns_33s_33_2_1_Adder_3_U.clk )
\add_33ns_33s_33_2_1_U6.top_add_33ns_33s_33_2_1_Adder_3_U.bin_s1  <= _174_;
always @(posedge \add_33ns_33s_33_2_1_U6.top_add_33ns_33s_33_2_1_Adder_3_U.clk )
\add_33ns_33s_33_2_1_U6.top_add_33ns_33s_33_2_1_Adder_3_U.ain_s1  <= _173_;
always @(posedge \add_33ns_33s_33_2_1_U6.top_add_33ns_33s_33_2_1_Adder_3_U.clk )
\add_33ns_33s_33_2_1_U6.top_add_33ns_33s_33_2_1_Adder_3_U.sum_s1  <= _176_;
always @(posedge \add_33ns_33s_33_2_1_U6.top_add_33ns_33s_33_2_1_Adder_3_U.clk )
\add_33ns_33s_33_2_1_U6.top_add_33ns_33s_33_2_1_Adder_3_U.carry_s1  <= _175_;
assign _174_ = \add_33ns_33s_33_2_1_U6.top_add_33ns_33s_33_2_1_Adder_3_U.ce  ? \add_33ns_33s_33_2_1_U6.top_add_33ns_33s_33_2_1_Adder_3_U.b [32:16] : \add_33ns_33s_33_2_1_U6.top_add_33ns_33s_33_2_1_Adder_3_U.bin_s1 ;
assign _173_ = \add_33ns_33s_33_2_1_U6.top_add_33ns_33s_33_2_1_Adder_3_U.ce  ? \add_33ns_33s_33_2_1_U6.top_add_33ns_33s_33_2_1_Adder_3_U.a [32:16] : \add_33ns_33s_33_2_1_U6.top_add_33ns_33s_33_2_1_Adder_3_U.ain_s1 ;
assign _175_ = \add_33ns_33s_33_2_1_U6.top_add_33ns_33s_33_2_1_Adder_3_U.ce  ? \add_33ns_33s_33_2_1_U6.top_add_33ns_33s_33_2_1_Adder_3_U.facout_s1  : \add_33ns_33s_33_2_1_U6.top_add_33ns_33s_33_2_1_Adder_3_U.carry_s1 ;
assign _176_ = \add_33ns_33s_33_2_1_U6.top_add_33ns_33s_33_2_1_Adder_3_U.ce  ? \add_33ns_33s_33_2_1_U6.top_add_33ns_33s_33_2_1_Adder_3_U.fas_s1  : \add_33ns_33s_33_2_1_U6.top_add_33ns_33s_33_2_1_Adder_3_U.sum_s1 ;
assign _177_ = \add_33ns_33s_33_2_1_U6.top_add_33ns_33s_33_2_1_Adder_3_U.u1.a  + \add_33ns_33s_33_2_1_U6.top_add_33ns_33s_33_2_1_Adder_3_U.u1.b ;
assign { \add_33ns_33s_33_2_1_U6.top_add_33ns_33s_33_2_1_Adder_3_U.u1.cout , \add_33ns_33s_33_2_1_U6.top_add_33ns_33s_33_2_1_Adder_3_U.u1.s  } = _177_ + \add_33ns_33s_33_2_1_U6.top_add_33ns_33s_33_2_1_Adder_3_U.u1.cin ;
assign _178_ = \add_33ns_33s_33_2_1_U6.top_add_33ns_33s_33_2_1_Adder_3_U.u2.a  + \add_33ns_33s_33_2_1_U6.top_add_33ns_33s_33_2_1_Adder_3_U.u2.b ;
assign { \add_33ns_33s_33_2_1_U6.top_add_33ns_33s_33_2_1_Adder_3_U.u2.cout , \add_33ns_33s_33_2_1_U6.top_add_33ns_33s_33_2_1_Adder_3_U.u2.s  } = _178_ + \add_33ns_33s_33_2_1_U6.top_add_33ns_33s_33_2_1_Adder_3_U.u2.cin ;
always @(posedge \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.clk )
\add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.bin_s1  <= _180_;
always @(posedge \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.clk )
\add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.ain_s1  <= _179_;
always @(posedge \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.clk )
\add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.sum_s1  <= _182_;
always @(posedge \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.clk )
\add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.carry_s1  <= _181_;
assign _180_ = \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.ce  ? \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.b [34:17] : \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.bin_s1 ;
assign _179_ = \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.ce  ? \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.a [34:17] : \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.ain_s1 ;
assign _181_ = \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.ce  ? \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.facout_s1  : \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.carry_s1 ;
assign _182_ = \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.ce  ? \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.fas_s1  : \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.sum_s1 ;
assign _183_ = \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.u1.a  + \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.u1.b ;
assign { \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.u1.cout , \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.u1.s  } = _183_ + \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.u1.cin ;
assign _184_ = \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.u2.a  + \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.u2.b ;
assign { \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.u2.cout , \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.u2.s  } = _184_ + \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.u2.cin ;
always @(posedge \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_8_U.clk )
\add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_8_U.bin_s1  <= _186_;
always @(posedge \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_8_U.clk )
\add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_8_U.ain_s1  <= _185_;
always @(posedge \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_8_U.clk )
\add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_8_U.sum_s1  <= _188_;
always @(posedge \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_8_U.clk )
\add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_8_U.carry_s1  <= _187_;
assign _186_ = \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_8_U.ce  ? \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_8_U.b [2:1] : \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_8_U.bin_s1 ;
assign _185_ = \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_8_U.ce  ? \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_8_U.a [2:1] : \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_8_U.ain_s1 ;
assign _187_ = \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_8_U.ce  ? \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_8_U.facout_s1  : \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_8_U.carry_s1 ;
assign _188_ = \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_8_U.ce  ? \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_8_U.fas_s1  : \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_8_U.sum_s1 ;
assign _189_ = \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_8_U.u1.a  + \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_8_U.u1.b ;
assign { \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_8_U.u1.cout , \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_8_U.u1.s  } = _189_ + \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_8_U.u1.cin ;
assign _190_ = \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_8_U.u2.a  + \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_8_U.u2.b ;
assign { \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_8_U.u2.cout , \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_8_U.u2.s  } = _190_ + \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_8_U.u2.cin ;
always @(posedge \add_46s_46s_46_2_1_U18.top_add_46s_46s_46_2_1_Adder_12_U.clk )
\add_46s_46s_46_2_1_U18.top_add_46s_46s_46_2_1_Adder_12_U.bin_s1  <= _192_;
always @(posedge \add_46s_46s_46_2_1_U18.top_add_46s_46s_46_2_1_Adder_12_U.clk )
\add_46s_46s_46_2_1_U18.top_add_46s_46s_46_2_1_Adder_12_U.ain_s1  <= _191_;
always @(posedge \add_46s_46s_46_2_1_U18.top_add_46s_46s_46_2_1_Adder_12_U.clk )
\add_46s_46s_46_2_1_U18.top_add_46s_46s_46_2_1_Adder_12_U.sum_s1  <= _194_;
always @(posedge \add_46s_46s_46_2_1_U18.top_add_46s_46s_46_2_1_Adder_12_U.clk )
\add_46s_46s_46_2_1_U18.top_add_46s_46s_46_2_1_Adder_12_U.carry_s1  <= _193_;
assign _192_ = \add_46s_46s_46_2_1_U18.top_add_46s_46s_46_2_1_Adder_12_U.ce  ? \add_46s_46s_46_2_1_U18.top_add_46s_46s_46_2_1_Adder_12_U.b [45:23] : \add_46s_46s_46_2_1_U18.top_add_46s_46s_46_2_1_Adder_12_U.bin_s1 ;
assign _191_ = \add_46s_46s_46_2_1_U18.top_add_46s_46s_46_2_1_Adder_12_U.ce  ? \add_46s_46s_46_2_1_U18.top_add_46s_46s_46_2_1_Adder_12_U.a [45:23] : \add_46s_46s_46_2_1_U18.top_add_46s_46s_46_2_1_Adder_12_U.ain_s1 ;
assign _193_ = \add_46s_46s_46_2_1_U18.top_add_46s_46s_46_2_1_Adder_12_U.ce  ? \add_46s_46s_46_2_1_U18.top_add_46s_46s_46_2_1_Adder_12_U.facout_s1  : \add_46s_46s_46_2_1_U18.top_add_46s_46s_46_2_1_Adder_12_U.carry_s1 ;
assign _194_ = \add_46s_46s_46_2_1_U18.top_add_46s_46s_46_2_1_Adder_12_U.ce  ? \add_46s_46s_46_2_1_U18.top_add_46s_46s_46_2_1_Adder_12_U.fas_s1  : \add_46s_46s_46_2_1_U18.top_add_46s_46s_46_2_1_Adder_12_U.sum_s1 ;
assign _195_ = \add_46s_46s_46_2_1_U18.top_add_46s_46s_46_2_1_Adder_12_U.u1.a  + \add_46s_46s_46_2_1_U18.top_add_46s_46s_46_2_1_Adder_12_U.u1.b ;
assign { \add_46s_46s_46_2_1_U18.top_add_46s_46s_46_2_1_Adder_12_U.u1.cout , \add_46s_46s_46_2_1_U18.top_add_46s_46s_46_2_1_Adder_12_U.u1.s  } = _195_ + \add_46s_46s_46_2_1_U18.top_add_46s_46s_46_2_1_Adder_12_U.u1.cin ;
assign _196_ = \add_46s_46s_46_2_1_U18.top_add_46s_46s_46_2_1_Adder_12_U.u2.a  + \add_46s_46s_46_2_1_U18.top_add_46s_46s_46_2_1_Adder_12_U.u2.b ;
assign { \add_46s_46s_46_2_1_U18.top_add_46s_46s_46_2_1_Adder_12_U.u2.cout , \add_46s_46s_46_2_1_U18.top_add_46s_46s_46_2_1_Adder_12_U.u2.s  } = _196_ + \add_46s_46s_46_2_1_U18.top_add_46s_46s_46_2_1_Adder_12_U.u2.cin ;
always @(posedge \add_4ns_4ns_4_2_1_U7.top_add_4ns_4ns_4_2_1_Adder_4_U.clk )
\add_4ns_4ns_4_2_1_U7.top_add_4ns_4ns_4_2_1_Adder_4_U.bin_s1  <= _198_;
always @(posedge \add_4ns_4ns_4_2_1_U7.top_add_4ns_4ns_4_2_1_Adder_4_U.clk )
\add_4ns_4ns_4_2_1_U7.top_add_4ns_4ns_4_2_1_Adder_4_U.ain_s1  <= _197_;
always @(posedge \add_4ns_4ns_4_2_1_U7.top_add_4ns_4ns_4_2_1_Adder_4_U.clk )
\add_4ns_4ns_4_2_1_U7.top_add_4ns_4ns_4_2_1_Adder_4_U.sum_s1  <= _200_;
always @(posedge \add_4ns_4ns_4_2_1_U7.top_add_4ns_4ns_4_2_1_Adder_4_U.clk )
\add_4ns_4ns_4_2_1_U7.top_add_4ns_4ns_4_2_1_Adder_4_U.carry_s1  <= _199_;
assign _198_ = \add_4ns_4ns_4_2_1_U7.top_add_4ns_4ns_4_2_1_Adder_4_U.ce  ? \add_4ns_4ns_4_2_1_U7.top_add_4ns_4ns_4_2_1_Adder_4_U.b [3:2] : \add_4ns_4ns_4_2_1_U7.top_add_4ns_4ns_4_2_1_Adder_4_U.bin_s1 ;
assign _197_ = \add_4ns_4ns_4_2_1_U7.top_add_4ns_4ns_4_2_1_Adder_4_U.ce  ? \add_4ns_4ns_4_2_1_U7.top_add_4ns_4ns_4_2_1_Adder_4_U.a [3:2] : \add_4ns_4ns_4_2_1_U7.top_add_4ns_4ns_4_2_1_Adder_4_U.ain_s1 ;
assign _199_ = \add_4ns_4ns_4_2_1_U7.top_add_4ns_4ns_4_2_1_Adder_4_U.ce  ? \add_4ns_4ns_4_2_1_U7.top_add_4ns_4ns_4_2_1_Adder_4_U.facout_s1  : \add_4ns_4ns_4_2_1_U7.top_add_4ns_4ns_4_2_1_Adder_4_U.carry_s1 ;
assign _200_ = \add_4ns_4ns_4_2_1_U7.top_add_4ns_4ns_4_2_1_Adder_4_U.ce  ? \add_4ns_4ns_4_2_1_U7.top_add_4ns_4ns_4_2_1_Adder_4_U.fas_s1  : \add_4ns_4ns_4_2_1_U7.top_add_4ns_4ns_4_2_1_Adder_4_U.sum_s1 ;
assign _201_ = \add_4ns_4ns_4_2_1_U7.top_add_4ns_4ns_4_2_1_Adder_4_U.u1.a  + \add_4ns_4ns_4_2_1_U7.top_add_4ns_4ns_4_2_1_Adder_4_U.u1.b ;
assign { \add_4ns_4ns_4_2_1_U7.top_add_4ns_4ns_4_2_1_Adder_4_U.u1.cout , \add_4ns_4ns_4_2_1_U7.top_add_4ns_4ns_4_2_1_Adder_4_U.u1.s  } = _201_ + \add_4ns_4ns_4_2_1_U7.top_add_4ns_4ns_4_2_1_Adder_4_U.u1.cin ;
assign _202_ = \add_4ns_4ns_4_2_1_U7.top_add_4ns_4ns_4_2_1_Adder_4_U.u2.a  + \add_4ns_4ns_4_2_1_U7.top_add_4ns_4ns_4_2_1_Adder_4_U.u2.b ;
assign { \add_4ns_4ns_4_2_1_U7.top_add_4ns_4ns_4_2_1_Adder_4_U.u2.cout , \add_4ns_4ns_4_2_1_U7.top_add_4ns_4ns_4_2_1_Adder_4_U.u2.s  } = _202_ + \add_4ns_4ns_4_2_1_U7.top_add_4ns_4ns_4_2_1_Adder_4_U.u2.cin ;
always @(posedge \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_4_U.clk )
\add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_4_U.bin_s1  <= _204_;
always @(posedge \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_4_U.clk )
\add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_4_U.ain_s1  <= _203_;
always @(posedge \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_4_U.clk )
\add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_4_U.sum_s1  <= _206_;
always @(posedge \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_4_U.clk )
\add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_4_U.carry_s1  <= _205_;
assign _204_ = \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_4_U.ce  ? \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_4_U.b [3:2] : \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_4_U.bin_s1 ;
assign _203_ = \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_4_U.ce  ? \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_4_U.a [3:2] : \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_4_U.ain_s1 ;
assign _205_ = \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_4_U.ce  ? \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_4_U.facout_s1  : \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_4_U.carry_s1 ;
assign _206_ = \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_4_U.ce  ? \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_4_U.fas_s1  : \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_4_U.sum_s1 ;
assign _207_ = \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_4_U.u1.a  + \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_4_U.u1.b ;
assign { \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_4_U.u1.cout , \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_4_U.u1.s  } = _207_ + \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_4_U.u1.cin ;
assign _208_ = \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_4_U.u2.a  + \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_4_U.u2.b ;
assign { \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_4_U.u2.cout , \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_4_U.u2.s  } = _208_ + \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_4_U.u2.cin ;
always @(posedge \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.clk )
\add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.bin_s1  <= _210_;
always @(posedge \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.clk )
\add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.ain_s1  <= _209_;
always @(posedge \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.clk )
\add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.sum_s1  <= _212_;
always @(posedge \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.clk )
\add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.carry_s1  <= _211_;
assign _210_ = \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.ce  ? \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.b [3:2] : \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.bin_s1 ;
assign _209_ = \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.ce  ? \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.a [3:2] : \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.ain_s1 ;
assign _211_ = \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.ce  ? \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.facout_s1  : \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.carry_s1 ;
assign _212_ = \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.ce  ? \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.fas_s1  : \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.sum_s1 ;
assign _213_ = \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.u1.a  + \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.u1.b ;
assign { \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.u1.cout , \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.u1.s  } = _213_ + \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.u1.cin ;
assign _214_ = \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.u2.a  + \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.u2.b ;
assign { \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.u2.cout , \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.u2.s  } = _214_ + \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.u2.cin ;
always @(posedge \add_5s_5s_5_2_1_U16.top_add_5s_5s_5_2_1_Adder_10_U.clk )
\add_5s_5s_5_2_1_U16.top_add_5s_5s_5_2_1_Adder_10_U.bin_s1  <= _216_;
always @(posedge \add_5s_5s_5_2_1_U16.top_add_5s_5s_5_2_1_Adder_10_U.clk )
\add_5s_5s_5_2_1_U16.top_add_5s_5s_5_2_1_Adder_10_U.ain_s1  <= _215_;
always @(posedge \add_5s_5s_5_2_1_U16.top_add_5s_5s_5_2_1_Adder_10_U.clk )
\add_5s_5s_5_2_1_U16.top_add_5s_5s_5_2_1_Adder_10_U.sum_s1  <= _218_;
always @(posedge \add_5s_5s_5_2_1_U16.top_add_5s_5s_5_2_1_Adder_10_U.clk )
\add_5s_5s_5_2_1_U16.top_add_5s_5s_5_2_1_Adder_10_U.carry_s1  <= _217_;
assign _216_ = \add_5s_5s_5_2_1_U16.top_add_5s_5s_5_2_1_Adder_10_U.ce  ? \add_5s_5s_5_2_1_U16.top_add_5s_5s_5_2_1_Adder_10_U.b [4:2] : \add_5s_5s_5_2_1_U16.top_add_5s_5s_5_2_1_Adder_10_U.bin_s1 ;
assign _215_ = \add_5s_5s_5_2_1_U16.top_add_5s_5s_5_2_1_Adder_10_U.ce  ? \add_5s_5s_5_2_1_U16.top_add_5s_5s_5_2_1_Adder_10_U.a [4:2] : \add_5s_5s_5_2_1_U16.top_add_5s_5s_5_2_1_Adder_10_U.ain_s1 ;
assign _217_ = \add_5s_5s_5_2_1_U16.top_add_5s_5s_5_2_1_Adder_10_U.ce  ? \add_5s_5s_5_2_1_U16.top_add_5s_5s_5_2_1_Adder_10_U.facout_s1  : \add_5s_5s_5_2_1_U16.top_add_5s_5s_5_2_1_Adder_10_U.carry_s1 ;
assign _218_ = \add_5s_5s_5_2_1_U16.top_add_5s_5s_5_2_1_Adder_10_U.ce  ? \add_5s_5s_5_2_1_U16.top_add_5s_5s_5_2_1_Adder_10_U.fas_s1  : \add_5s_5s_5_2_1_U16.top_add_5s_5s_5_2_1_Adder_10_U.sum_s1 ;
assign _219_ = \add_5s_5s_5_2_1_U16.top_add_5s_5s_5_2_1_Adder_10_U.u1.a  + \add_5s_5s_5_2_1_U16.top_add_5s_5s_5_2_1_Adder_10_U.u1.b ;
assign { \add_5s_5s_5_2_1_U16.top_add_5s_5s_5_2_1_Adder_10_U.u1.cout , \add_5s_5s_5_2_1_U16.top_add_5s_5s_5_2_1_Adder_10_U.u1.s  } = _219_ + \add_5s_5s_5_2_1_U16.top_add_5s_5s_5_2_1_Adder_10_U.u1.cin ;
assign _220_ = \add_5s_5s_5_2_1_U16.top_add_5s_5s_5_2_1_Adder_10_U.u2.a  + \add_5s_5s_5_2_1_U16.top_add_5s_5s_5_2_1_Adder_10_U.u2.b ;
assign { \add_5s_5s_5_2_1_U16.top_add_5s_5s_5_2_1_Adder_10_U.u2.cout , \add_5s_5s_5_2_1_U16.top_add_5s_5s_5_2_1_Adder_10_U.u2.s  } = _220_ + \add_5s_5s_5_2_1_U16.top_add_5s_5s_5_2_1_Adder_10_U.u2.cin ;
always @(posedge \add_6ns_6ns_6_2_1_U19.top_add_6ns_6ns_6_2_1_Adder_13_U.clk )
\add_6ns_6ns_6_2_1_U19.top_add_6ns_6ns_6_2_1_Adder_13_U.bin_s1  <= _222_;
always @(posedge \add_6ns_6ns_6_2_1_U19.top_add_6ns_6ns_6_2_1_Adder_13_U.clk )
\add_6ns_6ns_6_2_1_U19.top_add_6ns_6ns_6_2_1_Adder_13_U.ain_s1  <= _221_;
always @(posedge \add_6ns_6ns_6_2_1_U19.top_add_6ns_6ns_6_2_1_Adder_13_U.clk )
\add_6ns_6ns_6_2_1_U19.top_add_6ns_6ns_6_2_1_Adder_13_U.sum_s1  <= _224_;
always @(posedge \add_6ns_6ns_6_2_1_U19.top_add_6ns_6ns_6_2_1_Adder_13_U.clk )
\add_6ns_6ns_6_2_1_U19.top_add_6ns_6ns_6_2_1_Adder_13_U.carry_s1  <= _223_;
assign _222_ = \add_6ns_6ns_6_2_1_U19.top_add_6ns_6ns_6_2_1_Adder_13_U.ce  ? \add_6ns_6ns_6_2_1_U19.top_add_6ns_6ns_6_2_1_Adder_13_U.b [5:3] : \add_6ns_6ns_6_2_1_U19.top_add_6ns_6ns_6_2_1_Adder_13_U.bin_s1 ;
assign _221_ = \add_6ns_6ns_6_2_1_U19.top_add_6ns_6ns_6_2_1_Adder_13_U.ce  ? \add_6ns_6ns_6_2_1_U19.top_add_6ns_6ns_6_2_1_Adder_13_U.a [5:3] : \add_6ns_6ns_6_2_1_U19.top_add_6ns_6ns_6_2_1_Adder_13_U.ain_s1 ;
assign _223_ = \add_6ns_6ns_6_2_1_U19.top_add_6ns_6ns_6_2_1_Adder_13_U.ce  ? \add_6ns_6ns_6_2_1_U19.top_add_6ns_6ns_6_2_1_Adder_13_U.facout_s1  : \add_6ns_6ns_6_2_1_U19.top_add_6ns_6ns_6_2_1_Adder_13_U.carry_s1 ;
assign _224_ = \add_6ns_6ns_6_2_1_U19.top_add_6ns_6ns_6_2_1_Adder_13_U.ce  ? \add_6ns_6ns_6_2_1_U19.top_add_6ns_6ns_6_2_1_Adder_13_U.fas_s1  : \add_6ns_6ns_6_2_1_U19.top_add_6ns_6ns_6_2_1_Adder_13_U.sum_s1 ;
assign _225_ = \add_6ns_6ns_6_2_1_U19.top_add_6ns_6ns_6_2_1_Adder_13_U.u1.a  + \add_6ns_6ns_6_2_1_U19.top_add_6ns_6ns_6_2_1_Adder_13_U.u1.b ;
assign { \add_6ns_6ns_6_2_1_U19.top_add_6ns_6ns_6_2_1_Adder_13_U.u1.cout , \add_6ns_6ns_6_2_1_U19.top_add_6ns_6ns_6_2_1_Adder_13_U.u1.s  } = _225_ + \add_6ns_6ns_6_2_1_U19.top_add_6ns_6ns_6_2_1_Adder_13_U.u1.cin ;
assign _226_ = \add_6ns_6ns_6_2_1_U19.top_add_6ns_6ns_6_2_1_Adder_13_U.u2.a  + \add_6ns_6ns_6_2_1_U19.top_add_6ns_6ns_6_2_1_Adder_13_U.u2.b ;
assign { \add_6ns_6ns_6_2_1_U19.top_add_6ns_6ns_6_2_1_Adder_13_U.u2.cout , \add_6ns_6ns_6_2_1_U19.top_add_6ns_6ns_6_2_1_Adder_13_U.u2.s  } = _226_ + \add_6ns_6ns_6_2_1_U19.top_add_6ns_6ns_6_2_1_Adder_13_U.u2.cin ;
assign \mul_4ns_4s_8_7_1_U14.top_mul_4ns_4s_8_7_1_Mul_DSP_2_U.tmp_product  = $signed({ 1'h0, \mul_4ns_4s_8_7_1_U14.top_mul_4ns_4s_8_7_1_Mul_DSP_2_U.a_reg0  }) * $signed(\mul_4ns_4s_8_7_1_U14.top_mul_4ns_4s_8_7_1_Mul_DSP_2_U.b_reg0 );
always @(posedge \mul_4ns_4s_8_7_1_U14.top_mul_4ns_4s_8_7_1_Mul_DSP_2_U.clk )
\mul_4ns_4s_8_7_1_U14.top_mul_4ns_4s_8_7_1_Mul_DSP_2_U.a_reg0  <= _227_;
always @(posedge \mul_4ns_4s_8_7_1_U14.top_mul_4ns_4s_8_7_1_Mul_DSP_2_U.clk )
\mul_4ns_4s_8_7_1_U14.top_mul_4ns_4s_8_7_1_Mul_DSP_2_U.b_reg0  <= _228_;
always @(posedge \mul_4ns_4s_8_7_1_U14.top_mul_4ns_4s_8_7_1_Mul_DSP_2_U.clk )
\mul_4ns_4s_8_7_1_U14.top_mul_4ns_4s_8_7_1_Mul_DSP_2_U.buff0  <= _229_;
always @(posedge \mul_4ns_4s_8_7_1_U14.top_mul_4ns_4s_8_7_1_Mul_DSP_2_U.clk )
\mul_4ns_4s_8_7_1_U14.top_mul_4ns_4s_8_7_1_Mul_DSP_2_U.buff1  <= _230_;
always @(posedge \mul_4ns_4s_8_7_1_U14.top_mul_4ns_4s_8_7_1_Mul_DSP_2_U.clk )
\mul_4ns_4s_8_7_1_U14.top_mul_4ns_4s_8_7_1_Mul_DSP_2_U.buff2  <= _231_;
always @(posedge \mul_4ns_4s_8_7_1_U14.top_mul_4ns_4s_8_7_1_Mul_DSP_2_U.clk )
\mul_4ns_4s_8_7_1_U14.top_mul_4ns_4s_8_7_1_Mul_DSP_2_U.buff3  <= _232_;
always @(posedge \mul_4ns_4s_8_7_1_U14.top_mul_4ns_4s_8_7_1_Mul_DSP_2_U.clk )
\mul_4ns_4s_8_7_1_U14.top_mul_4ns_4s_8_7_1_Mul_DSP_2_U.buff4  <= _233_;
assign _233_ = \mul_4ns_4s_8_7_1_U14.top_mul_4ns_4s_8_7_1_Mul_DSP_2_U.ce  ? \mul_4ns_4s_8_7_1_U14.top_mul_4ns_4s_8_7_1_Mul_DSP_2_U.buff3  : \mul_4ns_4s_8_7_1_U14.top_mul_4ns_4s_8_7_1_Mul_DSP_2_U.buff4 ;
assign _232_ = \mul_4ns_4s_8_7_1_U14.top_mul_4ns_4s_8_7_1_Mul_DSP_2_U.ce  ? \mul_4ns_4s_8_7_1_U14.top_mul_4ns_4s_8_7_1_Mul_DSP_2_U.buff2  : \mul_4ns_4s_8_7_1_U14.top_mul_4ns_4s_8_7_1_Mul_DSP_2_U.buff3 ;
assign _231_ = \mul_4ns_4s_8_7_1_U14.top_mul_4ns_4s_8_7_1_Mul_DSP_2_U.ce  ? \mul_4ns_4s_8_7_1_U14.top_mul_4ns_4s_8_7_1_Mul_DSP_2_U.buff1  : \mul_4ns_4s_8_7_1_U14.top_mul_4ns_4s_8_7_1_Mul_DSP_2_U.buff2 ;
assign _230_ = \mul_4ns_4s_8_7_1_U14.top_mul_4ns_4s_8_7_1_Mul_DSP_2_U.ce  ? \mul_4ns_4s_8_7_1_U14.top_mul_4ns_4s_8_7_1_Mul_DSP_2_U.buff0  : \mul_4ns_4s_8_7_1_U14.top_mul_4ns_4s_8_7_1_Mul_DSP_2_U.buff1 ;
assign _229_ = \mul_4ns_4s_8_7_1_U14.top_mul_4ns_4s_8_7_1_Mul_DSP_2_U.ce  ? \mul_4ns_4s_8_7_1_U14.top_mul_4ns_4s_8_7_1_Mul_DSP_2_U.tmp_product  : \mul_4ns_4s_8_7_1_U14.top_mul_4ns_4s_8_7_1_Mul_DSP_2_U.buff0 ;
assign _228_ = \mul_4ns_4s_8_7_1_U14.top_mul_4ns_4s_8_7_1_Mul_DSP_2_U.ce  ? \mul_4ns_4s_8_7_1_U14.top_mul_4ns_4s_8_7_1_Mul_DSP_2_U.b  : \mul_4ns_4s_8_7_1_U14.top_mul_4ns_4s_8_7_1_Mul_DSP_2_U.b_reg0 ;
assign _227_ = \mul_4ns_4s_8_7_1_U14.top_mul_4ns_4s_8_7_1_Mul_DSP_2_U.ce  ? \mul_4ns_4s_8_7_1_U14.top_mul_4ns_4s_8_7_1_Mul_DSP_2_U.a  : \mul_4ns_4s_8_7_1_U14.top_mul_4ns_4s_8_7_1_Mul_DSP_2_U.a_reg0 ;
assign \mul_8ns_8s_16_7_1_U2.top_mul_8ns_8s_16_7_1_Mul_DSP_1_U.tmp_product  = $signed({ 1'h0, \mul_8ns_8s_16_7_1_U2.top_mul_8ns_8s_16_7_1_Mul_DSP_1_U.a_reg0  }) * $signed(\mul_8ns_8s_16_7_1_U2.top_mul_8ns_8s_16_7_1_Mul_DSP_1_U.b_reg0 );
always @(posedge \mul_8ns_8s_16_7_1_U2.top_mul_8ns_8s_16_7_1_Mul_DSP_1_U.clk )
\mul_8ns_8s_16_7_1_U2.top_mul_8ns_8s_16_7_1_Mul_DSP_1_U.a_reg0  <= _234_;
always @(posedge \mul_8ns_8s_16_7_1_U2.top_mul_8ns_8s_16_7_1_Mul_DSP_1_U.clk )
\mul_8ns_8s_16_7_1_U2.top_mul_8ns_8s_16_7_1_Mul_DSP_1_U.b_reg0  <= _235_;
always @(posedge \mul_8ns_8s_16_7_1_U2.top_mul_8ns_8s_16_7_1_Mul_DSP_1_U.clk )
\mul_8ns_8s_16_7_1_U2.top_mul_8ns_8s_16_7_1_Mul_DSP_1_U.buff0  <= _236_;
always @(posedge \mul_8ns_8s_16_7_1_U2.top_mul_8ns_8s_16_7_1_Mul_DSP_1_U.clk )
\mul_8ns_8s_16_7_1_U2.top_mul_8ns_8s_16_7_1_Mul_DSP_1_U.buff1  <= _237_;
always @(posedge \mul_8ns_8s_16_7_1_U2.top_mul_8ns_8s_16_7_1_Mul_DSP_1_U.clk )
\mul_8ns_8s_16_7_1_U2.top_mul_8ns_8s_16_7_1_Mul_DSP_1_U.buff2  <= _238_;
always @(posedge \mul_8ns_8s_16_7_1_U2.top_mul_8ns_8s_16_7_1_Mul_DSP_1_U.clk )
\mul_8ns_8s_16_7_1_U2.top_mul_8ns_8s_16_7_1_Mul_DSP_1_U.buff3  <= _239_;
always @(posedge \mul_8ns_8s_16_7_1_U2.top_mul_8ns_8s_16_7_1_Mul_DSP_1_U.clk )
\mul_8ns_8s_16_7_1_U2.top_mul_8ns_8s_16_7_1_Mul_DSP_1_U.buff4  <= _240_;
assign _240_ = \mul_8ns_8s_16_7_1_U2.top_mul_8ns_8s_16_7_1_Mul_DSP_1_U.ce  ? \mul_8ns_8s_16_7_1_U2.top_mul_8ns_8s_16_7_1_Mul_DSP_1_U.buff3  : \mul_8ns_8s_16_7_1_U2.top_mul_8ns_8s_16_7_1_Mul_DSP_1_U.buff4 ;
assign _239_ = \mul_8ns_8s_16_7_1_U2.top_mul_8ns_8s_16_7_1_Mul_DSP_1_U.ce  ? \mul_8ns_8s_16_7_1_U2.top_mul_8ns_8s_16_7_1_Mul_DSP_1_U.buff2  : \mul_8ns_8s_16_7_1_U2.top_mul_8ns_8s_16_7_1_Mul_DSP_1_U.buff3 ;
assign _238_ = \mul_8ns_8s_16_7_1_U2.top_mul_8ns_8s_16_7_1_Mul_DSP_1_U.ce  ? \mul_8ns_8s_16_7_1_U2.top_mul_8ns_8s_16_7_1_Mul_DSP_1_U.buff1  : \mul_8ns_8s_16_7_1_U2.top_mul_8ns_8s_16_7_1_Mul_DSP_1_U.buff2 ;
assign _237_ = \mul_8ns_8s_16_7_1_U2.top_mul_8ns_8s_16_7_1_Mul_DSP_1_U.ce  ? \mul_8ns_8s_16_7_1_U2.top_mul_8ns_8s_16_7_1_Mul_DSP_1_U.buff0  : \mul_8ns_8s_16_7_1_U2.top_mul_8ns_8s_16_7_1_Mul_DSP_1_U.buff1 ;
assign _236_ = \mul_8ns_8s_16_7_1_U2.top_mul_8ns_8s_16_7_1_Mul_DSP_1_U.ce  ? \mul_8ns_8s_16_7_1_U2.top_mul_8ns_8s_16_7_1_Mul_DSP_1_U.tmp_product  : \mul_8ns_8s_16_7_1_U2.top_mul_8ns_8s_16_7_1_Mul_DSP_1_U.buff0 ;
assign _235_ = \mul_8ns_8s_16_7_1_U2.top_mul_8ns_8s_16_7_1_Mul_DSP_1_U.ce  ? \mul_8ns_8s_16_7_1_U2.top_mul_8ns_8s_16_7_1_Mul_DSP_1_U.b  : \mul_8ns_8s_16_7_1_U2.top_mul_8ns_8s_16_7_1_Mul_DSP_1_U.b_reg0 ;
assign _234_ = \mul_8ns_8s_16_7_1_U2.top_mul_8ns_8s_16_7_1_Mul_DSP_1_U.ce  ? \mul_8ns_8s_16_7_1_U2.top_mul_8ns_8s_16_7_1_Mul_DSP_1_U.a  : \mul_8ns_8s_16_7_1_U2.top_mul_8ns_8s_16_7_1_Mul_DSP_1_U.a_reg0 ;
assign \mul_8s_3ns_11_7_1_U1.top_mul_8s_3ns_11_7_1_Mul_DSP_0_U.tmp_product  = $signed(\mul_8s_3ns_11_7_1_U1.top_mul_8s_3ns_11_7_1_Mul_DSP_0_U.a_reg0 ) * $signed({ 1'h0, \mul_8s_3ns_11_7_1_U1.top_mul_8s_3ns_11_7_1_Mul_DSP_0_U.b_reg0  });
always @(posedge \mul_8s_3ns_11_7_1_U1.top_mul_8s_3ns_11_7_1_Mul_DSP_0_U.clk )
\mul_8s_3ns_11_7_1_U1.top_mul_8s_3ns_11_7_1_Mul_DSP_0_U.a_reg0  <= _241_;
always @(posedge \mul_8s_3ns_11_7_1_U1.top_mul_8s_3ns_11_7_1_Mul_DSP_0_U.clk )
\mul_8s_3ns_11_7_1_U1.top_mul_8s_3ns_11_7_1_Mul_DSP_0_U.b_reg0  <= _242_;
always @(posedge \mul_8s_3ns_11_7_1_U1.top_mul_8s_3ns_11_7_1_Mul_DSP_0_U.clk )
\mul_8s_3ns_11_7_1_U1.top_mul_8s_3ns_11_7_1_Mul_DSP_0_U.buff0  <= _243_;
always @(posedge \mul_8s_3ns_11_7_1_U1.top_mul_8s_3ns_11_7_1_Mul_DSP_0_U.clk )
\mul_8s_3ns_11_7_1_U1.top_mul_8s_3ns_11_7_1_Mul_DSP_0_U.buff1  <= _244_;
always @(posedge \mul_8s_3ns_11_7_1_U1.top_mul_8s_3ns_11_7_1_Mul_DSP_0_U.clk )
\mul_8s_3ns_11_7_1_U1.top_mul_8s_3ns_11_7_1_Mul_DSP_0_U.buff2  <= _245_;
always @(posedge \mul_8s_3ns_11_7_1_U1.top_mul_8s_3ns_11_7_1_Mul_DSP_0_U.clk )
\mul_8s_3ns_11_7_1_U1.top_mul_8s_3ns_11_7_1_Mul_DSP_0_U.buff3  <= _246_;
always @(posedge \mul_8s_3ns_11_7_1_U1.top_mul_8s_3ns_11_7_1_Mul_DSP_0_U.clk )
\mul_8s_3ns_11_7_1_U1.top_mul_8s_3ns_11_7_1_Mul_DSP_0_U.buff4  <= _247_;
assign _247_ = \mul_8s_3ns_11_7_1_U1.top_mul_8s_3ns_11_7_1_Mul_DSP_0_U.ce  ? \mul_8s_3ns_11_7_1_U1.top_mul_8s_3ns_11_7_1_Mul_DSP_0_U.buff3  : \mul_8s_3ns_11_7_1_U1.top_mul_8s_3ns_11_7_1_Mul_DSP_0_U.buff4 ;
assign _246_ = \mul_8s_3ns_11_7_1_U1.top_mul_8s_3ns_11_7_1_Mul_DSP_0_U.ce  ? \mul_8s_3ns_11_7_1_U1.top_mul_8s_3ns_11_7_1_Mul_DSP_0_U.buff2  : \mul_8s_3ns_11_7_1_U1.top_mul_8s_3ns_11_7_1_Mul_DSP_0_U.buff3 ;
assign _245_ = \mul_8s_3ns_11_7_1_U1.top_mul_8s_3ns_11_7_1_Mul_DSP_0_U.ce  ? \mul_8s_3ns_11_7_1_U1.top_mul_8s_3ns_11_7_1_Mul_DSP_0_U.buff1  : \mul_8s_3ns_11_7_1_U1.top_mul_8s_3ns_11_7_1_Mul_DSP_0_U.buff2 ;
assign _244_ = \mul_8s_3ns_11_7_1_U1.top_mul_8s_3ns_11_7_1_Mul_DSP_0_U.ce  ? \mul_8s_3ns_11_7_1_U1.top_mul_8s_3ns_11_7_1_Mul_DSP_0_U.buff0  : \mul_8s_3ns_11_7_1_U1.top_mul_8s_3ns_11_7_1_Mul_DSP_0_U.buff1 ;
assign _243_ = \mul_8s_3ns_11_7_1_U1.top_mul_8s_3ns_11_7_1_Mul_DSP_0_U.ce  ? \mul_8s_3ns_11_7_1_U1.top_mul_8s_3ns_11_7_1_Mul_DSP_0_U.tmp_product  : \mul_8s_3ns_11_7_1_U1.top_mul_8s_3ns_11_7_1_Mul_DSP_0_U.buff0 ;
assign _242_ = \mul_8s_3ns_11_7_1_U1.top_mul_8s_3ns_11_7_1_Mul_DSP_0_U.ce  ? \mul_8s_3ns_11_7_1_U1.top_mul_8s_3ns_11_7_1_Mul_DSP_0_U.b  : \mul_8s_3ns_11_7_1_U1.top_mul_8s_3ns_11_7_1_Mul_DSP_0_U.b_reg0 ;
assign _241_ = \mul_8s_3ns_11_7_1_U1.top_mul_8s_3ns_11_7_1_Mul_DSP_0_U.ce  ? \mul_8s_3ns_11_7_1_U1.top_mul_8s_3ns_11_7_1_Mul_DSP_0_U.a  : \mul_8s_3ns_11_7_1_U1.top_mul_8s_3ns_11_7_1_Mul_DSP_0_U.a_reg0 ;
assign \sub_33s_33s_33_2_1_U3.top_sub_33s_33s_33_2_1_Adder_0_U.bin_s0  = ~ \sub_33s_33s_33_2_1_U3.top_sub_33s_33s_33_2_1_Adder_0_U.b ;
always @(posedge \sub_33s_33s_33_2_1_U3.top_sub_33s_33s_33_2_1_Adder_0_U.clk )
\sub_33s_33s_33_2_1_U3.top_sub_33s_33s_33_2_1_Adder_0_U.bin_s1  <= _249_;
always @(posedge \sub_33s_33s_33_2_1_U3.top_sub_33s_33s_33_2_1_Adder_0_U.clk )
\sub_33s_33s_33_2_1_U3.top_sub_33s_33s_33_2_1_Adder_0_U.ain_s1  <= _248_;
always @(posedge \sub_33s_33s_33_2_1_U3.top_sub_33s_33s_33_2_1_Adder_0_U.clk )
\sub_33s_33s_33_2_1_U3.top_sub_33s_33s_33_2_1_Adder_0_U.sum_s1  <= _251_;
always @(posedge \sub_33s_33s_33_2_1_U3.top_sub_33s_33s_33_2_1_Adder_0_U.clk )
\sub_33s_33s_33_2_1_U3.top_sub_33s_33s_33_2_1_Adder_0_U.carry_s1  <= _250_;
assign _249_ = \sub_33s_33s_33_2_1_U3.top_sub_33s_33s_33_2_1_Adder_0_U.ce  ? \sub_33s_33s_33_2_1_U3.top_sub_33s_33s_33_2_1_Adder_0_U.bin_s0 [32:16] : \sub_33s_33s_33_2_1_U3.top_sub_33s_33s_33_2_1_Adder_0_U.bin_s1 ;
assign _248_ = \sub_33s_33s_33_2_1_U3.top_sub_33s_33s_33_2_1_Adder_0_U.ce  ? \sub_33s_33s_33_2_1_U3.top_sub_33s_33s_33_2_1_Adder_0_U.a [32:16] : \sub_33s_33s_33_2_1_U3.top_sub_33s_33s_33_2_1_Adder_0_U.ain_s1 ;
assign _250_ = \sub_33s_33s_33_2_1_U3.top_sub_33s_33s_33_2_1_Adder_0_U.ce  ? \sub_33s_33s_33_2_1_U3.top_sub_33s_33s_33_2_1_Adder_0_U.facout_s1  : \sub_33s_33s_33_2_1_U3.top_sub_33s_33s_33_2_1_Adder_0_U.carry_s1 ;
assign _251_ = \sub_33s_33s_33_2_1_U3.top_sub_33s_33s_33_2_1_Adder_0_U.ce  ? \sub_33s_33s_33_2_1_U3.top_sub_33s_33s_33_2_1_Adder_0_U.fas_s1  : \sub_33s_33s_33_2_1_U3.top_sub_33s_33s_33_2_1_Adder_0_U.sum_s1 ;
assign _252_ = \sub_33s_33s_33_2_1_U3.top_sub_33s_33s_33_2_1_Adder_0_U.u1.a  + \sub_33s_33s_33_2_1_U3.top_sub_33s_33s_33_2_1_Adder_0_U.u1.b ;
assign { \sub_33s_33s_33_2_1_U3.top_sub_33s_33s_33_2_1_Adder_0_U.u1.cout , \sub_33s_33s_33_2_1_U3.top_sub_33s_33s_33_2_1_Adder_0_U.u1.s  } = _252_ + \sub_33s_33s_33_2_1_U3.top_sub_33s_33s_33_2_1_Adder_0_U.u1.cin ;
assign _253_ = \sub_33s_33s_33_2_1_U3.top_sub_33s_33s_33_2_1_Adder_0_U.u2.a  + \sub_33s_33s_33_2_1_U3.top_sub_33s_33s_33_2_1_Adder_0_U.u2.b ;
assign { \sub_33s_33s_33_2_1_U3.top_sub_33s_33s_33_2_1_Adder_0_U.u2.cout , \sub_33s_33s_33_2_1_U3.top_sub_33s_33s_33_2_1_Adder_0_U.u2.s  } = _253_ + \sub_33s_33s_33_2_1_U3.top_sub_33s_33s_33_2_1_Adder_0_U.u2.cin ;
assign \sub_7ns_7ns_7_2_1_U4.top_sub_7ns_7ns_7_2_1_Adder_1_U.bin_s0  = ~ \sub_7ns_7ns_7_2_1_U4.top_sub_7ns_7ns_7_2_1_Adder_1_U.b ;
always @(posedge \sub_7ns_7ns_7_2_1_U4.top_sub_7ns_7ns_7_2_1_Adder_1_U.clk )
\sub_7ns_7ns_7_2_1_U4.top_sub_7ns_7ns_7_2_1_Adder_1_U.bin_s1  <= _255_;
always @(posedge \sub_7ns_7ns_7_2_1_U4.top_sub_7ns_7ns_7_2_1_Adder_1_U.clk )
\sub_7ns_7ns_7_2_1_U4.top_sub_7ns_7ns_7_2_1_Adder_1_U.ain_s1  <= _254_;
always @(posedge \sub_7ns_7ns_7_2_1_U4.top_sub_7ns_7ns_7_2_1_Adder_1_U.clk )
\sub_7ns_7ns_7_2_1_U4.top_sub_7ns_7ns_7_2_1_Adder_1_U.sum_s1  <= _257_;
always @(posedge \sub_7ns_7ns_7_2_1_U4.top_sub_7ns_7ns_7_2_1_Adder_1_U.clk )
\sub_7ns_7ns_7_2_1_U4.top_sub_7ns_7ns_7_2_1_Adder_1_U.carry_s1  <= _256_;
assign _255_ = \sub_7ns_7ns_7_2_1_U4.top_sub_7ns_7ns_7_2_1_Adder_1_U.ce  ? \sub_7ns_7ns_7_2_1_U4.top_sub_7ns_7ns_7_2_1_Adder_1_U.bin_s0 [6:3] : \sub_7ns_7ns_7_2_1_U4.top_sub_7ns_7ns_7_2_1_Adder_1_U.bin_s1 ;
assign _254_ = \sub_7ns_7ns_7_2_1_U4.top_sub_7ns_7ns_7_2_1_Adder_1_U.ce  ? \sub_7ns_7ns_7_2_1_U4.top_sub_7ns_7ns_7_2_1_Adder_1_U.a [6:3] : \sub_7ns_7ns_7_2_1_U4.top_sub_7ns_7ns_7_2_1_Adder_1_U.ain_s1 ;
assign _256_ = \sub_7ns_7ns_7_2_1_U4.top_sub_7ns_7ns_7_2_1_Adder_1_U.ce  ? \sub_7ns_7ns_7_2_1_U4.top_sub_7ns_7ns_7_2_1_Adder_1_U.facout_s1  : \sub_7ns_7ns_7_2_1_U4.top_sub_7ns_7ns_7_2_1_Adder_1_U.carry_s1 ;
assign _257_ = \sub_7ns_7ns_7_2_1_U4.top_sub_7ns_7ns_7_2_1_Adder_1_U.ce  ? \sub_7ns_7ns_7_2_1_U4.top_sub_7ns_7ns_7_2_1_Adder_1_U.fas_s1  : \sub_7ns_7ns_7_2_1_U4.top_sub_7ns_7ns_7_2_1_Adder_1_U.sum_s1 ;
assign _258_ = \sub_7ns_7ns_7_2_1_U4.top_sub_7ns_7ns_7_2_1_Adder_1_U.u1.a  + \sub_7ns_7ns_7_2_1_U4.top_sub_7ns_7ns_7_2_1_Adder_1_U.u1.b ;
assign { \sub_7ns_7ns_7_2_1_U4.top_sub_7ns_7ns_7_2_1_Adder_1_U.u1.cout , \sub_7ns_7ns_7_2_1_U4.top_sub_7ns_7ns_7_2_1_Adder_1_U.u1.s  } = _258_ + \sub_7ns_7ns_7_2_1_U4.top_sub_7ns_7ns_7_2_1_Adder_1_U.u1.cin ;
assign _259_ = \sub_7ns_7ns_7_2_1_U4.top_sub_7ns_7ns_7_2_1_Adder_1_U.u2.a  + \sub_7ns_7ns_7_2_1_U4.top_sub_7ns_7ns_7_2_1_Adder_1_U.u2.b ;
assign { \sub_7ns_7ns_7_2_1_U4.top_sub_7ns_7ns_7_2_1_Adder_1_U.u2.cout , \sub_7ns_7ns_7_2_1_U4.top_sub_7ns_7ns_7_2_1_Adder_1_U.u2.s  } = _259_ + \sub_7ns_7ns_7_2_1_U4.top_sub_7ns_7ns_7_2_1_Adder_1_U.u2.cin ;
assign _260_ = $signed({ 1'h0, signbit_reg_1488, 7'h00 }) < $signed(op_6);
assign _261_ = $signed(op_1[15:1]) < $signed(2'h1);
assign _262_ = | { trunc_ln851_4_reg_1834, 3'h0 };
assign _263_ = | trunc_ln851_5_reg_1988;
assign _264_ = | op_15[12:0];
assign _265_ = ret_V_22_reg_1792 != op_8;
assign _266_ = | trunc_ln1115_reg_1531;
assign or_ln340_1_fu_967_p2 = overflow_1_fu_962_p2 | neg_src_4_fu_947_p2;
assign or_ln340_2_fu_1036_p2 = or_ln340_reg_1918 | and_ln786_reg_1880;
assign or_ln340_3_fu_1061_p2 = and_ln785_2_fu_1047_p2 | and_ln340_fu_1056_p2;
assign or_ln340_4_fu_1113_p2 = or_ln340_1_reg_1929 | and_ln786_1_reg_1900;
assign or_ln340_5_fu_1138_p2 = and_ln785_6_fu_1124_p2 | and_ln340_1_fu_1133_p2;
assign or_ln340_fu_917_p2 = overflow_fu_912_p2 | neg_src_fu_897_p2;
assign or_ln406_fu_580_p2 = r_V_3_reg_1595[0] | p_Result_21_reg_1602;
assign or_ln785_1_fu_957_p2 = xor_ln785_2_fu_952_p2 | p_Result_29_reg_1785;
assign or_ln785_2_fu_927_p2 = p_Result_21_reg_1602 | and_ln785_fu_923_p2;
assign or_ln785_3_fu_977_p2 = p_Result_26_reg_1536 | and_ln785_4_fu_973_p2;
assign or_ln785_fu_907_p2 = xor_ln785_fu_902_p2 | p_Result_24_reg_1769;
always @(posedge ap_clk)
trunc_ln728_reg_1478 <= _091_;
always @(posedge ap_clk)
signbit_reg_1488 <= _086_;
always @(posedge ap_clk)
select_ln353_1_reg_2065 <= _082_;
always @(posedge ap_clk)
select_ln340_reg_1947 <= _081_;
always @(posedge ap_clk)
select_ln340_1_reg_1957 <= _080_;
always @(posedge ap_clk)
sel_tmp11_reg_1952 <= _078_;
always @(posedge ap_clk)
sel_tmp25_reg_1962 <= _079_;
always @(posedge ap_clk)
ret_V_9_reg_2119 <= _075_;
always @(posedge ap_clk)
ret_V_26_reg_2033 <= _066_;
always @(posedge ap_clk)
ret_V_34_cast_reg_2038 <= _069_;
always @(posedge ap_clk)
ret_V_23_reg_2129 <= _063_;
always @(posedge ap_clk)
ret_V_28_reg_2134 <= _068_;
always @(posedge ap_clk)
ret_V_19_reg_1740 <= _060_;
always @(posedge ap_clk)
ret_V_6_reg_1755 <= _073_;
always @(posedge ap_clk)
ret_V_13_reg_1797 <= _058_;
always @(posedge ap_clk)
r_V_reg_2085 <= _056_;
always @(posedge ap_clk)
ret_V_7_reg_2090 <= _074_;
always @(posedge ap_clk)
trunc_ln851_2_reg_2097 <= _093_;
always @(posedge ap_clk)
ret_V_27_reg_2102 <= _067_;
always @(posedge ap_clk)
ret_V_36_cast_reg_2107 <= _070_;
always @(posedge ap_clk)
p_Val2_3_reg_1760 <= _050_;
always @(posedge ap_clk)
p_Result_24_reg_1769 <= _041_;
always @(posedge ap_clk)
p_Val2_7_reg_1776 <= _052_;
always @(posedge ap_clk)
p_Result_29_reg_1785 <= _046_;
always @(posedge ap_clk)
ret_V_22_reg_1792 <= _062_;
always @(posedge ap_clk)
op_14_V_reg_1972 <= _033_;
always @(posedge ap_clk)
op_9_V_reg_1977 <= _035_;
always @(posedge ap_clk)
select_ln353_reg_1983 <= _083_;
always @(posedge ap_clk)
trunc_ln851_5_reg_1988 <= _095_;
always @(posedge ap_clk)
ret_V_18_reg_1509 <= _059_;
always @(posedge ap_clk)
ret_V_cast_reg_1514 <= _076_;
always @(posedge ap_clk)
trunc_ln851_reg_1521 <= _096_;
always @(posedge ap_clk)
r_V_4_reg_1526 <= _055_;
always @(posedge ap_clk)
trunc_ln1115_reg_1531 <= _090_;
always @(posedge ap_clk)
p_Result_26_reg_1536 <= _043_;
always @(posedge ap_clk)
p_Val2_6_reg_1543 <= _051_;
always @(posedge ap_clk)
r_1_reg_1548 <= _053_;
always @(posedge ap_clk)
p_Result_28_reg_1553 <= _045_;
always @(posedge ap_clk)
p_Result_30_reg_1558 <= _047_;
always @(posedge ap_clk)
tmp_1_reg_1564 <= _087_;
always @(posedge ap_clk)
tmp_2_reg_1569 <= _088_;
always @(posedge ap_clk)
lhs_V_4_reg_1585 <= _032_;
always @(posedge ap_clk)
ret_V_3_reg_1802 <= _071_;
always @(posedge ap_clk)
xor_ln416_reg_1807 <= _098_;
always @(posedge ap_clk)
xor_ln416_1_reg_1813 <= _097_;
always @(posedge ap_clk)
_700_ <= _101_;
assign zext_ln1116_reg_1819[3:0] = _700_;
always @(posedge ap_clk)
icmp_ln874_reg_1824 <= _031_;
always @(posedge ap_clk)
select_ln850_5_reg_1829 <= _084_;
always @(posedge ap_clk)
trunc_ln851_4_reg_1834 <= _094_;
always @(posedge ap_clk)
icmp_ln851_6_reg_2080 <= _029_;
always @(posedge ap_clk)
icmp_ln851_2_reg_2114 <= _025_;
always @(posedge ap_clk)
icmp_ln1496_reg_1504 <= _023_;
always @(posedge ap_clk)
carry_1_reg_1839 <= _019_;
always @(posedge ap_clk)
carry_3_reg_1846 <= _020_;
always @(posedge ap_clk)
icmp_ln851_4_reg_1863 <= _027_;
always @(posedge ap_clk)
deleted_zeros_reg_1868 <= _022_;
always @(posedge ap_clk)
xor_ln785_1_reg_1874 <= _099_;
always @(posedge ap_clk)
and_ln786_reg_1880 <= _017_;
always @(posedge ap_clk)
deleted_zeros_1_reg_1888 <= _021_;
always @(posedge ap_clk)
xor_ln785_3_reg_1894 <= _100_;
always @(posedge ap_clk)
and_ln786_1_reg_1900 <= _016_;
always @(posedge ap_clk)
ret_V_25_reg_1908 <= _065_;
always @(posedge ap_clk)
tmp_3_reg_1913 <= _089_;
always @(posedge ap_clk)
or_ln340_reg_1918 <= _037_;
always @(posedge ap_clk)
and_ln785_1_reg_1924 <= _014_;
always @(posedge ap_clk)
or_ln340_1_reg_1929 <= _036_;
always @(posedge ap_clk)
and_ln785_5_reg_1935 <= _015_;
always @(posedge ap_clk)
sext_ln850_reg_1940 <= _085_;
always @(posedge ap_clk)
add_ln69_reg_2144 <= _011_;
always @(posedge ap_clk)
add_ln69_2_reg_2055 <= _010_;
always @(posedge ap_clk)
op_16_V_reg_2003 <= _034_;
always @(posedge ap_clk)
icmp_ln851_5_reg_2023 <= _028_;
always @(posedge ap_clk)
add_ln69_1_reg_2028 <= _009_;
always @(posedge ap_clk)
add_ln691_reg_1967 <= _008_;
always @(posedge ap_clk)
add_ln691_2_reg_2124 <= _007_;
always @(posedge ap_clk)
add_ln691_1_reg_2060 <= _006_;
always @(posedge ap_clk)
ret_V_reg_1691 <= _077_;
always @(posedge ap_clk)
and_ln406_reg_1696 <= _012_;
always @(posedge ap_clk)
Range2_all_ones_reg_1701 <= _005_;
always @(posedge ap_clk)
Range1_all_ones_reg_1706 <= _001_;
always @(posedge ap_clk)
Range1_all_zeros_reg_1713 <= _003_;
always @(posedge ap_clk)
and_ln408_reg_1718 <= _013_;
always @(posedge ap_clk)
icmp_ln851_1_reg_1723 <= _024_;
always @(posedge ap_clk)
ret_V_24_reg_1728 <= _064_;
always @(posedge ap_clk)
ret_V_12_reg_1733 <= _057_;
always @(posedge ap_clk)
icmp_ln851_reg_1590 <= _030_;
always @(posedge ap_clk)
r_V_3_reg_1595 <= _054_;
always @(posedge ap_clk)
p_Result_21_reg_1602 <= _039_;
always @(posedge ap_clk)
p_Val2_2_reg_1610 <= _049_;
always @(posedge ap_clk)
p_Result_23_reg_1615 <= _040_;
always @(posedge ap_clk)
p_Result_25_reg_1620 <= _042_;
always @(posedge ap_clk)
p_Result_s_22_reg_1626 <= _048_;
always @(posedge ap_clk)
p_Result_1_reg_1631 <= _038_;
always @(posedge ap_clk)
p_Result_27_reg_1637 <= _044_;
always @(posedge ap_clk)
Range2_all_ones_1_reg_1642 <= _004_;
always @(posedge ap_clk)
Range1_all_ones_1_reg_1647 <= _000_;
always @(posedge ap_clk)
Range1_all_zeros_1_reg_1654 <= _002_;
always @(posedge ap_clk)
ret_V_21_reg_1659 <= _061_;
always @(posedge ap_clk)
ret_V_6_cast_reg_1664 <= _072_;
always @(posedge ap_clk)
trunc_ln851_1_reg_1671 <= _092_;
always @(posedge ap_clk)
icmp_ln851_3_reg_1686 <= _026_;
always @(posedge ap_clk)
ap_CS_fsm <= _018_;
assign _102_ = _110_ ? 2'h2 : 2'h1;
assign _267_ = ap_CS_fsm == 1'h1;
function [30:0] _759_;
input [30:0] a;
input [960:0] b;
input [30:0] s;
case (s)
31'b0000000000000000000000000000001:
_759_ = b[30:0];
31'b0000000000000000000000000000010:
_759_ = b[61:31];
31'b0000000000000000000000000000100:
_759_ = b[92:62];
31'b0000000000000000000000000001000:
_759_ = b[123:93];
31'b0000000000000000000000000010000:
_759_ = b[154:124];
31'b0000000000000000000000000100000:
_759_ = b[185:155];
31'b0000000000000000000000001000000:
_759_ = b[216:186];
31'b0000000000000000000000010000000:
_759_ = b[247:217];
31'b0000000000000000000000100000000:
_759_ = b[278:248];
31'b0000000000000000000001000000000:
_759_ = b[309:279];
31'b0000000000000000000010000000000:
_759_ = b[340:310];
31'b0000000000000000000100000000000:
_759_ = b[371:341];
31'b0000000000000000001000000000000:
_759_ = b[402:372];
31'b0000000000000000010000000000000:
_759_ = b[433:403];
31'b0000000000000000100000000000000:
_759_ = b[464:434];
31'b0000000000000001000000000000000:
_759_ = b[495:465];
31'b0000000000000010000000000000000:
_759_ = b[526:496];
31'b0000000000000100000000000000000:
_759_ = b[557:527];
31'b0000000000001000000000000000000:
_759_ = b[588:558];
31'b0000000000010000000000000000000:
_759_ = b[619:589];
31'b0000000000100000000000000000000:
_759_ = b[650:620];
31'b0000000001000000000000000000000:
_759_ = b[681:651];
31'b0000000010000000000000000000000:
_759_ = b[712:682];
31'b0000000100000000000000000000000:
_759_ = b[743:713];
31'b0000001000000000000000000000000:
_759_ = b[774:744];
31'b0000010000000000000000000000000:
_759_ = b[805:775];
31'b0000100000000000000000000000000:
_759_ = b[836:806];
31'b0001000000000000000000000000000:
_759_ = b[867:837];
31'b0010000000000000000000000000000:
_759_ = b[898:868];
31'b0100000000000000000000000000000:
_759_ = b[929:899];
31'b1000000000000000000000000000000:
_759_ = b[960:930];
31'b0000000000000000000000000000000:
_759_ = a;
default:
_759_ = 31'bx;
endcase
endfunction
assign ap_NS_fsm = _759_(31'hxxxxxxxx, { 29'h00000000, _102_, 930'h00000002000000080000002000000080000002000000080000002000000080000002000000080000002000000080000002000000080000002000000080000002000000080000002000000080000002000000080000002000000080000002000000080000002000000080000002000000000000001 }, { _267_, _297_, _296_, _295_, _294_, _293_, _292_, _291_, _290_, _289_, _288_, _287_, _286_, _285_, _284_, _283_, _282_, _281_, _280_, _279_, _278_, _277_, _276_, _275_, _274_, _273_, _272_, _271_, _270_, _269_, _268_ });
assign _268_ = ap_CS_fsm == 31'h40000000;
assign _269_ = ap_CS_fsm == 30'h20000000;
assign _270_ = ap_CS_fsm == 29'h10000000;
assign _271_ = ap_CS_fsm == 28'h8000000;
assign _272_ = ap_CS_fsm == 27'h4000000;
assign _273_ = ap_CS_fsm == 26'h2000000;
assign _274_ = ap_CS_fsm == 25'h1000000;
assign _275_ = ap_CS_fsm == 24'h800000;
assign _276_ = ap_CS_fsm == 23'h400000;
assign _277_ = ap_CS_fsm == 22'h200000;
assign _278_ = ap_CS_fsm == 21'h100000;
assign _279_ = ap_CS_fsm == 20'h80000;
assign _280_ = ap_CS_fsm == 19'h40000;
assign _281_ = ap_CS_fsm == 18'h20000;
assign _282_ = ap_CS_fsm == 17'h10000;
assign _283_ = ap_CS_fsm == 16'h8000;
assign _284_ = ap_CS_fsm == 15'h4000;
assign _285_ = ap_CS_fsm == 14'h2000;
assign _286_ = ap_CS_fsm == 13'h1000;
assign _287_ = ap_CS_fsm == 12'h800;
assign _288_ = ap_CS_fsm == 11'h400;
assign _289_ = ap_CS_fsm == 10'h200;
assign _290_ = ap_CS_fsm == 9'h100;
assign _291_ = ap_CS_fsm == 8'h80;
assign _292_ = ap_CS_fsm == 7'h40;
assign _293_ = ap_CS_fsm == 6'h20;
assign _294_ = ap_CS_fsm == 5'h10;
assign _295_ = ap_CS_fsm == 4'h8;
assign _296_ = ap_CS_fsm == 3'h4;
assign _297_ = ap_CS_fsm == 2'h2;
assign op_28_ap_vld = ap_CS_fsm[30] ? 1'h1 : 1'h0;
assign ap_idle = _109_ ? 1'h1 : 1'h0;
assign _091_ = ap_CS_fsm[1] ? op_8[3:0] : trunc_ln728_reg_1478;
assign _086_ = ap_CS_fsm[4] ? signbit_fu_288_p2 : signbit_reg_1488;
assign _082_ = ap_CS_fsm[21] ? select_ln353_1_fu_1305_p3 : select_ln353_1_reg_2065;
assign _081_ = _108_ ? select_ln340_fu_1040_p3 : select_ln340_reg_1947;
assign _080_ = _107_ ? select_ln340_1_fu_1117_p3 : select_ln340_1_reg_1957;
assign _079_ = ap_CS_fsm[15] ? sel_tmp25_fu_1144_p2 : sel_tmp25_reg_1962;
assign _078_ = ap_CS_fsm[15] ? sel_tmp11_fu_1067_p2 : sel_tmp11_reg_1952;
assign _075_ = ap_CS_fsm[25] ? grp_fu_1372_p2 : ret_V_9_reg_2119;
assign _069_ = ap_CS_fsm[18] ? grp_fu_1255_p2[33:2] : ret_V_34_cast_reg_2038;
assign _066_ = ap_CS_fsm[18] ? grp_fu_1255_p2 : ret_V_26_reg_2033;
assign _068_ = ap_CS_fsm[26] ? ret_V_28_fu_1413_p3 : ret_V_28_reg_2134;
assign _063_ = ap_CS_fsm[26] ? ret_V_23_fu_1394_p3 : ret_V_23_reg_2129;
assign _073_ = ap_CS_fsm[9] ? grp_fu_615_p2 : ret_V_6_reg_1755;
assign _060_ = ap_CS_fsm[9] ? ret_V_19_fu_642_p3 : ret_V_19_reg_1740;
assign _058_ = _106_ ? grp_fu_665_p2 : ret_V_13_reg_1797;
assign _070_ = ap_CS_fsm[23] ? grp_fu_1327_p2[44:13] : ret_V_36_cast_reg_2107;
assign _067_ = ap_CS_fsm[23] ? grp_fu_1327_p2 : ret_V_27_reg_2102;
assign _093_ = ap_CS_fsm[23] ? grp_fu_1236_p2[1:0] : trunc_ln851_2_reg_2097;
assign _074_ = ap_CS_fsm[23] ? grp_fu_1236_p2[7:2] : ret_V_7_reg_2090;
assign _056_ = ap_CS_fsm[23] ? grp_fu_1236_p2 : r_V_reg_2085;
assign _062_ = ap_CS_fsm[10] ? ret_V_22_fu_698_p3 : ret_V_22_reg_1792;
assign _046_ = ap_CS_fsm[10] ? grp_fu_660_p2[3] : p_Result_29_reg_1785;
assign _052_ = ap_CS_fsm[10] ? grp_fu_660_p2 : p_Val2_7_reg_1776;
assign _041_ = ap_CS_fsm[10] ? grp_fu_652_p2[3] : p_Result_24_reg_1769;
assign _050_ = ap_CS_fsm[10] ? grp_fu_652_p2 : p_Val2_3_reg_1760;
assign _095_ = ap_CS_fsm[16] ? op_14_V_fu_1155_p3[1:0] : trunc_ln851_5_reg_1988;
assign _083_ = ap_CS_fsm[16] ? select_ln353_fu_1184_p3 : select_ln353_reg_1983;
assign _035_ = ap_CS_fsm[16] ? op_9_V_fu_1166_p3 : op_9_V_reg_1977;
assign _033_ = ap_CS_fsm[16] ? op_14_V_fu_1155_p3 : op_14_V_reg_1972;
assign _032_ = ap_CS_fsm[6] ? lhs_V_4_fu_436_p2 : lhs_V_4_reg_1585;
assign _088_ = ap_CS_fsm[6] ? grp_fu_255_p2[10:6] : tmp_2_reg_1569;
assign _087_ = ap_CS_fsm[6] ? grp_fu_255_p2[10:7] : tmp_1_reg_1564;
assign _047_ = ap_CS_fsm[6] ? grp_fu_255_p2[6] : p_Result_30_reg_1558;
assign _045_ = ap_CS_fsm[6] ? grp_fu_255_p2[5] : p_Result_28_reg_1553;
assign _053_ = ap_CS_fsm[6] ? grp_fu_255_p2[0] : r_1_reg_1548;
assign _051_ = ap_CS_fsm[6] ? grp_fu_255_p2[5:2] : p_Val2_6_reg_1543;
assign _043_ = ap_CS_fsm[6] ? grp_fu_255_p2[10] : p_Result_26_reg_1536;
assign _090_ = ap_CS_fsm[6] ? grp_fu_255_p2[1:0] : trunc_ln1115_reg_1531;
assign _055_ = ap_CS_fsm[6] ? grp_fu_255_p2 : r_V_4_reg_1526;
assign _096_ = ap_CS_fsm[6] ? grp_fu_309_p2[6:0] : trunc_ln851_reg_1521;
assign _076_ = ap_CS_fsm[6] ? grp_fu_309_p2[8:7] : ret_V_cast_reg_1514;
assign _059_ = ap_CS_fsm[6] ? grp_fu_309_p2 : ret_V_18_reg_1509;
assign _094_ = ap_CS_fsm[11] ? ret_V_3_fu_719_p2[3:0] : trunc_ln851_4_reg_1834;
assign _084_ = ap_CS_fsm[11] ? select_ln850_5_fu_755_p3 : select_ln850_5_reg_1829;
assign _031_ = ap_CS_fsm[11] ? icmp_ln874_fu_738_p2 : icmp_ln874_reg_1824;
assign _101_ = ap_CS_fsm[11] ? ret_V_22_reg_1792 : zext_ln1116_reg_1819[3:0];
assign _097_ = ap_CS_fsm[11] ? xor_ln416_1_fu_730_p2 : xor_ln416_1_reg_1813;
assign _098_ = ap_CS_fsm[11] ? xor_ln416_fu_725_p2 : xor_ln416_reg_1807;
assign _071_ = ap_CS_fsm[11] ? ret_V_3_fu_719_p2 : ret_V_3_reg_1802;
assign _029_ = ap_CS_fsm[22] ? icmp_ln851_6_fu_1337_p2 : icmp_ln851_6_reg_2080;
assign _025_ = ap_CS_fsm[24] ? icmp_ln851_2_fu_1367_p2 : icmp_ln851_2_reg_2114;
assign _023_ = ap_CS_fsm[5] ? icmp_ln1496_fu_326_p2 : icmp_ln1496_reg_1504;
assign _027_ = ap_CS_fsm[12] ? icmp_ln851_4_fu_809_p2 : icmp_ln851_4_reg_1863;
assign _020_ = ap_CS_fsm[12] ? carry_3_fu_777_p2 : carry_3_reg_1846;
assign _019_ = ap_CS_fsm[12] ? carry_1_fu_773_p2 : carry_1_reg_1839;
assign _089_ = ap_CS_fsm[13] ? grp_fu_796_p2[24:7] : tmp_3_reg_1913;
assign _065_ = ap_CS_fsm[13] ? grp_fu_796_p2 : ret_V_25_reg_1908;
assign _016_ = ap_CS_fsm[13] ? and_ln786_1_fu_872_p2 : and_ln786_1_reg_1900;
assign _100_ = ap_CS_fsm[13] ? xor_ln785_3_fu_867_p2 : xor_ln785_3_reg_1894;
assign _021_ = ap_CS_fsm[13] ? deleted_zeros_1_fu_846_p3 : deleted_zeros_1_reg_1888;
assign _017_ = ap_CS_fsm[13] ? and_ln786_fu_841_p2 : and_ln786_reg_1880;
assign _099_ = ap_CS_fsm[13] ? xor_ln785_1_fu_836_p2 : xor_ln785_1_reg_1874;
assign _022_ = ap_CS_fsm[13] ? deleted_zeros_fu_815_p3 : deleted_zeros_reg_1868;
assign _085_ = ap_CS_fsm[14] ? { tmp_3_reg_1913[17], tmp_3_reg_1913 } : sext_ln850_reg_1940;
assign _015_ = ap_CS_fsm[14] ? and_ln785_5_fu_982_p2 : and_ln785_5_reg_1935;
assign _036_ = ap_CS_fsm[14] ? or_ln340_1_fu_967_p2 : or_ln340_1_reg_1929;
assign _014_ = ap_CS_fsm[14] ? and_ln785_1_fu_932_p2 : and_ln785_1_reg_1924;
assign _037_ = ap_CS_fsm[14] ? or_ln340_fu_917_p2 : or_ln340_reg_1918;
assign _011_ = ap_CS_fsm[28] ? grp_fu_1427_p2 : add_ln69_reg_2144;
assign _010_ = ap_CS_fsm[19] ? grp_fu_1282_p2 : add_ln69_2_reg_2055;
assign _009_ = ap_CS_fsm[17] ? grp_fu_1201_p2 : add_ln69_1_reg_2028;
assign _028_ = ap_CS_fsm[17] ? icmp_ln851_5_fu_1261_p2 : icmp_ln851_5_reg_2023;
assign _034_ = ap_CS_fsm[17] ? ret_V_20_fu_1217_p2[5:2] : op_16_V_reg_2003;
assign _008_ = _105_ ? grp_fu_990_p2 : add_ln691_reg_1967;
assign _007_ = _104_ ? grp_fu_1377_p2 : add_ln691_2_reg_2124;
assign _006_ = _103_ ? grp_fu_1288_p2 : add_ln691_1_reg_2060;
assign _057_ = ap_CS_fsm[8] ? grp_fu_554_p2[32:16] : ret_V_12_reg_1733;
assign _064_ = ap_CS_fsm[8] ? grp_fu_554_p2 : ret_V_24_reg_1728;
assign _024_ = ap_CS_fsm[8] ? icmp_ln851_1_fu_610_p2 : icmp_ln851_1_reg_1723;
assign _013_ = ap_CS_fsm[8] ? and_ln408_fu_606_p2 : and_ln408_reg_1718;
assign _003_ = ap_CS_fsm[8] ? Range1_all_zeros_fu_601_p2 : Range1_all_zeros_reg_1713;
assign _001_ = ap_CS_fsm[8] ? Range1_all_ones_fu_596_p2 : Range1_all_ones_reg_1706;
assign _005_ = ap_CS_fsm[8] ? Range2_all_ones_fu_591_p2 : Range2_all_ones_reg_1701;
assign _012_ = ap_CS_fsm[8] ? and_ln406_fu_585_p2 : and_ln406_reg_1696;
assign _077_ = ap_CS_fsm[8] ? grp_fu_446_p2 : ret_V_reg_1691;
assign _026_ = ap_CS_fsm[7] ? icmp_ln851_3_fu_564_p2 : icmp_ln851_3_reg_1686;
assign _092_ = ap_CS_fsm[7] ? grp_fu_430_p2[2:0] : trunc_ln851_1_reg_1671;
assign _072_ = ap_CS_fsm[7] ? grp_fu_430_p2[6:3] : ret_V_6_cast_reg_1664;
assign _061_ = ap_CS_fsm[7] ? grp_fu_430_p2 : ret_V_21_reg_1659;
assign _002_ = ap_CS_fsm[7] ? Range1_all_zeros_1_fu_520_p2 : Range1_all_zeros_1_reg_1654;
assign _000_ = ap_CS_fsm[7] ? Range1_all_ones_1_fu_515_p2 : Range1_all_ones_1_reg_1647;
assign _004_ = ap_CS_fsm[7] ? Range2_all_ones_1_fu_510_p2 : Range2_all_ones_1_reg_1642;
assign _044_ = ap_CS_fsm[7] ? p_Result_27_fu_505_p2 : p_Result_27_reg_1637;
assign _038_ = ap_CS_fsm[7] ? grp_fu_268_p2[15:6] : p_Result_1_reg_1631;
assign _048_ = ap_CS_fsm[7] ? grp_fu_268_p2[15:7] : p_Result_s_22_reg_1626;
assign _042_ = ap_CS_fsm[7] ? grp_fu_268_p2[6] : p_Result_25_reg_1620;
assign _040_ = ap_CS_fsm[7] ? grp_fu_268_p2[5] : p_Result_23_reg_1615;
assign _049_ = ap_CS_fsm[7] ? grp_fu_268_p2[5:2] : p_Val2_2_reg_1610;
assign _039_ = ap_CS_fsm[7] ? grp_fu_268_p2[15] : p_Result_21_reg_1602;
assign _054_ = ap_CS_fsm[7] ? grp_fu_268_p2 : r_V_3_reg_1595;
assign _030_ = ap_CS_fsm[7] ? icmp_ln851_fu_441_p2 : icmp_ln851_reg_1590;
assign _018_ = ap_rst ? 31'h00000001 : ap_NS_fsm;
assign Range1_all_ones_1_fu_515_p2 = _115_ ? 1'h1 : 1'h0;
assign Range1_all_ones_fu_596_p2 = _116_ ? 1'h1 : 1'h0;
assign Range1_all_zeros_1_fu_520_p2 = _117_ ? 1'h1 : 1'h0;
assign Range1_all_zeros_fu_601_p2 = _118_ ? 1'h1 : 1'h0;
assign Range2_all_ones_1_fu_510_p2 = _119_ ? 1'h1 : 1'h0;
assign Range2_all_ones_fu_591_p2 = _120_ ? 1'h1 : 1'h0;
assign deleted_ones_1_fu_861_p3 = carry_3_reg_1846 ? and_ln780_1_fu_856_p2 : Range1_all_ones_1_reg_1647;
assign deleted_ones_fu_830_p3 = carry_1_reg_1839 ? and_ln780_fu_825_p2 : Range1_all_ones_reg_1706;
assign deleted_zeros_1_fu_846_p3 = carry_3_reg_1846 ? Range1_all_ones_1_reg_1647 : Range1_all_zeros_1_reg_1654;
assign deleted_zeros_fu_815_p3 = carry_1_reg_1839 ? Range1_all_ones_reg_1706 : Range1_all_zeros_reg_1713;
assign icmp_ln1496_fu_326_p2 = _260_ ? 1'h1 : 1'h0;
assign icmp_ln851_1_fu_610_p2 = _121_ ? 1'h1 : 1'h0;
assign icmp_ln851_2_fu_1367_p2 = _122_ ? 1'h1 : 1'h0;
assign icmp_ln851_3_fu_564_p2 = _123_ ? 1'h1 : 1'h0;
assign icmp_ln851_4_fu_809_p2 = _262_ ? 1'h1 : 1'h0;
assign icmp_ln851_5_fu_1261_p2 = _263_ ? 1'h1 : 1'h0;
assign icmp_ln851_6_fu_1337_p2 = _264_ ? 1'h1 : 1'h0;
assign icmp_ln851_fu_441_p2 = _124_ ? 1'h1 : 1'h0;
assign icmp_ln874_fu_738_p2 = _265_ ? 1'h1 : 1'h0;
assign op_14_V_fu_1155_p3 = sel_tmp11_reg_1952 ? p_Val2_3_reg_1760 : select_ln785_fu_1150_p3;
assign op_9_V_fu_1166_p3 = sel_tmp25_reg_1962 ? p_Val2_7_reg_1776 : select_ln785_1_fu_1161_p3;
assign p_Result_27_fu_505_p2 = _266_ ? 1'h1 : 1'h0;
assign ret_V_19_fu_642_p3 = ret_V_18_reg_1509[32] ? select_ln850_fu_637_p3 : ret_V_cast_reg_1514;
assign ret_V_22_fu_698_p3 = ret_V_21_reg_1659[6] ? select_ln850_1_fu_693_p3 : ret_V_6_cast_reg_1664;
assign ret_V_23_fu_1394_p3 = r_V_reg_2085[7] ? select_ln850_2_fu_1389_p3 : ret_V_7_reg_2090;
assign ret_V_28_fu_1413_p3 = ret_V_27_reg_2102[45] ? select_ln850_6_fu_1408_p3 : ret_V_36_cast_reg_2107;
assign select_ln340_1_fu_1117_p3 = or_ln340_4_fu_1113_p2 ? { p_Result_30_reg_1558, p_Val2_8_fu_1099_p2 } : p_Val2_7_reg_1776;
assign select_ln340_fu_1040_p3 = or_ln340_2_fu_1036_p2 ? { p_Result_25_reg_1620, p_Val2_4_fu_1022_p2 } : p_Val2_3_reg_1760;
assign select_ln353_1_fu_1305_p3 = ret_V_26_reg_2033[34] ? select_ln850_8_fu_1300_p3 : ret_V_34_cast_reg_2038;
assign select_ln353_fu_1184_p3 = ret_V_25_reg_1908[24] ? select_ln850_7_fu_1179_p3 : sext_ln850_reg_1940;
assign select_ln785_1_fu_1161_p3 = and_ln785_5_reg_1935 ? p_Val2_7_reg_1776 : select_ln340_1_reg_1957;
assign select_ln785_fu_1150_p3 = and_ln785_1_reg_1924 ? p_Val2_3_reg_1760 : select_ln340_reg_1947;
assign select_ln850_1_fu_693_p3 = icmp_ln851_1_reg_1723 ? ret_V_6_cast_reg_1664 : ret_V_6_reg_1755;
assign select_ln850_2_fu_1389_p3 = icmp_ln851_2_reg_2114 ? ret_V_7_reg_2090 : ret_V_9_reg_2119;
assign select_ln850_4_fu_750_p3 = icmp_ln851_3_reg_1686 ? ret_V_12_reg_1733 : ret_V_13_reg_1797;
assign select_ln850_5_fu_755_p3 = ret_V_24_reg_1728[32] ? select_ln850_4_fu_750_p3 : ret_V_12_reg_1733;
assign select_ln850_6_fu_1408_p3 = icmp_ln851_6_reg_2080 ? add_ln691_2_reg_2124 : ret_V_36_cast_reg_2107;
assign select_ln850_7_fu_1179_p3 = icmp_ln851_4_reg_1863 ? add_ln691_reg_1967 : sext_ln850_reg_1940;
assign select_ln850_8_fu_1300_p3 = icmp_ln851_5_reg_2023 ? add_ln691_1_reg_2060 : ret_V_34_cast_reg_2038;
assign select_ln850_fu_637_p3 = icmp_ln851_reg_1590 ? ret_V_cast_reg_1514 : ret_V_reg_1691;
assign signbit_fu_288_p2 = _261_ ? 1'h1 : 1'h0;
assign ret_V_3_fu_719_p2 = { op_8, 4'h0 } ^ { op_4[7], op_4[7], op_4[7], op_4[7], op_4[7], op_4 };
assign xor_ln365_2_fu_1087_p2 = p_Val2_7_reg_1776[3] ^ r_V_4_reg_1526[6];
assign xor_ln365_fu_1010_p2 = r_V_3_reg_1595[6] ^ p_Val2_3_reg_1760[3];
assign ap_CS_fsm_state1 = ap_CS_fsm[0];
assign ap_CS_fsm_state10 = ap_CS_fsm[9];
assign ap_CS_fsm_state11 = ap_CS_fsm[10];
assign ap_CS_fsm_state12 = ap_CS_fsm[11];
assign ap_CS_fsm_state13 = ap_CS_fsm[12];
assign ap_CS_fsm_state14 = ap_CS_fsm[13];
assign ap_CS_fsm_state15 = ap_CS_fsm[14];
assign ap_CS_fsm_state16 = ap_CS_fsm[15];
assign ap_CS_fsm_state17 = ap_CS_fsm[16];
assign ap_CS_fsm_state18 = ap_CS_fsm[17];
assign ap_CS_fsm_state19 = ap_CS_fsm[18];
assign ap_CS_fsm_state2 = ap_CS_fsm[1];
assign ap_CS_fsm_state20 = ap_CS_fsm[19];
assign ap_CS_fsm_state21 = ap_CS_fsm[20];
assign ap_CS_fsm_state22 = ap_CS_fsm[21];
assign ap_CS_fsm_state23 = ap_CS_fsm[22];
assign ap_CS_fsm_state24 = ap_CS_fsm[23];
assign ap_CS_fsm_state25 = ap_CS_fsm[24];
assign ap_CS_fsm_state26 = ap_CS_fsm[25];
assign ap_CS_fsm_state27 = ap_CS_fsm[26];
assign ap_CS_fsm_state28 = ap_CS_fsm[27];
assign ap_CS_fsm_state29 = ap_CS_fsm[28];
assign ap_CS_fsm_state30 = ap_CS_fsm[29];
assign ap_CS_fsm_state31 = ap_CS_fsm[30];
assign ap_CS_fsm_state5 = ap_CS_fsm[4];
assign ap_CS_fsm_state6 = ap_CS_fsm[5];
assign ap_CS_fsm_state7 = ap_CS_fsm[6];
assign ap_CS_fsm_state8 = ap_CS_fsm[7];
assign ap_CS_fsm_state9 = ap_CS_fsm[8];
assign ap_done = op_28_ap_vld;
assign ap_ready = op_28_ap_vld;
assign grp_fu_1201_p0 = { ret_V_19_reg_1740[1], ret_V_19_reg_1740 };
assign grp_fu_1201_p1 = { 2'h0, icmp_ln874_reg_1824 };
assign grp_fu_1236_p0 = zext_ln1116_reg_1819[3:0];
assign grp_fu_1255_p0 = { select_ln353_reg_1983[18], select_ln353_reg_1983[18], select_ln353_reg_1983[18], select_ln353_reg_1983[18], select_ln353_reg_1983[18], select_ln353_reg_1983[18], select_ln353_reg_1983[18], select_ln353_reg_1983[18], select_ln353_reg_1983[18], select_ln353_reg_1983[18], select_ln353_reg_1983[18], select_ln353_reg_1983[18], select_ln353_reg_1983[18], select_ln353_reg_1983[18], select_ln353_reg_1983, 2'h0 };
assign grp_fu_1255_p1 = { op_14_V_reg_1972[3], op_14_V_reg_1972[3], op_14_V_reg_1972[3], op_14_V_reg_1972[3], op_14_V_reg_1972[3], op_14_V_reg_1972[3], op_14_V_reg_1972[3], op_14_V_reg_1972[3], op_14_V_reg_1972[3], op_14_V_reg_1972[3], op_14_V_reg_1972[3], op_14_V_reg_1972[3], op_14_V_reg_1972[3], op_14_V_reg_1972[3], op_14_V_reg_1972[3], op_14_V_reg_1972[3], op_14_V_reg_1972[3], op_14_V_reg_1972[3], op_14_V_reg_1972[3], op_14_V_reg_1972[3], op_14_V_reg_1972[3], op_14_V_reg_1972[3], op_14_V_reg_1972[3], op_14_V_reg_1972[3], op_14_V_reg_1972[3], op_14_V_reg_1972[3], op_14_V_reg_1972[3], op_14_V_reg_1972[3], op_14_V_reg_1972[3], op_14_V_reg_1972[3], op_14_V_reg_1972[3], op_14_V_reg_1972 };
assign grp_fu_1282_p0 = { add_ln69_1_reg_2028[2], add_ln69_1_reg_2028[2], add_ln69_1_reg_2028 };
assign grp_fu_1282_p1 = { op_16_V_reg_2003[3], op_16_V_reg_2003 };
assign grp_fu_1327_p0 = { select_ln353_1_reg_2065[31], select_ln353_1_reg_2065, 13'h0000 };
assign grp_fu_1327_p1 = { op_15[15], op_15[15], op_15[15], op_15[15], op_15[15], op_15[15], op_15[15], op_15[15], op_15[15], op_15[15], op_15[15], op_15[15], op_15[15], op_15[15], op_15[15], op_15[15], op_15[15], op_15[15], op_15[15], op_15[15], op_15[15], op_15[15], op_15[15], op_15[15], op_15[15], op_15[15], op_15[15], op_15[15], op_15[15], op_15[15], op_15 };
assign grp_fu_1427_p1 = { 16'h0000, ret_V_23_reg_2129[5], ret_V_23_reg_2129[5], ret_V_23_reg_2129[5], ret_V_23_reg_2129[5], ret_V_23_reg_2129[5], ret_V_23_reg_2129[5], ret_V_23_reg_2129[5], ret_V_23_reg_2129[5], ret_V_23_reg_2129[5], ret_V_23_reg_2129[5], ret_V_23_reg_2129 };
assign grp_fu_1435_p0 = { add_ln69_2_reg_2055[4], add_ln69_2_reg_2055[4], add_ln69_2_reg_2055[4], add_ln69_2_reg_2055[4], add_ln69_2_reg_2055[4], add_ln69_2_reg_2055[4], add_ln69_2_reg_2055[4], add_ln69_2_reg_2055[4], add_ln69_2_reg_2055[4], add_ln69_2_reg_2055[4], add_ln69_2_reg_2055[4], add_ln69_2_reg_2055[4], add_ln69_2_reg_2055[4], add_ln69_2_reg_2055[4], add_ln69_2_reg_2055[4], add_ln69_2_reg_2055[4], add_ln69_2_reg_2055[4], add_ln69_2_reg_2055[4], add_ln69_2_reg_2055[4], add_ln69_2_reg_2055[4], add_ln69_2_reg_2055[4], add_ln69_2_reg_2055[4], add_ln69_2_reg_2055[4], add_ln69_2_reg_2055[4], add_ln69_2_reg_2055[4], add_ln69_2_reg_2055[4], add_ln69_2_reg_2055[4], add_ln69_2_reg_2055 };
assign grp_fu_255_p1 = { op_0, 1'h0 };
assign grp_fu_255_p10 = { 8'h00, op_0, 1'h0 };
assign grp_fu_268_p0 = op_8;
assign grp_fu_268_p00 = { 8'h00, op_8 };
assign grp_fu_309_p0 = { op_1[15], op_1[15], op_1[15], op_1[15], op_1[15], op_1[15], op_1[15], op_1[15], op_1[15], op_1[15], op_1[15], op_1, 6'h00 };
assign grp_fu_309_p1 = { op_6[31], op_6 };
assign grp_fu_430_p0 = { 1'h0, op_0, 4'h0 };
assign grp_fu_430_p1 = { 3'h0, signbit_reg_1488, 3'h0 };
assign grp_fu_554_p0 = { 16'h0000, lhs_V_4_reg_1585, 16'h0000 };
assign grp_fu_554_p1 = { op_11[31], op_11 };
assign grp_fu_652_p1 = { 3'h0, and_ln406_reg_1696 };
assign grp_fu_660_p1 = { 3'h0, and_ln408_reg_1718 };
assign grp_fu_796_p0 = { select_ln850_5_reg_1829[16], select_ln850_5_reg_1829, 7'h00 };
assign grp_fu_796_p1 = { ret_V_3_reg_1802[12], ret_V_3_reg_1802[12], ret_V_3_reg_1802[12], ret_V_3_reg_1802[12], ret_V_3_reg_1802[12], ret_V_3_reg_1802[12], ret_V_3_reg_1802[12], ret_V_3_reg_1802[12], ret_V_3_reg_1802[12], ret_V_3_reg_1802, 3'h0 };
assign grp_fu_990_p0 = { tmp_3_reg_1913[17], tmp_3_reg_1913 };
assign icmp_ln1496_fu_326_p1 = op_6;
assign lhs_V_2_fu_415_p3 = { op_0, 4'h0 };
assign lhs_V_5_fu_539_p3 = { lhs_V_4_reg_1585, 16'h0000 };
assign lhs_V_fu_1207_p3 = { trunc_ln728_reg_1478, 2'h0 };
assign lhs_fu_294_p3 = { op_1, 6'h00 };
assign op_12_V_fu_766_p3 = { ret_V_3_reg_1802, 3'h0 };
assign op_28 = grp_fu_1435_p2;
assign op_5_V_fu_408_p3 = { signbit_reg_1488, 3'h0 };
assign p_Result_14_fu_1104_p4 = { p_Result_30_reg_1558, p_Val2_8_fu_1099_p2 };
assign p_Result_15_fu_686_p3 = ret_V_21_reg_1659[6];
assign p_Result_16_fu_1382_p3 = r_V_reg_2085[7];
assign p_Result_17_fu_743_p3 = ret_V_24_reg_1728[32];
assign p_Result_18_fu_1172_p3 = ret_V_25_reg_1908[24];
assign p_Result_19_fu_1293_p3 = ret_V_26_reg_2033[34];
assign p_Result_20_fu_1401_p3 = ret_V_27_reg_2102[45];
assign p_Result_22_fu_570_p3 = r_V_3_reg_1595[1];
assign p_Result_5_fu_802_p3 = { trunc_ln851_4_reg_1834, 3'h0 };
assign p_Result_8_fu_1027_p4 = { p_Result_25_reg_1620, p_Val2_4_fu_1022_p2 };
assign p_Result_s_fu_630_p3 = ret_V_18_reg_1509[32];
assign r_1_fu_368_p1 = grp_fu_255_p2[0];
assign r_fu_577_p1 = r_V_3_reg_1595[0];
assign ret_fu_239_p3 = { op_0, 1'h0 };
assign rhs_3_fu_785_p3 = { select_ln850_5_reg_1829, 7'h00 };
assign rhs_4_fu_1316_p3 = { select_ln353_1_reg_2065, 13'h0000 };
assign rhs_fu_708_p3 = { op_8, 4'h0 };
assign sext_ln1194_fu_1214_p1 = { op_9_V_reg_1977[3], op_9_V_reg_1977[3], op_9_V_reg_1977 };
assign sext_ln69_1_fu_1420_p1 = { ret_V_23_reg_2129[5], ret_V_23_reg_2129[5], ret_V_23_reg_2129[5], ret_V_23_reg_2129[5], ret_V_23_reg_2129[5], ret_V_23_reg_2129[5], ret_V_23_reg_2129[5], ret_V_23_reg_2129[5], ret_V_23_reg_2129[5], ret_V_23_reg_2129[5], ret_V_23_reg_2129 };
assign sext_ln703_1_fu_705_p0 = op_4;
assign sext_ln703_1_fu_705_p1 = { op_4[7], op_4[7], op_4[7], op_4[7], op_4[7], op_4 };
assign sext_ln703_2_fu_550_p0 = op_11;
assign sext_ln703_4_fu_1312_p0 = op_15;
assign sext_ln703_fu_305_p0 = op_6;
assign sext_ln850_fu_987_p1 = { tmp_3_reg_1913[17], tmp_3_reg_1913 };
assign shl_ln_fu_315_p3 = { signbit_reg_1488, 7'h00 };
assign tmp_10_fu_1073_p3 = r_V_4_reg_1526[6];
assign tmp_11_fu_1080_p3 = p_Val2_7_reg_1776[3];
assign tmp_13_fu_278_p4 = op_1[15:1];
assign tmp_18_fu_1244_p3 = { select_ln353_reg_1983, 2'h0 };
assign tmp_4_fu_1003_p3 = p_Val2_3_reg_1760[3];
assign tmp_fu_996_p3 = r_V_3_reg_1595[6];
assign trunc_ln1115_fu_346_p1 = grp_fu_255_p2[1:0];
assign trunc_ln728_fu_274_p1 = op_8[3:0];
assign trunc_ln851_1_fu_535_p1 = grp_fu_430_p2[2:0];
assign trunc_ln851_2_fu_1353_p1 = grp_fu_1236_p2[1:0];
assign trunc_ln851_3_fu_560_p0 = op_11;
assign trunc_ln851_3_fu_560_p1 = op_11[15:0];
assign trunc_ln851_4_fu_762_p1 = ret_V_3_fu_719_p2[3:0];
assign trunc_ln851_5_fu_1191_p1 = op_14_V_fu_1155_p3[1:0];
assign trunc_ln851_6_fu_1333_p0 = op_15;
assign trunc_ln851_6_fu_1333_p1 = op_15[12:0];
assign trunc_ln851_fu_342_p1 = grp_fu_309_p2[6:0];
assign zext_ln1116_fu_735_p1 = { 4'h0, ret_V_22_reg_1792 };
assign zext_ln1196_fu_715_p1 = { 1'h0, op_8, 4'h0 };
assign zext_ln1496_fu_322_p1 = { 24'h000000, signbit_reg_1488, 7'h00 };
assign \sub_7ns_7ns_7_2_1_U4.top_sub_7ns_7ns_7_2_1_Adder_1_U.ain_s0  = \sub_7ns_7ns_7_2_1_U4.top_sub_7ns_7ns_7_2_1_Adder_1_U.a ;
assign \sub_7ns_7ns_7_2_1_U4.top_sub_7ns_7ns_7_2_1_Adder_1_U.s  = { \sub_7ns_7ns_7_2_1_U4.top_sub_7ns_7ns_7_2_1_Adder_1_U.fas_s2 , \sub_7ns_7ns_7_2_1_U4.top_sub_7ns_7ns_7_2_1_Adder_1_U.sum_s1  };
assign \sub_7ns_7ns_7_2_1_U4.top_sub_7ns_7ns_7_2_1_Adder_1_U.u2.a  = \sub_7ns_7ns_7_2_1_U4.top_sub_7ns_7ns_7_2_1_Adder_1_U.ain_s1 ;
assign \sub_7ns_7ns_7_2_1_U4.top_sub_7ns_7ns_7_2_1_Adder_1_U.u2.b  = \sub_7ns_7ns_7_2_1_U4.top_sub_7ns_7ns_7_2_1_Adder_1_U.bin_s1 ;
assign \sub_7ns_7ns_7_2_1_U4.top_sub_7ns_7ns_7_2_1_Adder_1_U.u2.cin  = \sub_7ns_7ns_7_2_1_U4.top_sub_7ns_7ns_7_2_1_Adder_1_U.carry_s1 ;
assign \sub_7ns_7ns_7_2_1_U4.top_sub_7ns_7ns_7_2_1_Adder_1_U.facout_s2  = \sub_7ns_7ns_7_2_1_U4.top_sub_7ns_7ns_7_2_1_Adder_1_U.u2.cout ;
assign \sub_7ns_7ns_7_2_1_U4.top_sub_7ns_7ns_7_2_1_Adder_1_U.fas_s2  = \sub_7ns_7ns_7_2_1_U4.top_sub_7ns_7ns_7_2_1_Adder_1_U.u2.s ;
assign \sub_7ns_7ns_7_2_1_U4.top_sub_7ns_7ns_7_2_1_Adder_1_U.u1.a  = \sub_7ns_7ns_7_2_1_U4.top_sub_7ns_7ns_7_2_1_Adder_1_U.a [2:0];
assign \sub_7ns_7ns_7_2_1_U4.top_sub_7ns_7ns_7_2_1_Adder_1_U.u1.b  = \sub_7ns_7ns_7_2_1_U4.top_sub_7ns_7ns_7_2_1_Adder_1_U.bin_s0 [2:0];
assign \sub_7ns_7ns_7_2_1_U4.top_sub_7ns_7ns_7_2_1_Adder_1_U.u1.cin  = 1'h1;
assign \sub_7ns_7ns_7_2_1_U4.top_sub_7ns_7ns_7_2_1_Adder_1_U.facout_s1  = \sub_7ns_7ns_7_2_1_U4.top_sub_7ns_7ns_7_2_1_Adder_1_U.u1.cout ;
assign \sub_7ns_7ns_7_2_1_U4.top_sub_7ns_7ns_7_2_1_Adder_1_U.fas_s1  = \sub_7ns_7ns_7_2_1_U4.top_sub_7ns_7ns_7_2_1_Adder_1_U.u1.s ;
assign \sub_7ns_7ns_7_2_1_U4.top_sub_7ns_7ns_7_2_1_Adder_1_U.a  = \sub_7ns_7ns_7_2_1_U4.din0 ;
assign \sub_7ns_7ns_7_2_1_U4.top_sub_7ns_7ns_7_2_1_Adder_1_U.b  = \sub_7ns_7ns_7_2_1_U4.din1 ;
assign \sub_7ns_7ns_7_2_1_U4.top_sub_7ns_7ns_7_2_1_Adder_1_U.ce  = \sub_7ns_7ns_7_2_1_U4.ce ;
assign \sub_7ns_7ns_7_2_1_U4.top_sub_7ns_7ns_7_2_1_Adder_1_U.clk  = \sub_7ns_7ns_7_2_1_U4.clk ;
assign \sub_7ns_7ns_7_2_1_U4.top_sub_7ns_7ns_7_2_1_Adder_1_U.reset  = \sub_7ns_7ns_7_2_1_U4.reset ;
assign \sub_7ns_7ns_7_2_1_U4.dout  = \sub_7ns_7ns_7_2_1_U4.top_sub_7ns_7ns_7_2_1_Adder_1_U.s ;
assign \sub_7ns_7ns_7_2_1_U4.ce  = 1'h1;
assign \sub_7ns_7ns_7_2_1_U4.clk  = ap_clk;
assign \sub_7ns_7ns_7_2_1_U4.din0  = { 1'h0, op_0, 4'h0 };
assign \sub_7ns_7ns_7_2_1_U4.din1  = { 3'h0, signbit_reg_1488, 3'h0 };
assign grp_fu_430_p2 = \sub_7ns_7ns_7_2_1_U4.dout ;
assign \sub_7ns_7ns_7_2_1_U4.reset  = ap_rst;
assign \sub_33s_33s_33_2_1_U3.top_sub_33s_33s_33_2_1_Adder_0_U.ain_s0  = \sub_33s_33s_33_2_1_U3.top_sub_33s_33s_33_2_1_Adder_0_U.a ;
assign \sub_33s_33s_33_2_1_U3.top_sub_33s_33s_33_2_1_Adder_0_U.s  = { \sub_33s_33s_33_2_1_U3.top_sub_33s_33s_33_2_1_Adder_0_U.fas_s2 , \sub_33s_33s_33_2_1_U3.top_sub_33s_33s_33_2_1_Adder_0_U.sum_s1  };
assign \sub_33s_33s_33_2_1_U3.top_sub_33s_33s_33_2_1_Adder_0_U.u2.a  = \sub_33s_33s_33_2_1_U3.top_sub_33s_33s_33_2_1_Adder_0_U.ain_s1 ;
assign \sub_33s_33s_33_2_1_U3.top_sub_33s_33s_33_2_1_Adder_0_U.u2.b  = \sub_33s_33s_33_2_1_U3.top_sub_33s_33s_33_2_1_Adder_0_U.bin_s1 ;
assign \sub_33s_33s_33_2_1_U3.top_sub_33s_33s_33_2_1_Adder_0_U.u2.cin  = \sub_33s_33s_33_2_1_U3.top_sub_33s_33s_33_2_1_Adder_0_U.carry_s1 ;
assign \sub_33s_33s_33_2_1_U3.top_sub_33s_33s_33_2_1_Adder_0_U.facout_s2  = \sub_33s_33s_33_2_1_U3.top_sub_33s_33s_33_2_1_Adder_0_U.u2.cout ;
assign \sub_33s_33s_33_2_1_U3.top_sub_33s_33s_33_2_1_Adder_0_U.fas_s2  = \sub_33s_33s_33_2_1_U3.top_sub_33s_33s_33_2_1_Adder_0_U.u2.s ;
assign \sub_33s_33s_33_2_1_U3.top_sub_33s_33s_33_2_1_Adder_0_U.u1.a  = \sub_33s_33s_33_2_1_U3.top_sub_33s_33s_33_2_1_Adder_0_U.a [15:0];
assign \sub_33s_33s_33_2_1_U3.top_sub_33s_33s_33_2_1_Adder_0_U.u1.b  = \sub_33s_33s_33_2_1_U3.top_sub_33s_33s_33_2_1_Adder_0_U.bin_s0 [15:0];
assign \sub_33s_33s_33_2_1_U3.top_sub_33s_33s_33_2_1_Adder_0_U.u1.cin  = 1'h1;
assign \sub_33s_33s_33_2_1_U3.top_sub_33s_33s_33_2_1_Adder_0_U.facout_s1  = \sub_33s_33s_33_2_1_U3.top_sub_33s_33s_33_2_1_Adder_0_U.u1.cout ;
assign \sub_33s_33s_33_2_1_U3.top_sub_33s_33s_33_2_1_Adder_0_U.fas_s1  = \sub_33s_33s_33_2_1_U3.top_sub_33s_33s_33_2_1_Adder_0_U.u1.s ;
assign \sub_33s_33s_33_2_1_U3.top_sub_33s_33s_33_2_1_Adder_0_U.a  = \sub_33s_33s_33_2_1_U3.din0 ;
assign \sub_33s_33s_33_2_1_U3.top_sub_33s_33s_33_2_1_Adder_0_U.b  = \sub_33s_33s_33_2_1_U3.din1 ;
assign \sub_33s_33s_33_2_1_U3.top_sub_33s_33s_33_2_1_Adder_0_U.ce  = \sub_33s_33s_33_2_1_U3.ce ;
assign \sub_33s_33s_33_2_1_U3.top_sub_33s_33s_33_2_1_Adder_0_U.clk  = \sub_33s_33s_33_2_1_U3.clk ;
assign \sub_33s_33s_33_2_1_U3.top_sub_33s_33s_33_2_1_Adder_0_U.reset  = \sub_33s_33s_33_2_1_U3.reset ;
assign \sub_33s_33s_33_2_1_U3.dout  = \sub_33s_33s_33_2_1_U3.top_sub_33s_33s_33_2_1_Adder_0_U.s ;
assign \sub_33s_33s_33_2_1_U3.ce  = 1'h1;
assign \sub_33s_33s_33_2_1_U3.clk  = ap_clk;
assign \sub_33s_33s_33_2_1_U3.din0  = { op_1[15], op_1[15], op_1[15], op_1[15], op_1[15], op_1[15], op_1[15], op_1[15], op_1[15], op_1[15], op_1[15], op_1, 6'h00 };
assign \sub_33s_33s_33_2_1_U3.din1  = { op_6[31], op_6 };
assign grp_fu_309_p2 = \sub_33s_33s_33_2_1_U3.dout ;
assign \sub_33s_33s_33_2_1_U3.reset  = ap_rst;
assign \mul_8s_3ns_11_7_1_U1.top_mul_8s_3ns_11_7_1_Mul_DSP_0_U.p  = \mul_8s_3ns_11_7_1_U1.top_mul_8s_3ns_11_7_1_Mul_DSP_0_U.buff4 ;
assign \mul_8s_3ns_11_7_1_U1.top_mul_8s_3ns_11_7_1_Mul_DSP_0_U.a  = \mul_8s_3ns_11_7_1_U1.din0 ;
assign \mul_8s_3ns_11_7_1_U1.top_mul_8s_3ns_11_7_1_Mul_DSP_0_U.b  = \mul_8s_3ns_11_7_1_U1.din1 ;
assign \mul_8s_3ns_11_7_1_U1.top_mul_8s_3ns_11_7_1_Mul_DSP_0_U.ce  = \mul_8s_3ns_11_7_1_U1.ce ;
assign \mul_8s_3ns_11_7_1_U1.top_mul_8s_3ns_11_7_1_Mul_DSP_0_U.clk  = \mul_8s_3ns_11_7_1_U1.clk ;
assign \mul_8s_3ns_11_7_1_U1.dout  = \mul_8s_3ns_11_7_1_U1.top_mul_8s_3ns_11_7_1_Mul_DSP_0_U.p ;
assign \mul_8s_3ns_11_7_1_U1.ce  = 1'h1;
assign \mul_8s_3ns_11_7_1_U1.clk  = ap_clk;
assign \mul_8s_3ns_11_7_1_U1.din0  = op_4;
assign \mul_8s_3ns_11_7_1_U1.din1  = { op_0, 1'h0 };
assign grp_fu_255_p2 = \mul_8s_3ns_11_7_1_U1.dout ;
assign \mul_8s_3ns_11_7_1_U1.reset  = ap_rst;
assign \mul_8ns_8s_16_7_1_U2.top_mul_8ns_8s_16_7_1_Mul_DSP_1_U.p  = \mul_8ns_8s_16_7_1_U2.top_mul_8ns_8s_16_7_1_Mul_DSP_1_U.buff4 ;
assign \mul_8ns_8s_16_7_1_U2.top_mul_8ns_8s_16_7_1_Mul_DSP_1_U.a  = \mul_8ns_8s_16_7_1_U2.din0 ;
assign \mul_8ns_8s_16_7_1_U2.top_mul_8ns_8s_16_7_1_Mul_DSP_1_U.b  = \mul_8ns_8s_16_7_1_U2.din1 ;
assign \mul_8ns_8s_16_7_1_U2.top_mul_8ns_8s_16_7_1_Mul_DSP_1_U.ce  = \mul_8ns_8s_16_7_1_U2.ce ;
assign \mul_8ns_8s_16_7_1_U2.top_mul_8ns_8s_16_7_1_Mul_DSP_1_U.clk  = \mul_8ns_8s_16_7_1_U2.clk ;
assign \mul_8ns_8s_16_7_1_U2.dout  = \mul_8ns_8s_16_7_1_U2.top_mul_8ns_8s_16_7_1_Mul_DSP_1_U.p ;
assign \mul_8ns_8s_16_7_1_U2.ce  = 1'h1;
assign \mul_8ns_8s_16_7_1_U2.clk  = ap_clk;
assign \mul_8ns_8s_16_7_1_U2.din0  = op_8;
assign \mul_8ns_8s_16_7_1_U2.din1  = op_4;
assign grp_fu_268_p2 = \mul_8ns_8s_16_7_1_U2.dout ;
assign \mul_8ns_8s_16_7_1_U2.reset  = ap_rst;
assign \mul_4ns_4s_8_7_1_U14.top_mul_4ns_4s_8_7_1_Mul_DSP_2_U.p  = \mul_4ns_4s_8_7_1_U14.top_mul_4ns_4s_8_7_1_Mul_DSP_2_U.buff4 ;
assign \mul_4ns_4s_8_7_1_U14.top_mul_4ns_4s_8_7_1_Mul_DSP_2_U.a  = \mul_4ns_4s_8_7_1_U14.din0 ;
assign \mul_4ns_4s_8_7_1_U14.top_mul_4ns_4s_8_7_1_Mul_DSP_2_U.b  = \mul_4ns_4s_8_7_1_U14.din1 ;
assign \mul_4ns_4s_8_7_1_U14.top_mul_4ns_4s_8_7_1_Mul_DSP_2_U.ce  = \mul_4ns_4s_8_7_1_U14.ce ;
assign \mul_4ns_4s_8_7_1_U14.top_mul_4ns_4s_8_7_1_Mul_DSP_2_U.clk  = \mul_4ns_4s_8_7_1_U14.clk ;
assign \mul_4ns_4s_8_7_1_U14.dout  = \mul_4ns_4s_8_7_1_U14.top_mul_4ns_4s_8_7_1_Mul_DSP_2_U.p ;
assign \mul_4ns_4s_8_7_1_U14.ce  = 1'h1;
assign \mul_4ns_4s_8_7_1_U14.clk  = ap_clk;
assign \mul_4ns_4s_8_7_1_U14.din0  = zext_ln1116_reg_1819[3:0];
assign \mul_4ns_4s_8_7_1_U14.din1  = op_9_V_reg_1977;
assign grp_fu_1236_p2 = \mul_4ns_4s_8_7_1_U14.dout ;
assign \mul_4ns_4s_8_7_1_U14.reset  = ap_rst;
assign \add_6ns_6ns_6_2_1_U19.top_add_6ns_6ns_6_2_1_Adder_13_U.ain_s0  = \add_6ns_6ns_6_2_1_U19.top_add_6ns_6ns_6_2_1_Adder_13_U.a ;
assign \add_6ns_6ns_6_2_1_U19.top_add_6ns_6ns_6_2_1_Adder_13_U.bin_s0  = \add_6ns_6ns_6_2_1_U19.top_add_6ns_6ns_6_2_1_Adder_13_U.b ;
assign \add_6ns_6ns_6_2_1_U19.top_add_6ns_6ns_6_2_1_Adder_13_U.s  = { \add_6ns_6ns_6_2_1_U19.top_add_6ns_6ns_6_2_1_Adder_13_U.fas_s2 , \add_6ns_6ns_6_2_1_U19.top_add_6ns_6ns_6_2_1_Adder_13_U.sum_s1  };
assign \add_6ns_6ns_6_2_1_U19.top_add_6ns_6ns_6_2_1_Adder_13_U.u2.a  = \add_6ns_6ns_6_2_1_U19.top_add_6ns_6ns_6_2_1_Adder_13_U.ain_s1 ;
assign \add_6ns_6ns_6_2_1_U19.top_add_6ns_6ns_6_2_1_Adder_13_U.u2.b  = \add_6ns_6ns_6_2_1_U19.top_add_6ns_6ns_6_2_1_Adder_13_U.bin_s1 ;
assign \add_6ns_6ns_6_2_1_U19.top_add_6ns_6ns_6_2_1_Adder_13_U.u2.cin  = \add_6ns_6ns_6_2_1_U19.top_add_6ns_6ns_6_2_1_Adder_13_U.carry_s1 ;
assign \add_6ns_6ns_6_2_1_U19.top_add_6ns_6ns_6_2_1_Adder_13_U.facout_s2  = \add_6ns_6ns_6_2_1_U19.top_add_6ns_6ns_6_2_1_Adder_13_U.u2.cout ;
assign \add_6ns_6ns_6_2_1_U19.top_add_6ns_6ns_6_2_1_Adder_13_U.fas_s2  = \add_6ns_6ns_6_2_1_U19.top_add_6ns_6ns_6_2_1_Adder_13_U.u2.s ;
assign \add_6ns_6ns_6_2_1_U19.top_add_6ns_6ns_6_2_1_Adder_13_U.u1.a  = \add_6ns_6ns_6_2_1_U19.top_add_6ns_6ns_6_2_1_Adder_13_U.a [2:0];
assign \add_6ns_6ns_6_2_1_U19.top_add_6ns_6ns_6_2_1_Adder_13_U.u1.b  = \add_6ns_6ns_6_2_1_U19.top_add_6ns_6ns_6_2_1_Adder_13_U.b [2:0];
assign \add_6ns_6ns_6_2_1_U19.top_add_6ns_6ns_6_2_1_Adder_13_U.u1.cin  = 1'h0;
assign \add_6ns_6ns_6_2_1_U19.top_add_6ns_6ns_6_2_1_Adder_13_U.facout_s1  = \add_6ns_6ns_6_2_1_U19.top_add_6ns_6ns_6_2_1_Adder_13_U.u1.cout ;
assign \add_6ns_6ns_6_2_1_U19.top_add_6ns_6ns_6_2_1_Adder_13_U.fas_s1  = \add_6ns_6ns_6_2_1_U19.top_add_6ns_6ns_6_2_1_Adder_13_U.u1.s ;
assign \add_6ns_6ns_6_2_1_U19.top_add_6ns_6ns_6_2_1_Adder_13_U.a  = \add_6ns_6ns_6_2_1_U19.din0 ;
assign \add_6ns_6ns_6_2_1_U19.top_add_6ns_6ns_6_2_1_Adder_13_U.b  = \add_6ns_6ns_6_2_1_U19.din1 ;
assign \add_6ns_6ns_6_2_1_U19.top_add_6ns_6ns_6_2_1_Adder_13_U.ce  = \add_6ns_6ns_6_2_1_U19.ce ;
assign \add_6ns_6ns_6_2_1_U19.top_add_6ns_6ns_6_2_1_Adder_13_U.clk  = \add_6ns_6ns_6_2_1_U19.clk ;
assign \add_6ns_6ns_6_2_1_U19.top_add_6ns_6ns_6_2_1_Adder_13_U.reset  = \add_6ns_6ns_6_2_1_U19.reset ;
assign \add_6ns_6ns_6_2_1_U19.dout  = \add_6ns_6ns_6_2_1_U19.top_add_6ns_6ns_6_2_1_Adder_13_U.s ;
assign \add_6ns_6ns_6_2_1_U19.ce  = 1'h1;
assign \add_6ns_6ns_6_2_1_U19.clk  = ap_clk;
assign \add_6ns_6ns_6_2_1_U19.din0  = ret_V_7_reg_2090;
assign \add_6ns_6ns_6_2_1_U19.din1  = 6'h01;
assign grp_fu_1372_p2 = \add_6ns_6ns_6_2_1_U19.dout ;
assign \add_6ns_6ns_6_2_1_U19.reset  = ap_rst;
assign \add_5s_5s_5_2_1_U16.top_add_5s_5s_5_2_1_Adder_10_U.ain_s0  = \add_5s_5s_5_2_1_U16.top_add_5s_5s_5_2_1_Adder_10_U.a ;
assign \add_5s_5s_5_2_1_U16.top_add_5s_5s_5_2_1_Adder_10_U.bin_s0  = \add_5s_5s_5_2_1_U16.top_add_5s_5s_5_2_1_Adder_10_U.b ;
assign \add_5s_5s_5_2_1_U16.top_add_5s_5s_5_2_1_Adder_10_U.s  = { \add_5s_5s_5_2_1_U16.top_add_5s_5s_5_2_1_Adder_10_U.fas_s2 , \add_5s_5s_5_2_1_U16.top_add_5s_5s_5_2_1_Adder_10_U.sum_s1  };
assign \add_5s_5s_5_2_1_U16.top_add_5s_5s_5_2_1_Adder_10_U.u2.a  = \add_5s_5s_5_2_1_U16.top_add_5s_5s_5_2_1_Adder_10_U.ain_s1 ;
assign \add_5s_5s_5_2_1_U16.top_add_5s_5s_5_2_1_Adder_10_U.u2.b  = \add_5s_5s_5_2_1_U16.top_add_5s_5s_5_2_1_Adder_10_U.bin_s1 ;
assign \add_5s_5s_5_2_1_U16.top_add_5s_5s_5_2_1_Adder_10_U.u2.cin  = \add_5s_5s_5_2_1_U16.top_add_5s_5s_5_2_1_Adder_10_U.carry_s1 ;
assign \add_5s_5s_5_2_1_U16.top_add_5s_5s_5_2_1_Adder_10_U.facout_s2  = \add_5s_5s_5_2_1_U16.top_add_5s_5s_5_2_1_Adder_10_U.u2.cout ;
assign \add_5s_5s_5_2_1_U16.top_add_5s_5s_5_2_1_Adder_10_U.fas_s2  = \add_5s_5s_5_2_1_U16.top_add_5s_5s_5_2_1_Adder_10_U.u2.s ;
assign \add_5s_5s_5_2_1_U16.top_add_5s_5s_5_2_1_Adder_10_U.u1.a  = \add_5s_5s_5_2_1_U16.top_add_5s_5s_5_2_1_Adder_10_U.a [1:0];
assign \add_5s_5s_5_2_1_U16.top_add_5s_5s_5_2_1_Adder_10_U.u1.b  = \add_5s_5s_5_2_1_U16.top_add_5s_5s_5_2_1_Adder_10_U.b [1:0];
assign \add_5s_5s_5_2_1_U16.top_add_5s_5s_5_2_1_Adder_10_U.u1.cin  = 1'h0;
assign \add_5s_5s_5_2_1_U16.top_add_5s_5s_5_2_1_Adder_10_U.facout_s1  = \add_5s_5s_5_2_1_U16.top_add_5s_5s_5_2_1_Adder_10_U.u1.cout ;
assign \add_5s_5s_5_2_1_U16.top_add_5s_5s_5_2_1_Adder_10_U.fas_s1  = \add_5s_5s_5_2_1_U16.top_add_5s_5s_5_2_1_Adder_10_U.u1.s ;
assign \add_5s_5s_5_2_1_U16.top_add_5s_5s_5_2_1_Adder_10_U.a  = \add_5s_5s_5_2_1_U16.din0 ;
assign \add_5s_5s_5_2_1_U16.top_add_5s_5s_5_2_1_Adder_10_U.b  = \add_5s_5s_5_2_1_U16.din1 ;
assign \add_5s_5s_5_2_1_U16.top_add_5s_5s_5_2_1_Adder_10_U.ce  = \add_5s_5s_5_2_1_U16.ce ;
assign \add_5s_5s_5_2_1_U16.top_add_5s_5s_5_2_1_Adder_10_U.clk  = \add_5s_5s_5_2_1_U16.clk ;
assign \add_5s_5s_5_2_1_U16.top_add_5s_5s_5_2_1_Adder_10_U.reset  = \add_5s_5s_5_2_1_U16.reset ;
assign \add_5s_5s_5_2_1_U16.dout  = \add_5s_5s_5_2_1_U16.top_add_5s_5s_5_2_1_Adder_10_U.s ;
assign \add_5s_5s_5_2_1_U16.ce  = 1'h1;
assign \add_5s_5s_5_2_1_U16.clk  = ap_clk;
assign \add_5s_5s_5_2_1_U16.din0  = { add_ln69_1_reg_2028[2], add_ln69_1_reg_2028[2], add_ln69_1_reg_2028 };
assign \add_5s_5s_5_2_1_U16.din1  = { op_16_V_reg_2003[3], op_16_V_reg_2003 };
assign grp_fu_1282_p2 = \add_5s_5s_5_2_1_U16.dout ;
assign \add_5s_5s_5_2_1_U16.reset  = ap_rst;
assign \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.ain_s0  = \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.a ;
assign \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.bin_s0  = \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.b ;
assign \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.s  = { \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.fas_s2 , \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.sum_s1  };
assign \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.u2.a  = \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.ain_s1 ;
assign \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.u2.b  = \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.bin_s1 ;
assign \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.u2.cin  = \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.carry_s1 ;
assign \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.facout_s2  = \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.u2.cout ;
assign \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.fas_s2  = \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.u2.s ;
assign \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.u1.a  = \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.a [1:0];
assign \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.u1.b  = \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.b [1:0];
assign \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.u1.cin  = 1'h0;
assign \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.facout_s1  = \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.u1.cout ;
assign \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.fas_s1  = \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.u1.s ;
assign \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.a  = \add_4ns_4ns_4_2_1_U9.din0 ;
assign \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.b  = \add_4ns_4ns_4_2_1_U9.din1 ;
assign \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.ce  = \add_4ns_4ns_4_2_1_U9.ce ;
assign \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.clk  = \add_4ns_4ns_4_2_1_U9.clk ;
assign \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.reset  = \add_4ns_4ns_4_2_1_U9.reset ;
assign \add_4ns_4ns_4_2_1_U9.dout  = \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.s ;
assign \add_4ns_4ns_4_2_1_U9.ce  = 1'h1;
assign \add_4ns_4ns_4_2_1_U9.clk  = ap_clk;
assign \add_4ns_4ns_4_2_1_U9.din0  = p_Val2_6_reg_1543;
assign \add_4ns_4ns_4_2_1_U9.din1  = { 3'h0, and_ln408_reg_1718 };
assign grp_fu_660_p2 = \add_4ns_4ns_4_2_1_U9.dout ;
assign \add_4ns_4ns_4_2_1_U9.reset  = ap_rst;
assign \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_4_U.ain_s0  = \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_4_U.a ;
assign \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_4_U.bin_s0  = \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_4_U.b ;
assign \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_4_U.s  = { \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_4_U.fas_s2 , \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_4_U.sum_s1  };
assign \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_4_U.u2.a  = \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_4_U.ain_s1 ;
assign \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_4_U.u2.b  = \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_4_U.bin_s1 ;
assign \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_4_U.u2.cin  = \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_4_U.carry_s1 ;
assign \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_4_U.facout_s2  = \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_4_U.u2.cout ;
assign \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_4_U.fas_s2  = \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_4_U.u2.s ;
assign \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_4_U.u1.a  = \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_4_U.a [1:0];
assign \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_4_U.u1.b  = \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_4_U.b [1:0];
assign \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_4_U.u1.cin  = 1'h0;
assign \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_4_U.facout_s1  = \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_4_U.u1.cout ;
assign \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_4_U.fas_s1  = \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_4_U.u1.s ;
assign \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_4_U.a  = \add_4ns_4ns_4_2_1_U8.din0 ;
assign \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_4_U.b  = \add_4ns_4ns_4_2_1_U8.din1 ;
assign \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_4_U.ce  = \add_4ns_4ns_4_2_1_U8.ce ;
assign \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_4_U.clk  = \add_4ns_4ns_4_2_1_U8.clk ;
assign \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_4_U.reset  = \add_4ns_4ns_4_2_1_U8.reset ;
assign \add_4ns_4ns_4_2_1_U8.dout  = \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_4_U.s ;
assign \add_4ns_4ns_4_2_1_U8.ce  = 1'h1;
assign \add_4ns_4ns_4_2_1_U8.clk  = ap_clk;
assign \add_4ns_4ns_4_2_1_U8.din0  = p_Val2_2_reg_1610;
assign \add_4ns_4ns_4_2_1_U8.din1  = { 3'h0, and_ln406_reg_1696 };
assign grp_fu_652_p2 = \add_4ns_4ns_4_2_1_U8.dout ;
assign \add_4ns_4ns_4_2_1_U8.reset  = ap_rst;
assign \add_4ns_4ns_4_2_1_U7.top_add_4ns_4ns_4_2_1_Adder_4_U.ain_s0  = \add_4ns_4ns_4_2_1_U7.top_add_4ns_4ns_4_2_1_Adder_4_U.a ;
assign \add_4ns_4ns_4_2_1_U7.top_add_4ns_4ns_4_2_1_Adder_4_U.bin_s0  = \add_4ns_4ns_4_2_1_U7.top_add_4ns_4ns_4_2_1_Adder_4_U.b ;
assign \add_4ns_4ns_4_2_1_U7.top_add_4ns_4ns_4_2_1_Adder_4_U.s  = { \add_4ns_4ns_4_2_1_U7.top_add_4ns_4ns_4_2_1_Adder_4_U.fas_s2 , \add_4ns_4ns_4_2_1_U7.top_add_4ns_4ns_4_2_1_Adder_4_U.sum_s1  };
assign \add_4ns_4ns_4_2_1_U7.top_add_4ns_4ns_4_2_1_Adder_4_U.u2.a  = \add_4ns_4ns_4_2_1_U7.top_add_4ns_4ns_4_2_1_Adder_4_U.ain_s1 ;
assign \add_4ns_4ns_4_2_1_U7.top_add_4ns_4ns_4_2_1_Adder_4_U.u2.b  = \add_4ns_4ns_4_2_1_U7.top_add_4ns_4ns_4_2_1_Adder_4_U.bin_s1 ;
assign \add_4ns_4ns_4_2_1_U7.top_add_4ns_4ns_4_2_1_Adder_4_U.u2.cin  = \add_4ns_4ns_4_2_1_U7.top_add_4ns_4ns_4_2_1_Adder_4_U.carry_s1 ;
assign \add_4ns_4ns_4_2_1_U7.top_add_4ns_4ns_4_2_1_Adder_4_U.facout_s2  = \add_4ns_4ns_4_2_1_U7.top_add_4ns_4ns_4_2_1_Adder_4_U.u2.cout ;
assign \add_4ns_4ns_4_2_1_U7.top_add_4ns_4ns_4_2_1_Adder_4_U.fas_s2  = \add_4ns_4ns_4_2_1_U7.top_add_4ns_4ns_4_2_1_Adder_4_U.u2.s ;
assign \add_4ns_4ns_4_2_1_U7.top_add_4ns_4ns_4_2_1_Adder_4_U.u1.a  = \add_4ns_4ns_4_2_1_U7.top_add_4ns_4ns_4_2_1_Adder_4_U.a [1:0];
assign \add_4ns_4ns_4_2_1_U7.top_add_4ns_4ns_4_2_1_Adder_4_U.u1.b  = \add_4ns_4ns_4_2_1_U7.top_add_4ns_4ns_4_2_1_Adder_4_U.b [1:0];
assign \add_4ns_4ns_4_2_1_U7.top_add_4ns_4ns_4_2_1_Adder_4_U.u1.cin  = 1'h0;
assign \add_4ns_4ns_4_2_1_U7.top_add_4ns_4ns_4_2_1_Adder_4_U.facout_s1  = \add_4ns_4ns_4_2_1_U7.top_add_4ns_4ns_4_2_1_Adder_4_U.u1.cout ;
assign \add_4ns_4ns_4_2_1_U7.top_add_4ns_4ns_4_2_1_Adder_4_U.fas_s1  = \add_4ns_4ns_4_2_1_U7.top_add_4ns_4ns_4_2_1_Adder_4_U.u1.s ;
assign \add_4ns_4ns_4_2_1_U7.top_add_4ns_4ns_4_2_1_Adder_4_U.a  = \add_4ns_4ns_4_2_1_U7.din0 ;
assign \add_4ns_4ns_4_2_1_U7.top_add_4ns_4ns_4_2_1_Adder_4_U.b  = \add_4ns_4ns_4_2_1_U7.din1 ;
assign \add_4ns_4ns_4_2_1_U7.top_add_4ns_4ns_4_2_1_Adder_4_U.ce  = \add_4ns_4ns_4_2_1_U7.ce ;
assign \add_4ns_4ns_4_2_1_U7.top_add_4ns_4ns_4_2_1_Adder_4_U.clk  = \add_4ns_4ns_4_2_1_U7.clk ;
assign \add_4ns_4ns_4_2_1_U7.top_add_4ns_4ns_4_2_1_Adder_4_U.reset  = \add_4ns_4ns_4_2_1_U7.reset ;
assign \add_4ns_4ns_4_2_1_U7.dout  = \add_4ns_4ns_4_2_1_U7.top_add_4ns_4ns_4_2_1_Adder_4_U.s ;
assign \add_4ns_4ns_4_2_1_U7.ce  = 1'h1;
assign \add_4ns_4ns_4_2_1_U7.clk  = ap_clk;
assign \add_4ns_4ns_4_2_1_U7.din0  = ret_V_6_cast_reg_1664;
assign \add_4ns_4ns_4_2_1_U7.din1  = 4'h1;
assign grp_fu_615_p2 = \add_4ns_4ns_4_2_1_U7.dout ;
assign \add_4ns_4ns_4_2_1_U7.reset  = ap_rst;
assign \add_46s_46s_46_2_1_U18.top_add_46s_46s_46_2_1_Adder_12_U.ain_s0  = \add_46s_46s_46_2_1_U18.top_add_46s_46s_46_2_1_Adder_12_U.a ;
assign \add_46s_46s_46_2_1_U18.top_add_46s_46s_46_2_1_Adder_12_U.bin_s0  = \add_46s_46s_46_2_1_U18.top_add_46s_46s_46_2_1_Adder_12_U.b ;
assign \add_46s_46s_46_2_1_U18.top_add_46s_46s_46_2_1_Adder_12_U.s  = { \add_46s_46s_46_2_1_U18.top_add_46s_46s_46_2_1_Adder_12_U.fas_s2 , \add_46s_46s_46_2_1_U18.top_add_46s_46s_46_2_1_Adder_12_U.sum_s1  };
assign \add_46s_46s_46_2_1_U18.top_add_46s_46s_46_2_1_Adder_12_U.u2.a  = \add_46s_46s_46_2_1_U18.top_add_46s_46s_46_2_1_Adder_12_U.ain_s1 ;
assign \add_46s_46s_46_2_1_U18.top_add_46s_46s_46_2_1_Adder_12_U.u2.b  = \add_46s_46s_46_2_1_U18.top_add_46s_46s_46_2_1_Adder_12_U.bin_s1 ;
assign \add_46s_46s_46_2_1_U18.top_add_46s_46s_46_2_1_Adder_12_U.u2.cin  = \add_46s_46s_46_2_1_U18.top_add_46s_46s_46_2_1_Adder_12_U.carry_s1 ;
assign \add_46s_46s_46_2_1_U18.top_add_46s_46s_46_2_1_Adder_12_U.facout_s2  = \add_46s_46s_46_2_1_U18.top_add_46s_46s_46_2_1_Adder_12_U.u2.cout ;
assign \add_46s_46s_46_2_1_U18.top_add_46s_46s_46_2_1_Adder_12_U.fas_s2  = \add_46s_46s_46_2_1_U18.top_add_46s_46s_46_2_1_Adder_12_U.u2.s ;
assign \add_46s_46s_46_2_1_U18.top_add_46s_46s_46_2_1_Adder_12_U.u1.a  = \add_46s_46s_46_2_1_U18.top_add_46s_46s_46_2_1_Adder_12_U.a [22:0];
assign \add_46s_46s_46_2_1_U18.top_add_46s_46s_46_2_1_Adder_12_U.u1.b  = \add_46s_46s_46_2_1_U18.top_add_46s_46s_46_2_1_Adder_12_U.b [22:0];
assign \add_46s_46s_46_2_1_U18.top_add_46s_46s_46_2_1_Adder_12_U.u1.cin  = 1'h0;
assign \add_46s_46s_46_2_1_U18.top_add_46s_46s_46_2_1_Adder_12_U.facout_s1  = \add_46s_46s_46_2_1_U18.top_add_46s_46s_46_2_1_Adder_12_U.u1.cout ;
assign \add_46s_46s_46_2_1_U18.top_add_46s_46s_46_2_1_Adder_12_U.fas_s1  = \add_46s_46s_46_2_1_U18.top_add_46s_46s_46_2_1_Adder_12_U.u1.s ;
assign \add_46s_46s_46_2_1_U18.top_add_46s_46s_46_2_1_Adder_12_U.a  = \add_46s_46s_46_2_1_U18.din0 ;
assign \add_46s_46s_46_2_1_U18.top_add_46s_46s_46_2_1_Adder_12_U.b  = \add_46s_46s_46_2_1_U18.din1 ;
assign \add_46s_46s_46_2_1_U18.top_add_46s_46s_46_2_1_Adder_12_U.ce  = \add_46s_46s_46_2_1_U18.ce ;
assign \add_46s_46s_46_2_1_U18.top_add_46s_46s_46_2_1_Adder_12_U.clk  = \add_46s_46s_46_2_1_U18.clk ;
assign \add_46s_46s_46_2_1_U18.top_add_46s_46s_46_2_1_Adder_12_U.reset  = \add_46s_46s_46_2_1_U18.reset ;
assign \add_46s_46s_46_2_1_U18.dout  = \add_46s_46s_46_2_1_U18.top_add_46s_46s_46_2_1_Adder_12_U.s ;
assign \add_46s_46s_46_2_1_U18.ce  = 1'h1;
assign \add_46s_46s_46_2_1_U18.clk  = ap_clk;
assign \add_46s_46s_46_2_1_U18.din0  = { select_ln353_1_reg_2065[31], select_ln353_1_reg_2065, 13'h0000 };
assign \add_46s_46s_46_2_1_U18.din1  = { op_15[15], op_15[15], op_15[15], op_15[15], op_15[15], op_15[15], op_15[15], op_15[15], op_15[15], op_15[15], op_15[15], op_15[15], op_15[15], op_15[15], op_15[15], op_15[15], op_15[15], op_15[15], op_15[15], op_15[15], op_15[15], op_15[15], op_15[15], op_15[15], op_15[15], op_15[15], op_15[15], op_15[15], op_15[15], op_15[15], op_15 };
assign grp_fu_1327_p2 = \add_46s_46s_46_2_1_U18.dout ;
assign \add_46s_46s_46_2_1_U18.reset  = ap_rst;
assign \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_8_U.ain_s0  = \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_8_U.a ;
assign \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_8_U.bin_s0  = \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_8_U.b ;
assign \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_8_U.s  = { \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_8_U.fas_s2 , \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_8_U.sum_s1  };
assign \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_8_U.u2.a  = \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_8_U.ain_s1 ;
assign \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_8_U.u2.b  = \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_8_U.bin_s1 ;
assign \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_8_U.u2.cin  = \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_8_U.carry_s1 ;
assign \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_8_U.facout_s2  = \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_8_U.u2.cout ;
assign \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_8_U.fas_s2  = \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_8_U.u2.s ;
assign \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_8_U.u1.a  = \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_8_U.a [0];
assign \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_8_U.u1.b  = \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_8_U.b [0];
assign \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_8_U.u1.cin  = 1'h0;
assign \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_8_U.facout_s1  = \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_8_U.u1.cout ;
assign \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_8_U.fas_s1  = \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_8_U.u1.s ;
assign \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_8_U.a  = \add_3s_3ns_3_2_1_U13.din0 ;
assign \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_8_U.b  = \add_3s_3ns_3_2_1_U13.din1 ;
assign \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_8_U.ce  = \add_3s_3ns_3_2_1_U13.ce ;
assign \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_8_U.clk  = \add_3s_3ns_3_2_1_U13.clk ;
assign \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_8_U.reset  = \add_3s_3ns_3_2_1_U13.reset ;
assign \add_3s_3ns_3_2_1_U13.dout  = \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_8_U.s ;
assign \add_3s_3ns_3_2_1_U13.ce  = 1'h1;
assign \add_3s_3ns_3_2_1_U13.clk  = ap_clk;
assign \add_3s_3ns_3_2_1_U13.din0  = { ret_V_19_reg_1740[1], ret_V_19_reg_1740 };
assign \add_3s_3ns_3_2_1_U13.din1  = { 2'h0, icmp_ln874_reg_1824 };
assign grp_fu_1201_p2 = \add_3s_3ns_3_2_1_U13.dout ;
assign \add_3s_3ns_3_2_1_U13.reset  = ap_rst;
assign \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.ain_s0  = \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.a ;
assign \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.bin_s0  = \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.b ;
assign \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.s  = { \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.fas_s2 , \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.sum_s1  };
assign \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.u2.a  = \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.ain_s1 ;
assign \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.u2.b  = \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.bin_s1 ;
assign \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.u2.cin  = \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.carry_s1 ;
assign \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.facout_s2  = \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.u2.cout ;
assign \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.fas_s2  = \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.u2.s ;
assign \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.u1.a  = \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.a [16:0];
assign \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.u1.b  = \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.b [16:0];
assign \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.u1.cin  = 1'h0;
assign \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.facout_s1  = \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.u1.cout ;
assign \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.fas_s1  = \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.u1.s ;
assign \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.a  = \add_35s_35s_35_2_1_U15.din0 ;
assign \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.b  = \add_35s_35s_35_2_1_U15.din1 ;
assign \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.ce  = \add_35s_35s_35_2_1_U15.ce ;
assign \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.clk  = \add_35s_35s_35_2_1_U15.clk ;
assign \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.reset  = \add_35s_35s_35_2_1_U15.reset ;
assign \add_35s_35s_35_2_1_U15.dout  = \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.s ;
assign \add_35s_35s_35_2_1_U15.ce  = 1'h1;
assign \add_35s_35s_35_2_1_U15.clk  = ap_clk;
assign \add_35s_35s_35_2_1_U15.din0  = { select_ln353_reg_1983[18], select_ln353_reg_1983[18], select_ln353_reg_1983[18], select_ln353_reg_1983[18], select_ln353_reg_1983[18], select_ln353_reg_1983[18], select_ln353_reg_1983[18], select_ln353_reg_1983[18], select_ln353_reg_1983[18], select_ln353_reg_1983[18], select_ln353_reg_1983[18], select_ln353_reg_1983[18], select_ln353_reg_1983[18], select_ln353_reg_1983[18], select_ln353_reg_1983, 2'h0 };
assign \add_35s_35s_35_2_1_U15.din1  = { op_14_V_reg_1972[3], op_14_V_reg_1972[3], op_14_V_reg_1972[3], op_14_V_reg_1972[3], op_14_V_reg_1972[3], op_14_V_reg_1972[3], op_14_V_reg_1972[3], op_14_V_reg_1972[3], op_14_V_reg_1972[3], op_14_V_reg_1972[3], op_14_V_reg_1972[3], op_14_V_reg_1972[3], op_14_V_reg_1972[3], op_14_V_reg_1972[3], op_14_V_reg_1972[3], op_14_V_reg_1972[3], op_14_V_reg_1972[3], op_14_V_reg_1972[3], op_14_V_reg_1972[3], op_14_V_reg_1972[3], op_14_V_reg_1972[3], op_14_V_reg_1972[3], op_14_V_reg_1972[3], op_14_V_reg_1972[3], op_14_V_reg_1972[3], op_14_V_reg_1972[3], op_14_V_reg_1972[3], op_14_V_reg_1972[3], op_14_V_reg_1972[3], op_14_V_reg_1972[3], op_14_V_reg_1972[3], op_14_V_reg_1972 };
assign grp_fu_1255_p2 = \add_35s_35s_35_2_1_U15.dout ;
assign \add_35s_35s_35_2_1_U15.reset  = ap_rst;
assign \add_33ns_33s_33_2_1_U6.top_add_33ns_33s_33_2_1_Adder_3_U.ain_s0  = \add_33ns_33s_33_2_1_U6.top_add_33ns_33s_33_2_1_Adder_3_U.a ;
assign \add_33ns_33s_33_2_1_U6.top_add_33ns_33s_33_2_1_Adder_3_U.bin_s0  = \add_33ns_33s_33_2_1_U6.top_add_33ns_33s_33_2_1_Adder_3_U.b ;
assign \add_33ns_33s_33_2_1_U6.top_add_33ns_33s_33_2_1_Adder_3_U.s  = { \add_33ns_33s_33_2_1_U6.top_add_33ns_33s_33_2_1_Adder_3_U.fas_s2 , \add_33ns_33s_33_2_1_U6.top_add_33ns_33s_33_2_1_Adder_3_U.sum_s1  };
assign \add_33ns_33s_33_2_1_U6.top_add_33ns_33s_33_2_1_Adder_3_U.u2.a  = \add_33ns_33s_33_2_1_U6.top_add_33ns_33s_33_2_1_Adder_3_U.ain_s1 ;
assign \add_33ns_33s_33_2_1_U6.top_add_33ns_33s_33_2_1_Adder_3_U.u2.b  = \add_33ns_33s_33_2_1_U6.top_add_33ns_33s_33_2_1_Adder_3_U.bin_s1 ;
assign \add_33ns_33s_33_2_1_U6.top_add_33ns_33s_33_2_1_Adder_3_U.u2.cin  = \add_33ns_33s_33_2_1_U6.top_add_33ns_33s_33_2_1_Adder_3_U.carry_s1 ;
assign \add_33ns_33s_33_2_1_U6.top_add_33ns_33s_33_2_1_Adder_3_U.facout_s2  = \add_33ns_33s_33_2_1_U6.top_add_33ns_33s_33_2_1_Adder_3_U.u2.cout ;
assign \add_33ns_33s_33_2_1_U6.top_add_33ns_33s_33_2_1_Adder_3_U.fas_s2  = \add_33ns_33s_33_2_1_U6.top_add_33ns_33s_33_2_1_Adder_3_U.u2.s ;
assign \add_33ns_33s_33_2_1_U6.top_add_33ns_33s_33_2_1_Adder_3_U.u1.a  = \add_33ns_33s_33_2_1_U6.top_add_33ns_33s_33_2_1_Adder_3_U.a [15:0];
assign \add_33ns_33s_33_2_1_U6.top_add_33ns_33s_33_2_1_Adder_3_U.u1.b  = \add_33ns_33s_33_2_1_U6.top_add_33ns_33s_33_2_1_Adder_3_U.b [15:0];
assign \add_33ns_33s_33_2_1_U6.top_add_33ns_33s_33_2_1_Adder_3_U.u1.cin  = 1'h0;
assign \add_33ns_33s_33_2_1_U6.top_add_33ns_33s_33_2_1_Adder_3_U.facout_s1  = \add_33ns_33s_33_2_1_U6.top_add_33ns_33s_33_2_1_Adder_3_U.u1.cout ;
assign \add_33ns_33s_33_2_1_U6.top_add_33ns_33s_33_2_1_Adder_3_U.fas_s1  = \add_33ns_33s_33_2_1_U6.top_add_33ns_33s_33_2_1_Adder_3_U.u1.s ;
assign \add_33ns_33s_33_2_1_U6.top_add_33ns_33s_33_2_1_Adder_3_U.a  = \add_33ns_33s_33_2_1_U6.din0 ;
assign \add_33ns_33s_33_2_1_U6.top_add_33ns_33s_33_2_1_Adder_3_U.b  = \add_33ns_33s_33_2_1_U6.din1 ;
assign \add_33ns_33s_33_2_1_U6.top_add_33ns_33s_33_2_1_Adder_3_U.ce  = \add_33ns_33s_33_2_1_U6.ce ;
assign \add_33ns_33s_33_2_1_U6.top_add_33ns_33s_33_2_1_Adder_3_U.clk  = \add_33ns_33s_33_2_1_U6.clk ;
assign \add_33ns_33s_33_2_1_U6.top_add_33ns_33s_33_2_1_Adder_3_U.reset  = \add_33ns_33s_33_2_1_U6.reset ;
assign \add_33ns_33s_33_2_1_U6.dout  = \add_33ns_33s_33_2_1_U6.top_add_33ns_33s_33_2_1_Adder_3_U.s ;
assign \add_33ns_33s_33_2_1_U6.ce  = 1'h1;
assign \add_33ns_33s_33_2_1_U6.clk  = ap_clk;
assign \add_33ns_33s_33_2_1_U6.din0  = { 16'h0000, lhs_V_4_reg_1585, 16'h0000 };
assign \add_33ns_33s_33_2_1_U6.din1  = { op_11[31], op_11 };
assign grp_fu_554_p2 = \add_33ns_33s_33_2_1_U6.dout ;
assign \add_33ns_33s_33_2_1_U6.reset  = ap_rst;
assign \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_14_U.ain_s0  = \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_14_U.a ;
assign \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_14_U.bin_s0  = \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_14_U.b ;
assign \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_14_U.s  = { \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_14_U.fas_s2 , \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_14_U.sum_s1  };
assign \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_14_U.u2.a  = \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_14_U.ain_s1 ;
assign \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_14_U.u2.b  = \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_14_U.bin_s1 ;
assign \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_14_U.u2.cin  = \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_14_U.carry_s1 ;
assign \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_14_U.facout_s2  = \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_14_U.u2.cout ;
assign \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_14_U.fas_s2  = \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_14_U.u2.s ;
assign \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_14_U.u1.a  = \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_14_U.a [15:0];
assign \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_14_U.u1.b  = \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_14_U.b [15:0];
assign \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_14_U.u1.cin  = 1'h0;
assign \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_14_U.facout_s1  = \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_14_U.u1.cout ;
assign \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_14_U.fas_s1  = \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_14_U.u1.s ;
assign \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_14_U.a  = \add_32s_32ns_32_2_1_U22.din0 ;
assign \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_14_U.b  = \add_32s_32ns_32_2_1_U22.din1 ;
assign \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_14_U.ce  = \add_32s_32ns_32_2_1_U22.ce ;
assign \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_14_U.clk  = \add_32s_32ns_32_2_1_U22.clk ;
assign \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_14_U.reset  = \add_32s_32ns_32_2_1_U22.reset ;
assign \add_32s_32ns_32_2_1_U22.dout  = \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_14_U.s ;
assign \add_32s_32ns_32_2_1_U22.ce  = 1'h1;
assign \add_32s_32ns_32_2_1_U22.clk  = ap_clk;
assign \add_32s_32ns_32_2_1_U22.din0  = { add_ln69_2_reg_2055[4], add_ln69_2_reg_2055[4], add_ln69_2_reg_2055[4], add_ln69_2_reg_2055[4], add_ln69_2_reg_2055[4], add_ln69_2_reg_2055[4], add_ln69_2_reg_2055[4], add_ln69_2_reg_2055[4], add_ln69_2_reg_2055[4], add_ln69_2_reg_2055[4], add_ln69_2_reg_2055[4], add_ln69_2_reg_2055[4], add_ln69_2_reg_2055[4], add_ln69_2_reg_2055[4], add_ln69_2_reg_2055[4], add_ln69_2_reg_2055[4], add_ln69_2_reg_2055[4], add_ln69_2_reg_2055[4], add_ln69_2_reg_2055[4], add_ln69_2_reg_2055[4], add_ln69_2_reg_2055[4], add_ln69_2_reg_2055[4], add_ln69_2_reg_2055[4], add_ln69_2_reg_2055[4], add_ln69_2_reg_2055[4], add_ln69_2_reg_2055[4], add_ln69_2_reg_2055[4], add_ln69_2_reg_2055 };
assign \add_32s_32ns_32_2_1_U22.din1  = add_ln69_reg_2144;
assign grp_fu_1435_p2 = \add_32s_32ns_32_2_1_U22.dout ;
assign \add_32s_32ns_32_2_1_U22.reset  = ap_rst;
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.ain_s0  = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.a ;
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.bin_s0  = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.b ;
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.s  = { \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.fas_s2 , \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.sum_s1  };
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.a  = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.ain_s1 ;
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.b  = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.bin_s1 ;
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.cin  = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.carry_s1 ;
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.facout_s2  = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.cout ;
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.fas_s2  = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.s ;
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.a  = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.a [15:0];
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.b  = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.b [15:0];
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.cin  = 1'h0;
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.facout_s1  = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.cout ;
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.fas_s1  = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.s ;
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.a  = \add_32ns_32ns_32_2_1_U21.din0 ;
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.b  = \add_32ns_32ns_32_2_1_U21.din1 ;
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.ce  = \add_32ns_32ns_32_2_1_U21.ce ;
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.clk  = \add_32ns_32ns_32_2_1_U21.clk ;
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.reset  = \add_32ns_32ns_32_2_1_U21.reset ;
assign \add_32ns_32ns_32_2_1_U21.dout  = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.s ;
assign \add_32ns_32ns_32_2_1_U21.ce  = 1'h1;
assign \add_32ns_32ns_32_2_1_U21.clk  = ap_clk;
assign \add_32ns_32ns_32_2_1_U21.din0  = ret_V_28_reg_2134;
assign \add_32ns_32ns_32_2_1_U21.din1  = { 16'h0000, ret_V_23_reg_2129[5], ret_V_23_reg_2129[5], ret_V_23_reg_2129[5], ret_V_23_reg_2129[5], ret_V_23_reg_2129[5], ret_V_23_reg_2129[5], ret_V_23_reg_2129[5], ret_V_23_reg_2129[5], ret_V_23_reg_2129[5], ret_V_23_reg_2129[5], ret_V_23_reg_2129 };
assign grp_fu_1427_p2 = \add_32ns_32ns_32_2_1_U21.dout ;
assign \add_32ns_32ns_32_2_1_U21.reset  = ap_rst;
assign \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.ain_s0  = \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.a ;
assign \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.bin_s0  = \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.b ;
assign \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.s  = { \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.fas_s2 , \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.sum_s1  };
assign \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.a  = \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.ain_s1 ;
assign \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.b  = \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.bin_s1 ;
assign \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.cin  = \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.carry_s1 ;
assign \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.facout_s2  = \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.cout ;
assign \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.fas_s2  = \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.s ;
assign \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.a  = \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.a [15:0];
assign \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.b  = \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.b [15:0];
assign \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.cin  = 1'h0;
assign \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.facout_s1  = \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.cout ;
assign \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.fas_s1  = \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.s ;
assign \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.a  = \add_32ns_32ns_32_2_1_U20.din0 ;
assign \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.b  = \add_32ns_32ns_32_2_1_U20.din1 ;
assign \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.ce  = \add_32ns_32ns_32_2_1_U20.ce ;
assign \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.clk  = \add_32ns_32ns_32_2_1_U20.clk ;
assign \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.reset  = \add_32ns_32ns_32_2_1_U20.reset ;
assign \add_32ns_32ns_32_2_1_U20.dout  = \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.s ;
assign \add_32ns_32ns_32_2_1_U20.ce  = 1'h1;
assign \add_32ns_32ns_32_2_1_U20.clk  = ap_clk;
assign \add_32ns_32ns_32_2_1_U20.din0  = ret_V_36_cast_reg_2107;
assign \add_32ns_32ns_32_2_1_U20.din1  = 32'd1;
assign grp_fu_1377_p2 = \add_32ns_32ns_32_2_1_U20.dout ;
assign \add_32ns_32ns_32_2_1_U20.reset  = ap_rst;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.ain_s0  = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.a ;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.bin_s0  = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.b ;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.s  = { \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.fas_s2 , \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.sum_s1  };
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.a  = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.ain_s1 ;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.b  = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.bin_s1 ;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.cin  = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.carry_s1 ;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.facout_s2  = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.cout ;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.fas_s2  = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.s ;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.a  = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.a [15:0];
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.b  = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.b [15:0];
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.cin  = 1'h0;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.facout_s1  = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.cout ;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.fas_s1  = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.s ;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.a  = \add_32ns_32ns_32_2_1_U17.din0 ;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.b  = \add_32ns_32ns_32_2_1_U17.din1 ;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.ce  = \add_32ns_32ns_32_2_1_U17.ce ;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.clk  = \add_32ns_32ns_32_2_1_U17.clk ;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.reset  = \add_32ns_32ns_32_2_1_U17.reset ;
assign \add_32ns_32ns_32_2_1_U17.dout  = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.s ;
assign \add_32ns_32ns_32_2_1_U17.ce  = 1'h1;
assign \add_32ns_32ns_32_2_1_U17.clk  = ap_clk;
assign \add_32ns_32ns_32_2_1_U17.din0  = ret_V_34_cast_reg_2038;
assign \add_32ns_32ns_32_2_1_U17.din1  = 32'd1;
assign grp_fu_1288_p2 = \add_32ns_32ns_32_2_1_U17.dout ;
assign \add_32ns_32ns_32_2_1_U17.reset  = ap_rst;
assign \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_2_U.ain_s0  = \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_2_U.a ;
assign \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_2_U.bin_s0  = \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_2_U.b ;
assign \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_2_U.s  = { \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_2_U.fas_s2 , \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_2_U.sum_s1  };
assign \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_2_U.u2.a  = \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_2_U.ain_s1 ;
assign \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_2_U.u2.b  = \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_2_U.bin_s1 ;
assign \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_2_U.u2.cin  = \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_2_U.carry_s1 ;
assign \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_2_U.facout_s2  = \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_2_U.u2.cout ;
assign \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_2_U.fas_s2  = \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_2_U.u2.s ;
assign \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_2_U.u1.a  = \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_2_U.a [0];
assign \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_2_U.u1.b  = \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_2_U.b [0];
assign \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_2_U.u1.cin  = 1'h0;
assign \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_2_U.facout_s1  = \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_2_U.u1.cout ;
assign \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_2_U.fas_s1  = \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_2_U.u1.s ;
assign \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_2_U.a  = \add_2ns_2ns_2_2_1_U5.din0 ;
assign \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_2_U.b  = \add_2ns_2ns_2_2_1_U5.din1 ;
assign \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_2_U.ce  = \add_2ns_2ns_2_2_1_U5.ce ;
assign \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_2_U.clk  = \add_2ns_2ns_2_2_1_U5.clk ;
assign \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_2_U.reset  = \add_2ns_2ns_2_2_1_U5.reset ;
assign \add_2ns_2ns_2_2_1_U5.dout  = \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_2_U.s ;
assign \add_2ns_2ns_2_2_1_U5.ce  = 1'h1;
assign \add_2ns_2ns_2_2_1_U5.clk  = ap_clk;
assign \add_2ns_2ns_2_2_1_U5.din0  = ret_V_cast_reg_1514;
assign \add_2ns_2ns_2_2_1_U5.din1  = 2'h1;
assign grp_fu_446_p2 = \add_2ns_2ns_2_2_1_U5.dout ;
assign \add_2ns_2ns_2_2_1_U5.reset  = ap_rst;
assign \add_25s_25s_25_2_1_U11.top_add_25s_25s_25_2_1_Adder_6_U.ain_s0  = \add_25s_25s_25_2_1_U11.top_add_25s_25s_25_2_1_Adder_6_U.a ;
assign \add_25s_25s_25_2_1_U11.top_add_25s_25s_25_2_1_Adder_6_U.bin_s0  = \add_25s_25s_25_2_1_U11.top_add_25s_25s_25_2_1_Adder_6_U.b ;
assign \add_25s_25s_25_2_1_U11.top_add_25s_25s_25_2_1_Adder_6_U.s  = { \add_25s_25s_25_2_1_U11.top_add_25s_25s_25_2_1_Adder_6_U.fas_s2 , \add_25s_25s_25_2_1_U11.top_add_25s_25s_25_2_1_Adder_6_U.sum_s1  };
assign \add_25s_25s_25_2_1_U11.top_add_25s_25s_25_2_1_Adder_6_U.u2.a  = \add_25s_25s_25_2_1_U11.top_add_25s_25s_25_2_1_Adder_6_U.ain_s1 ;
assign \add_25s_25s_25_2_1_U11.top_add_25s_25s_25_2_1_Adder_6_U.u2.b  = \add_25s_25s_25_2_1_U11.top_add_25s_25s_25_2_1_Adder_6_U.bin_s1 ;
assign \add_25s_25s_25_2_1_U11.top_add_25s_25s_25_2_1_Adder_6_U.u2.cin  = \add_25s_25s_25_2_1_U11.top_add_25s_25s_25_2_1_Adder_6_U.carry_s1 ;
assign \add_25s_25s_25_2_1_U11.top_add_25s_25s_25_2_1_Adder_6_U.facout_s2  = \add_25s_25s_25_2_1_U11.top_add_25s_25s_25_2_1_Adder_6_U.u2.cout ;
assign \add_25s_25s_25_2_1_U11.top_add_25s_25s_25_2_1_Adder_6_U.fas_s2  = \add_25s_25s_25_2_1_U11.top_add_25s_25s_25_2_1_Adder_6_U.u2.s ;
assign \add_25s_25s_25_2_1_U11.top_add_25s_25s_25_2_1_Adder_6_U.u1.a  = \add_25s_25s_25_2_1_U11.top_add_25s_25s_25_2_1_Adder_6_U.a [11:0];
assign \add_25s_25s_25_2_1_U11.top_add_25s_25s_25_2_1_Adder_6_U.u1.b  = \add_25s_25s_25_2_1_U11.top_add_25s_25s_25_2_1_Adder_6_U.b [11:0];
assign \add_25s_25s_25_2_1_U11.top_add_25s_25s_25_2_1_Adder_6_U.u1.cin  = 1'h0;
assign \add_25s_25s_25_2_1_U11.top_add_25s_25s_25_2_1_Adder_6_U.facout_s1  = \add_25s_25s_25_2_1_U11.top_add_25s_25s_25_2_1_Adder_6_U.u1.cout ;
assign \add_25s_25s_25_2_1_U11.top_add_25s_25s_25_2_1_Adder_6_U.fas_s1  = \add_25s_25s_25_2_1_U11.top_add_25s_25s_25_2_1_Adder_6_U.u1.s ;
assign \add_25s_25s_25_2_1_U11.top_add_25s_25s_25_2_1_Adder_6_U.a  = \add_25s_25s_25_2_1_U11.din0 ;
assign \add_25s_25s_25_2_1_U11.top_add_25s_25s_25_2_1_Adder_6_U.b  = \add_25s_25s_25_2_1_U11.din1 ;
assign \add_25s_25s_25_2_1_U11.top_add_25s_25s_25_2_1_Adder_6_U.ce  = \add_25s_25s_25_2_1_U11.ce ;
assign \add_25s_25s_25_2_1_U11.top_add_25s_25s_25_2_1_Adder_6_U.clk  = \add_25s_25s_25_2_1_U11.clk ;
assign \add_25s_25s_25_2_1_U11.top_add_25s_25s_25_2_1_Adder_6_U.reset  = \add_25s_25s_25_2_1_U11.reset ;
assign \add_25s_25s_25_2_1_U11.dout  = \add_25s_25s_25_2_1_U11.top_add_25s_25s_25_2_1_Adder_6_U.s ;
assign \add_25s_25s_25_2_1_U11.ce  = 1'h1;
assign \add_25s_25s_25_2_1_U11.clk  = ap_clk;
assign \add_25s_25s_25_2_1_U11.din0  = { select_ln850_5_reg_1829[16], select_ln850_5_reg_1829, 7'h00 };
assign \add_25s_25s_25_2_1_U11.din1  = { ret_V_3_reg_1802[12], ret_V_3_reg_1802[12], ret_V_3_reg_1802[12], ret_V_3_reg_1802[12], ret_V_3_reg_1802[12], ret_V_3_reg_1802[12], ret_V_3_reg_1802[12], ret_V_3_reg_1802[12], ret_V_3_reg_1802[12], ret_V_3_reg_1802, 3'h0 };
assign grp_fu_796_p2 = \add_25s_25s_25_2_1_U11.dout ;
assign \add_25s_25s_25_2_1_U11.reset  = ap_rst;
assign \add_19s_19ns_19_2_1_U12.top_add_19s_19ns_19_2_1_Adder_7_U.ain_s0  = \add_19s_19ns_19_2_1_U12.top_add_19s_19ns_19_2_1_Adder_7_U.a ;
assign \add_19s_19ns_19_2_1_U12.top_add_19s_19ns_19_2_1_Adder_7_U.bin_s0  = \add_19s_19ns_19_2_1_U12.top_add_19s_19ns_19_2_1_Adder_7_U.b ;
assign \add_19s_19ns_19_2_1_U12.top_add_19s_19ns_19_2_1_Adder_7_U.s  = { \add_19s_19ns_19_2_1_U12.top_add_19s_19ns_19_2_1_Adder_7_U.fas_s2 , \add_19s_19ns_19_2_1_U12.top_add_19s_19ns_19_2_1_Adder_7_U.sum_s1  };
assign \add_19s_19ns_19_2_1_U12.top_add_19s_19ns_19_2_1_Adder_7_U.u2.a  = \add_19s_19ns_19_2_1_U12.top_add_19s_19ns_19_2_1_Adder_7_U.ain_s1 ;
assign \add_19s_19ns_19_2_1_U12.top_add_19s_19ns_19_2_1_Adder_7_U.u2.b  = \add_19s_19ns_19_2_1_U12.top_add_19s_19ns_19_2_1_Adder_7_U.bin_s1 ;
assign \add_19s_19ns_19_2_1_U12.top_add_19s_19ns_19_2_1_Adder_7_U.u2.cin  = \add_19s_19ns_19_2_1_U12.top_add_19s_19ns_19_2_1_Adder_7_U.carry_s1 ;
assign \add_19s_19ns_19_2_1_U12.top_add_19s_19ns_19_2_1_Adder_7_U.facout_s2  = \add_19s_19ns_19_2_1_U12.top_add_19s_19ns_19_2_1_Adder_7_U.u2.cout ;
assign \add_19s_19ns_19_2_1_U12.top_add_19s_19ns_19_2_1_Adder_7_U.fas_s2  = \add_19s_19ns_19_2_1_U12.top_add_19s_19ns_19_2_1_Adder_7_U.u2.s ;
assign \add_19s_19ns_19_2_1_U12.top_add_19s_19ns_19_2_1_Adder_7_U.u1.a  = \add_19s_19ns_19_2_1_U12.top_add_19s_19ns_19_2_1_Adder_7_U.a [8:0];
assign \add_19s_19ns_19_2_1_U12.top_add_19s_19ns_19_2_1_Adder_7_U.u1.b  = \add_19s_19ns_19_2_1_U12.top_add_19s_19ns_19_2_1_Adder_7_U.b [8:0];
assign \add_19s_19ns_19_2_1_U12.top_add_19s_19ns_19_2_1_Adder_7_U.u1.cin  = 1'h0;
assign \add_19s_19ns_19_2_1_U12.top_add_19s_19ns_19_2_1_Adder_7_U.facout_s1  = \add_19s_19ns_19_2_1_U12.top_add_19s_19ns_19_2_1_Adder_7_U.u1.cout ;
assign \add_19s_19ns_19_2_1_U12.top_add_19s_19ns_19_2_1_Adder_7_U.fas_s1  = \add_19s_19ns_19_2_1_U12.top_add_19s_19ns_19_2_1_Adder_7_U.u1.s ;
assign \add_19s_19ns_19_2_1_U12.top_add_19s_19ns_19_2_1_Adder_7_U.a  = \add_19s_19ns_19_2_1_U12.din0 ;
assign \add_19s_19ns_19_2_1_U12.top_add_19s_19ns_19_2_1_Adder_7_U.b  = \add_19s_19ns_19_2_1_U12.din1 ;
assign \add_19s_19ns_19_2_1_U12.top_add_19s_19ns_19_2_1_Adder_7_U.ce  = \add_19s_19ns_19_2_1_U12.ce ;
assign \add_19s_19ns_19_2_1_U12.top_add_19s_19ns_19_2_1_Adder_7_U.clk  = \add_19s_19ns_19_2_1_U12.clk ;
assign \add_19s_19ns_19_2_1_U12.top_add_19s_19ns_19_2_1_Adder_7_U.reset  = \add_19s_19ns_19_2_1_U12.reset ;
assign \add_19s_19ns_19_2_1_U12.dout  = \add_19s_19ns_19_2_1_U12.top_add_19s_19ns_19_2_1_Adder_7_U.s ;
assign \add_19s_19ns_19_2_1_U12.ce  = 1'h1;
assign \add_19s_19ns_19_2_1_U12.clk  = ap_clk;
assign \add_19s_19ns_19_2_1_U12.din0  = { tmp_3_reg_1913[17], tmp_3_reg_1913 };
assign \add_19s_19ns_19_2_1_U12.din1  = 19'h00001;
assign grp_fu_990_p2 = \add_19s_19ns_19_2_1_U12.dout ;
assign \add_19s_19ns_19_2_1_U12.reset  = ap_rst;
assign \add_17ns_17ns_17_2_1_U10.top_add_17ns_17ns_17_2_1_Adder_5_U.ain_s0  = \add_17ns_17ns_17_2_1_U10.top_add_17ns_17ns_17_2_1_Adder_5_U.a ;
assign \add_17ns_17ns_17_2_1_U10.top_add_17ns_17ns_17_2_1_Adder_5_U.bin_s0  = \add_17ns_17ns_17_2_1_U10.top_add_17ns_17ns_17_2_1_Adder_5_U.b ;
assign \add_17ns_17ns_17_2_1_U10.top_add_17ns_17ns_17_2_1_Adder_5_U.s  = { \add_17ns_17ns_17_2_1_U10.top_add_17ns_17ns_17_2_1_Adder_5_U.fas_s2 , \add_17ns_17ns_17_2_1_U10.top_add_17ns_17ns_17_2_1_Adder_5_U.sum_s1  };
assign \add_17ns_17ns_17_2_1_U10.top_add_17ns_17ns_17_2_1_Adder_5_U.u2.a  = \add_17ns_17ns_17_2_1_U10.top_add_17ns_17ns_17_2_1_Adder_5_U.ain_s1 ;
assign \add_17ns_17ns_17_2_1_U10.top_add_17ns_17ns_17_2_1_Adder_5_U.u2.b  = \add_17ns_17ns_17_2_1_U10.top_add_17ns_17ns_17_2_1_Adder_5_U.bin_s1 ;
assign \add_17ns_17ns_17_2_1_U10.top_add_17ns_17ns_17_2_1_Adder_5_U.u2.cin  = \add_17ns_17ns_17_2_1_U10.top_add_17ns_17ns_17_2_1_Adder_5_U.carry_s1 ;
assign \add_17ns_17ns_17_2_1_U10.top_add_17ns_17ns_17_2_1_Adder_5_U.facout_s2  = \add_17ns_17ns_17_2_1_U10.top_add_17ns_17ns_17_2_1_Adder_5_U.u2.cout ;
assign \add_17ns_17ns_17_2_1_U10.top_add_17ns_17ns_17_2_1_Adder_5_U.fas_s2  = \add_17ns_17ns_17_2_1_U10.top_add_17ns_17ns_17_2_1_Adder_5_U.u2.s ;
assign \add_17ns_17ns_17_2_1_U10.top_add_17ns_17ns_17_2_1_Adder_5_U.u1.a  = \add_17ns_17ns_17_2_1_U10.top_add_17ns_17ns_17_2_1_Adder_5_U.a [7:0];
assign \add_17ns_17ns_17_2_1_U10.top_add_17ns_17ns_17_2_1_Adder_5_U.u1.b  = \add_17ns_17ns_17_2_1_U10.top_add_17ns_17ns_17_2_1_Adder_5_U.b [7:0];
assign \add_17ns_17ns_17_2_1_U10.top_add_17ns_17ns_17_2_1_Adder_5_U.u1.cin  = 1'h0;
assign \add_17ns_17ns_17_2_1_U10.top_add_17ns_17ns_17_2_1_Adder_5_U.facout_s1  = \add_17ns_17ns_17_2_1_U10.top_add_17ns_17ns_17_2_1_Adder_5_U.u1.cout ;
assign \add_17ns_17ns_17_2_1_U10.top_add_17ns_17ns_17_2_1_Adder_5_U.fas_s1  = \add_17ns_17ns_17_2_1_U10.top_add_17ns_17ns_17_2_1_Adder_5_U.u1.s ;
assign \add_17ns_17ns_17_2_1_U10.top_add_17ns_17ns_17_2_1_Adder_5_U.a  = \add_17ns_17ns_17_2_1_U10.din0 ;
assign \add_17ns_17ns_17_2_1_U10.top_add_17ns_17ns_17_2_1_Adder_5_U.b  = \add_17ns_17ns_17_2_1_U10.din1 ;
assign \add_17ns_17ns_17_2_1_U10.top_add_17ns_17ns_17_2_1_Adder_5_U.ce  = \add_17ns_17ns_17_2_1_U10.ce ;
assign \add_17ns_17ns_17_2_1_U10.top_add_17ns_17ns_17_2_1_Adder_5_U.clk  = \add_17ns_17ns_17_2_1_U10.clk ;
assign \add_17ns_17ns_17_2_1_U10.top_add_17ns_17ns_17_2_1_Adder_5_U.reset  = \add_17ns_17ns_17_2_1_U10.reset ;
assign \add_17ns_17ns_17_2_1_U10.dout  = \add_17ns_17ns_17_2_1_U10.top_add_17ns_17ns_17_2_1_Adder_5_U.s ;
assign \add_17ns_17ns_17_2_1_U10.ce  = 1'h1;
assign \add_17ns_17ns_17_2_1_U10.clk  = ap_clk;
assign \add_17ns_17ns_17_2_1_U10.din0  = ret_V_12_reg_1733;
assign \add_17ns_17ns_17_2_1_U10.din1  = 17'h00001;
assign grp_fu_665_p2 = \add_17ns_17ns_17_2_1_U10.dout ;
assign \add_17ns_17ns_17_2_1_U10.reset  = ap_rst;
endmodule


// Machine B:
// Processed by function `add_clk_enable_signal` in `verilog_tricks.py`.
// Processed by function `remove_reset_signal` in `verilog_tricks.py`.
module top_B (
  ap_clk,
  ap_start,
  ap_done,
  ap_idle,
  ap_ready,
  op_0,
  op_1,
  op_4,
  op_6,
  op_8,
  op_11,
  op_15,
  op_28,
  op_28_ap_vld,
clk_enable
);
input clk_enable;


input ap_clk;
wire ap_rst;
assign ap_rst = op_28_ap_vld;
input ap_start;
input [1:0] op_0;
input [15:0] op_1;
input [31:0] op_11;
input [15:0] op_15;
input [7:0] op_4;
input [31:0] op_6;
input [7:0] op_8;
output ap_done;
output ap_idle;
output ap_ready;
output [31:0] op_28;
output op_28_ap_vld;


reg Range1_all_ones_1_reg_1669;
reg Range1_all_ones_reg_1740;
reg Range1_all_zeros_1_reg_1676;
reg Range1_all_zeros_reg_1747;
reg Range2_all_ones_1_reg_1664;
reg Range2_all_ones_reg_1735;
reg [31:0] add_ln691_1_reg_1841;
reg [2:0] add_ln69_1_reg_1703;
reg [4:0] add_ln69_2_reg_1814;
reg and_ln785_5_reg_1757;
reg [9:0] ap_CS_fsm = 10'h001;
reg carry_1_reg_1728;
reg icmp_ln1496_reg_1594;
reg icmp_ln851_1_reg_1584;
reg icmp_ln851_2_reg_1789;
reg icmp_ln851_3_reg_1698;
reg icmp_ln851_4_reg_1804;
reg icmp_ln851_5_reg_1836;
reg icmp_ln851_6_reg_1858;
reg icmp_ln851_reg_1527;
reg [3:0] op_14_V_reg_1772;
reg [9:0] p_Result_1_reg_1637;
reg p_Result_21_reg_1613;
reg p_Result_23_reg_1621;
reg p_Result_24_reg_1717;
reg p_Result_25_reg_1626;
reg p_Result_26_reg_1544;
reg p_Result_28_reg_1551;
reg p_Result_29_reg_1652;
reg p_Result_30_reg_1556;
reg [8:0] p_Result_s_22_reg_1632;
reg [3:0] p_Val2_3_reg_1708;
reg [3:0] p_Val2_7_reg_1643;
reg [15:0] r_V_3_reg_1605;
reg [10:0] r_V_4_reg_1532;
reg [7:0] r_V_reg_1777;
reg [16:0] ret_V_12_reg_1691;
reg [16:0] ret_V_13_reg_1767;
reg [32:0] ret_V_18_reg_1515;
reg [5:0] ret_V_23_reg_1819;
reg [32:0] ret_V_24_reg_1686;
reg [34:0] ret_V_26_reg_1824;
reg [45:0] ret_V_27_reg_1846;
reg [31:0] ret_V_28_reg_1863;
reg [31:0] ret_V_34_cast_reg_1829;
reg [31:0] ret_V_36_cast_reg_1851;
reg [3:0] ret_V_6_cast_reg_1578;
reg [3:0] ret_V_6_reg_1589;
reg [5:0] ret_V_7_reg_1782;
reg [1:0] ret_V_cast_reg_1520;
reg sel_tmp25_reg_1762;
reg [3:0] select_ln340_1_reg_1752;
reg signbit_reg_1503;
reg [3:0] tmp_1_reg_1562;
reg [4:0] tmp_2_reg_1567;
reg [17:0] tmp_3_reg_1799;
reg [1:0] trunc_ln1115_reg_1539;
reg [1:0] trunc_ln851_5_reg_1809;
reg xor_ln416_1_reg_1658;
reg xor_ln416_reg_1723;
reg [3:0] _213_;
reg [21:0] _222_;
reg [3:0] _250_;
wire _000_;
wire _001_;
wire _002_;
wire _003_;
wire _004_;
wire _005_;
wire [31:0] _006_;
wire [2:0] _007_;
wire [4:0] _008_;
wire _009_;
wire [9:0] _010_;
wire _011_;
wire _012_;
wire _013_;
wire _014_;
wire _015_;
wire _016_;
wire _017_;
wire _018_;
wire _019_;
wire [3:0] _020_;
wire [9:0] _021_;
wire _022_;
wire _023_;
wire _024_;
wire _025_;
wire _026_;
wire _027_;
wire _028_;
wire _029_;
wire [8:0] _030_;
wire [3:0] _031_;
wire [3:0] _032_;
wire [15:0] _033_;
wire [10:0] _034_;
wire [7:0] _035_;
wire [16:0] _036_;
wire [16:0] _037_;
wire [32:0] _038_;
wire [3:0] _039_;
wire [5:0] _040_;
wire [32:0] _041_;
wire [21:0] _042_;
wire [34:0] _043_;
wire [45:0] _044_;
wire [31:0] _045_;
wire [31:0] _046_;
wire [31:0] _047_;
wire [3:0] _048_;
wire [3:0] _049_;
wire [5:0] _050_;
wire [1:0] _051_;
wire _052_;
wire [3:0] _053_;
wire _054_;
wire [3:0] _055_;
wire [4:0] _056_;
wire [17:0] _057_;
wire [1:0] _058_;
wire [1:0] _059_;
wire _060_;
wire _061_;
wire [3:0] _062_;
wire [1:0] _063_;
wire _064_;
wire _065_;
wire _066_;
wire _067_;
wire _068_;
wire _069_;
wire _070_;
wire _071_;
wire _072_;
wire _073_;
wire _074_;
wire _075_;
wire _076_;
wire _077_;
wire _078_;
wire _079_;
wire _080_;
wire _081_;
wire _082_;
wire _083_;
wire _084_;
wire _085_;
wire _086_;
wire _087_;
wire _088_;
wire _089_;
wire _090_;
wire _091_;
wire _092_;
wire _093_;
wire _094_;
wire _095_;
wire _096_;
wire Range1_all_ones_1_fu_572_p2;
wire Range1_all_ones_fu_736_p2;
wire Range1_all_zeros_1_fu_577_p2;
wire Range1_all_zeros_fu_741_p2;
wire Range2_all_ones_1_fu_567_p2;
wire Range2_all_ones_fu_731_p2;
wire [31:0] add_ln691_1_fu_1385_p2;
wire [31:0] add_ln691_2_fu_1458_p2;
wire [18:0] add_ln691_fu_1328_p2;
wire [2:0] add_ln69_1_fu_666_p2;
wire [4:0] add_ln69_2_fu_1287_p2;
wire [31:0] add_ln69_fu_1483_p2;
wire and_ln340_1_fu_903_p2;
wire and_ln340_fu_1111_p2;
wire and_ln406_fu_696_p2;
wire and_ln408_fu_537_p2;
wire and_ln780_1_fu_761_p2;
wire and_ln780_fu_964_p2;
wire and_ln781_1_fu_773_p2;
wire and_ln781_fu_975_p2;
wire and_ln785_1_fu_1086_p2;
wire and_ln785_2_fu_1099_p2;
wire and_ln785_4_fu_875_p2;
wire and_ln785_5_fu_885_p2;
wire and_ln785_6_fu_891_p2;
wire and_ln785_fu_1076_p2;
wire and_ln786_1_fu_811_p2;
wire and_ln786_fu_1012_p2;
wire ap_CS_fsm_state1;
wire ap_CS_fsm_state10;
wire ap_CS_fsm_state2;
wire ap_CS_fsm_state3;
wire ap_CS_fsm_state4;
wire ap_CS_fsm_state5;
wire ap_CS_fsm_state6;
wire ap_CS_fsm_state7;
wire ap_CS_fsm_state8;
wire ap_CS_fsm_state9;
wire [9:0] ap_NS_fsm;
wire ap_clk;
wire ap_done;
wire ap_idle;
wire ap_ready;
wire ap_rst;
wire ap_start;
wire carry_1_fu_726_p2;
wire carry_3_fu_746_p2;
wire deleted_ones_1_fu_766_p3;
wire deleted_ones_fu_969_p3;
wire deleted_zeros_1_fu_750_p3;
wire deleted_zeros_fu_954_p3;
wire [31:0] icmp_ln1496_fu_432_p1;
wire icmp_ln1496_fu_432_p2;
wire icmp_ln851_1_fu_409_p2;
wire icmp_ln851_2_fu_1201_p2;
wire icmp_ln851_3_fu_652_p2;
wire icmp_ln851_4_fu_1270_p2;
wire icmp_ln851_5_fu_1380_p2;
wire icmp_ln851_6_fu_1445_p2;
wire icmp_ln851_fu_298_p2;
wire icmp_ln874_fu_610_p2;
wire [5:0] lhs_V_2_fu_373_p3;
wire lhs_V_4_fu_601_p2;
wire [16:0] lhs_V_5_fu_616_p3;
wire [5:0] lhs_V_fu_1150_p3;
wire [21:0] lhs_fu_263_p3;
wire [3:0] \mul_4ns_4s_8_1_1_U3.din0 ;
wire [3:0] \mul_4ns_4s_8_1_1_U3.din1 ;
wire [7:0] \mul_4ns_4s_8_1_1_U3.dout ;
wire [3:0] \mul_4ns_4s_8_1_1_U3.top_mul_4ns_4s_8_1_1_Multiplier_2_U.a ;
wire [3:0] \mul_4ns_4s_8_1_1_U3.top_mul_4ns_4s_8_1_1_Multiplier_2_U.b ;
wire [7:0] \mul_4ns_4s_8_1_1_U3.top_mul_4ns_4s_8_1_1_Multiplier_2_U.p ;
wire [7:0] \mul_8ns_8s_16_1_1_U2.din0 ;
wire [7:0] \mul_8ns_8s_16_1_1_U2.din1 ;
wire [15:0] \mul_8ns_8s_16_1_1_U2.dout ;
wire [7:0] \mul_8ns_8s_16_1_1_U2.top_mul_8ns_8s_16_1_1_Multiplier_1_U.a ;
wire [7:0] \mul_8ns_8s_16_1_1_U2.top_mul_8ns_8s_16_1_1_Multiplier_1_U.b ;
wire [15:0] \mul_8ns_8s_16_1_1_U2.top_mul_8ns_8s_16_1_1_Multiplier_1_U.p ;
wire [7:0] \mul_8s_3ns_11_1_1_U1.din0 ;
wire [2:0] \mul_8s_3ns_11_1_1_U1.din1 ;
wire [10:0] \mul_8s_3ns_11_1_1_U1.dout ;
wire [7:0] \mul_8s_3ns_11_1_1_U1.top_mul_8s_3ns_11_1_1_Multiplier_0_U.a ;
wire [2:0] \mul_8s_3ns_11_1_1_U1.top_mul_8s_3ns_11_1_1_Multiplier_0_U.b ;
wire [10:0] \mul_8s_3ns_11_1_1_U1.top_mul_8s_3ns_11_1_1_Multiplier_0_U.p ;
wire neg_src_4_fu_784_p2;
wire neg_src_fu_985_p2;
wire [1:0] op_0;
wire [15:0] op_1;
wire [31:0] op_11;
wire [15:0] op_12_V_fu_946_p3;
wire [3:0] op_14_V_fu_1129_p3;
wire [15:0] op_15;
wire [3:0] op_16_V_fu_1168_p4;
wire [31:0] op_28;
wire op_28_ap_vld;
wire [7:0] op_4;
wire [3:0] op_5_V_fu_366_p3;
wire [31:0] op_6;
wire [7:0] op_8;
wire [3:0] op_9_V_fu_1141_p3;
wire or_ln340_1_fu_816_p2;
wire or_ln340_2_fu_1063_p2;
wire or_ln340_3_fu_1117_p2;
wire or_ln340_4_fu_862_p2;
wire or_ln340_5_fu_909_p2;
wire or_ln340_fu_1017_p2;
wire or_ln406_fu_691_p2;
wire or_ln785_1_fu_795_p2;
wire or_ln785_2_fu_1081_p2;
wire or_ln785_3_fu_880_p2;
wire or_ln785_fu_996_p2;
wire overflow_1_fu_805_p2;
wire overflow_fu_1006_p2;
wire [3:0] p_Result_14_fu_853_p4;
wire p_Result_15_fu_582_p3;
wire p_Result_16_fu_1293_p3;
wire p_Result_17_fu_1207_p3;
wire p_Result_18_fu_1321_p3;
wire p_Result_19_fu_1390_p3;
wire p_Result_20_fu_1451_p3;
wire p_Result_22_fu_681_p3;
wire p_Result_24_fu_712_p3;
wire p_Result_27_fu_529_p2;
wire p_Result_29_fu_553_p3;
wire [6:0] p_Result_5_fu_1262_p3;
wire [3:0] p_Result_8_fu_1054_p4;
wire p_Result_s_fu_438_p3;
wire [3:0] p_Val2_2_fu_672_p4;
wire [3:0] p_Val2_3_fu_706_p2;
wire [2:0] p_Val2_4_fu_1049_p2;
wire [3:0] p_Val2_6_fu_520_p4;
wire [3:0] p_Val2_7_fu_547_p2;
wire [2:0] p_Val2_8_fu_848_p2;
wire r_1_fu_534_p1;
wire [7:0] r_V_3_fu_470_p0;
wire [15:0] r_V_3_fu_470_p00;
wire [15:0] r_V_3_fu_470_p2;
wire [2:0] r_V_4_fu_312_p1;
wire [10:0] r_V_4_fu_312_p10;
wire [10:0] r_V_4_fu_312_p2;
wire [3:0] r_V_fu_1182_p0;
wire [7:0] r_V_fu_1182_p2;
wire r_fu_688_p1;
wire [16:0] ret_V_13_fu_921_p2;
wire [32:0] ret_V_18_fu_278_p2;
wire [1:0] ret_V_19_fu_456_p3;
wire [5:0] ret_V_20_fu_1162_p2;
wire [6:0] ret_V_21_fu_389_p2;
wire [6:0] ret_V_21_reg_1573;
wire [3:0] ret_V_22_fu_594_p3;
wire [5:0] ret_V_23_fu_1311_p3;
wire [32:0] ret_V_24_fu_632_p2;
wire [24:0] ret_V_25_fu_1242_p2;
wire [24:0] ret_V_25_reg_1794;
wire [34:0] ret_V_26_fu_1364_p2;
wire [45:0] ret_V_27_fu_1425_p2;
wire [31:0] ret_V_28_fu_1469_p3;
wire [12:0] ret_V_3_fu_940_p2;
wire [3:0] ret_V_6_cast_fu_395_p4;
wire [3:0] ret_V_6_fu_415_p2;
wire [5:0] ret_V_9_fu_1300_p2;
wire [1:0] ret_V_fu_445_p2;
wire [2:0] ret_fu_255_p3;
wire [23:0] rhs_3_fu_1230_p3;
wire [44:0] rhs_4_fu_1413_p3;
wire [11:0] rhs_fu_929_p3;
wire sel_tmp11_fu_1123_p2;
wire sel_tmp25_fu_915_p2;
wire [3:0] select_ln340_1_fu_868_p3;
wire [3:0] select_ln340_fu_1069_p3;
wire [31:0] select_ln353_1_fu_1406_p3;
wire [18:0] select_ln353_fu_1344_p3;
wire [3:0] select_ln785_1_fu_1136_p3;
wire [3:0] select_ln785_fu_1092_p3;
wire [3:0] select_ln850_1_fu_589_p3;
wire [5:0] select_ln850_2_fu_1305_p3;
wire [16:0] select_ln850_4_fu_1218_p3;
wire [16:0] select_ln850_5_fu_1223_p3;
wire [31:0] select_ln850_6_fu_1463_p3;
wire [18:0] select_ln850_7_fu_1337_p3;
wire [31:0] select_ln850_8_fu_1401_p3;
wire [1:0] select_ln850_fu_450_p3;
wire [24:0] sext_ln1192_1_fu_1238_p1;
wire [34:0] sext_ln1192_2_fu_1360_p1;
wire [45:0] sext_ln1192_3_fu_1421_p1;
wire [24:0] sext_ln1192_fu_1214_p1;
wire [32:0] sext_ln1193_fu_270_p1;
wire [5:0] sext_ln1194_fu_1158_p1;
wire [15:0] sext_ln69_1_fu_1476_p1;
wire [2:0] sext_ln69_2_fu_658_p1;
wire [4:0] sext_ln69_3_fu_1284_p1;
wire [31:0] sext_ln69_4_fu_1488_p1;
wire [4:0] sext_ln69_fu_1280_p1;
wire [7:0] sext_ln703_1_fu_926_p0;
wire [12:0] sext_ln703_1_fu_926_p1;
wire [31:0] sext_ln703_2_fu_628_p0;
wire [32:0] sext_ln703_2_fu_628_p1;
wire [34:0] sext_ln703_3_fu_1334_p1;
wire [15:0] sext_ln703_4_fu_1397_p0;
wire [45:0] sext_ln703_4_fu_1397_p1;
wire [31:0] sext_ln703_fu_274_p0;
wire [32:0] sext_ln703_fu_274_p1;
wire [18:0] sext_ln850_fu_1318_p1;
wire [7:0] shl_ln_fu_421_p3;
wire signbit_fu_249_p2;
wire tmp_10_fu_822_p3;
wire tmp_11_fu_829_p3;
wire [14:0] tmp_13_fu_239_p4;
wire [20:0] tmp_18_fu_1352_p3;
wire tmp_4_fu_1030_p3;
wire tmp_fu_1023_p3;
wire [1:0] trunc_ln1115_fu_318_p1;
wire [3:0] trunc_ln728_fu_1147_p1;
wire [2:0] trunc_ln851_1_fu_405_p1;
wire [1:0] trunc_ln851_2_fu_1197_p1;
wire [31:0] trunc_ln851_3_fu_648_p0;
wire [15:0] trunc_ln851_3_fu_648_p1;
wire [3:0] trunc_ln851_4_fu_1258_p1;
wire [1:0] trunc_ln851_5_fu_1276_p1;
wire [15:0] trunc_ln851_6_fu_1441_p0;
wire [12:0] trunc_ln851_6_fu_1441_p1;
wire [6:0] trunc_ln851_fu_294_p1;
wire xor_ln365_1_fu_1043_p2;
wire xor_ln365_2_fu_836_p2;
wire xor_ln365_3_fu_842_p2;
wire xor_ln365_fu_1037_p2;
wire xor_ln416_1_fu_561_p2;
wire xor_ln416_fu_720_p2;
wire xor_ln780_1_fu_756_p2;
wire xor_ln780_fu_959_p2;
wire xor_ln781_1_fu_778_p2;
wire xor_ln781_fu_979_p2;
wire xor_ln785_1_fu_1001_p2;
wire xor_ln785_2_fu_789_p2;
wire xor_ln785_3_fu_800_p2;
wire xor_ln785_fu_990_p2;
wire xor_ln786_1_fu_897_p2;
wire xor_ln786_fu_1105_p2;
wire [7:0] zext_ln1116_fu_606_p1;
wire [7:0] zext_ln1116_reg_1681;
wire [32:0] zext_ln1192_fu_624_p1;
wire [6:0] zext_ln1193_1_fu_385_p1;
wire [6:0] zext_ln1193_fu_381_p1;
wire [12:0] zext_ln1196_fu_936_p1;
wire [31:0] zext_ln1496_fu_428_p1;
wire [3:0] zext_ln415_1_fu_543_p1;
wire [3:0] zext_ln415_fu_702_p1;
wire [2:0] zext_ln69_1_fu_662_p1;
wire [31:0] zext_ln69_fu_1479_p1;


assign add_ln691_1_fu_1385_p2 = ret_V_34_cast_reg_1829 + 1'h1;
assign add_ln691_2_fu_1458_p2 = ret_V_36_cast_reg_1851 + 1'h1;
assign add_ln691_fu_1328_p2 = $signed(tmp_3_reg_1799) + $signed(2'h1);
assign add_ln69_1_fu_666_p2 = $signed(ret_V_19_fu_456_p3) + $signed({ 1'h0, icmp_ln874_fu_610_p2 });
assign add_ln69_2_fu_1287_p2 = $signed(add_ln69_1_reg_1703) + $signed(ret_V_20_fu_1162_p2[5:2]);
assign add_ln69_fu_1483_p2 = ret_V_28_reg_1863 + { ret_V_23_reg_1819[5], ret_V_23_reg_1819[5], ret_V_23_reg_1819[5], ret_V_23_reg_1819[5], ret_V_23_reg_1819[5], ret_V_23_reg_1819[5], ret_V_23_reg_1819[5], ret_V_23_reg_1819[5], ret_V_23_reg_1819[5], ret_V_23_reg_1819[5], ret_V_23_reg_1819 };
assign op_28 = $signed(add_ln69_2_reg_1814) + $signed(add_ln69_fu_1483_p2);
assign p_Val2_3_fu_706_p2 = r_V_3_reg_1605[5:2] + and_ln406_fu_696_p2;
assign p_Val2_7_fu_547_p2 = r_V_4_reg_1532[5:2] + and_ln408_fu_537_p2;
assign ret_V_13_fu_921_p2 = ret_V_12_reg_1691 + 1'h1;
assign ret_V_24_fu_632_p2 = $signed({ 1'h0, lhs_V_4_fu_601_p2, 16'h0000 }) + $signed(op_11);
assign ret_V_25_fu_1242_p2 = $signed({ select_ln850_5_fu_1223_p3, 7'h00 }) + $signed({ ret_V_3_fu_940_p2, 3'h0 });
assign { ret_V_26_fu_1364_p2[34], ret_V_26_fu_1364_p2[20:0] } = $signed({ select_ln353_fu_1344_p3, 2'h0 }) + $signed(op_14_V_reg_1772);
assign ret_V_27_fu_1425_p2 = $signed({ select_ln353_1_fu_1406_p3, 13'h0000 }) + $signed(op_15);
assign ret_V_6_fu_415_p2 = ret_V_21_fu_389_p2[6:3] + 1'h1;
assign ret_V_9_fu_1300_p2 = ret_V_7_reg_1782 + 1'h1;
assign ret_V_fu_445_p2 = ret_V_cast_reg_1520 + 1'h1;
assign _064_ = ap_CS_fsm[6] & icmp_ln851_5_reg_1836;
assign _065_ = ap_CS_fsm[3] & _068_;
assign _066_ = ap_CS_fsm[0] & _069_;
assign _067_ = ap_CS_fsm[0] & ap_start;
assign and_ln340_1_fu_903_p2 = xor_ln786_1_fu_897_p2 & or_ln340_1_fu_816_p2;
assign and_ln340_fu_1111_p2 = xor_ln786_fu_1105_p2 & or_ln340_fu_1017_p2;
assign and_ln406_fu_696_p2 = r_V_3_reg_1605[1] & or_ln406_fu_691_p2;
assign and_ln408_fu_537_p2 = r_V_4_reg_1532[0] & p_Result_27_fu_529_p2;
assign and_ln780_1_fu_761_p2 = xor_ln780_1_fu_756_p2 & Range2_all_ones_1_reg_1664;
assign and_ln780_fu_964_p2 = xor_ln780_fu_959_p2 & Range2_all_ones_reg_1735;
assign and_ln781_1_fu_773_p2 = carry_3_fu_746_p2 & Range1_all_ones_1_reg_1669;
assign and_ln781_fu_975_p2 = carry_1_reg_1728 & Range1_all_ones_reg_1740;
assign and_ln785_1_fu_1086_p2 = or_ln785_2_fu_1081_p2 & and_ln786_fu_1012_p2;
assign and_ln785_2_fu_1099_p2 = xor_ln785_1_fu_1001_p2 & and_ln786_fu_1012_p2;
assign and_ln785_4_fu_875_p2 = xor_ln416_1_reg_1658 & deleted_zeros_1_fu_750_p3;
assign and_ln785_5_fu_885_p2 = or_ln785_3_fu_880_p2 & and_ln786_1_fu_811_p2;
assign and_ln785_6_fu_891_p2 = xor_ln785_3_fu_800_p2 & and_ln786_1_fu_811_p2;
assign and_ln785_fu_1076_p2 = xor_ln416_reg_1723 & deleted_zeros_fu_954_p3;
assign and_ln786_1_fu_811_p2 = p_Result_29_reg_1652 & deleted_ones_1_fu_766_p3;
assign and_ln786_fu_1012_p2 = p_Result_24_reg_1717 & deleted_ones_fu_969_p3;
assign carry_1_fu_726_p2 = xor_ln416_fu_720_p2 & p_Result_23_reg_1621;
assign carry_3_fu_746_p2 = xor_ln416_1_reg_1658 & p_Result_28_reg_1551;
assign neg_src_4_fu_784_p2 = xor_ln781_1_fu_778_p2 & p_Result_26_reg_1544;
assign neg_src_fu_985_p2 = xor_ln781_fu_979_p2 & p_Result_21_reg_1613;
assign overflow_1_fu_805_p2 = xor_ln785_3_fu_800_p2 & or_ln785_1_fu_795_p2;
assign overflow_fu_1006_p2 = xor_ln785_1_fu_1001_p2 & or_ln785_fu_996_p2;
assign ret_V_20_fu_1162_p2 = { op_9_V_fu_1141_p3[3], op_9_V_fu_1141_p3[3], op_9_V_fu_1141_p3 } & { op_8[3:0], 2'h0 };
assign sel_tmp11_fu_1123_p2 = xor_ln365_1_fu_1043_p2 & or_ln340_3_fu_1117_p2;
assign sel_tmp25_fu_915_p2 = xor_ln365_3_fu_842_p2 & or_ln340_5_fu_909_p2;
assign xor_ln781_1_fu_778_p2 = ~ and_ln781_1_fu_773_p2;
assign xor_ln785_2_fu_789_p2 = ~ deleted_zeros_1_fu_750_p3;
assign xor_ln785_3_fu_800_p2 = ~ p_Result_26_reg_1544;
assign xor_ln780_1_fu_756_p2 = ~ p_Result_30_reg_1556;
assign xor_ln786_1_fu_897_p2 = ~ and_ln786_1_fu_811_p2;
assign xor_ln781_fu_979_p2 = ~ and_ln781_fu_975_p2;
assign xor_ln785_fu_990_p2 = ~ deleted_zeros_fu_954_p3;
assign xor_ln785_1_fu_1001_p2 = ~ p_Result_21_reg_1613;
assign xor_ln780_fu_959_p2 = ~ p_Result_25_reg_1626;
assign xor_ln786_fu_1105_p2 = ~ and_ln786_fu_1012_p2;
assign xor_ln416_fu_720_p2 = ~ p_Val2_3_fu_706_p2[3];
assign lhs_V_4_fu_601_p2 = ~ icmp_ln1496_reg_1594;
assign xor_ln365_1_fu_1043_p2 = ~ xor_ln365_fu_1037_p2;
assign xor_ln365_3_fu_842_p2 = ~ xor_ln365_2_fu_836_p2;
assign xor_ln416_1_fu_561_p2 = ~ p_Val2_7_fu_547_p2[3];
assign p_Val2_4_fu_1049_p2 = ~ p_Val2_3_reg_1708[2:0];
assign p_Val2_8_fu_848_p2 = ~ p_Val2_7_reg_1643[2:0];
assign _068_ = ~ icmp_ln851_3_reg_1698;
assign _069_ = ~ ap_start;
assign _070_ = tmp_2_reg_1567 == 5'h1f;
assign _071_ = p_Result_1_reg_1637 == 10'h3ff;
assign _072_ = ! tmp_2_reg_1567;
assign _073_ = ! p_Result_1_reg_1637;
assign _074_ = tmp_1_reg_1562 == 4'hf;
assign _075_ = p_Result_s_22_reg_1632 == 9'h1ff;
assign _076_ = ! ret_V_21_fu_389_p2[2:0];
assign _077_ = ! r_V_fu_1182_p2[1:0];
assign _078_ = ! op_11[15:0];
assign _079_ = ! ret_V_18_fu_278_p2[6:0];
assign \mul_4ns_4s_8_1_1_U3.top_mul_4ns_4s_8_1_1_Multiplier_2_U.p  = $signed({ 1'h0, \mul_4ns_4s_8_1_1_U3.top_mul_4ns_4s_8_1_1_Multiplier_2_U.a  }) * $signed(\mul_4ns_4s_8_1_1_U3.top_mul_4ns_4s_8_1_1_Multiplier_2_U.b );
assign \mul_8ns_8s_16_1_1_U2.top_mul_8ns_8s_16_1_1_Multiplier_1_U.p  = $signed({ 1'h0, \mul_8ns_8s_16_1_1_U2.top_mul_8ns_8s_16_1_1_Multiplier_1_U.a  }) * $signed(\mul_8ns_8s_16_1_1_U2.top_mul_8ns_8s_16_1_1_Multiplier_1_U.b );
assign \mul_8s_3ns_11_1_1_U1.top_mul_8s_3ns_11_1_1_Multiplier_0_U.p  = $signed(\mul_8s_3ns_11_1_1_U1.top_mul_8s_3ns_11_1_1_Multiplier_0_U.a ) * $signed({ 1'h0, \mul_8s_3ns_11_1_1_U1.top_mul_8s_3ns_11_1_1_Multiplier_0_U.b  });
assign _080_ = $signed({ 1'h0, signbit_reg_1503, 7'h00 }) < $signed(op_6);
assign _081_ = $signed(op_1[15:1]) < $signed(2'h1);
assign _082_ = | { ret_V_3_fu_940_p2[3:0], 3'h0 };
assign _083_ = | trunc_ln851_5_reg_1809;
assign _084_ = | op_15[12:0];
assign _085_ = ret_V_22_fu_594_p3 != op_8;
assign _086_ = | trunc_ln1115_reg_1539;
assign or_ln340_1_fu_816_p2 = overflow_1_fu_805_p2 | neg_src_4_fu_784_p2;
assign or_ln340_2_fu_1063_p2 = or_ln340_fu_1017_p2 | and_ln786_fu_1012_p2;
assign or_ln340_3_fu_1117_p2 = and_ln785_2_fu_1099_p2 | and_ln340_fu_1111_p2;
assign or_ln340_4_fu_862_p2 = or_ln340_1_fu_816_p2 | and_ln786_1_fu_811_p2;
assign or_ln340_5_fu_909_p2 = and_ln785_6_fu_891_p2 | and_ln340_1_fu_903_p2;
assign or_ln340_fu_1017_p2 = overflow_fu_1006_p2 | neg_src_fu_985_p2;
assign or_ln406_fu_691_p2 = r_V_3_reg_1605[0] | p_Result_21_reg_1613;
assign or_ln785_1_fu_795_p2 = xor_ln785_2_fu_789_p2 | p_Result_29_reg_1652;
assign or_ln785_2_fu_1081_p2 = p_Result_21_reg_1613 | and_ln785_fu_1076_p2;
assign or_ln785_3_fu_880_p2 = p_Result_26_reg_1544 | and_ln785_4_fu_875_p2;
assign or_ln785_fu_996_p2 = xor_ln785_fu_990_p2 | p_Result_24_reg_1717;
always @(posedge ap_clk)
signbit_reg_1503 <= _054_;
always @(posedge ap_clk)
ret_V_28_reg_1863 <= _045_;
always @(posedge ap_clk)
ret_V_13_reg_1767 <= _037_;
always @(posedge ap_clk)
ret_V_27_reg_1846 <= _044_;
always @(posedge ap_clk)
ret_V_36_cast_reg_1851 <= _047_;
always @(posedge ap_clk)
icmp_ln851_6_reg_1858 <= _018_;
always @(posedge ap_clk)
ret_V_23_reg_1819 <= _040_;
always @(posedge ap_clk)
ret_V_26_reg_1824 <= _043_;
always @(posedge ap_clk)
ret_V_34_cast_reg_1829 <= _046_;
always @(posedge ap_clk)
icmp_ln851_5_reg_1836 <= _017_;
always @(posedge ap_clk)
ret_V_18_reg_1515 <= _038_;
always @(posedge ap_clk)
ret_V_cast_reg_1520 <= _051_;
always @(posedge ap_clk)
icmp_ln851_reg_1527 <= _019_;
always @(posedge ap_clk)
r_V_4_reg_1532 <= _034_;
always @(posedge ap_clk)
trunc_ln1115_reg_1539 <= _058_;
always @(posedge ap_clk)
p_Result_26_reg_1544 <= _026_;
always @(posedge ap_clk)
p_Result_28_reg_1551 <= _027_;
always @(posedge ap_clk)
p_Result_30_reg_1556 <= _029_;
always @(posedge ap_clk)
tmp_1_reg_1562 <= _055_;
always @(posedge ap_clk)
tmp_2_reg_1567 <= _056_;
always @(posedge ap_clk)
_213_ <= _039_;
assign ret_V_21_reg_1573[6:3] = _213_;
always @(posedge ap_clk)
ret_V_6_cast_reg_1578 <= _048_;
always @(posedge ap_clk)
icmp_ln851_1_reg_1584 <= _013_;
always @(posedge ap_clk)
ret_V_6_reg_1589 <= _049_;
always @(posedge ap_clk)
icmp_ln1496_reg_1594 <= _012_;
always @(posedge ap_clk)
op_14_V_reg_1772 <= _020_;
always @(posedge ap_clk)
r_V_reg_1777 <= _035_;
always @(posedge ap_clk)
ret_V_7_reg_1782 <= _050_;
always @(posedge ap_clk)
icmp_ln851_2_reg_1789 <= _014_;
always @(posedge ap_clk)
_222_ <= _042_;
assign ret_V_25_reg_1794[24:3] = _222_;
always @(posedge ap_clk)
tmp_3_reg_1799 <= _057_;
always @(posedge ap_clk)
icmp_ln851_4_reg_1804 <= _016_;
always @(posedge ap_clk)
trunc_ln851_5_reg_1809 <= _059_;
always @(posedge ap_clk)
add_ln69_2_reg_1814 <= _008_;
always @(posedge ap_clk)
add_ln691_1_reg_1841 <= _006_;
always @(posedge ap_clk)
p_Val2_3_reg_1708 <= _031_;
always @(posedge ap_clk)
p_Result_24_reg_1717 <= _024_;
always @(posedge ap_clk)
xor_ln416_reg_1723 <= _061_;
always @(posedge ap_clk)
carry_1_reg_1728 <= _011_;
always @(posedge ap_clk)
Range2_all_ones_reg_1735 <= _005_;
always @(posedge ap_clk)
Range1_all_ones_reg_1740 <= _001_;
always @(posedge ap_clk)
Range1_all_zeros_reg_1747 <= _003_;
always @(posedge ap_clk)
select_ln340_1_reg_1752 <= _053_;
always @(posedge ap_clk)
and_ln785_5_reg_1757 <= _009_;
always @(posedge ap_clk)
sel_tmp25_reg_1762 <= _052_;
always @(posedge ap_clk)
r_V_3_reg_1605 <= _033_;
always @(posedge ap_clk)
p_Result_21_reg_1613 <= _022_;
always @(posedge ap_clk)
p_Result_23_reg_1621 <= _023_;
always @(posedge ap_clk)
p_Result_25_reg_1626 <= _025_;
always @(posedge ap_clk)
p_Result_s_22_reg_1632 <= _030_;
always @(posedge ap_clk)
p_Result_1_reg_1637 <= _021_;
always @(posedge ap_clk)
p_Val2_7_reg_1643 <= _032_;
always @(posedge ap_clk)
p_Result_29_reg_1652 <= _028_;
always @(posedge ap_clk)
xor_ln416_1_reg_1658 <= _060_;
always @(posedge ap_clk)
Range2_all_ones_1_reg_1664 <= _004_;
always @(posedge ap_clk)
Range1_all_ones_1_reg_1669 <= _000_;
always @(posedge ap_clk)
Range1_all_zeros_1_reg_1676 <= _002_;
always @(posedge ap_clk)
_250_ <= _062_;
assign zext_ln1116_reg_1681[3:0] = _250_;
always @(posedge ap_clk)
ret_V_24_reg_1686 <= _041_;
always @(posedge ap_clk)
ret_V_12_reg_1691 <= _036_;
always @(posedge ap_clk)
icmp_ln851_3_reg_1698 <= _015_;
always @(posedge ap_clk)
add_ln69_1_reg_1703 <= _007_;
always @(posedge ap_clk)
ap_CS_fsm <= _010_;
assign _063_ = _067_ ? 2'h2 : 2'h1;
assign _087_ = ap_CS_fsm == 1'h1;
function [9:0] _258_;
input [9:0] a;
input [99:0] b;
input [9:0] s;
case (s)
10'b0000000001:
_258_ = b[9:0];
10'b0000000010:
_258_ = b[19:10];
10'b0000000100:
_258_ = b[29:20];
10'b0000001000:
_258_ = b[39:30];
10'b0000010000:
_258_ = b[49:40];
10'b0000100000:
_258_ = b[59:50];
10'b0001000000:
_258_ = b[69:60];
10'b0010000000:
_258_ = b[79:70];
10'b0100000000:
_258_ = b[89:80];
10'b1000000000:
_258_ = b[99:90];
10'b0000000000:
_258_ = a;
default:
_258_ = 10'bx;
endcase
endfunction
assign ap_NS_fsm = _258_(10'hxxx, { 8'h00, _063_, 90'h00402010080402010080001 }, { _087_, _096_, _095_, _094_, _093_, _092_, _091_, _090_, _089_, _088_ });
assign _088_ = ap_CS_fsm == 10'h200;
assign _089_ = ap_CS_fsm == 9'h100;
assign _090_ = ap_CS_fsm == 8'h80;
assign _091_ = ap_CS_fsm == 7'h40;
assign _092_ = ap_CS_fsm == 6'h20;
assign _093_ = ap_CS_fsm == 5'h10;
assign _094_ = ap_CS_fsm == 4'h8;
assign _095_ = ap_CS_fsm == 3'h4;
assign _096_ = ap_CS_fsm == 2'h2;
assign op_28_ap_vld = ap_CS_fsm[9] ? 1'h1 : 1'h0;
assign ap_idle = _066_ ? 1'h1 : 1'h0;
assign _054_ = ap_CS_fsm[0] ? signbit_fu_249_p2 : signbit_reg_1503;
assign _045_ = ap_CS_fsm[8] ? ret_V_28_fu_1469_p3 : ret_V_28_reg_1863;
assign _037_ = _065_ ? ret_V_13_fu_921_p2 : ret_V_13_reg_1767;
assign _018_ = ap_CS_fsm[7] ? icmp_ln851_6_fu_1445_p2 : icmp_ln851_6_reg_1858;
assign _047_ = ap_CS_fsm[7] ? ret_V_27_fu_1425_p2[44:13] : ret_V_36_cast_reg_1851;
assign _044_ = ap_CS_fsm[7] ? ret_V_27_fu_1425_p2 : ret_V_27_reg_1846;
assign _017_ = ap_CS_fsm[5] ? icmp_ln851_5_fu_1380_p2 : icmp_ln851_5_reg_1836;
assign _046_ = ap_CS_fsm[5] ? { ret_V_26_fu_1364_p2[34], ret_V_26_fu_1364_p2[34], ret_V_26_fu_1364_p2[34], ret_V_26_fu_1364_p2[34], ret_V_26_fu_1364_p2[34], ret_V_26_fu_1364_p2[34], ret_V_26_fu_1364_p2[34], ret_V_26_fu_1364_p2[34], ret_V_26_fu_1364_p2[34], ret_V_26_fu_1364_p2[34], ret_V_26_fu_1364_p2[34], ret_V_26_fu_1364_p2[34], ret_V_26_fu_1364_p2[34], ret_V_26_fu_1364_p2[20:2] } : ret_V_34_cast_reg_1829;
assign _043_ = ap_CS_fsm[5] ? { ret_V_26_fu_1364_p2[34], ret_V_26_fu_1364_p2[34], ret_V_26_fu_1364_p2[34], ret_V_26_fu_1364_p2[34], ret_V_26_fu_1364_p2[34], ret_V_26_fu_1364_p2[34], ret_V_26_fu_1364_p2[34], ret_V_26_fu_1364_p2[34], ret_V_26_fu_1364_p2[34], ret_V_26_fu_1364_p2[34], ret_V_26_fu_1364_p2[34], ret_V_26_fu_1364_p2[34], ret_V_26_fu_1364_p2[34], ret_V_26_fu_1364_p2[34], ret_V_26_fu_1364_p2[20:0] } : ret_V_26_reg_1824;
assign _040_ = ap_CS_fsm[5] ? ret_V_23_fu_1311_p3 : ret_V_23_reg_1819;
assign _012_ = ap_CS_fsm[1] ? icmp_ln1496_fu_432_p2 : icmp_ln1496_reg_1594;
assign _049_ = ap_CS_fsm[1] ? ret_V_6_fu_415_p2 : ret_V_6_reg_1589;
assign _013_ = ap_CS_fsm[1] ? icmp_ln851_1_fu_409_p2 : icmp_ln851_1_reg_1584;
assign _048_ = ap_CS_fsm[1] ? ret_V_21_fu_389_p2[6:3] : ret_V_6_cast_reg_1578;
assign _039_ = ap_CS_fsm[1] ? ret_V_21_fu_389_p2[6:3] : ret_V_21_reg_1573[6:3];
assign _056_ = ap_CS_fsm[1] ? r_V_4_fu_312_p2[10:6] : tmp_2_reg_1567;
assign _055_ = ap_CS_fsm[1] ? r_V_4_fu_312_p2[10:7] : tmp_1_reg_1562;
assign _029_ = ap_CS_fsm[1] ? r_V_4_fu_312_p2[6] : p_Result_30_reg_1556;
assign _027_ = ap_CS_fsm[1] ? r_V_4_fu_312_p2[5] : p_Result_28_reg_1551;
assign _026_ = ap_CS_fsm[1] ? r_V_4_fu_312_p2[10] : p_Result_26_reg_1544;
assign _058_ = ap_CS_fsm[1] ? r_V_4_fu_312_p2[1:0] : trunc_ln1115_reg_1539;
assign _034_ = ap_CS_fsm[1] ? r_V_4_fu_312_p2 : r_V_4_reg_1532;
assign _019_ = ap_CS_fsm[1] ? icmp_ln851_fu_298_p2 : icmp_ln851_reg_1527;
assign _051_ = ap_CS_fsm[1] ? ret_V_18_fu_278_p2[8:7] : ret_V_cast_reg_1520;
assign _038_ = ap_CS_fsm[1] ? ret_V_18_fu_278_p2 : ret_V_18_reg_1515;
assign _008_ = ap_CS_fsm[4] ? add_ln69_2_fu_1287_p2 : add_ln69_2_reg_1814;
assign _059_ = ap_CS_fsm[4] ? op_14_V_fu_1129_p3[1:0] : trunc_ln851_5_reg_1809;
assign _016_ = ap_CS_fsm[4] ? icmp_ln851_4_fu_1270_p2 : icmp_ln851_4_reg_1804;
assign _057_ = ap_CS_fsm[4] ? ret_V_25_fu_1242_p2[24:7] : tmp_3_reg_1799;
assign _042_ = ap_CS_fsm[4] ? ret_V_25_fu_1242_p2[24:3] : ret_V_25_reg_1794[24:3];
assign _014_ = ap_CS_fsm[4] ? icmp_ln851_2_fu_1201_p2 : icmp_ln851_2_reg_1789;
assign _050_ = ap_CS_fsm[4] ? r_V_fu_1182_p2[7:2] : ret_V_7_reg_1782;
assign _035_ = ap_CS_fsm[4] ? r_V_fu_1182_p2 : r_V_reg_1777;
assign _020_ = ap_CS_fsm[4] ? op_14_V_fu_1129_p3 : op_14_V_reg_1772;
assign _006_ = _064_ ? add_ln691_1_fu_1385_p2 : add_ln691_1_reg_1841;
assign _052_ = ap_CS_fsm[3] ? sel_tmp25_fu_915_p2 : sel_tmp25_reg_1762;
assign _009_ = ap_CS_fsm[3] ? and_ln785_5_fu_885_p2 : and_ln785_5_reg_1757;
assign _053_ = ap_CS_fsm[3] ? select_ln340_1_fu_868_p3 : select_ln340_1_reg_1752;
assign _003_ = ap_CS_fsm[3] ? Range1_all_zeros_fu_741_p2 : Range1_all_zeros_reg_1747;
assign _001_ = ap_CS_fsm[3] ? Range1_all_ones_fu_736_p2 : Range1_all_ones_reg_1740;
assign _005_ = ap_CS_fsm[3] ? Range2_all_ones_fu_731_p2 : Range2_all_ones_reg_1735;
assign _011_ = ap_CS_fsm[3] ? carry_1_fu_726_p2 : carry_1_reg_1728;
assign _061_ = ap_CS_fsm[3] ? xor_ln416_fu_720_p2 : xor_ln416_reg_1723;
assign _024_ = ap_CS_fsm[3] ? p_Val2_3_fu_706_p2[3] : p_Result_24_reg_1717;
assign _031_ = ap_CS_fsm[3] ? p_Val2_3_fu_706_p2 : p_Val2_3_reg_1708;
assign _007_ = ap_CS_fsm[2] ? add_ln69_1_fu_666_p2 : add_ln69_1_reg_1703;
assign _015_ = ap_CS_fsm[2] ? icmp_ln851_3_fu_652_p2 : icmp_ln851_3_reg_1698;
assign _036_ = ap_CS_fsm[2] ? ret_V_24_fu_632_p2[32:16] : ret_V_12_reg_1691;
assign _041_ = ap_CS_fsm[2] ? ret_V_24_fu_632_p2 : ret_V_24_reg_1686;
assign _062_ = ap_CS_fsm[2] ? ret_V_22_fu_594_p3 : zext_ln1116_reg_1681[3:0];
assign _002_ = ap_CS_fsm[2] ? Range1_all_zeros_1_fu_577_p2 : Range1_all_zeros_1_reg_1676;
assign _000_ = ap_CS_fsm[2] ? Range1_all_ones_1_fu_572_p2 : Range1_all_ones_1_reg_1669;
assign _004_ = ap_CS_fsm[2] ? Range2_all_ones_1_fu_567_p2 : Range2_all_ones_1_reg_1664;
assign _060_ = ap_CS_fsm[2] ? xor_ln416_1_fu_561_p2 : xor_ln416_1_reg_1658;
assign _028_ = ap_CS_fsm[2] ? p_Val2_7_fu_547_p2[3] : p_Result_29_reg_1652;
assign _032_ = ap_CS_fsm[2] ? p_Val2_7_fu_547_p2 : p_Val2_7_reg_1643;
assign _021_ = ap_CS_fsm[2] ? r_V_3_fu_470_p2[15:6] : p_Result_1_reg_1637;
assign _030_ = ap_CS_fsm[2] ? r_V_3_fu_470_p2[15:7] : p_Result_s_22_reg_1632;
assign _025_ = ap_CS_fsm[2] ? r_V_3_fu_470_p2[6] : p_Result_25_reg_1626;
assign _023_ = ap_CS_fsm[2] ? r_V_3_fu_470_p2[5] : p_Result_23_reg_1621;
assign _022_ = ap_CS_fsm[2] ? r_V_3_fu_470_p2[15] : p_Result_21_reg_1613;
assign _033_ = ap_CS_fsm[2] ? r_V_3_fu_470_p2 : r_V_3_reg_1605;
assign _010_ = ap_rst ? 10'h001 : ap_NS_fsm;
assign ret_V_18_fu_278_p2 = $signed({ op_1, 6'h00 }) - $signed(op_6);
assign ret_V_21_fu_389_p2 = { op_0, 4'h0 } - { signbit_reg_1503, 3'h0 };
assign Range1_all_ones_1_fu_572_p2 = _070_ ? 1'h1 : 1'h0;
assign Range1_all_ones_fu_736_p2 = _071_ ? 1'h1 : 1'h0;
assign Range1_all_zeros_1_fu_577_p2 = _072_ ? 1'h1 : 1'h0;
assign Range1_all_zeros_fu_741_p2 = _073_ ? 1'h1 : 1'h0;
assign Range2_all_ones_1_fu_567_p2 = _074_ ? 1'h1 : 1'h0;
assign Range2_all_ones_fu_731_p2 = _075_ ? 1'h1 : 1'h0;
assign deleted_ones_1_fu_766_p3 = carry_3_fu_746_p2 ? and_ln780_1_fu_761_p2 : Range1_all_ones_1_reg_1669;
assign deleted_ones_fu_969_p3 = carry_1_reg_1728 ? and_ln780_fu_964_p2 : Range1_all_ones_reg_1740;
assign deleted_zeros_1_fu_750_p3 = carry_3_fu_746_p2 ? Range1_all_ones_1_reg_1669 : Range1_all_zeros_1_reg_1676;
assign deleted_zeros_fu_954_p3 = carry_1_reg_1728 ? Range1_all_ones_reg_1740 : Range1_all_zeros_reg_1747;
assign icmp_ln1496_fu_432_p2 = _080_ ? 1'h1 : 1'h0;
assign icmp_ln851_1_fu_409_p2 = _076_ ? 1'h1 : 1'h0;
assign icmp_ln851_2_fu_1201_p2 = _077_ ? 1'h1 : 1'h0;
assign icmp_ln851_3_fu_652_p2 = _078_ ? 1'h1 : 1'h0;
assign icmp_ln851_4_fu_1270_p2 = _082_ ? 1'h1 : 1'h0;
assign icmp_ln851_5_fu_1380_p2 = _083_ ? 1'h1 : 1'h0;
assign icmp_ln851_6_fu_1445_p2 = _084_ ? 1'h1 : 1'h0;
assign icmp_ln851_fu_298_p2 = _079_ ? 1'h1 : 1'h0;
assign icmp_ln874_fu_610_p2 = _085_ ? 1'h1 : 1'h0;
assign op_14_V_fu_1129_p3 = sel_tmp11_fu_1123_p2 ? p_Val2_3_reg_1708 : select_ln785_fu_1092_p3;
assign op_9_V_fu_1141_p3 = sel_tmp25_reg_1762 ? p_Val2_7_reg_1643 : select_ln785_1_fu_1136_p3;
assign p_Result_27_fu_529_p2 = _086_ ? 1'h1 : 1'h0;
assign ret_V_19_fu_456_p3 = ret_V_18_reg_1515[32] ? select_ln850_fu_450_p3 : ret_V_cast_reg_1520;
assign ret_V_22_fu_594_p3 = ret_V_21_reg_1573[6] ? select_ln850_1_fu_589_p3 : ret_V_6_cast_reg_1578;
assign ret_V_23_fu_1311_p3 = r_V_reg_1777[7] ? select_ln850_2_fu_1305_p3 : ret_V_7_reg_1782;
assign ret_V_28_fu_1469_p3 = ret_V_27_reg_1846[45] ? select_ln850_6_fu_1463_p3 : ret_V_36_cast_reg_1851;
assign select_ln340_1_fu_868_p3 = or_ln340_4_fu_862_p2 ? { p_Result_30_reg_1556, p_Val2_8_fu_848_p2 } : p_Val2_7_reg_1643;
assign select_ln340_fu_1069_p3 = or_ln340_2_fu_1063_p2 ? { p_Result_25_reg_1626, p_Val2_4_fu_1049_p2 } : p_Val2_3_reg_1708;
assign select_ln353_1_fu_1406_p3 = ret_V_26_reg_1824[34] ? select_ln850_8_fu_1401_p3 : ret_V_34_cast_reg_1829;
assign select_ln353_fu_1344_p3 = ret_V_25_reg_1794[24] ? select_ln850_7_fu_1337_p3 : { tmp_3_reg_1799[17], tmp_3_reg_1799 };
assign select_ln785_1_fu_1136_p3 = and_ln785_5_reg_1757 ? p_Val2_7_reg_1643 : select_ln340_1_reg_1752;
assign select_ln785_fu_1092_p3 = and_ln785_1_fu_1086_p2 ? p_Val2_3_reg_1708 : select_ln340_fu_1069_p3;
assign select_ln850_1_fu_589_p3 = icmp_ln851_1_reg_1584 ? ret_V_6_cast_reg_1578 : ret_V_6_reg_1589;
assign select_ln850_2_fu_1305_p3 = icmp_ln851_2_reg_1789 ? ret_V_7_reg_1782 : ret_V_9_fu_1300_p2;
assign select_ln850_4_fu_1218_p3 = icmp_ln851_3_reg_1698 ? ret_V_12_reg_1691 : ret_V_13_reg_1767;
assign select_ln850_5_fu_1223_p3 = ret_V_24_reg_1686[32] ? select_ln850_4_fu_1218_p3 : ret_V_12_reg_1691;
assign select_ln850_6_fu_1463_p3 = icmp_ln851_6_reg_1858 ? add_ln691_2_fu_1458_p2 : ret_V_36_cast_reg_1851;
assign select_ln850_7_fu_1337_p3 = icmp_ln851_4_reg_1804 ? add_ln691_fu_1328_p2 : { tmp_3_reg_1799[17], tmp_3_reg_1799 };
assign select_ln850_8_fu_1401_p3 = icmp_ln851_5_reg_1836 ? add_ln691_1_reg_1841 : ret_V_34_cast_reg_1829;
assign select_ln850_fu_450_p3 = icmp_ln851_reg_1527 ? ret_V_cast_reg_1520 : ret_V_fu_445_p2;
assign signbit_fu_249_p2 = _081_ ? 1'h1 : 1'h0;
assign xor_ln365_2_fu_836_p2 = p_Val2_7_reg_1643[3] ^ r_V_4_reg_1532[6];
assign xor_ln365_fu_1037_p2 = r_V_3_reg_1605[6] ^ p_Val2_3_reg_1708[3];
assign ret_V_3_fu_940_p2 = { op_8, 4'h0 } ^ { op_4[7], op_4[7], op_4[7], op_4[7], op_4[7], op_4 };
assign ap_CS_fsm_state1 = ap_CS_fsm[0];
assign ap_CS_fsm_state10 = ap_CS_fsm[9];
assign ap_CS_fsm_state2 = ap_CS_fsm[1];
assign ap_CS_fsm_state3 = ap_CS_fsm[2];
assign ap_CS_fsm_state4 = ap_CS_fsm[3];
assign ap_CS_fsm_state5 = ap_CS_fsm[4];
assign ap_CS_fsm_state6 = ap_CS_fsm[5];
assign ap_CS_fsm_state7 = ap_CS_fsm[6];
assign ap_CS_fsm_state8 = ap_CS_fsm[7];
assign ap_CS_fsm_state9 = ap_CS_fsm[8];
assign ap_done = op_28_ap_vld;
assign ap_ready = op_28_ap_vld;
assign icmp_ln1496_fu_432_p1 = op_6;
assign lhs_V_2_fu_373_p3 = { op_0, 4'h0 };
assign lhs_V_5_fu_616_p3 = { lhs_V_4_fu_601_p2, 16'h0000 };
assign lhs_V_fu_1150_p3 = { op_8[3:0], 2'h0 };
assign lhs_fu_263_p3 = { op_1, 6'h00 };
assign op_12_V_fu_946_p3 = { ret_V_3_fu_940_p2, 3'h0 };
assign op_16_V_fu_1168_p4 = ret_V_20_fu_1162_p2[5:2];
assign op_5_V_fu_366_p3 = { signbit_reg_1503, 3'h0 };
assign p_Result_14_fu_853_p4 = { p_Result_30_reg_1556, p_Val2_8_fu_848_p2 };
assign p_Result_15_fu_582_p3 = ret_V_21_reg_1573[6];
assign p_Result_16_fu_1293_p3 = r_V_reg_1777[7];
assign p_Result_17_fu_1207_p3 = ret_V_24_reg_1686[32];
assign p_Result_18_fu_1321_p3 = ret_V_25_reg_1794[24];
assign p_Result_19_fu_1390_p3 = ret_V_26_reg_1824[34];
assign p_Result_20_fu_1451_p3 = ret_V_27_reg_1846[45];
assign p_Result_22_fu_681_p3 = r_V_3_reg_1605[1];
assign p_Result_24_fu_712_p3 = p_Val2_3_fu_706_p2[3];
assign p_Result_29_fu_553_p3 = p_Val2_7_fu_547_p2[3];
assign p_Result_5_fu_1262_p3 = { ret_V_3_fu_940_p2[3:0], 3'h0 };
assign p_Result_8_fu_1054_p4 = { p_Result_25_reg_1626, p_Val2_4_fu_1049_p2 };
assign p_Result_s_fu_438_p3 = ret_V_18_reg_1515[32];
assign p_Val2_2_fu_672_p4 = r_V_3_reg_1605[5:2];
assign p_Val2_6_fu_520_p4 = r_V_4_reg_1532[5:2];
assign r_1_fu_534_p1 = r_V_4_reg_1532[0];
assign r_V_3_fu_470_p0 = op_8;
assign r_V_3_fu_470_p00 = { 8'h00, op_8 };
assign r_V_4_fu_312_p1 = { op_0, 1'h0 };
assign r_V_4_fu_312_p10 = { 8'h00, op_0, 1'h0 };
assign r_V_fu_1182_p0 = zext_ln1116_reg_1681[3:0];
assign r_fu_688_p1 = r_V_3_reg_1605[0];
assign ret_V_26_fu_1364_p2[33:21] = { ret_V_26_fu_1364_p2[34], ret_V_26_fu_1364_p2[34], ret_V_26_fu_1364_p2[34], ret_V_26_fu_1364_p2[34], ret_V_26_fu_1364_p2[34], ret_V_26_fu_1364_p2[34], ret_V_26_fu_1364_p2[34], ret_V_26_fu_1364_p2[34], ret_V_26_fu_1364_p2[34], ret_V_26_fu_1364_p2[34], ret_V_26_fu_1364_p2[34], ret_V_26_fu_1364_p2[34], ret_V_26_fu_1364_p2[34] };
assign ret_V_6_cast_fu_395_p4 = ret_V_21_fu_389_p2[6:3];
assign ret_fu_255_p3 = { op_0, 1'h0 };
assign rhs_3_fu_1230_p3 = { select_ln850_5_fu_1223_p3, 7'h00 };
assign rhs_4_fu_1413_p3 = { select_ln353_1_fu_1406_p3, 13'h0000 };
assign rhs_fu_929_p3 = { op_8, 4'h0 };
assign sext_ln1192_1_fu_1238_p1 = { select_ln850_5_fu_1223_p3[16], select_ln850_5_fu_1223_p3, 7'h00 };
assign sext_ln1192_2_fu_1360_p1 = { select_ln353_fu_1344_p3[18], select_ln353_fu_1344_p3[18], select_ln353_fu_1344_p3[18], select_ln353_fu_1344_p3[18], select_ln353_fu_1344_p3[18], select_ln353_fu_1344_p3[18], select_ln353_fu_1344_p3[18], select_ln353_fu_1344_p3[18], select_ln353_fu_1344_p3[18], select_ln353_fu_1344_p3[18], select_ln353_fu_1344_p3[18], select_ln353_fu_1344_p3[18], select_ln353_fu_1344_p3[18], select_ln353_fu_1344_p3[18], select_ln353_fu_1344_p3, 2'h0 };
assign sext_ln1192_3_fu_1421_p1 = { select_ln353_1_fu_1406_p3[31], select_ln353_1_fu_1406_p3, 13'h0000 };
assign sext_ln1192_fu_1214_p1 = { ret_V_3_fu_940_p2[12], ret_V_3_fu_940_p2[12], ret_V_3_fu_940_p2[12], ret_V_3_fu_940_p2[12], ret_V_3_fu_940_p2[12], ret_V_3_fu_940_p2[12], ret_V_3_fu_940_p2[12], ret_V_3_fu_940_p2[12], ret_V_3_fu_940_p2[12], ret_V_3_fu_940_p2, 3'h0 };
assign sext_ln1193_fu_270_p1 = { op_1[15], op_1[15], op_1[15], op_1[15], op_1[15], op_1[15], op_1[15], op_1[15], op_1[15], op_1[15], op_1[15], op_1, 6'h00 };
assign sext_ln1194_fu_1158_p1 = { op_9_V_fu_1141_p3[3], op_9_V_fu_1141_p3[3], op_9_V_fu_1141_p3 };
assign sext_ln69_1_fu_1476_p1 = { ret_V_23_reg_1819[5], ret_V_23_reg_1819[5], ret_V_23_reg_1819[5], ret_V_23_reg_1819[5], ret_V_23_reg_1819[5], ret_V_23_reg_1819[5], ret_V_23_reg_1819[5], ret_V_23_reg_1819[5], ret_V_23_reg_1819[5], ret_V_23_reg_1819[5], ret_V_23_reg_1819 };
assign sext_ln69_2_fu_658_p1 = { ret_V_19_fu_456_p3[1], ret_V_19_fu_456_p3 };
assign sext_ln69_3_fu_1284_p1 = { add_ln69_1_reg_1703[2], add_ln69_1_reg_1703[2], add_ln69_1_reg_1703 };
assign sext_ln69_4_fu_1488_p1 = { add_ln69_2_reg_1814[4], add_ln69_2_reg_1814[4], add_ln69_2_reg_1814[4], add_ln69_2_reg_1814[4], add_ln69_2_reg_1814[4], add_ln69_2_reg_1814[4], add_ln69_2_reg_1814[4], add_ln69_2_reg_1814[4], add_ln69_2_reg_1814[4], add_ln69_2_reg_1814[4], add_ln69_2_reg_1814[4], add_ln69_2_reg_1814[4], add_ln69_2_reg_1814[4], add_ln69_2_reg_1814[4], add_ln69_2_reg_1814[4], add_ln69_2_reg_1814[4], add_ln69_2_reg_1814[4], add_ln69_2_reg_1814[4], add_ln69_2_reg_1814[4], add_ln69_2_reg_1814[4], add_ln69_2_reg_1814[4], add_ln69_2_reg_1814[4], add_ln69_2_reg_1814[4], add_ln69_2_reg_1814[4], add_ln69_2_reg_1814[4], add_ln69_2_reg_1814[4], add_ln69_2_reg_1814[4], add_ln69_2_reg_1814 };
assign sext_ln69_fu_1280_p1 = { ret_V_20_fu_1162_p2[5], ret_V_20_fu_1162_p2[5:2] };
assign sext_ln703_1_fu_926_p0 = op_4;
assign sext_ln703_1_fu_926_p1 = { op_4[7], op_4[7], op_4[7], op_4[7], op_4[7], op_4 };
assign sext_ln703_2_fu_628_p0 = op_11;
assign sext_ln703_2_fu_628_p1 = { op_11[31], op_11 };
assign sext_ln703_3_fu_1334_p1 = { op_14_V_reg_1772[3], op_14_V_reg_1772[3], op_14_V_reg_1772[3], op_14_V_reg_1772[3], op_14_V_reg_1772[3], op_14_V_reg_1772[3], op_14_V_reg_1772[3], op_14_V_reg_1772[3], op_14_V_reg_1772[3], op_14_V_reg_1772[3], op_14_V_reg_1772[3], op_14_V_reg_1772[3], op_14_V_reg_1772[3], op_14_V_reg_1772[3], op_14_V_reg_1772[3], op_14_V_reg_1772[3], op_14_V_reg_1772[3], op_14_V_reg_1772[3], op_14_V_reg_1772[3], op_14_V_reg_1772[3], op_14_V_reg_1772[3], op_14_V_reg_1772[3], op_14_V_reg_1772[3], op_14_V_reg_1772[3], op_14_V_reg_1772[3], op_14_V_reg_1772[3], op_14_V_reg_1772[3], op_14_V_reg_1772[3], op_14_V_reg_1772[3], op_14_V_reg_1772[3], op_14_V_reg_1772[3], op_14_V_reg_1772 };
assign sext_ln703_4_fu_1397_p0 = op_15;
assign sext_ln703_4_fu_1397_p1 = { op_15[15], op_15[15], op_15[15], op_15[15], op_15[15], op_15[15], op_15[15], op_15[15], op_15[15], op_15[15], op_15[15], op_15[15], op_15[15], op_15[15], op_15[15], op_15[15], op_15[15], op_15[15], op_15[15], op_15[15], op_15[15], op_15[15], op_15[15], op_15[15], op_15[15], op_15[15], op_15[15], op_15[15], op_15[15], op_15[15], op_15 };
assign sext_ln703_fu_274_p0 = op_6;
assign sext_ln703_fu_274_p1 = { op_6[31], op_6 };
assign sext_ln850_fu_1318_p1 = { tmp_3_reg_1799[17], tmp_3_reg_1799 };
assign shl_ln_fu_421_p3 = { signbit_reg_1503, 7'h00 };
assign tmp_10_fu_822_p3 = r_V_4_reg_1532[6];
assign tmp_11_fu_829_p3 = p_Val2_7_reg_1643[3];
assign tmp_13_fu_239_p4 = op_1[15:1];
assign tmp_18_fu_1352_p3 = { select_ln353_fu_1344_p3, 2'h0 };
assign tmp_4_fu_1030_p3 = p_Val2_3_reg_1708[3];
assign tmp_fu_1023_p3 = r_V_3_reg_1605[6];
assign trunc_ln1115_fu_318_p1 = r_V_4_fu_312_p2[1:0];
assign trunc_ln728_fu_1147_p1 = op_8[3:0];
assign trunc_ln851_1_fu_405_p1 = ret_V_21_fu_389_p2[2:0];
assign trunc_ln851_2_fu_1197_p1 = r_V_fu_1182_p2[1:0];
assign trunc_ln851_3_fu_648_p0 = op_11;
assign trunc_ln851_3_fu_648_p1 = op_11[15:0];
assign trunc_ln851_4_fu_1258_p1 = ret_V_3_fu_940_p2[3:0];
assign trunc_ln851_5_fu_1276_p1 = op_14_V_fu_1129_p3[1:0];
assign trunc_ln851_6_fu_1441_p0 = op_15;
assign trunc_ln851_6_fu_1441_p1 = op_15[12:0];
assign trunc_ln851_fu_294_p1 = ret_V_18_fu_278_p2[6:0];
assign zext_ln1116_fu_606_p1 = { 4'h0, ret_V_22_fu_594_p3 };
assign zext_ln1192_fu_624_p1 = { 16'h0000, lhs_V_4_fu_601_p2, 16'h0000 };
assign zext_ln1193_1_fu_385_p1 = { 3'h0, signbit_reg_1503, 3'h0 };
assign zext_ln1193_fu_381_p1 = { 1'h0, op_0, 4'h0 };
assign zext_ln1196_fu_936_p1 = { 1'h0, op_8, 4'h0 };
assign zext_ln1496_fu_428_p1 = { 24'h000000, signbit_reg_1503, 7'h00 };
assign zext_ln415_1_fu_543_p1 = { 3'h0, and_ln408_fu_537_p2 };
assign zext_ln415_fu_702_p1 = { 3'h0, and_ln406_fu_696_p2 };
assign zext_ln69_1_fu_662_p1 = { 2'h0, icmp_ln874_fu_610_p2 };
assign zext_ln69_fu_1479_p1 = { 16'h0000, ret_V_23_reg_1819[5], ret_V_23_reg_1819[5], ret_V_23_reg_1819[5], ret_V_23_reg_1819[5], ret_V_23_reg_1819[5], ret_V_23_reg_1819[5], ret_V_23_reg_1819[5], ret_V_23_reg_1819[5], ret_V_23_reg_1819[5], ret_V_23_reg_1819[5], ret_V_23_reg_1819 };
assign \mul_8s_3ns_11_1_1_U1.top_mul_8s_3ns_11_1_1_Multiplier_0_U.a  = \mul_8s_3ns_11_1_1_U1.din0 ;
assign \mul_8s_3ns_11_1_1_U1.top_mul_8s_3ns_11_1_1_Multiplier_0_U.b  = \mul_8s_3ns_11_1_1_U1.din1 ;
assign \mul_8s_3ns_11_1_1_U1.dout  = \mul_8s_3ns_11_1_1_U1.top_mul_8s_3ns_11_1_1_Multiplier_0_U.p ;
assign \mul_8s_3ns_11_1_1_U1.din0  = op_4;
assign \mul_8s_3ns_11_1_1_U1.din1  = { op_0, 1'h0 };
assign r_V_4_fu_312_p2 = \mul_8s_3ns_11_1_1_U1.dout ;
assign \mul_8ns_8s_16_1_1_U2.top_mul_8ns_8s_16_1_1_Multiplier_1_U.a  = \mul_8ns_8s_16_1_1_U2.din0 ;
assign \mul_8ns_8s_16_1_1_U2.top_mul_8ns_8s_16_1_1_Multiplier_1_U.b  = \mul_8ns_8s_16_1_1_U2.din1 ;
assign \mul_8ns_8s_16_1_1_U2.dout  = \mul_8ns_8s_16_1_1_U2.top_mul_8ns_8s_16_1_1_Multiplier_1_U.p ;
assign \mul_8ns_8s_16_1_1_U2.din0  = op_8;
assign \mul_8ns_8s_16_1_1_U2.din1  = op_4;
assign r_V_3_fu_470_p2 = \mul_8ns_8s_16_1_1_U2.dout ;
assign \mul_4ns_4s_8_1_1_U3.top_mul_4ns_4s_8_1_1_Multiplier_2_U.a  = \mul_4ns_4s_8_1_1_U3.din0 ;
assign \mul_4ns_4s_8_1_1_U3.top_mul_4ns_4s_8_1_1_Multiplier_2_U.b  = \mul_4ns_4s_8_1_1_U3.din1 ;
assign \mul_4ns_4s_8_1_1_U3.dout  = \mul_4ns_4s_8_1_1_U3.top_mul_4ns_4s_8_1_1_Multiplier_2_U.p ;
assign \mul_4ns_4s_8_1_1_U3.din0  = zext_ln1116_reg_1681[3:0];
assign \mul_4ns_4s_8_1_1_U3.din1  = op_9_V_fu_1141_p3;
assign r_V_fu_1182_p2 = \mul_4ns_4s_8_1_1_U3.dout ;
endmodule


// Product machine:
module top_A_times_top_B (ap_start, op_0, op_1, op_11, op_15, op_4, op_6, op_8, ap_clk, unsafe_signal);
input ap_start;
input [1:0] op_0;
input [15:0] op_1;
input [31:0] op_11;
input [15:0] op_15;
input [7:0] op_4;
input [31:0] op_6;
input [7:0] op_8;
input ap_clk;
output unsafe_signal;
reg _setup;
initial _setup = 1'b0;
always @ (posedge ap_clk) _setup <= 1'b1;
reg ap_start_internal;
always @ (posedge ap_clk) if (!_setup) ap_start_internal <= ap_start;
reg [1:0] op_0_internal;
always @ (posedge ap_clk) if (!_setup) op_0_internal <= op_0;
reg [15:0] op_1_internal;
always @ (posedge ap_clk) if (!_setup) op_1_internal <= op_1;
reg [31:0] op_11_internal;
always @ (posedge ap_clk) if (!_setup) op_11_internal <= op_11;
reg [15:0] op_15_internal;
always @ (posedge ap_clk) if (!_setup) op_15_internal <= op_15;
reg [7:0] op_4_internal;
always @ (posedge ap_clk) if (!_setup) op_4_internal <= op_4;
reg [31:0] op_6_internal;
always @ (posedge ap_clk) if (!_setup) op_6_internal <= op_6;
reg [7:0] op_8_internal;
always @ (posedge ap_clk) if (!_setup) op_8_internal <= op_8;
wire ap_done_A;
wire ap_done_B;
wire ap_done_eq;
assign ap_done_eq = ap_done_A == ap_done_B;
wire ap_idle_A;
wire ap_idle_B;
wire ap_idle_eq;
assign ap_idle_eq = ap_idle_A == ap_idle_B;
wire ap_ready_A;
wire ap_ready_B;
wire ap_ready_eq;
assign ap_ready_eq = ap_ready_A == ap_ready_B;
wire [31:0] op_28_A;
wire [31:0] op_28_B;
wire op_28_eq;
assign op_28_eq = op_28_A == op_28_B;
wire op_28_ap_vld_A;
wire op_28_ap_vld_B;
wire clk_enable_A;
wire clk_enable_B;
assign clk_enable_A = _setup & (~op_28_ap_vld_A | op_28_ap_vld_B);
assign clk_enable_B = _setup;
wire divergent;
assign divergent = ~(ap_done_eq & ap_idle_eq & ap_ready_eq & op_28_eq);
assign unsafe_signal = op_28_ap_vld_A & op_28_ap_vld_B & divergent;
top_A instance_A (
    .ap_clk(ap_clk),
    .clk_enable(clk_enable_A),
    .ap_start(ap_start_internal),
    .op_0(op_0_internal),
    .op_1(op_1_internal),
    .op_11(op_11_internal),
    .op_15(op_15_internal),
    .op_4(op_4_internal),
    .op_6(op_6_internal),
    .op_8(op_8_internal),
    .ap_done(ap_done_A),
    .ap_idle(ap_idle_A),
    .ap_ready(ap_ready_A),
    .op_28(op_28_A),
    .op_28_ap_vld(op_28_ap_vld_A)
);
top_B instance_B (
    .ap_clk(ap_clk),
    .clk_enable(clk_enable_B),
    .ap_start(ap_start_internal),
    .op_0(op_0_internal),
    .op_1(op_1_internal),
    .op_11(op_11_internal),
    .op_15(op_15_internal),
    .op_4(op_4_internal),
    .op_6(op_6_internal),
    .op_8(op_8_internal),
    .ap_done(ap_done_B),
    .ap_idle(ap_idle_B),
    .ap_ready(ap_ready_B),
    .op_28(op_28_B),
    .op_28_ap_vld(op_28_ap_vld_B)
);
endmodule
