// Processed by function `construct_kairos` in `verilog_tricks.py`.
// Machine A:
// Processed by function `add_clk_enable_signal` in `verilog_tricks.py`.
// Processed by function `remove_reset_signal` in `verilog_tricks.py`.
module top_A (
  ap_clk,
  ap_start,
  ap_done,
  ap_idle,
  ap_ready,
  op_0,
  op_2,
  op_3,
  op_5,
  op_6,
  op_7,
  op_8,
  op_12,
  op_13,
  op_15,
  op_16,
  op_17,
  op_19,
  op_30,
  op_30_ap_vld,
clk_enable
);
input clk_enable;


input ap_clk;
wire ap_rst;
assign ap_rst = op_30_ap_vld;
input ap_start;
input [7:0] op_0;
input op_12;
input [3:0] op_13;
input [3:0] op_15;
input [1:0] op_16;
input [7:0] op_17;
input [3:0] op_19;
input [7:0] op_2;
input [3:0] op_3;
input op_5;
input [1:0] op_6;
input [31:0] op_7;
input [7:0] op_8;
output ap_done;
output ap_idle;
output ap_ready;
output [31:0] op_30;
output op_30_ap_vld;


reg [4:0] add_ln69_3_reg_533;
reg [4:0] ap_CS_fsm = 5'h01;
reg [31:0] op_21_V_reg_513;
reg [31:0] op_27_V_reg_538;
reg [8:0] ret_2_reg_508;
reg [31:0] ret_V_10_reg_528;
reg [31:0] ret_V_12_reg_543;
reg [7:0] ret_V_9_reg_523;
wire [4:0] _00_;
wire [4:0] _01_;
wire [31:0] _02_;
wire [31:0] _03_;
wire [8:0] _04_;
wire [31:0] _05_;
wire [31:0] _06_;
wire [7:0] _07_;
wire [1:0] _08_;
wire _09_;
wire _10_;
wire _11_;
wire _12_;
wire _13_;
wire _14_;
wire _15_;
wire _16_;
wire _17_;
wire _18_;
wire [31:0] add_ln691_fu_452_p2;
wire [31:0] add_ln69_2_fu_379_p2;
wire [4:0] add_ln69_3_fu_366_p2;
wire [5:0] add_ln69_4_fu_387_p2;
wire [8:0] add_ln69_fu_219_p2;
wire ap_CS_fsm_state1;
wire ap_CS_fsm_state2;
wire ap_CS_fsm_state3;
wire ap_CS_fsm_state4;
wire ap_CS_fsm_state5;
wire [4:0] ap_NS_fsm;
wire ap_clk;
wire ap_done;
wire ap_idle;
wire ap_ready;
wire ap_rst;
wire ap_start;
wire icmp_ln851_1_fu_446_p2;
wire icmp_ln851_fu_289_p2;
wire [21:0] lhs_fu_249_p3;
wire [7:0] op_0;
wire [1:0] op_10_V_fu_205_p2;
wire [2:0] op_11_V_fu_242_p3;
wire op_12;
wire [3:0] op_13;
wire [3:0] op_15;
wire [1:0] op_16;
wire [7:0] op_17;
wire [3:0] op_19;
wire [7:0] op_2;
wire [31:0] op_21_V_fu_229_p2;
wire [31:0] op_22_V_fu_334_p4;
wire [31:0] op_27_V_fu_397_p2;
wire [31:0] op_29_V_fu_487_p2;
wire [3:0] op_3;
wire [31:0] op_30;
wire op_30_ap_vld;
wire op_5;
wire [1:0] op_6;
wire [31:0] op_7;
wire [7:0] op_8;
wire [28:0] op_9_V_fu_235_p3;
wire p_Result_1_fu_434_p3;
wire p_Result_s_fu_277_p3;
wire [32:0] p_Val2_2_fu_328_p2;
wire [8:0] ret_2_fu_191_p2;
wire [31:0] ret_V_10_fu_352_p2;
wire [36:0] ret_V_11_fu_418_p2;
wire [31:0] ret_V_12_fu_466_p3;
wire [31:0] ret_V_6_cast_fu_424_p4;
wire [28:0] ret_V_8_fu_261_p2;
wire [7:0] ret_V_9_fu_309_p3;
wire [7:0] ret_V_cast_fu_267_p4;
wire [7:0] ret_V_fu_295_p2;
wire [2:0] ret_fu_477_p2;
wire [32:0] rhs_2_fu_321_p3;
wire [35:0] rhs_5_fu_407_p3;
wire [31:0] select_ln1192_fu_344_p3;
wire [31:0] select_ln850_1_fu_458_p3;
wire [7:0] select_ln850_fu_301_p3;
wire [31:0] sext_ln1192_1_fu_492_p1;
wire [36:0] sext_ln1192_fu_414_p1;
wire [7:0] sext_ln1346_fu_183_p0;
wire [8:0] sext_ln1346_fu_183_p1;
wire [31:0] sext_ln69_1_fu_225_p1;
wire [4:0] sext_ln69_2_fu_358_p1;
wire [31:0] sext_ln69_3_fu_372_p1;
wire [5:0] sext_ln69_4_fu_375_p1;
wire [4:0] sext_ln69_5_fu_362_p1;
wire [31:0] sext_ln69_6_fu_483_p1;
wire [5:0] sext_ln69_7_fu_384_p1;
wire [31:0] sext_ln69_8_fu_393_p1;
wire [8:0] sext_ln69_fu_215_p1;
wire [7:0] sext_ln703_fu_403_p0;
wire [36:0] sext_ln703_fu_403_p1;
wire [8:0] sext_ln727_fu_211_p1;
wire [7:0] trunc_ln69_fu_197_p0;
wire [1:0] trunc_ln69_fu_197_p1;
wire [7:0] trunc_ln851_1_fu_442_p0;
wire [3:0] trunc_ln851_1_fu_442_p1;
wire [19:0] trunc_ln851_fu_285_p1;
wire [32:0] zext_ln1192_fu_317_p1;
wire [28:0] zext_ln1193_fu_257_p1;
wire [8:0] zext_ln1346_fu_187_p1;
wire [2:0] zext_ln215_fu_474_p1;
wire [1:0] zext_ln69_fu_201_p1;


assign add_ln691_fu_452_p2 = ret_V_11_fu_418_p2[35:4] + 1'h1;
assign add_ln69_2_fu_379_p2 = $signed(ret_V_10_reg_528) + $signed(ret_V_9_reg_523);
assign add_ln69_3_fu_366_p2 = $signed(op_13) + $signed(op_16);
assign add_ln69_4_fu_387_p2 = $signed(add_ln69_3_reg_533) + $signed(op_15);
assign add_ln69_fu_219_p2 = $signed(op_8) + $signed(op_10_V_fu_205_p2);
assign op_10_V_fu_205_p2 = op_2[1:0] + op_5;
assign op_21_V_fu_229_p2 = $signed(add_ln69_fu_219_p2) + $signed(op_7);
assign op_27_V_fu_397_p2 = $signed(add_ln69_4_fu_387_p2) + $signed(add_ln69_2_fu_379_p2);
assign op_29_V_fu_487_p2 = $signed(ret_V_12_reg_543) + $signed(ret_fu_477_p2);
assign op_30 = $signed(op_29_V_fu_487_p2) + $signed(op_19);
assign p_Val2_2_fu_328_p2 = { op_21_V_reg_513, 1'h0 } + { op_5, 2'h0 };
assign ret_2_fu_191_p2 = $signed(op_2) + $signed({ 1'h0, op_3 });
assign ret_V_10_fu_352_p2 = p_Val2_2_fu_328_p2[32:1] + select_ln1192_fu_344_p3;
assign ret_V_11_fu_418_p2 = $signed({ op_27_V_reg_538, 4'h0 }) + $signed(op_17);
assign ret_V_fu_295_p2 = ret_V_8_fu_261_p2[27:20] + 1'h1;
assign _09_ = ap_CS_fsm[0] & _11_;
assign _10_ = ap_CS_fsm[0] & ap_start;
assign _11_ = ~ ap_start;
assign _12_ = ! ret_V_8_fu_261_p2[19:0];
assign _13_ = | op_17[3:0];
always @(posedge ap_clk)
ret_V_12_reg_543 <= _06_;
always @(posedge ap_clk)
op_27_V_reg_538 <= _03_;
always @(posedge ap_clk)
ret_2_reg_508 <= _04_;
always @(posedge ap_clk)
op_21_V_reg_513 <= _02_;
always @(posedge ap_clk)
ret_V_9_reg_523 <= _07_;
always @(posedge ap_clk)
ret_V_10_reg_528 <= _05_;
always @(posedge ap_clk)
add_ln69_3_reg_533 <= _00_;
always @(posedge ap_clk)
ap_CS_fsm <= _01_;
assign _01_ = ap_rst ? 5'h01 : ap_NS_fsm;
assign _08_ = _10_ ? 2'h2 : 2'h1;
assign _14_ = ap_CS_fsm == 1'h1;
function [4:0] _50_;
input [4:0] a;
input [24:0] b;
input [4:0] s;
case (s)
5'b00001:
_50_ = b[4:0];
5'b00010:
_50_ = b[9:5];
5'b00100:
_50_ = b[14:10];
5'b01000:
_50_ = b[19:15];
5'b10000:
_50_ = b[24:20];
5'b00000:
_50_ = a;
default:
_50_ = 5'bx;
endcase
endfunction
assign ap_NS_fsm = _50_(5'hxx, { 3'h0, _08_, 20'h22201 }, { _14_, _18_, _17_, _16_, _15_ });
assign _15_ = ap_CS_fsm == 5'h10;
assign _16_ = ap_CS_fsm == 4'h8;
assign _17_ = ap_CS_fsm == 3'h4;
assign _18_ = ap_CS_fsm == 2'h2;
assign op_30_ap_vld = ap_CS_fsm[4] ? 1'h1 : 1'h0;
assign ap_idle = _09_ ? 1'h1 : 1'h0;
assign _06_ = ap_CS_fsm[3] ? ret_V_12_fu_466_p3 : ret_V_12_reg_543;
assign _03_ = ap_CS_fsm[2] ? op_27_V_fu_397_p2 : op_27_V_reg_538;
assign _02_ = ap_CS_fsm[0] ? op_21_V_fu_229_p2 : op_21_V_reg_513;
assign _04_ = ap_CS_fsm[0] ? ret_2_fu_191_p2 : ret_2_reg_508;
assign _00_ = ap_CS_fsm[1] ? add_ln69_3_fu_366_p2 : add_ln69_3_reg_533;
assign _05_ = ap_CS_fsm[1] ? ret_V_10_fu_352_p2 : ret_V_10_reg_528;
assign _07_ = ap_CS_fsm[1] ? ret_V_9_fu_309_p3 : ret_V_9_reg_523;
assign ret_V_8_fu_261_p2 = { op_6, 20'h00000 } - { ret_2_reg_508, 20'h00000 };
assign ret_fu_477_p2 = 1'h0 - op_6;
assign icmp_ln851_1_fu_446_p2 = _13_ ? 1'h1 : 1'h0;
assign icmp_ln851_fu_289_p2 = _12_ ? 1'h1 : 1'h0;
assign ret_V_12_fu_466_p3 = ret_V_11_fu_418_p2[36] ? select_ln850_1_fu_458_p3 : ret_V_11_fu_418_p2[35:4];
assign ret_V_9_fu_309_p3 = ret_V_8_fu_261_p2[28] ? select_ln850_fu_301_p3 : ret_V_8_fu_261_p2[27:20];
assign select_ln1192_fu_344_p3 = op_12 ? 32'd4294967295 : 32'd0;
assign select_ln850_1_fu_458_p3 = icmp_ln851_1_fu_446_p2 ? add_ln691_fu_452_p2 : ret_V_11_fu_418_p2[35:4];
assign select_ln850_fu_301_p3 = icmp_ln851_fu_289_p2 ? ret_V_8_fu_261_p2[27:20] : ret_V_fu_295_p2;
assign ap_CS_fsm_state1 = ap_CS_fsm[0];
assign ap_CS_fsm_state2 = ap_CS_fsm[1];
assign ap_CS_fsm_state3 = ap_CS_fsm[2];
assign ap_CS_fsm_state4 = ap_CS_fsm[3];
assign ap_CS_fsm_state5 = ap_CS_fsm[4];
assign ap_done = op_30_ap_vld;
assign ap_ready = op_30_ap_vld;
assign lhs_fu_249_p3 = { op_6, 20'h00000 };
assign op_11_V_fu_242_p3 = { op_5, 2'h0 };
assign op_22_V_fu_334_p4 = p_Val2_2_fu_328_p2[32:1];
assign op_9_V_fu_235_p3 = { ret_2_reg_508, 20'h00000 };
assign p_Result_1_fu_434_p3 = ret_V_11_fu_418_p2[36];
assign p_Result_s_fu_277_p3 = ret_V_8_fu_261_p2[28];
assign ret_V_6_cast_fu_424_p4 = ret_V_11_fu_418_p2[35:4];
assign ret_V_cast_fu_267_p4 = ret_V_8_fu_261_p2[27:20];
assign rhs_2_fu_321_p3 = { op_21_V_reg_513, 1'h0 };
assign rhs_5_fu_407_p3 = { op_27_V_reg_538, 4'h0 };
assign sext_ln1192_1_fu_492_p1 = { op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19 };
assign sext_ln1192_fu_414_p1 = { op_27_V_reg_538[31], op_27_V_reg_538, 4'h0 };
assign sext_ln1346_fu_183_p0 = op_2;
assign sext_ln1346_fu_183_p1 = { op_2[7], op_2 };
assign sext_ln69_1_fu_225_p1 = { add_ln69_fu_219_p2[8], add_ln69_fu_219_p2[8], add_ln69_fu_219_p2[8], add_ln69_fu_219_p2[8], add_ln69_fu_219_p2[8], add_ln69_fu_219_p2[8], add_ln69_fu_219_p2[8], add_ln69_fu_219_p2[8], add_ln69_fu_219_p2[8], add_ln69_fu_219_p2[8], add_ln69_fu_219_p2[8], add_ln69_fu_219_p2[8], add_ln69_fu_219_p2[8], add_ln69_fu_219_p2[8], add_ln69_fu_219_p2[8], add_ln69_fu_219_p2[8], add_ln69_fu_219_p2[8], add_ln69_fu_219_p2[8], add_ln69_fu_219_p2[8], add_ln69_fu_219_p2[8], add_ln69_fu_219_p2[8], add_ln69_fu_219_p2[8], add_ln69_fu_219_p2[8], add_ln69_fu_219_p2 };
assign sext_ln69_2_fu_358_p1 = { op_13[3], op_13 };
assign sext_ln69_3_fu_372_p1 = { ret_V_9_reg_523[7], ret_V_9_reg_523[7], ret_V_9_reg_523[7], ret_V_9_reg_523[7], ret_V_9_reg_523[7], ret_V_9_reg_523[7], ret_V_9_reg_523[7], ret_V_9_reg_523[7], ret_V_9_reg_523[7], ret_V_9_reg_523[7], ret_V_9_reg_523[7], ret_V_9_reg_523[7], ret_V_9_reg_523[7], ret_V_9_reg_523[7], ret_V_9_reg_523[7], ret_V_9_reg_523[7], ret_V_9_reg_523[7], ret_V_9_reg_523[7], ret_V_9_reg_523[7], ret_V_9_reg_523[7], ret_V_9_reg_523[7], ret_V_9_reg_523[7], ret_V_9_reg_523[7], ret_V_9_reg_523[7], ret_V_9_reg_523 };
assign sext_ln69_4_fu_375_p1 = { op_15[3], op_15[3], op_15 };
assign sext_ln69_5_fu_362_p1 = { op_16[1], op_16[1], op_16[1], op_16 };
assign sext_ln69_6_fu_483_p1 = { ret_fu_477_p2[2], ret_fu_477_p2[2], ret_fu_477_p2[2], ret_fu_477_p2[2], ret_fu_477_p2[2], ret_fu_477_p2[2], ret_fu_477_p2[2], ret_fu_477_p2[2], ret_fu_477_p2[2], ret_fu_477_p2[2], ret_fu_477_p2[2], ret_fu_477_p2[2], ret_fu_477_p2[2], ret_fu_477_p2[2], ret_fu_477_p2[2], ret_fu_477_p2[2], ret_fu_477_p2[2], ret_fu_477_p2[2], ret_fu_477_p2[2], ret_fu_477_p2[2], ret_fu_477_p2[2], ret_fu_477_p2[2], ret_fu_477_p2[2], ret_fu_477_p2[2], ret_fu_477_p2[2], ret_fu_477_p2[2], ret_fu_477_p2[2], ret_fu_477_p2[2], ret_fu_477_p2[2], ret_fu_477_p2 };
assign sext_ln69_7_fu_384_p1 = { add_ln69_3_reg_533[4], add_ln69_3_reg_533 };
assign sext_ln69_8_fu_393_p1 = { add_ln69_4_fu_387_p2[5], add_ln69_4_fu_387_p2[5], add_ln69_4_fu_387_p2[5], add_ln69_4_fu_387_p2[5], add_ln69_4_fu_387_p2[5], add_ln69_4_fu_387_p2[5], add_ln69_4_fu_387_p2[5], add_ln69_4_fu_387_p2[5], add_ln69_4_fu_387_p2[5], add_ln69_4_fu_387_p2[5], add_ln69_4_fu_387_p2[5], add_ln69_4_fu_387_p2[5], add_ln69_4_fu_387_p2[5], add_ln69_4_fu_387_p2[5], add_ln69_4_fu_387_p2[5], add_ln69_4_fu_387_p2[5], add_ln69_4_fu_387_p2[5], add_ln69_4_fu_387_p2[5], add_ln69_4_fu_387_p2[5], add_ln69_4_fu_387_p2[5], add_ln69_4_fu_387_p2[5], add_ln69_4_fu_387_p2[5], add_ln69_4_fu_387_p2[5], add_ln69_4_fu_387_p2[5], add_ln69_4_fu_387_p2[5], add_ln69_4_fu_387_p2[5], add_ln69_4_fu_387_p2 };
assign sext_ln69_fu_215_p1 = { op_10_V_fu_205_p2[1], op_10_V_fu_205_p2[1], op_10_V_fu_205_p2[1], op_10_V_fu_205_p2[1], op_10_V_fu_205_p2[1], op_10_V_fu_205_p2[1], op_10_V_fu_205_p2[1], op_10_V_fu_205_p2 };
assign sext_ln703_fu_403_p0 = op_17;
assign sext_ln703_fu_403_p1 = { op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17 };
assign sext_ln727_fu_211_p1 = { op_8[7], op_8 };
assign trunc_ln69_fu_197_p0 = op_2;
assign trunc_ln69_fu_197_p1 = op_2[1:0];
assign trunc_ln851_1_fu_442_p0 = op_17;
assign trunc_ln851_1_fu_442_p1 = op_17[3:0];
assign trunc_ln851_fu_285_p1 = ret_V_8_fu_261_p2[19:0];
assign zext_ln1192_fu_317_p1 = { 30'h00000000, op_5, 2'h0 };
assign zext_ln1193_fu_257_p1 = { 7'h00, op_6, 20'h00000 };
assign zext_ln1346_fu_187_p1 = { 5'h00, op_3 };
assign zext_ln215_fu_474_p1 = { 1'h0, op_6 };
assign zext_ln69_fu_201_p1 = { 1'h0, op_5 };
endmodule


// Machine B:
// Processed by function `add_clk_enable_signal` in `verilog_tricks.py`.
// Processed by function `remove_reset_signal` in `verilog_tricks.py`.
module top_B (
  ap_clk,
  ap_start,
  ap_done,
  ap_idle,
  ap_ready,
  op_0,
  op_2,
  op_3,
  op_5,
  op_6,
  op_7,
  op_8,
  op_12,
  op_13,
  op_15,
  op_16,
  op_17,
  op_19,
  op_30,
  op_30_ap_vld,
clk_enable
);
input clk_enable;


input ap_clk;
wire ap_rst;
assign ap_rst = op_30_ap_vld;
input ap_start;
input [7:0] op_0;
input op_12;
input [3:0] op_13;
input [3:0] op_15;
input [1:0] op_16;
input [7:0] op_17;
input [3:0] op_19;
input [7:0] op_2;
input [3:0] op_3;
input op_5;
input [1:0] op_6;
input [31:0] op_7;
input [7:0] op_8;
output ap_done;
output ap_idle;
output ap_ready;
output [31:0] op_30;
output op_30_ap_vld;


reg [31:0] add_ln691_reg_598;
reg [31:0] add_ln69_2_reg_561;
reg [4:0] add_ln69_3_reg_556;
reg [5:0] add_ln69_4_reg_566;
reg [8:0] add_ln69_reg_499;
reg [10:0] ap_CS_fsm = 11'h001;
reg icmp_ln851_1_reg_588;
reg icmp_ln851_reg_541;
reg [1:0] op_10_V_reg_494;
reg [31:0] op_21_V_reg_509;
reg [31:0] op_27_V_reg_571;
reg [31:0] op_29_V_reg_603;
reg [8:0] ret_2_reg_504;
reg [31:0] ret_V_10_reg_551;
reg [36:0] ret_V_11_reg_576;
reg [31:0] ret_V_6_cast_reg_581;
reg [7:0] ret_V_cast_reg_524;
reg [7:0] ret_V_reg_546;
reg [2:0] ret_reg_593;
reg [19:0] trunc_ln851_reg_531;
reg [8:0] _062_;
reg [31:0] _064_;
wire [31:0] _000_;
wire [31:0] _001_;
wire [4:0] _002_;
wire [5:0] _003_;
wire [8:0] _004_;
wire [10:0] _005_;
wire _006_;
wire _007_;
wire [1:0] _008_;
wire [31:0] _009_;
wire [31:0] _010_;
wire [31:0] _011_;
wire [31:0] _012_;
wire [8:0] _013_;
wire [31:0] _014_;
wire [36:0] _015_;
wire [31:0] _016_;
wire [8:0] _017_;
wire [7:0] _018_;
wire [7:0] _019_;
wire [2:0] _020_;
wire [1:0] _021_;
wire _022_;
wire _023_;
wire _024_;
wire _025_;
wire _026_;
wire _027_;
wire _028_;
wire _029_;
wire _030_;
wire _031_;
wire _032_;
wire _033_;
wire _034_;
wire _035_;
wire _036_;
wire _037_;
wire _038_;
wire [31:0] add_ln691_fu_441_p2;
wire [31:0] add_ln69_2_fu_369_p2;
wire [4:0] add_ln69_3_fu_336_p2;
wire [5:0] add_ln69_4_fu_377_p2;
wire [8:0] add_ln69_fu_204_p2;
wire ap_CS_fsm_state1;
wire ap_CS_fsm_state10;
wire ap_CS_fsm_state11;
wire ap_CS_fsm_state2;
wire ap_CS_fsm_state3;
wire ap_CS_fsm_state4;
wire ap_CS_fsm_state5;
wire ap_CS_fsm_state6;
wire ap_CS_fsm_state7;
wire ap_CS_fsm_state8;
wire ap_CS_fsm_state9;
wire [10:0] ap_NS_fsm;
wire ap_clk;
wire ap_done;
wire ap_idle;
wire ap_ready;
wire ap_rst;
wire ap_start;
wire icmp_ln851_1_fu_426_p2;
wire icmp_ln851_fu_295_p2;
wire [21:0] lhs_fu_246_p3;
wire [7:0] op_0;
wire [1:0] op_10_V_fu_191_p2;
wire [2:0] op_11_V_fu_239_p3;
wire op_12;
wire [3:0] op_13;
wire [3:0] op_15;
wire [1:0] op_16;
wire [7:0] op_17;
wire [3:0] op_19;
wire [7:0] op_2;
wire [31:0] op_21_V_fu_226_p2;
wire [31:0] op_22_V_fu_305_p4;
wire [31:0] op_27_V_fu_386_p2;
wire [31:0] op_29_V_fu_468_p2;
wire [3:0] op_3;
wire [31:0] op_30;
wire op_30_ap_vld;
wire op_5;
wire [1:0] op_6;
wire [31:0] op_7;
wire [7:0] op_8;
wire [28:0] op_9_V_fu_232_p3;
wire p_Result_1_fu_446_p3;
wire p_Result_s_fu_342_p3;
wire [32:0] p_Val2_2_fu_289_p2;
wire [32:0] p_Val2_2_reg_536;
wire [8:0] ret_2_fu_217_p2;
wire [31:0] ret_V_10_fu_322_p2;
wire [36:0] ret_V_11_fu_406_p2;
wire [31:0] ret_V_12_fu_458_p3;
wire [28:0] ret_V_8_fu_258_p2;
wire [28:0] ret_V_8_reg_519;
wire [7:0] ret_V_9_fu_354_p3;
wire [7:0] ret_V_fu_300_p2;
wire [2:0] ret_fu_435_p2;
wire [32:0] rhs_2_fu_282_p3;
wire [35:0] rhs_5_fu_395_p3;
wire [31:0] select_ln1192_fu_314_p3;
wire [31:0] select_ln850_1_fu_453_p3;
wire [7:0] select_ln850_fu_349_p3;
wire [31:0] sext_ln1192_1_fu_474_p1;
wire [36:0] sext_ln1192_fu_402_p1;
wire [7:0] sext_ln1346_fu_210_p0;
wire [8:0] sext_ln1346_fu_210_p1;
wire [31:0] sext_ln69_1_fu_223_p1;
wire [4:0] sext_ln69_2_fu_328_p1;
wire [31:0] sext_ln69_3_fu_361_p1;
wire [5:0] sext_ln69_4_fu_365_p1;
wire [4:0] sext_ln69_5_fu_332_p1;
wire [31:0] sext_ln69_6_fu_465_p1;
wire [5:0] sext_ln69_7_fu_374_p1;
wire [31:0] sext_ln69_8_fu_383_p1;
wire [8:0] sext_ln69_fu_201_p1;
wire [7:0] sext_ln703_fu_391_p0;
wire [36:0] sext_ln703_fu_391_p1;
wire [8:0] sext_ln727_fu_197_p1;
wire [7:0] trunc_ln69_fu_183_p0;
wire [1:0] trunc_ln69_fu_183_p1;
wire [7:0] trunc_ln851_1_fu_422_p0;
wire [3:0] trunc_ln851_1_fu_422_p1;
wire [19:0] trunc_ln851_fu_274_p1;
wire [32:0] zext_ln1192_fu_278_p1;
wire [28:0] zext_ln1193_fu_254_p1;
wire [8:0] zext_ln1346_fu_213_p1;
wire [2:0] zext_ln215_fu_432_p1;
wire [1:0] zext_ln69_fu_187_p1;


assign add_ln691_fu_441_p2 = ret_V_6_cast_reg_581 + 1'h1;
assign add_ln69_2_fu_369_p2 = $signed(ret_V_10_reg_551) + $signed(ret_V_9_fu_354_p3);
assign add_ln69_3_fu_336_p2 = $signed(op_13) + $signed(op_16);
assign add_ln69_4_fu_377_p2 = $signed(add_ln69_3_reg_556) + $signed(op_15);
assign add_ln69_fu_204_p2 = $signed(op_8) + $signed(op_10_V_reg_494);
assign op_10_V_fu_191_p2 = op_2[1:0] + op_5;
assign op_21_V_fu_226_p2 = $signed(add_ln69_reg_499) + $signed(op_7);
assign op_27_V_fu_386_p2 = $signed(add_ln69_4_reg_566) + $signed(add_ln69_2_reg_561);
assign op_29_V_fu_468_p2 = $signed(ret_V_12_fu_458_p3) + $signed(ret_reg_593);
assign op_30 = $signed(op_29_V_reg_603) + $signed(op_19);
assign p_Val2_2_fu_289_p2 = { op_21_V_reg_509, 1'h0 } + { op_5, 2'h0 };
assign ret_2_fu_217_p2 = $signed(op_2) + $signed({ 1'h0, op_3 });
assign ret_V_10_fu_322_p2 = p_Val2_2_reg_536[32:1] + select_ln1192_fu_314_p3;
assign ret_V_11_fu_406_p2 = $signed({ op_27_V_reg_571, 4'h0 }) + $signed(op_17);
assign ret_V_fu_300_p2 = ret_V_cast_reg_524 + 1'h1;
assign _022_ = ap_CS_fsm[8] & icmp_ln851_1_reg_588;
assign _023_ = ap_CS_fsm[0] & _025_;
assign _024_ = ap_CS_fsm[0] & ap_start;
assign _025_ = ~ ap_start;
assign _026_ = ! trunc_ln851_reg_531;
assign _027_ = | op_17[3:0];
always @(posedge ap_clk)
trunc_ln851_reg_531 <= 20'h00000;
always @(posedge ap_clk)
ret_reg_593 <= _020_;
always @(posedge ap_clk)
_062_ <= _017_;
assign ret_V_8_reg_519[28:20] = _062_;
always @(posedge ap_clk)
ret_V_cast_reg_524 <= _018_;
always @(posedge ap_clk)
_064_ <= _012_;
assign p_Val2_2_reg_536[32:1] = _064_;
always @(posedge ap_clk)
op_29_V_reg_603 <= _011_;
always @(posedge ap_clk)
op_27_V_reg_571 <= _010_;
always @(posedge ap_clk)
ret_2_reg_504 <= _013_;
always @(posedge ap_clk)
op_21_V_reg_509 <= _009_;
always @(posedge ap_clk)
op_10_V_reg_494 <= _008_;
always @(posedge ap_clk)
ret_V_11_reg_576 <= _015_;
always @(posedge ap_clk)
ret_V_6_cast_reg_581 <= _016_;
always @(posedge ap_clk)
icmp_ln851_1_reg_588 <= _006_;
always @(posedge ap_clk)
add_ln69_reg_499 <= _004_;
always @(posedge ap_clk)
icmp_ln851_reg_541 <= _007_;
always @(posedge ap_clk)
ret_V_reg_546 <= _019_;
always @(posedge ap_clk)
ret_V_10_reg_551 <= _014_;
always @(posedge ap_clk)
add_ln69_3_reg_556 <= _002_;
always @(posedge ap_clk)
add_ln69_2_reg_561 <= _001_;
always @(posedge ap_clk)
add_ln69_4_reg_566 <= _003_;
always @(posedge ap_clk)
add_ln691_reg_598 <= _000_;
always @(posedge ap_clk)
ap_CS_fsm <= _005_;
assign _028_ = ap_CS_fsm == 3'h4;
assign _029_ = ap_CS_fsm == 2'h2;
assign _030_ = ap_CS_fsm == 1'h1;
assign op_30_ap_vld = ap_CS_fsm[10] ? 1'h1 : 1'h0;
assign ap_idle = _023_ ? 1'h1 : 1'h0;
assign _020_ = ap_CS_fsm[8] ? ret_fu_435_p2 : ret_reg_593;
assign _012_ = ap_CS_fsm[3] ? p_Val2_2_fu_289_p2[32:1] : p_Val2_2_reg_536[32:1];
assign _018_ = ap_CS_fsm[3] ? ret_V_8_fu_258_p2[27:20] : ret_V_cast_reg_524;
assign _017_ = ap_CS_fsm[3] ? ret_V_8_fu_258_p2[28:20] : ret_V_8_reg_519[28:20];
assign _011_ = ap_CS_fsm[9] ? op_29_V_fu_468_p2 : op_29_V_reg_603;
assign _010_ = ap_CS_fsm[6] ? op_27_V_fu_386_p2 : op_27_V_reg_571;
assign _009_ = ap_CS_fsm[2] ? op_21_V_fu_226_p2 : op_21_V_reg_509;
assign _013_ = ap_CS_fsm[2] ? ret_2_fu_217_p2 : ret_2_reg_504;
assign _008_ = ap_CS_fsm[0] ? op_10_V_fu_191_p2 : op_10_V_reg_494;
assign _006_ = ap_CS_fsm[7] ? icmp_ln851_1_fu_426_p2 : icmp_ln851_1_reg_588;
assign _016_ = ap_CS_fsm[7] ? ret_V_11_fu_406_p2[35:4] : ret_V_6_cast_reg_581;
assign _015_ = ap_CS_fsm[7] ? ret_V_11_fu_406_p2 : ret_V_11_reg_576;
assign _004_ = ap_CS_fsm[1] ? add_ln69_fu_204_p2 : add_ln69_reg_499;
assign _002_ = ap_CS_fsm[4] ? add_ln69_3_fu_336_p2 : add_ln69_3_reg_556;
assign _014_ = ap_CS_fsm[4] ? ret_V_10_fu_322_p2 : ret_V_10_reg_551;
assign _019_ = ap_CS_fsm[4] ? ret_V_fu_300_p2 : ret_V_reg_546;
assign _007_ = ap_CS_fsm[4] ? icmp_ln851_fu_295_p2 : icmp_ln851_reg_541;
assign _003_ = ap_CS_fsm[5] ? add_ln69_4_fu_377_p2 : add_ln69_4_reg_566;
assign _001_ = ap_CS_fsm[5] ? add_ln69_2_fu_369_p2 : add_ln69_2_reg_561;
assign _000_ = _022_ ? add_ln691_fu_441_p2 : add_ln691_reg_598;
assign _005_ = ap_rst ? 11'h001 : ap_NS_fsm;
assign _021_ = _024_ ? 2'h2 : 2'h1;
function [10:0] _109_;
input [10:0] a;
input [120:0] b;
input [10:0] s;
case (s)
11'b00000000001:
_109_ = b[10:0];
11'b00000000010:
_109_ = b[21:11];
11'b00000000100:
_109_ = b[32:22];
11'b00000001000:
_109_ = b[43:33];
11'b00000010000:
_109_ = b[54:44];
11'b00000100000:
_109_ = b[65:55];
11'b00001000000:
_109_ = b[76:66];
11'b00010000000:
_109_ = b[87:77];
11'b00100000000:
_109_ = b[98:88];
11'b01000000000:
_109_ = b[109:99];
11'b10000000000:
_109_ = b[120:110];
11'b00000000000:
_109_ = a;
default:
_109_ = 11'bx;
endcase
endfunction
assign ap_NS_fsm = _109_(11'hxxx, { 9'h000, _021_, 110'h0020080200802008020080200001 }, { _030_, _029_, _028_, _038_, _037_, _036_, _035_, _034_, _033_, _032_, _031_ });
assign _031_ = ap_CS_fsm == 11'h400;
assign _032_ = ap_CS_fsm == 10'h200;
assign _033_ = ap_CS_fsm == 9'h100;
assign _034_ = ap_CS_fsm == 8'h80;
assign _035_ = ap_CS_fsm == 7'h40;
assign _036_ = ap_CS_fsm == 6'h20;
assign _037_ = ap_CS_fsm == 5'h10;
assign _038_ = ap_CS_fsm == 4'h8;
assign ret_V_8_fu_258_p2 = { op_6, 20'h00000 } - { ret_2_reg_504, 20'h00000 };
assign ret_fu_435_p2 = 1'h0 - op_6;
assign icmp_ln851_1_fu_426_p2 = _027_ ? 1'h1 : 1'h0;
assign icmp_ln851_fu_295_p2 = _026_ ? 1'h1 : 1'h0;
assign ret_V_12_fu_458_p3 = ret_V_11_reg_576[36] ? select_ln850_1_fu_453_p3 : ret_V_6_cast_reg_581;
assign ret_V_9_fu_354_p3 = ret_V_8_reg_519[28] ? select_ln850_fu_349_p3 : ret_V_cast_reg_524;
assign select_ln1192_fu_314_p3 = op_12 ? 32'd4294967295 : 32'd0;
assign select_ln850_1_fu_453_p3 = icmp_ln851_1_reg_588 ? add_ln691_reg_598 : ret_V_6_cast_reg_581;
assign select_ln850_fu_349_p3 = icmp_ln851_reg_541 ? ret_V_cast_reg_524 : ret_V_reg_546;
assign ap_CS_fsm_state1 = ap_CS_fsm[0];
assign ap_CS_fsm_state10 = ap_CS_fsm[9];
assign ap_CS_fsm_state11 = ap_CS_fsm[10];
assign ap_CS_fsm_state2 = ap_CS_fsm[1];
assign ap_CS_fsm_state3 = ap_CS_fsm[2];
assign ap_CS_fsm_state4 = ap_CS_fsm[3];
assign ap_CS_fsm_state5 = ap_CS_fsm[4];
assign ap_CS_fsm_state6 = ap_CS_fsm[5];
assign ap_CS_fsm_state7 = ap_CS_fsm[6];
assign ap_CS_fsm_state8 = ap_CS_fsm[7];
assign ap_CS_fsm_state9 = ap_CS_fsm[8];
assign ap_done = op_30_ap_vld;
assign ap_ready = op_30_ap_vld;
assign lhs_fu_246_p3 = { op_6, 20'h00000 };
assign op_11_V_fu_239_p3 = { op_5, 2'h0 };
assign op_22_V_fu_305_p4 = p_Val2_2_reg_536[32:1];
assign op_9_V_fu_232_p3 = { ret_2_reg_504, 20'h00000 };
assign p_Result_1_fu_446_p3 = ret_V_11_reg_576[36];
assign p_Result_s_fu_342_p3 = ret_V_8_reg_519[28];
assign rhs_2_fu_282_p3 = { op_21_V_reg_509, 1'h0 };
assign rhs_5_fu_395_p3 = { op_27_V_reg_571, 4'h0 };
assign sext_ln1192_1_fu_474_p1 = { op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19 };
assign sext_ln1192_fu_402_p1 = { op_27_V_reg_571[31], op_27_V_reg_571, 4'h0 };
assign sext_ln1346_fu_210_p0 = op_2;
assign sext_ln1346_fu_210_p1 = { op_2[7], op_2 };
assign sext_ln69_1_fu_223_p1 = { add_ln69_reg_499[8], add_ln69_reg_499[8], add_ln69_reg_499[8], add_ln69_reg_499[8], add_ln69_reg_499[8], add_ln69_reg_499[8], add_ln69_reg_499[8], add_ln69_reg_499[8], add_ln69_reg_499[8], add_ln69_reg_499[8], add_ln69_reg_499[8], add_ln69_reg_499[8], add_ln69_reg_499[8], add_ln69_reg_499[8], add_ln69_reg_499[8], add_ln69_reg_499[8], add_ln69_reg_499[8], add_ln69_reg_499[8], add_ln69_reg_499[8], add_ln69_reg_499[8], add_ln69_reg_499[8], add_ln69_reg_499[8], add_ln69_reg_499[8], add_ln69_reg_499 };
assign sext_ln69_2_fu_328_p1 = { op_13[3], op_13 };
assign sext_ln69_3_fu_361_p1 = { ret_V_9_fu_354_p3[7], ret_V_9_fu_354_p3[7], ret_V_9_fu_354_p3[7], ret_V_9_fu_354_p3[7], ret_V_9_fu_354_p3[7], ret_V_9_fu_354_p3[7], ret_V_9_fu_354_p3[7], ret_V_9_fu_354_p3[7], ret_V_9_fu_354_p3[7], ret_V_9_fu_354_p3[7], ret_V_9_fu_354_p3[7], ret_V_9_fu_354_p3[7], ret_V_9_fu_354_p3[7], ret_V_9_fu_354_p3[7], ret_V_9_fu_354_p3[7], ret_V_9_fu_354_p3[7], ret_V_9_fu_354_p3[7], ret_V_9_fu_354_p3[7], ret_V_9_fu_354_p3[7], ret_V_9_fu_354_p3[7], ret_V_9_fu_354_p3[7], ret_V_9_fu_354_p3[7], ret_V_9_fu_354_p3[7], ret_V_9_fu_354_p3[7], ret_V_9_fu_354_p3 };
assign sext_ln69_4_fu_365_p1 = { op_15[3], op_15[3], op_15 };
assign sext_ln69_5_fu_332_p1 = { op_16[1], op_16[1], op_16[1], op_16 };
assign sext_ln69_6_fu_465_p1 = { ret_reg_593[2], ret_reg_593[2], ret_reg_593[2], ret_reg_593[2], ret_reg_593[2], ret_reg_593[2], ret_reg_593[2], ret_reg_593[2], ret_reg_593[2], ret_reg_593[2], ret_reg_593[2], ret_reg_593[2], ret_reg_593[2], ret_reg_593[2], ret_reg_593[2], ret_reg_593[2], ret_reg_593[2], ret_reg_593[2], ret_reg_593[2], ret_reg_593[2], ret_reg_593[2], ret_reg_593[2], ret_reg_593[2], ret_reg_593[2], ret_reg_593[2], ret_reg_593[2], ret_reg_593[2], ret_reg_593[2], ret_reg_593[2], ret_reg_593 };
assign sext_ln69_7_fu_374_p1 = { add_ln69_3_reg_556[4], add_ln69_3_reg_556 };
assign sext_ln69_8_fu_383_p1 = { add_ln69_4_reg_566[5], add_ln69_4_reg_566[5], add_ln69_4_reg_566[5], add_ln69_4_reg_566[5], add_ln69_4_reg_566[5], add_ln69_4_reg_566[5], add_ln69_4_reg_566[5], add_ln69_4_reg_566[5], add_ln69_4_reg_566[5], add_ln69_4_reg_566[5], add_ln69_4_reg_566[5], add_ln69_4_reg_566[5], add_ln69_4_reg_566[5], add_ln69_4_reg_566[5], add_ln69_4_reg_566[5], add_ln69_4_reg_566[5], add_ln69_4_reg_566[5], add_ln69_4_reg_566[5], add_ln69_4_reg_566[5], add_ln69_4_reg_566[5], add_ln69_4_reg_566[5], add_ln69_4_reg_566[5], add_ln69_4_reg_566[5], add_ln69_4_reg_566[5], add_ln69_4_reg_566[5], add_ln69_4_reg_566[5], add_ln69_4_reg_566 };
assign sext_ln69_fu_201_p1 = { op_10_V_reg_494[1], op_10_V_reg_494[1], op_10_V_reg_494[1], op_10_V_reg_494[1], op_10_V_reg_494[1], op_10_V_reg_494[1], op_10_V_reg_494[1], op_10_V_reg_494 };
assign sext_ln703_fu_391_p0 = op_17;
assign sext_ln703_fu_391_p1 = { op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17 };
assign sext_ln727_fu_197_p1 = { op_8[7], op_8 };
assign trunc_ln69_fu_183_p0 = op_2;
assign trunc_ln69_fu_183_p1 = op_2[1:0];
assign trunc_ln851_1_fu_422_p0 = op_17;
assign trunc_ln851_1_fu_422_p1 = op_17[3:0];
assign trunc_ln851_fu_274_p1 = ret_V_8_fu_258_p2[19:0];
assign zext_ln1192_fu_278_p1 = { 30'h00000000, op_5, 2'h0 };
assign zext_ln1193_fu_254_p1 = { 7'h00, op_6, 20'h00000 };
assign zext_ln1346_fu_213_p1 = { 5'h00, op_3 };
assign zext_ln215_fu_432_p1 = { 1'h0, op_6 };
assign zext_ln69_fu_187_p1 = { 1'h0, op_5 };
endmodule


// Product machine:
module top_A_times_top_B (ap_start, op_0, op_12, op_13, op_15, op_16, op_17, op_19, op_2, op_3, op_5, op_6, op_7, op_8, ap_clk, unsafe_signal);
input ap_start;
input [7:0] op_0;
input op_12;
input [3:0] op_13;
input [3:0] op_15;
input [1:0] op_16;
input [7:0] op_17;
input [3:0] op_19;
input [7:0] op_2;
input [3:0] op_3;
input op_5;
input [1:0] op_6;
input [31:0] op_7;
input [7:0] op_8;
input ap_clk;
output unsafe_signal;
reg _setup;
initial _setup = 1'b0;
always @ (posedge ap_clk) _setup <= 1'b1;
reg ap_start_internal;
always @ (posedge ap_clk) if (!_setup) ap_start_internal <= ap_start;
reg [7:0] op_0_internal;
always @ (posedge ap_clk) if (!_setup) op_0_internal <= op_0;
reg op_12_internal;
always @ (posedge ap_clk) if (!_setup) op_12_internal <= op_12;
reg [3:0] op_13_internal;
always @ (posedge ap_clk) if (!_setup) op_13_internal <= op_13;
reg [3:0] op_15_internal;
always @ (posedge ap_clk) if (!_setup) op_15_internal <= op_15;
reg [1:0] op_16_internal;
always @ (posedge ap_clk) if (!_setup) op_16_internal <= op_16;
reg [7:0] op_17_internal;
always @ (posedge ap_clk) if (!_setup) op_17_internal <= op_17;
reg [3:0] op_19_internal;
always @ (posedge ap_clk) if (!_setup) op_19_internal <= op_19;
reg [7:0] op_2_internal;
always @ (posedge ap_clk) if (!_setup) op_2_internal <= op_2;
reg [3:0] op_3_internal;
always @ (posedge ap_clk) if (!_setup) op_3_internal <= op_3;
reg op_5_internal;
always @ (posedge ap_clk) if (!_setup) op_5_internal <= op_5;
reg [1:0] op_6_internal;
always @ (posedge ap_clk) if (!_setup) op_6_internal <= op_6;
reg [31:0] op_7_internal;
always @ (posedge ap_clk) if (!_setup) op_7_internal <= op_7;
reg [7:0] op_8_internal;
always @ (posedge ap_clk) if (!_setup) op_8_internal <= op_8;
wire ap_done_A;
wire ap_done_B;
wire ap_done_eq;
assign ap_done_eq = ap_done_A == ap_done_B;
wire ap_idle_A;
wire ap_idle_B;
wire ap_idle_eq;
assign ap_idle_eq = ap_idle_A == ap_idle_B;
wire ap_ready_A;
wire ap_ready_B;
wire ap_ready_eq;
assign ap_ready_eq = ap_ready_A == ap_ready_B;
wire [31:0] op_30_A;
wire [31:0] op_30_B;
wire op_30_eq;
assign op_30_eq = op_30_A == op_30_B;
wire op_30_ap_vld_A;
wire op_30_ap_vld_B;
wire clk_enable_A;
wire clk_enable_B;
assign clk_enable_A = _setup & (~op_30_ap_vld_A | op_30_ap_vld_B);
assign clk_enable_B = _setup;
wire divergent;
assign divergent = ~(ap_done_eq & ap_idle_eq & ap_ready_eq & op_30_eq);
assign unsafe_signal = op_30_ap_vld_A & op_30_ap_vld_B & divergent;
top_A instance_A (
    .ap_clk(ap_clk),
    .clk_enable(clk_enable_A),
    .ap_start(ap_start_internal),
    .op_0(op_0_internal),
    .op_12(op_12_internal),
    .op_13(op_13_internal),
    .op_15(op_15_internal),
    .op_16(op_16_internal),
    .op_17(op_17_internal),
    .op_19(op_19_internal),
    .op_2(op_2_internal),
    .op_3(op_3_internal),
    .op_5(op_5_internal),
    .op_6(op_6_internal),
    .op_7(op_7_internal),
    .op_8(op_8_internal),
    .ap_done(ap_done_A),
    .ap_idle(ap_idle_A),
    .ap_ready(ap_ready_A),
    .op_30(op_30_A),
    .op_30_ap_vld(op_30_ap_vld_A)
);
top_B instance_B (
    .ap_clk(ap_clk),
    .clk_enable(clk_enable_B),
    .ap_start(ap_start_internal),
    .op_0(op_0_internal),
    .op_12(op_12_internal),
    .op_13(op_13_internal),
    .op_15(op_15_internal),
    .op_16(op_16_internal),
    .op_17(op_17_internal),
    .op_19(op_19_internal),
    .op_2(op_2_internal),
    .op_3(op_3_internal),
    .op_5(op_5_internal),
    .op_6(op_6_internal),
    .op_7(op_7_internal),
    .op_8(op_8_internal),
    .ap_done(ap_done_B),
    .ap_idle(ap_idle_B),
    .ap_ready(ap_ready_B),
    .op_30(op_30_B),
    .op_30_ap_vld(op_30_ap_vld_B)
);
endmodule
