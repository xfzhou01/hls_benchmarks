// Processed by function `construct_kairos` in `verilog_tricks.py`.
// Machine A:
// Processed by function `add_clk_enable_signal` in `verilog_tricks.py`.
// Processed by function `remove_reset_signal` in `verilog_tricks.py`.
module top_A (
  ap_clk,
  ap_start,
  ap_done,
  ap_idle,
  ap_ready,
  op_0,
  op_2,
  op_3,
  op_5,
  op_8,
  op_10,
  op_11,
  op_14,
  op_16,
  op_18,
  op_19,
  op_30,
  op_30_ap_vld,
clk_enable
);
input clk_enable;


input ap_clk;
wire ap_rst;
assign ap_rst = op_30_ap_vld;
input ap_start;
input [3:0] op_0;
input [7:0] op_10;
input [7:0] op_11;
input [3:0] op_14;
input [7:0] op_16;
input [31:0] op_18;
input op_19;
input [3:0] op_2;
input [31:0] op_3;
input [15:0] op_5;
input [3:0] op_8;
output ap_done;
output ap_idle;
output ap_ready;
output [31:0] op_30;
output op_30_ap_vld;


reg [31:0] add_ln691_4_reg_883;
reg [4:0] add_ln69_1_reg_792;
reg [11:0] ap_CS_fsm = 12'h001;
reg icmp_ln851_1_reg_824;
reg icmp_ln851_2_reg_878;
reg [31:0] op_13_V_reg_797;
reg [1:0] op_15_V_reg_787;
reg [24:0] op_23_V_reg_802;
reg [31:0] op_28_V_reg_861;
reg [1:0] ret_V_15_reg_751;
reg [32:0] ret_V_16_reg_756;
reg [24:0] ret_V_17_reg_782;
reg [31:0] ret_V_19_cast_reg_849;
reg [55:0] ret_V_19_reg_812;
reg [31:0] ret_V_20_reg_829;
reg [31:0] ret_V_21_cast_reg_871;
reg [31:0] ret_V_22_reg_834;
reg [33:0] ret_V_23_reg_844;
reg [31:0] ret_V_24_reg_856;
reg [38:0] ret_V_25_reg_866;
reg [31:0] ret_V_8_cast_reg_817;
reg [3:0] ret_reg_776;
reg [23:0] tmp_1_reg_761;
reg [8:0] trunc_ln851_1_reg_766;
reg [22:0] trunc_ln851_2_reg_807;
wire [31:0] _000_;
wire [4:0] _001_;
wire [11:0] _002_;
wire _003_;
wire _004_;
wire [31:0] _005_;
wire [1:0] _006_;
wire [24:0] _007_;
wire [31:0] _008_;
wire [1:0] _009_;
wire [32:0] _010_;
wire [24:0] _011_;
wire [31:0] _012_;
wire [55:0] _013_;
wire [31:0] _014_;
wire [31:0] _015_;
wire [31:0] _016_;
wire [33:0] _017_;
wire [31:0] _018_;
wire [38:0] _019_;
wire [31:0] _020_;
wire [3:0] _021_;
wire [23:0] _022_;
wire [8:0] _023_;
wire [22:0] _024_;
wire [1:0] _025_;
wire _026_;
wire _027_;
wire _028_;
wire _029_;
wire _030_;
wire _031_;
wire _032_;
wire _033_;
wire _034_;
wire _035_;
wire _036_;
wire _037_;
wire _038_;
wire _039_;
wire _040_;
wire _041_;
wire _042_;
wire _043_;
wire _044_;
wire [24:0] add_ln691_1_fu_343_p2;
wire [31:0] add_ln691_2_fu_553_p2;
wire [31:0] add_ln691_3_fu_630_p2;
wire [31:0] add_ln691_4_fu_712_p2;
wire [1:0] add_ln691_fu_255_p2;
wire [4:0] add_ln69_1_fu_397_p2;
wire [24:0] add_ln69_fu_493_p2;
wire ap_CS_fsm_state1;
wire ap_CS_fsm_state10;
wire ap_CS_fsm_state11;
wire ap_CS_fsm_state12;
wire ap_CS_fsm_state2;
wire ap_CS_fsm_state3;
wire ap_CS_fsm_state4;
wire ap_CS_fsm_state5;
wire ap_CS_fsm_state6;
wire ap_CS_fsm_state7;
wire ap_CS_fsm_state8;
wire ap_CS_fsm_state9;
wire [11:0] ap_NS_fsm;
wire ap_clk;
wire ap_done;
wire ap_idle;
wire ap_ready;
wire ap_rst;
wire ap_start;
wire [15:0] empty_16_fu_301_p0;
wire [9:0] empty_16_fu_301_p1;
wire [2:0] empty_fu_223_p1;
wire icmp_ln851_1_fu_541_p2;
wire icmp_ln851_2_fu_706_p2;
wire icmp_ln851_fu_338_p2;
wire [20:0] lhs_V_fu_369_p3;
wire [1:0] \mul_2s_2s_4_1_1_U1.din0 ;
wire [1:0] \mul_2s_2s_4_1_1_U1.din1 ;
wire [3:0] \mul_2s_2s_4_1_1_U1.dout ;
wire [1:0] \mul_2s_2s_4_1_1_U1.top_mul_2s_2s_4_1_1_Multiplier_0_U.a ;
wire [1:0] \mul_2s_2s_4_1_1_U1.top_mul_2s_2s_4_1_1_Multiplier_0_U.b ;
wire [3:0] \mul_2s_2s_4_1_1_U1.top_mul_2s_2s_4_1_1_Multiplier_0_U.p ;
wire [3:0] op_0;
wire [7:0] op_10;
wire [7:0] op_11;
wire [20:0] op_12_V_fu_311_p3;
wire [31:0] op_13_V_fu_481_p3;
wire [3:0] op_14;
wire [7:0] op_16;
wire op_17_V_fu_656_p2;
wire [31:0] op_18;
wire op_19;
wire [3:0] op_2;
wire [24:0] op_23_V_fu_501_p2;
wire [31:0] op_28_V_fu_666_p2;
wire [31:0] op_3;
wire [31:0] op_30;
wire op_30_ap_vld;
wire [15:0] op_5;
wire [3:0] op_8;
wire overflow_fu_461_p2;
wire p_Result_1_fu_331_p3;
wire p_Result_4_fu_546_p3;
wire p_Result_5_fu_620_p3;
wire p_Result_6_fu_717_p3;
wire p_Result_7_fu_427_p3;
wire p_Result_8_fu_447_p3;
wire p_Result_s_fu_243_p3;
wire [31:0] p_Val2_3_fu_439_p3;
wire [9:0] r_fu_305_p2;
wire [2:0] ret_V_14_fu_227_p2;
wire [1:0] ret_V_15_fu_269_p3;
wire [32:0] ret_V_16_fu_281_p2;
wire [24:0] ret_V_17_fu_357_p3;
wire [17:0] ret_V_18_fu_421_p2;
wire [55:0] ret_V_19_fu_525_p2;
wire [31:0] ret_V_20_fu_564_p3;
wire [31:0] ret_V_21_fu_575_p2;
wire [31:0] ret_V_22_fu_583_p2;
wire [33:0] ret_V_23_fu_604_p2;
wire [31:0] ret_V_24_fu_642_p3;
wire [38:0] ret_V_25_fu_686_p2;
wire [31:0] ret_V_26_fu_729_p3;
wire [1:0] ret_V_cast_fu_233_p4;
wire [20:0] ret_V_fu_377_p2;
wire [1:0] ret_fu_322_p0;
wire [1:0] ret_fu_322_p1;
wire [3:0] ret_fu_322_p2;
wire [11:0] rhs_1_fu_406_p3;
wire [32:0] rhs_7_fu_593_p3;
wire [37:0] rhs_9_fu_675_p3;
wire [31:0] select_ln384_fu_473_p3;
wire [31:0] select_ln69_fu_736_p3;
wire [24:0] select_ln850_1_fu_349_p3;
wire [31:0] select_ln850_2_fu_558_p3;
wire [31:0] select_ln850_3_fu_635_p3;
wire [31:0] select_ln850_4_fu_724_p3;
wire [1:0] select_ln850_fu_261_p3;
wire [55:0] sext_ln1192_1_fu_521_p1;
wire [31:0] sext_ln1192_2_fu_571_p1;
wire [31:0] sext_ln1192_3_fu_580_p1;
wire [33:0] sext_ln1192_4_fu_600_p1;
wire [38:0] sext_ln1192_5_fu_682_p1;
wire [15:0] sext_ln1192_6_fu_413_p1;
wire [32:0] sext_ln1192_fu_277_p1;
wire [3:0] sext_ln1345_fu_319_p1;
wire [24:0] sext_ln69_1_fu_489_p1;
wire [24:0] sext_ln69_3_fu_498_p1;
wire [4:0] sext_ln69_fu_393_p1;
wire [55:0] sext_ln703_1_fu_511_p1;
wire [7:0] sext_ln703_2_fu_589_p0;
wire [33:0] sext_ln703_2_fu_589_p1;
wire [31:0] sext_ln703_3_fu_671_p0;
wire [38:0] sext_ln703_3_fu_671_p1;
wire [15:0] sext_ln703_fu_403_p0;
wire [17:0] sext_ln703_fu_403_p1;
wire [24:0] sext_ln850_fu_328_p1;
wire [47:0] tmp_fu_514_p3;
wire trunc_ln213_1_fu_652_p1;
wire trunc_ln213_fu_649_p1;
wire [1:0] trunc_ln728_1_fu_365_p1;
wire [16:0] trunc_ln728_fu_435_p1;
wire [8:0] trunc_ln851_1_fu_297_p1;
wire [22:0] trunc_ln851_2_fu_507_p1;
wire [7:0] trunc_ln851_3_fu_627_p0;
wire trunc_ln851_3_fu_627_p1;
wire [31:0] trunc_ln851_4_fu_702_p0;
wire [5:0] trunc_ln851_4_fu_702_p1;
wire trunc_ln851_fu_251_p1;
wire xor_ln340_fu_467_p2;
wire xor_ln785_fu_455_p2;
wire [17:0] zext_ln1192_fu_417_p1;
wire [31:0] zext_ln69_fu_662_p1;


assign add_ln691_1_fu_343_p2 = $signed(tmp_1_reg_761) + $signed(2'h1);
assign add_ln691_2_fu_553_p2 = ret_V_8_cast_reg_817 + 1'h1;
assign add_ln691_3_fu_630_p2 = ret_V_19_cast_reg_849 + 1'h1;
assign add_ln691_4_fu_712_p2 = ret_V_21_cast_reg_871 + 1'h1;
assign add_ln691_fu_255_p2 = { op_2[2], 1'h1 } + 1'h1;
assign add_ln69_1_fu_397_p2 = $signed(op_8) + $signed(2'h1);
assign add_ln69_fu_493_p2 = $signed(ret_V_17_reg_782) + $signed(op_11);
assign op_23_V_fu_501_p2 = $signed(add_ln69_1_reg_792) + $signed(add_ln69_fu_493_p2);
assign op_28_V_fu_666_p2 = ret_V_24_reg_856 + op_17_V_fu_656_p2;
assign op_30 = ret_V_26_fu_729_p3 + select_ln69_fu_736_p3;
assign ret_V_16_fu_281_p2 = $signed(op_3) + $signed(11'h200);
assign ret_V_18_fu_421_p2 = $signed({ 1'h0, ret_reg_776[3], ret_reg_776[3], ret_reg_776[3], ret_reg_776[3], ret_reg_776, 8'h00 }) + $signed(op_5);
assign { ret_V_19_fu_525_p2[55], ret_V_19_fu_525_p2[47:0] } = $signed({ op_23_V_reg_802, 23'h000000 }) + $signed(op_13_V_reg_797);
assign ret_V_21_fu_575_p2 = $signed(ret_V_20_reg_829) + $signed(op_14);
assign ret_V_22_fu_583_p2 = $signed(ret_V_21_fu_575_p2) + $signed(op_15_V_reg_787);
assign ret_V_23_fu_604_p2 = $signed({ ret_V_22_reg_834, 1'h0 }) + $signed(op_16);
assign ret_V_25_fu_686_p2 = $signed({ op_28_V_reg_861, 6'h00 }) + $signed(op_18);
assign _026_ = ap_CS_fsm[10] & icmp_ln851_2_reg_878;
assign _027_ = ap_CS_fsm[0] & _029_;
assign _028_ = ap_CS_fsm[0] & ap_start;
assign overflow_fu_461_p2 = xor_ln785_fu_455_p2 & ret_V_18_fu_421_p2[16];
assign ret_V_fu_377_p2 = { op_12_V_fu_311_p3[20:19], op_5[7:0], 11'h000 } & { ret_fu_322_p2[1:0], 19'h00000 };
assign xor_ln785_fu_455_p2 = ~ ret_V_18_fu_421_p2[17];
assign op_12_V_fu_311_p3[20:19] = ~ op_5[9:8];
assign _029_ = ~ ap_start;
assign \mul_2s_2s_4_1_1_U1.top_mul_2s_2s_4_1_1_Multiplier_0_U.p  = $signed(\mul_2s_2s_4_1_1_U1.top_mul_2s_2s_4_1_1_Multiplier_0_U.a ) * $signed(\mul_2s_2s_4_1_1_U1.top_mul_2s_2s_4_1_1_Multiplier_0_U.b );
assign _030_ = | trunc_ln851_2_reg_807;
assign _031_ = | op_18[5:0];
assign _032_ = | trunc_ln851_1_reg_766;
always @(posedge ap_clk)
ret_V_24_reg_856 <= _018_;
always @(posedge ap_clk)
ret_V_22_reg_834 <= _016_;
always @(posedge ap_clk)
ret_V_20_reg_829 <= _014_;
always @(posedge ap_clk)
ret_V_23_reg_844 <= _017_;
always @(posedge ap_clk)
ret_V_19_cast_reg_849 <= _012_;
always @(posedge ap_clk)
ret_V_15_reg_751 <= _009_;
always @(posedge ap_clk)
ret_V_16_reg_756 <= _010_;
always @(posedge ap_clk)
tmp_1_reg_761 <= _022_;
always @(posedge ap_clk)
trunc_ln851_1_reg_766 <= _023_;
always @(posedge ap_clk)
op_28_V_reg_861 <= _008_;
always @(posedge ap_clk)
op_13_V_reg_797 <= _005_;
always @(posedge ap_clk)
op_23_V_reg_802 <= _007_;
always @(posedge ap_clk)
trunc_ln851_2_reg_807 <= _024_;
always @(posedge ap_clk)
ret_V_25_reg_866 <= _019_;
always @(posedge ap_clk)
ret_V_21_cast_reg_871 <= _015_;
always @(posedge ap_clk)
icmp_ln851_2_reg_878 <= _004_;
always @(posedge ap_clk)
ret_V_19_reg_812 <= _013_;
always @(posedge ap_clk)
ret_V_8_cast_reg_817 <= _020_;
always @(posedge ap_clk)
icmp_ln851_1_reg_824 <= _003_;
always @(posedge ap_clk)
ret_reg_776 <= _021_;
always @(posedge ap_clk)
ret_V_17_reg_782 <= _011_;
always @(posedge ap_clk)
op_15_V_reg_787 <= _006_;
always @(posedge ap_clk)
add_ln69_1_reg_792 <= _001_;
always @(posedge ap_clk)
add_ln691_4_reg_883 <= _000_;
always @(posedge ap_clk)
ap_CS_fsm <= _002_;
assign _025_ = _028_ ? 2'h2 : 2'h1;
assign _033_ = ap_CS_fsm == 1'h1;
function [11:0] _101_;
input [11:0] a;
input [143:0] b;
input [11:0] s;
case (s)
12'b000000000001:
_101_ = b[11:0];
12'b000000000010:
_101_ = b[23:12];
12'b000000000100:
_101_ = b[35:24];
12'b000000001000:
_101_ = b[47:36];
12'b000000010000:
_101_ = b[59:48];
12'b000000100000:
_101_ = b[71:60];
12'b000001000000:
_101_ = b[83:72];
12'b000010000000:
_101_ = b[95:84];
12'b000100000000:
_101_ = b[107:96];
12'b001000000000:
_101_ = b[119:108];
12'b010000000000:
_101_ = b[131:120];
12'b100000000000:
_101_ = b[143:132];
12'b000000000000:
_101_ = a;
default:
_101_ = 12'bx;
endcase
endfunction
assign ap_NS_fsm = _101_(12'hxxx, { 10'h000, _025_, 132'h004008010020040080100200400800001 }, { _033_, _044_, _043_, _042_, _041_, _040_, _039_, _038_, _037_, _036_, _035_, _034_ });
assign _034_ = ap_CS_fsm == 12'h800;
assign _035_ = ap_CS_fsm == 11'h400;
assign _036_ = ap_CS_fsm == 10'h200;
assign _037_ = ap_CS_fsm == 9'h100;
assign _038_ = ap_CS_fsm == 8'h80;
assign _039_ = ap_CS_fsm == 7'h40;
assign _040_ = ap_CS_fsm == 6'h20;
assign _041_ = ap_CS_fsm == 5'h10;
assign _042_ = ap_CS_fsm == 4'h8;
assign _043_ = ap_CS_fsm == 3'h4;
assign _044_ = ap_CS_fsm == 2'h2;
assign op_30_ap_vld = ap_CS_fsm[11] ? 1'h1 : 1'h0;
assign ap_idle = _027_ ? 1'h1 : 1'h0;
assign _018_ = ap_CS_fsm[7] ? ret_V_24_fu_642_p3 : ret_V_24_reg_856;
assign _016_ = ap_CS_fsm[5] ? ret_V_22_fu_583_p2 : ret_V_22_reg_834;
assign _014_ = ap_CS_fsm[4] ? ret_V_20_fu_564_p3 : ret_V_20_reg_829;
assign _012_ = ap_CS_fsm[6] ? ret_V_23_fu_604_p2[32:1] : ret_V_19_cast_reg_849;
assign _017_ = ap_CS_fsm[6] ? ret_V_23_fu_604_p2 : ret_V_23_reg_844;
assign _023_ = ap_CS_fsm[0] ? ret_V_16_fu_281_p2[8:0] : trunc_ln851_1_reg_766;
assign _022_ = ap_CS_fsm[0] ? ret_V_16_fu_281_p2[32:9] : tmp_1_reg_761;
assign _010_ = ap_CS_fsm[0] ? ret_V_16_fu_281_p2 : ret_V_16_reg_756;
assign _009_ = ap_CS_fsm[0] ? ret_V_15_fu_269_p3 : ret_V_15_reg_751;
assign _008_ = ap_CS_fsm[8] ? op_28_V_fu_666_p2 : op_28_V_reg_861;
assign _024_ = ap_CS_fsm[2] ? op_13_V_fu_481_p3[22:0] : trunc_ln851_2_reg_807;
assign _007_ = ap_CS_fsm[2] ? op_23_V_fu_501_p2 : op_23_V_reg_802;
assign _005_ = ap_CS_fsm[2] ? op_13_V_fu_481_p3 : op_13_V_reg_797;
assign _004_ = ap_CS_fsm[9] ? icmp_ln851_2_fu_706_p2 : icmp_ln851_2_reg_878;
assign _015_ = ap_CS_fsm[9] ? ret_V_25_fu_686_p2[37:6] : ret_V_21_cast_reg_871;
assign _019_ = ap_CS_fsm[9] ? ret_V_25_fu_686_p2 : ret_V_25_reg_866;
assign _003_ = ap_CS_fsm[3] ? icmp_ln851_1_fu_541_p2 : icmp_ln851_1_reg_824;
assign _020_ = ap_CS_fsm[3] ? { ret_V_19_fu_525_p2[55], ret_V_19_fu_525_p2[55], ret_V_19_fu_525_p2[55], ret_V_19_fu_525_p2[55], ret_V_19_fu_525_p2[55], ret_V_19_fu_525_p2[55], ret_V_19_fu_525_p2[55], ret_V_19_fu_525_p2[47:23] } : ret_V_8_cast_reg_817;
assign _013_ = ap_CS_fsm[3] ? { ret_V_19_fu_525_p2[55], ret_V_19_fu_525_p2[55], ret_V_19_fu_525_p2[55], ret_V_19_fu_525_p2[55], ret_V_19_fu_525_p2[55], ret_V_19_fu_525_p2[55], ret_V_19_fu_525_p2[55], ret_V_19_fu_525_p2[55], ret_V_19_fu_525_p2[47:0] } : ret_V_19_reg_812;
assign _001_ = ap_CS_fsm[1] ? add_ln69_1_fu_397_p2 : add_ln69_1_reg_792;
assign _006_ = ap_CS_fsm[1] ? ret_V_fu_377_p2[20:19] : op_15_V_reg_787;
assign _011_ = ap_CS_fsm[1] ? ret_V_17_fu_357_p3 : ret_V_17_reg_782;
assign _021_ = ap_CS_fsm[1] ? ret_fu_322_p2 : ret_reg_776;
assign _000_ = _026_ ? add_ln691_4_fu_712_p2 : add_ln691_4_reg_883;
assign _002_ = ap_rst ? 12'h001 : ap_NS_fsm;
assign icmp_ln851_1_fu_541_p2 = _030_ ? 1'h1 : 1'h0;
assign icmp_ln851_2_fu_706_p2 = _031_ ? 1'h1 : 1'h0;
assign icmp_ln851_fu_338_p2 = _032_ ? 1'h1 : 1'h0;
assign op_13_V_fu_481_p3 = xor_ln340_fu_467_p2 ? select_ln384_fu_473_p3 : { ret_V_18_fu_421_p2[16:0], 15'h0000 };
assign ret_V_15_fu_269_p3 = op_2[3] ? select_ln850_fu_261_p3 : { op_2[2], 1'h1 };
assign ret_V_17_fu_357_p3 = ret_V_16_reg_756[32] ? select_ln850_1_fu_349_p3 : { tmp_1_reg_761[23], tmp_1_reg_761 };
assign ret_V_20_fu_564_p3 = ret_V_19_reg_812[55] ? select_ln850_2_fu_558_p3 : ret_V_8_cast_reg_817;
assign ret_V_24_fu_642_p3 = ret_V_23_reg_844[33] ? select_ln850_3_fu_635_p3 : ret_V_19_cast_reg_849;
assign ret_V_26_fu_729_p3 = ret_V_25_reg_866[38] ? select_ln850_4_fu_724_p3 : ret_V_21_cast_reg_871;
assign select_ln384_fu_473_p3 = overflow_fu_461_p2 ? 32'd2147483647 : 32'd2147483648;
assign select_ln69_fu_736_p3 = op_19 ? 32'd4294967295 : 32'd0;
assign select_ln850_1_fu_349_p3 = icmp_ln851_fu_338_p2 ? add_ln691_1_fu_343_p2 : { tmp_1_reg_761[23], tmp_1_reg_761 };
assign select_ln850_2_fu_558_p3 = icmp_ln851_1_reg_824 ? add_ln691_2_fu_553_p2 : ret_V_8_cast_reg_817;
assign select_ln850_3_fu_635_p3 = op_16[0] ? add_ln691_3_fu_630_p2 : ret_V_19_cast_reg_849;
assign select_ln850_4_fu_724_p3 = icmp_ln851_2_reg_878 ? add_ln691_4_reg_883 : ret_V_21_cast_reg_871;
assign select_ln850_fu_261_p3 = op_2[0] ? add_ln691_fu_255_p2 : { op_2[2], 1'h1 };
assign op_17_V_fu_656_p2 = ret_reg_776[0] ^ op_10[0];
assign xor_ln340_fu_467_p2 = ret_V_18_fu_421_p2[16] ^ ret_V_18_fu_421_p2[17];
assign ap_CS_fsm_state1 = ap_CS_fsm[0];
assign ap_CS_fsm_state10 = ap_CS_fsm[9];
assign ap_CS_fsm_state11 = ap_CS_fsm[10];
assign ap_CS_fsm_state12 = ap_CS_fsm[11];
assign ap_CS_fsm_state2 = ap_CS_fsm[1];
assign ap_CS_fsm_state3 = ap_CS_fsm[2];
assign ap_CS_fsm_state4 = ap_CS_fsm[3];
assign ap_CS_fsm_state5 = ap_CS_fsm[4];
assign ap_CS_fsm_state6 = ap_CS_fsm[5];
assign ap_CS_fsm_state7 = ap_CS_fsm[6];
assign ap_CS_fsm_state8 = ap_CS_fsm[7];
assign ap_CS_fsm_state9 = ap_CS_fsm[8];
assign ap_done = op_30_ap_vld;
assign ap_ready = op_30_ap_vld;
assign empty_16_fu_301_p0 = op_5;
assign empty_16_fu_301_p1 = op_5[9:0];
assign empty_fu_223_p1 = op_2[2:0];
assign lhs_V_fu_369_p3 = { ret_fu_322_p2[1:0], 19'h00000 };
assign op_12_V_fu_311_p3[18:0] = { op_5[7:0], 11'h000 };
assign p_Result_1_fu_331_p3 = ret_V_16_reg_756[32];
assign p_Result_4_fu_546_p3 = ret_V_19_reg_812[55];
assign p_Result_5_fu_620_p3 = ret_V_23_reg_844[33];
assign p_Result_6_fu_717_p3 = ret_V_25_reg_866[38];
assign p_Result_7_fu_427_p3 = ret_V_18_fu_421_p2[17];
assign p_Result_8_fu_447_p3 = ret_V_18_fu_421_p2[16];
assign p_Result_s_fu_243_p3 = op_2[3];
assign p_Val2_3_fu_439_p3 = { ret_V_18_fu_421_p2[16:0], 15'h0000 };
assign r_fu_305_p2 = { op_12_V_fu_311_p3[20:19], op_5[7:0] };
assign ret_V_14_fu_227_p2 = { op_2[2], 1'h1, op_2[0] };
assign ret_V_19_fu_525_p2[54:48] = { ret_V_19_fu_525_p2[55], ret_V_19_fu_525_p2[55], ret_V_19_fu_525_p2[55], ret_V_19_fu_525_p2[55], ret_V_19_fu_525_p2[55], ret_V_19_fu_525_p2[55], ret_V_19_fu_525_p2[55] };
assign ret_V_cast_fu_233_p4 = { op_2[2], 1'h1 };
assign ret_fu_322_p0 = ret_V_15_reg_751;
assign ret_fu_322_p1 = ret_V_15_reg_751;
assign rhs_1_fu_406_p3 = { ret_reg_776, 8'h00 };
assign rhs_7_fu_593_p3 = { ret_V_22_reg_834, 1'h0 };
assign rhs_9_fu_675_p3 = { op_28_V_reg_861, 6'h00 };
assign sext_ln1192_1_fu_521_p1 = { op_23_V_reg_802[24], op_23_V_reg_802[24], op_23_V_reg_802[24], op_23_V_reg_802[24], op_23_V_reg_802[24], op_23_V_reg_802[24], op_23_V_reg_802[24], op_23_V_reg_802[24], op_23_V_reg_802, 23'h000000 };
assign sext_ln1192_2_fu_571_p1 = { op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14 };
assign sext_ln1192_3_fu_580_p1 = { op_15_V_reg_787[1], op_15_V_reg_787[1], op_15_V_reg_787[1], op_15_V_reg_787[1], op_15_V_reg_787[1], op_15_V_reg_787[1], op_15_V_reg_787[1], op_15_V_reg_787[1], op_15_V_reg_787[1], op_15_V_reg_787[1], op_15_V_reg_787[1], op_15_V_reg_787[1], op_15_V_reg_787[1], op_15_V_reg_787[1], op_15_V_reg_787[1], op_15_V_reg_787[1], op_15_V_reg_787[1], op_15_V_reg_787[1], op_15_V_reg_787[1], op_15_V_reg_787[1], op_15_V_reg_787[1], op_15_V_reg_787[1], op_15_V_reg_787[1], op_15_V_reg_787[1], op_15_V_reg_787[1], op_15_V_reg_787[1], op_15_V_reg_787[1], op_15_V_reg_787[1], op_15_V_reg_787[1], op_15_V_reg_787[1], op_15_V_reg_787 };
assign sext_ln1192_4_fu_600_p1 = { ret_V_22_reg_834[31], ret_V_22_reg_834, 1'h0 };
assign sext_ln1192_5_fu_682_p1 = { op_28_V_reg_861[31], op_28_V_reg_861, 6'h00 };
assign sext_ln1192_6_fu_413_p1 = { ret_reg_776[3], ret_reg_776[3], ret_reg_776[3], ret_reg_776[3], ret_reg_776, 8'h00 };
assign sext_ln1192_fu_277_p1 = { op_3[31], op_3 };
assign sext_ln1345_fu_319_p1 = { ret_V_15_reg_751[1], ret_V_15_reg_751[1], ret_V_15_reg_751 };
assign sext_ln69_1_fu_489_p1 = { op_11[7], op_11[7], op_11[7], op_11[7], op_11[7], op_11[7], op_11[7], op_11[7], op_11[7], op_11[7], op_11[7], op_11[7], op_11[7], op_11[7], op_11[7], op_11[7], op_11[7], op_11 };
assign sext_ln69_3_fu_498_p1 = { add_ln69_1_reg_792[4], add_ln69_1_reg_792[4], add_ln69_1_reg_792[4], add_ln69_1_reg_792[4], add_ln69_1_reg_792[4], add_ln69_1_reg_792[4], add_ln69_1_reg_792[4], add_ln69_1_reg_792[4], add_ln69_1_reg_792[4], add_ln69_1_reg_792[4], add_ln69_1_reg_792[4], add_ln69_1_reg_792[4], add_ln69_1_reg_792[4], add_ln69_1_reg_792[4], add_ln69_1_reg_792[4], add_ln69_1_reg_792[4], add_ln69_1_reg_792[4], add_ln69_1_reg_792[4], add_ln69_1_reg_792[4], add_ln69_1_reg_792[4], add_ln69_1_reg_792 };
assign sext_ln69_fu_393_p1 = { op_8[3], op_8 };
assign sext_ln703_1_fu_511_p1 = { op_13_V_reg_797[31], op_13_V_reg_797[31], op_13_V_reg_797[31], op_13_V_reg_797[31], op_13_V_reg_797[31], op_13_V_reg_797[31], op_13_V_reg_797[31], op_13_V_reg_797[31], op_13_V_reg_797[31], op_13_V_reg_797[31], op_13_V_reg_797[31], op_13_V_reg_797[31], op_13_V_reg_797[31], op_13_V_reg_797[31], op_13_V_reg_797[31], op_13_V_reg_797[31], op_13_V_reg_797[31], op_13_V_reg_797[31], op_13_V_reg_797[31], op_13_V_reg_797[31], op_13_V_reg_797[31], op_13_V_reg_797[31], op_13_V_reg_797[31], op_13_V_reg_797[31], op_13_V_reg_797 };
assign sext_ln703_2_fu_589_p0 = op_16;
assign sext_ln703_2_fu_589_p1 = { op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16 };
assign sext_ln703_3_fu_671_p0 = op_18;
assign sext_ln703_3_fu_671_p1 = { op_18[31], op_18[31], op_18[31], op_18[31], op_18[31], op_18[31], op_18[31], op_18 };
assign sext_ln703_fu_403_p0 = op_5;
assign sext_ln703_fu_403_p1 = { op_5[15], op_5[15], op_5 };
assign sext_ln850_fu_328_p1 = { tmp_1_reg_761[23], tmp_1_reg_761 };
assign tmp_fu_514_p3 = { op_23_V_reg_802, 23'h000000 };
assign trunc_ln213_1_fu_652_p1 = op_10[0];
assign trunc_ln213_fu_649_p1 = ret_reg_776[0];
assign trunc_ln728_1_fu_365_p1 = ret_fu_322_p2[1:0];
assign trunc_ln728_fu_435_p1 = ret_V_18_fu_421_p2[16:0];
assign trunc_ln851_1_fu_297_p1 = ret_V_16_fu_281_p2[8:0];
assign trunc_ln851_2_fu_507_p1 = op_13_V_fu_481_p3[22:0];
assign trunc_ln851_3_fu_627_p0 = op_16;
assign trunc_ln851_3_fu_627_p1 = op_16[0];
assign trunc_ln851_4_fu_702_p0 = op_18;
assign trunc_ln851_4_fu_702_p1 = op_18[5:0];
assign trunc_ln851_fu_251_p1 = op_2[0];
assign zext_ln1192_fu_417_p1 = { 2'h0, ret_reg_776[3], ret_reg_776[3], ret_reg_776[3], ret_reg_776[3], ret_reg_776, 8'h00 };
assign zext_ln69_fu_662_p1 = { 31'h00000000, op_17_V_fu_656_p2 };
assign \mul_2s_2s_4_1_1_U1.top_mul_2s_2s_4_1_1_Multiplier_0_U.a  = \mul_2s_2s_4_1_1_U1.din0 ;
assign \mul_2s_2s_4_1_1_U1.top_mul_2s_2s_4_1_1_Multiplier_0_U.b  = \mul_2s_2s_4_1_1_U1.din1 ;
assign \mul_2s_2s_4_1_1_U1.dout  = \mul_2s_2s_4_1_1_U1.top_mul_2s_2s_4_1_1_Multiplier_0_U.p ;
assign \mul_2s_2s_4_1_1_U1.din0  = ret_V_15_reg_751;
assign \mul_2s_2s_4_1_1_U1.din1  = ret_V_15_reg_751;
assign ret_fu_322_p2 = \mul_2s_2s_4_1_1_U1.dout ;
endmodule


// Machine B:
// Processed by function `add_clk_enable_signal` in `verilog_tricks.py`.
// Processed by function `remove_reset_signal` in `verilog_tricks.py`.
module top_B (
  ap_clk,
  ap_start,
  ap_done,
  ap_idle,
  ap_ready,
  op_0,
  op_2,
  op_3,
  op_5,
  op_8,
  op_10,
  op_11,
  op_14,
  op_16,
  op_18,
  op_19,
  op_30,
  op_30_ap_vld,
clk_enable
);
input clk_enable;


input ap_clk;
wire ap_rst;
assign ap_rst = op_30_ap_vld;
input ap_start;
input [3:0] op_0;
input [7:0] op_10;
input [7:0] op_11;
input [3:0] op_14;
input [7:0] op_16;
input [31:0] op_18;
input op_19;
input [3:0] op_2;
input [31:0] op_3;
input [15:0] op_5;
input [3:0] op_8;
output ap_done;
output ap_idle;
output ap_ready;
output [31:0] op_30;
output op_30_ap_vld;


reg [8:0] \add_18ns_18s_18_2_1_U7.top_add_18ns_18s_18_2_1_Adder_5_U.ain_s1 ;
reg [8:0] \add_18ns_18s_18_2_1_U7.top_add_18ns_18s_18_2_1_Adder_5_U.bin_s1 ;
reg \add_18ns_18s_18_2_1_U7.top_add_18ns_18s_18_2_1_Adder_5_U.carry_s1 ;
reg [8:0] \add_18ns_18s_18_2_1_U7.top_add_18ns_18s_18_2_1_Adder_5_U.sum_s1 ;
reg [12:0] \add_25ns_25s_25_2_1_U5.top_add_25ns_25s_25_2_1_Adder_3_U.ain_s1 ;
reg [12:0] \add_25ns_25s_25_2_1_U5.top_add_25ns_25s_25_2_1_Adder_3_U.bin_s1 ;
reg \add_25ns_25s_25_2_1_U5.top_add_25ns_25s_25_2_1_Adder_3_U.carry_s1 ;
reg [11:0] \add_25ns_25s_25_2_1_U5.top_add_25ns_25s_25_2_1_Adder_3_U.sum_s1 ;
reg [12:0] \add_25s_25ns_25_2_1_U3.top_add_25s_25ns_25_2_1_Adder_2_U.ain_s1 ;
reg [12:0] \add_25s_25ns_25_2_1_U3.top_add_25s_25ns_25_2_1_Adder_2_U.bin_s1 ;
reg \add_25s_25ns_25_2_1_U3.top_add_25s_25ns_25_2_1_Adder_2_U.carry_s1 ;
reg [11:0] \add_25s_25ns_25_2_1_U3.top_add_25s_25ns_25_2_1_Adder_2_U.sum_s1 ;
reg [12:0] \add_25s_25ns_25_2_1_U8.top_add_25s_25ns_25_2_1_Adder_2_U.ain_s1 ;
reg [12:0] \add_25s_25ns_25_2_1_U8.top_add_25s_25ns_25_2_1_Adder_2_U.bin_s1 ;
reg \add_25s_25ns_25_2_1_U8.top_add_25s_25ns_25_2_1_Adder_2_U.carry_s1 ;
reg [11:0] \add_25s_25ns_25_2_1_U8.top_add_25s_25ns_25_2_1_Adder_2_U.sum_s1 ;
reg \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.ain_s1 ;
reg \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.bin_s1 ;
reg \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.carry_s1 ;
reg \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.sum_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s1 ;
reg \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.carry_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.sum_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s1 ;
reg \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.carry_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.sum_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s1 ;
reg \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.carry_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.sum_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s1 ;
reg \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_7_U.carry_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_7_U.sum_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s1 ;
reg \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.carry_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.sum_s1 ;
reg [15:0] \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.ain_s1 ;
reg [15:0] \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.bin_s1 ;
reg \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.carry_s1 ;
reg [15:0] \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.sum_s1 ;
reg [15:0] \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.ain_s1 ;
reg [15:0] \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.bin_s1 ;
reg \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.carry_s1 ;
reg [15:0] \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.sum_s1 ;
reg [16:0] \add_33s_33ns_33_2_1_U1.top_add_33s_33ns_33_2_1_Adder_0_U.ain_s1 ;
reg [16:0] \add_33s_33ns_33_2_1_U1.top_add_33s_33ns_33_2_1_Adder_0_U.bin_s1 ;
reg \add_33s_33ns_33_2_1_U1.top_add_33s_33ns_33_2_1_Adder_0_U.carry_s1 ;
reg [15:0] \add_33s_33ns_33_2_1_U1.top_add_33s_33ns_33_2_1_Adder_0_U.sum_s1 ;
reg [16:0] \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_9_U.ain_s1 ;
reg [16:0] \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_9_U.bin_s1 ;
reg \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_9_U.carry_s1 ;
reg [16:0] \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_9_U.sum_s1 ;
reg [19:0] \add_39s_39s_39_2_1_U16.top_add_39s_39s_39_2_1_Adder_10_U.ain_s1 ;
reg [19:0] \add_39s_39s_39_2_1_U16.top_add_39s_39s_39_2_1_Adder_10_U.bin_s1 ;
reg \add_39s_39s_39_2_1_U16.top_add_39s_39s_39_2_1_Adder_10_U.carry_s1 ;
reg [18:0] \add_39s_39s_39_2_1_U16.top_add_39s_39s_39_2_1_Adder_10_U.sum_s1 ;
reg [27:0] \add_56s_56s_56_2_1_U9.top_add_56s_56s_56_2_1_Adder_6_U.ain_s1 ;
reg [27:0] \add_56s_56s_56_2_1_U9.top_add_56s_56s_56_2_1_Adder_6_U.bin_s1 ;
reg \add_56s_56s_56_2_1_U9.top_add_56s_56s_56_2_1_Adder_6_U.carry_s1 ;
reg [27:0] \add_56s_56s_56_2_1_U9.top_add_56s_56s_56_2_1_Adder_6_U.sum_s1 ;
reg [2:0] \add_5s_5ns_5_2_1_U6.top_add_5s_5ns_5_2_1_Adder_4_U.ain_s1 ;
reg [2:0] \add_5s_5ns_5_2_1_U6.top_add_5s_5ns_5_2_1_Adder_4_U.bin_s1 ;
reg \add_5s_5ns_5_2_1_U6.top_add_5s_5ns_5_2_1_Adder_4_U.carry_s1 ;
reg [1:0] \add_5s_5ns_5_2_1_U6.top_add_5s_5ns_5_2_1_Adder_4_U.sum_s1 ;
reg [24:0] add_ln691_1_reg_780;
reg [31:0] add_ln691_2_reg_905;
reg [31:0] add_ln691_3_reg_962;
reg [31:0] add_ln691_4_reg_1014;
reg [1:0] add_ln691_reg_775;
reg [4:0] add_ln69_1_reg_836;
reg [24:0] add_ln69_reg_831;
reg [31:0] ap_CS_fsm = 32'd1;
reg icmp_ln851_1_reg_888;
reg icmp_ln851_2_reg_997;
reg icmp_ln851_reg_770;
reg [31:0] op_13_V_reg_863;
reg [1:0] op_15_V_reg_826;
reg op_17_V_reg_967;
reg [24:0] op_23_V_reg_868;
reg [31:0] op_28_V_reg_982;
reg p_Result_7_reg_846;
reg p_Result_8_reg_852;
reg [1:0] ret_V_15_reg_785;
reg [32:0] ret_V_16_reg_735;
reg [24:0] ret_V_17_reg_790;
reg [17:0] ret_V_18_reg_841;
reg [31:0] ret_V_19_cast_reg_955;
reg [55:0] ret_V_19_reg_893;
reg [31:0] ret_V_20_reg_910;
reg [31:0] ret_V_21_cast_reg_1007;
reg [31:0] ret_V_21_reg_920;
reg [31:0] ret_V_22_reg_930;
reg [33:0] ret_V_23_reg_950;
reg [31:0] ret_V_24_reg_972;
reg [38:0] ret_V_25_reg_1002;
reg [31:0] ret_V_26_reg_1019;
reg [31:0] ret_V_8_cast_reg_898;
reg [1:0] ret_V_cast_reg_756;
reg [3:0] ret_reg_795;
reg [31:0] select_ln69_reg_1024;
reg [24:0] sext_ln850_reg_763;
reg [23:0] tmp_1_reg_740;
reg trunc_ln213_reg_801;
reg [8:0] trunc_ln851_1_reg_745;
reg [22:0] trunc_ln851_2_reg_873;
wire [24:0] _000_;
wire [31:0] _001_;
wire [31:0] _002_;
wire [31:0] _003_;
wire [1:0] _004_;
wire [4:0] _005_;
wire [24:0] _006_;
wire [31:0] _007_;
wire _008_;
wire _009_;
wire _010_;
wire [31:0] _011_;
wire [1:0] _012_;
wire _013_;
wire [24:0] _014_;
wire [31:0] _015_;
wire _016_;
wire _017_;
wire [1:0] _018_;
wire [32:0] _019_;
wire [24:0] _020_;
wire [17:0] _021_;
wire [31:0] _022_;
wire [55:0] _023_;
wire [31:0] _024_;
wire [31:0] _025_;
wire [31:0] _026_;
wire [31:0] _027_;
wire [33:0] _028_;
wire [31:0] _029_;
wire [38:0] _030_;
wire [31:0] _031_;
wire [31:0] _032_;
wire [1:0] _033_;
wire [3:0] _034_;
wire [31:0] _035_;
wire [24:0] _036_;
wire [23:0] _037_;
wire _038_;
wire [8:0] _039_;
wire [22:0] _040_;
wire [1:0] _041_;
wire _042_;
wire _043_;
wire _044_;
wire _045_;
wire _046_;
wire [8:0] _047_;
wire [8:0] _048_;
wire _049_;
wire [8:0] _050_;
wire [9:0] _051_;
wire [9:0] _052_;
wire [12:0] _053_;
wire [12:0] _054_;
wire _055_;
wire [11:0] _056_;
wire [12:0] _057_;
wire [13:0] _058_;
wire [12:0] _059_;
wire [12:0] _060_;
wire _061_;
wire [11:0] _062_;
wire [12:0] _063_;
wire [13:0] _064_;
wire [12:0] _065_;
wire [12:0] _066_;
wire _067_;
wire [11:0] _068_;
wire [12:0] _069_;
wire [13:0] _070_;
wire _071_;
wire _072_;
wire _073_;
wire _074_;
wire [1:0] _075_;
wire [1:0] _076_;
wire [15:0] _077_;
wire [15:0] _078_;
wire _079_;
wire [15:0] _080_;
wire [16:0] _081_;
wire [16:0] _082_;
wire [15:0] _083_;
wire [15:0] _084_;
wire _085_;
wire [15:0] _086_;
wire [16:0] _087_;
wire [16:0] _088_;
wire [15:0] _089_;
wire [15:0] _090_;
wire _091_;
wire [15:0] _092_;
wire [16:0] _093_;
wire [16:0] _094_;
wire [15:0] _095_;
wire [15:0] _096_;
wire _097_;
wire [15:0] _098_;
wire [16:0] _099_;
wire [16:0] _100_;
wire [15:0] _101_;
wire [15:0] _102_;
wire _103_;
wire [15:0] _104_;
wire [16:0] _105_;
wire [16:0] _106_;
wire [15:0] _107_;
wire [15:0] _108_;
wire _109_;
wire [15:0] _110_;
wire [16:0] _111_;
wire [16:0] _112_;
wire [15:0] _113_;
wire [15:0] _114_;
wire _115_;
wire [15:0] _116_;
wire [16:0] _117_;
wire [16:0] _118_;
wire [16:0] _119_;
wire [16:0] _120_;
wire _121_;
wire [15:0] _122_;
wire [16:0] _123_;
wire [17:0] _124_;
wire [16:0] _125_;
wire [16:0] _126_;
wire _127_;
wire [16:0] _128_;
wire [17:0] _129_;
wire [17:0] _130_;
wire [19:0] _131_;
wire [19:0] _132_;
wire _133_;
wire [18:0] _134_;
wire [19:0] _135_;
wire [20:0] _136_;
wire [27:0] _137_;
wire [27:0] _138_;
wire _139_;
wire [27:0] _140_;
wire [28:0] _141_;
wire [28:0] _142_;
wire [2:0] _143_;
wire [2:0] _144_;
wire _145_;
wire [1:0] _146_;
wire [2:0] _147_;
wire [3:0] _148_;
wire _149_;
wire _150_;
wire _151_;
wire _152_;
wire _153_;
wire _154_;
wire _155_;
wire _156_;
wire _157_;
wire _158_;
wire _159_;
wire _160_;
wire _161_;
wire _162_;
wire _163_;
wire _164_;
wire _165_;
wire _166_;
wire _167_;
wire _168_;
wire _169_;
wire _170_;
wire _171_;
wire _172_;
wire _173_;
wire _174_;
wire _175_;
wire _176_;
wire _177_;
wire _178_;
wire _179_;
wire _180_;
wire _181_;
wire _182_;
wire _183_;
wire \add_18ns_18s_18_2_1_U7.ce ;
wire \add_18ns_18s_18_2_1_U7.clk ;
wire [17:0] \add_18ns_18s_18_2_1_U7.din0 ;
wire [17:0] \add_18ns_18s_18_2_1_U7.din1 ;
wire [17:0] \add_18ns_18s_18_2_1_U7.dout ;
wire \add_18ns_18s_18_2_1_U7.reset ;
wire [17:0] \add_18ns_18s_18_2_1_U7.top_add_18ns_18s_18_2_1_Adder_5_U.a ;
wire [17:0] \add_18ns_18s_18_2_1_U7.top_add_18ns_18s_18_2_1_Adder_5_U.ain_s0 ;
wire [17:0] \add_18ns_18s_18_2_1_U7.top_add_18ns_18s_18_2_1_Adder_5_U.b ;
wire [17:0] \add_18ns_18s_18_2_1_U7.top_add_18ns_18s_18_2_1_Adder_5_U.bin_s0 ;
wire \add_18ns_18s_18_2_1_U7.top_add_18ns_18s_18_2_1_Adder_5_U.ce ;
wire \add_18ns_18s_18_2_1_U7.top_add_18ns_18s_18_2_1_Adder_5_U.clk ;
wire \add_18ns_18s_18_2_1_U7.top_add_18ns_18s_18_2_1_Adder_5_U.facout_s1 ;
wire \add_18ns_18s_18_2_1_U7.top_add_18ns_18s_18_2_1_Adder_5_U.facout_s2 ;
wire [8:0] \add_18ns_18s_18_2_1_U7.top_add_18ns_18s_18_2_1_Adder_5_U.fas_s1 ;
wire [8:0] \add_18ns_18s_18_2_1_U7.top_add_18ns_18s_18_2_1_Adder_5_U.fas_s2 ;
wire \add_18ns_18s_18_2_1_U7.top_add_18ns_18s_18_2_1_Adder_5_U.reset ;
wire [17:0] \add_18ns_18s_18_2_1_U7.top_add_18ns_18s_18_2_1_Adder_5_U.s ;
wire [8:0] \add_18ns_18s_18_2_1_U7.top_add_18ns_18s_18_2_1_Adder_5_U.u1.a ;
wire [8:0] \add_18ns_18s_18_2_1_U7.top_add_18ns_18s_18_2_1_Adder_5_U.u1.b ;
wire \add_18ns_18s_18_2_1_U7.top_add_18ns_18s_18_2_1_Adder_5_U.u1.cin ;
wire \add_18ns_18s_18_2_1_U7.top_add_18ns_18s_18_2_1_Adder_5_U.u1.cout ;
wire [8:0] \add_18ns_18s_18_2_1_U7.top_add_18ns_18s_18_2_1_Adder_5_U.u1.s ;
wire [8:0] \add_18ns_18s_18_2_1_U7.top_add_18ns_18s_18_2_1_Adder_5_U.u2.a ;
wire [8:0] \add_18ns_18s_18_2_1_U7.top_add_18ns_18s_18_2_1_Adder_5_U.u2.b ;
wire \add_18ns_18s_18_2_1_U7.top_add_18ns_18s_18_2_1_Adder_5_U.u2.cin ;
wire \add_18ns_18s_18_2_1_U7.top_add_18ns_18s_18_2_1_Adder_5_U.u2.cout ;
wire [8:0] \add_18ns_18s_18_2_1_U7.top_add_18ns_18s_18_2_1_Adder_5_U.u2.s ;
wire \add_25ns_25s_25_2_1_U5.ce ;
wire \add_25ns_25s_25_2_1_U5.clk ;
wire [24:0] \add_25ns_25s_25_2_1_U5.din0 ;
wire [24:0] \add_25ns_25s_25_2_1_U5.din1 ;
wire [24:0] \add_25ns_25s_25_2_1_U5.dout ;
wire \add_25ns_25s_25_2_1_U5.reset ;
wire [24:0] \add_25ns_25s_25_2_1_U5.top_add_25ns_25s_25_2_1_Adder_3_U.a ;
wire [24:0] \add_25ns_25s_25_2_1_U5.top_add_25ns_25s_25_2_1_Adder_3_U.ain_s0 ;
wire [24:0] \add_25ns_25s_25_2_1_U5.top_add_25ns_25s_25_2_1_Adder_3_U.b ;
wire [24:0] \add_25ns_25s_25_2_1_U5.top_add_25ns_25s_25_2_1_Adder_3_U.bin_s0 ;
wire \add_25ns_25s_25_2_1_U5.top_add_25ns_25s_25_2_1_Adder_3_U.ce ;
wire \add_25ns_25s_25_2_1_U5.top_add_25ns_25s_25_2_1_Adder_3_U.clk ;
wire \add_25ns_25s_25_2_1_U5.top_add_25ns_25s_25_2_1_Adder_3_U.facout_s1 ;
wire \add_25ns_25s_25_2_1_U5.top_add_25ns_25s_25_2_1_Adder_3_U.facout_s2 ;
wire [11:0] \add_25ns_25s_25_2_1_U5.top_add_25ns_25s_25_2_1_Adder_3_U.fas_s1 ;
wire [12:0] \add_25ns_25s_25_2_1_U5.top_add_25ns_25s_25_2_1_Adder_3_U.fas_s2 ;
wire \add_25ns_25s_25_2_1_U5.top_add_25ns_25s_25_2_1_Adder_3_U.reset ;
wire [24:0] \add_25ns_25s_25_2_1_U5.top_add_25ns_25s_25_2_1_Adder_3_U.s ;
wire [11:0] \add_25ns_25s_25_2_1_U5.top_add_25ns_25s_25_2_1_Adder_3_U.u1.a ;
wire [11:0] \add_25ns_25s_25_2_1_U5.top_add_25ns_25s_25_2_1_Adder_3_U.u1.b ;
wire \add_25ns_25s_25_2_1_U5.top_add_25ns_25s_25_2_1_Adder_3_U.u1.cin ;
wire \add_25ns_25s_25_2_1_U5.top_add_25ns_25s_25_2_1_Adder_3_U.u1.cout ;
wire [11:0] \add_25ns_25s_25_2_1_U5.top_add_25ns_25s_25_2_1_Adder_3_U.u1.s ;
wire [12:0] \add_25ns_25s_25_2_1_U5.top_add_25ns_25s_25_2_1_Adder_3_U.u2.a ;
wire [12:0] \add_25ns_25s_25_2_1_U5.top_add_25ns_25s_25_2_1_Adder_3_U.u2.b ;
wire \add_25ns_25s_25_2_1_U5.top_add_25ns_25s_25_2_1_Adder_3_U.u2.cin ;
wire \add_25ns_25s_25_2_1_U5.top_add_25ns_25s_25_2_1_Adder_3_U.u2.cout ;
wire [12:0] \add_25ns_25s_25_2_1_U5.top_add_25ns_25s_25_2_1_Adder_3_U.u2.s ;
wire \add_25s_25ns_25_2_1_U3.ce ;
wire \add_25s_25ns_25_2_1_U3.clk ;
wire [24:0] \add_25s_25ns_25_2_1_U3.din0 ;
wire [24:0] \add_25s_25ns_25_2_1_U3.din1 ;
wire [24:0] \add_25s_25ns_25_2_1_U3.dout ;
wire \add_25s_25ns_25_2_1_U3.reset ;
wire [24:0] \add_25s_25ns_25_2_1_U3.top_add_25s_25ns_25_2_1_Adder_2_U.a ;
wire [24:0] \add_25s_25ns_25_2_1_U3.top_add_25s_25ns_25_2_1_Adder_2_U.ain_s0 ;
wire [24:0] \add_25s_25ns_25_2_1_U3.top_add_25s_25ns_25_2_1_Adder_2_U.b ;
wire [24:0] \add_25s_25ns_25_2_1_U3.top_add_25s_25ns_25_2_1_Adder_2_U.bin_s0 ;
wire \add_25s_25ns_25_2_1_U3.top_add_25s_25ns_25_2_1_Adder_2_U.ce ;
wire \add_25s_25ns_25_2_1_U3.top_add_25s_25ns_25_2_1_Adder_2_U.clk ;
wire \add_25s_25ns_25_2_1_U3.top_add_25s_25ns_25_2_1_Adder_2_U.facout_s1 ;
wire \add_25s_25ns_25_2_1_U3.top_add_25s_25ns_25_2_1_Adder_2_U.facout_s2 ;
wire [11:0] \add_25s_25ns_25_2_1_U3.top_add_25s_25ns_25_2_1_Adder_2_U.fas_s1 ;
wire [12:0] \add_25s_25ns_25_2_1_U3.top_add_25s_25ns_25_2_1_Adder_2_U.fas_s2 ;
wire \add_25s_25ns_25_2_1_U3.top_add_25s_25ns_25_2_1_Adder_2_U.reset ;
wire [24:0] \add_25s_25ns_25_2_1_U3.top_add_25s_25ns_25_2_1_Adder_2_U.s ;
wire [11:0] \add_25s_25ns_25_2_1_U3.top_add_25s_25ns_25_2_1_Adder_2_U.u1.a ;
wire [11:0] \add_25s_25ns_25_2_1_U3.top_add_25s_25ns_25_2_1_Adder_2_U.u1.b ;
wire \add_25s_25ns_25_2_1_U3.top_add_25s_25ns_25_2_1_Adder_2_U.u1.cin ;
wire \add_25s_25ns_25_2_1_U3.top_add_25s_25ns_25_2_1_Adder_2_U.u1.cout ;
wire [11:0] \add_25s_25ns_25_2_1_U3.top_add_25s_25ns_25_2_1_Adder_2_U.u1.s ;
wire [12:0] \add_25s_25ns_25_2_1_U3.top_add_25s_25ns_25_2_1_Adder_2_U.u2.a ;
wire [12:0] \add_25s_25ns_25_2_1_U3.top_add_25s_25ns_25_2_1_Adder_2_U.u2.b ;
wire \add_25s_25ns_25_2_1_U3.top_add_25s_25ns_25_2_1_Adder_2_U.u2.cin ;
wire \add_25s_25ns_25_2_1_U3.top_add_25s_25ns_25_2_1_Adder_2_U.u2.cout ;
wire [12:0] \add_25s_25ns_25_2_1_U3.top_add_25s_25ns_25_2_1_Adder_2_U.u2.s ;
wire \add_25s_25ns_25_2_1_U8.ce ;
wire \add_25s_25ns_25_2_1_U8.clk ;
wire [24:0] \add_25s_25ns_25_2_1_U8.din0 ;
wire [24:0] \add_25s_25ns_25_2_1_U8.din1 ;
wire [24:0] \add_25s_25ns_25_2_1_U8.dout ;
wire \add_25s_25ns_25_2_1_U8.reset ;
wire [24:0] \add_25s_25ns_25_2_1_U8.top_add_25s_25ns_25_2_1_Adder_2_U.a ;
wire [24:0] \add_25s_25ns_25_2_1_U8.top_add_25s_25ns_25_2_1_Adder_2_U.ain_s0 ;
wire [24:0] \add_25s_25ns_25_2_1_U8.top_add_25s_25ns_25_2_1_Adder_2_U.b ;
wire [24:0] \add_25s_25ns_25_2_1_U8.top_add_25s_25ns_25_2_1_Adder_2_U.bin_s0 ;
wire \add_25s_25ns_25_2_1_U8.top_add_25s_25ns_25_2_1_Adder_2_U.ce ;
wire \add_25s_25ns_25_2_1_U8.top_add_25s_25ns_25_2_1_Adder_2_U.clk ;
wire \add_25s_25ns_25_2_1_U8.top_add_25s_25ns_25_2_1_Adder_2_U.facout_s1 ;
wire \add_25s_25ns_25_2_1_U8.top_add_25s_25ns_25_2_1_Adder_2_U.facout_s2 ;
wire [11:0] \add_25s_25ns_25_2_1_U8.top_add_25s_25ns_25_2_1_Adder_2_U.fas_s1 ;
wire [12:0] \add_25s_25ns_25_2_1_U8.top_add_25s_25ns_25_2_1_Adder_2_U.fas_s2 ;
wire \add_25s_25ns_25_2_1_U8.top_add_25s_25ns_25_2_1_Adder_2_U.reset ;
wire [24:0] \add_25s_25ns_25_2_1_U8.top_add_25s_25ns_25_2_1_Adder_2_U.s ;
wire [11:0] \add_25s_25ns_25_2_1_U8.top_add_25s_25ns_25_2_1_Adder_2_U.u1.a ;
wire [11:0] \add_25s_25ns_25_2_1_U8.top_add_25s_25ns_25_2_1_Adder_2_U.u1.b ;
wire \add_25s_25ns_25_2_1_U8.top_add_25s_25ns_25_2_1_Adder_2_U.u1.cin ;
wire \add_25s_25ns_25_2_1_U8.top_add_25s_25ns_25_2_1_Adder_2_U.u1.cout ;
wire [11:0] \add_25s_25ns_25_2_1_U8.top_add_25s_25ns_25_2_1_Adder_2_U.u1.s ;
wire [12:0] \add_25s_25ns_25_2_1_U8.top_add_25s_25ns_25_2_1_Adder_2_U.u2.a ;
wire [12:0] \add_25s_25ns_25_2_1_U8.top_add_25s_25ns_25_2_1_Adder_2_U.u2.b ;
wire \add_25s_25ns_25_2_1_U8.top_add_25s_25ns_25_2_1_Adder_2_U.u2.cin ;
wire \add_25s_25ns_25_2_1_U8.top_add_25s_25ns_25_2_1_Adder_2_U.u2.cout ;
wire [12:0] \add_25s_25ns_25_2_1_U8.top_add_25s_25ns_25_2_1_Adder_2_U.u2.s ;
wire \add_2ns_2ns_2_2_1_U2.ce ;
wire \add_2ns_2ns_2_2_1_U2.clk ;
wire [1:0] \add_2ns_2ns_2_2_1_U2.din0 ;
wire [1:0] \add_2ns_2ns_2_2_1_U2.din1 ;
wire [1:0] \add_2ns_2ns_2_2_1_U2.dout ;
wire \add_2ns_2ns_2_2_1_U2.reset ;
wire [1:0] \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.a ;
wire [1:0] \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.ain_s0 ;
wire [1:0] \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.b ;
wire [1:0] \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.bin_s0 ;
wire \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.ce ;
wire \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.clk ;
wire \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.facout_s1 ;
wire \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.facout_s2 ;
wire \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.fas_s1 ;
wire \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.fas_s2 ;
wire \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.reset ;
wire [1:0] \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.s ;
wire \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.a ;
wire \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.b ;
wire \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.cin ;
wire \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.cout ;
wire \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.s ;
wire \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.a ;
wire \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.b ;
wire \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.cin ;
wire \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.cout ;
wire \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.s ;
wire \add_32ns_32ns_32_2_1_U10.ce ;
wire \add_32ns_32ns_32_2_1_U10.clk ;
wire [31:0] \add_32ns_32ns_32_2_1_U10.din0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U10.din1 ;
wire [31:0] \add_32ns_32ns_32_2_1_U10.dout ;
wire \add_32ns_32ns_32_2_1_U10.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.a ;
wire [31:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.b ;
wire [31:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s0 ;
wire \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.ce ;
wire \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.clk ;
wire \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.facout_s1 ;
wire \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.facout_s2 ;
wire [15:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s1 ;
wire [15:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s2 ;
wire \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.b ;
wire \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cin ;
wire \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.b ;
wire \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cin ;
wire \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.s ;
wire \add_32ns_32ns_32_2_1_U14.ce ;
wire \add_32ns_32ns_32_2_1_U14.clk ;
wire [31:0] \add_32ns_32ns_32_2_1_U14.din0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U14.din1 ;
wire [31:0] \add_32ns_32ns_32_2_1_U14.dout ;
wire \add_32ns_32ns_32_2_1_U14.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.a ;
wire [31:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.b ;
wire [31:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s0 ;
wire \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.ce ;
wire \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.clk ;
wire \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.facout_s1 ;
wire \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.facout_s2 ;
wire [15:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s1 ;
wire [15:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s2 ;
wire \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.b ;
wire \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cin ;
wire \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.b ;
wire \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cin ;
wire \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.s ;
wire \add_32ns_32ns_32_2_1_U15.ce ;
wire \add_32ns_32ns_32_2_1_U15.clk ;
wire [31:0] \add_32ns_32ns_32_2_1_U15.din0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U15.din1 ;
wire [31:0] \add_32ns_32ns_32_2_1_U15.dout ;
wire \add_32ns_32ns_32_2_1_U15.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.a ;
wire [31:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.b ;
wire [31:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s0 ;
wire \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.ce ;
wire \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.clk ;
wire \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.facout_s1 ;
wire \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.facout_s2 ;
wire [15:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s1 ;
wire [15:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s2 ;
wire \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.b ;
wire \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cin ;
wire \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.b ;
wire \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cin ;
wire \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.s ;
wire \add_32ns_32ns_32_2_1_U17.ce ;
wire \add_32ns_32ns_32_2_1_U17.clk ;
wire [31:0] \add_32ns_32ns_32_2_1_U17.din0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U17.din1 ;
wire [31:0] \add_32ns_32ns_32_2_1_U17.dout ;
wire \add_32ns_32ns_32_2_1_U17.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_7_U.a ;
wire [31:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_7_U.b ;
wire [31:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s0 ;
wire \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_7_U.ce ;
wire \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_7_U.clk ;
wire \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_7_U.facout_s1 ;
wire \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_7_U.facout_s2 ;
wire [15:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s1 ;
wire [15:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s2 ;
wire \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_7_U.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_7_U.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.b ;
wire \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cin ;
wire \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.b ;
wire \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cin ;
wire \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.s ;
wire \add_32ns_32ns_32_2_1_U18.ce ;
wire \add_32ns_32ns_32_2_1_U18.clk ;
wire [31:0] \add_32ns_32ns_32_2_1_U18.din0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U18.din1 ;
wire [31:0] \add_32ns_32ns_32_2_1_U18.dout ;
wire \add_32ns_32ns_32_2_1_U18.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.a ;
wire [31:0] \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.b ;
wire [31:0] \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s0 ;
wire \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.ce ;
wire \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.clk ;
wire \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.facout_s1 ;
wire \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.facout_s2 ;
wire [15:0] \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s1 ;
wire [15:0] \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s2 ;
wire \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.b ;
wire \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cin ;
wire \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.b ;
wire \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cin ;
wire \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.s ;
wire \add_32ns_32s_32_2_1_U11.ce ;
wire \add_32ns_32s_32_2_1_U11.clk ;
wire [31:0] \add_32ns_32s_32_2_1_U11.din0 ;
wire [31:0] \add_32ns_32s_32_2_1_U11.din1 ;
wire [31:0] \add_32ns_32s_32_2_1_U11.dout ;
wire \add_32ns_32s_32_2_1_U11.reset ;
wire [31:0] \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.a ;
wire [31:0] \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.ain_s0 ;
wire [31:0] \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.b ;
wire [31:0] \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.bin_s0 ;
wire \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.ce ;
wire \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.clk ;
wire \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.facout_s1 ;
wire \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.facout_s2 ;
wire [15:0] \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.fas_s1 ;
wire [15:0] \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.fas_s2 ;
wire \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.reset ;
wire [31:0] \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.s ;
wire [15:0] \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.u1.a ;
wire [15:0] \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.u1.b ;
wire \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.u1.cin ;
wire \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.u1.cout ;
wire [15:0] \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.u1.s ;
wire [15:0] \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.u2.a ;
wire [15:0] \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.u2.b ;
wire \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.u2.cin ;
wire \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.u2.cout ;
wire [15:0] \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.u2.s ;
wire \add_32ns_32s_32_2_1_U12.ce ;
wire \add_32ns_32s_32_2_1_U12.clk ;
wire [31:0] \add_32ns_32s_32_2_1_U12.din0 ;
wire [31:0] \add_32ns_32s_32_2_1_U12.din1 ;
wire [31:0] \add_32ns_32s_32_2_1_U12.dout ;
wire \add_32ns_32s_32_2_1_U12.reset ;
wire [31:0] \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.a ;
wire [31:0] \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.ain_s0 ;
wire [31:0] \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.b ;
wire [31:0] \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.bin_s0 ;
wire \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.ce ;
wire \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.clk ;
wire \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.facout_s1 ;
wire \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.facout_s2 ;
wire [15:0] \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.fas_s1 ;
wire [15:0] \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.fas_s2 ;
wire \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.reset ;
wire [31:0] \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.s ;
wire [15:0] \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.u1.a ;
wire [15:0] \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.u1.b ;
wire \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.u1.cin ;
wire \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.u1.cout ;
wire [15:0] \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.u1.s ;
wire [15:0] \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.u2.a ;
wire [15:0] \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.u2.b ;
wire \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.u2.cin ;
wire \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.u2.cout ;
wire [15:0] \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.u2.s ;
wire \add_33s_33ns_33_2_1_U1.ce ;
wire \add_33s_33ns_33_2_1_U1.clk ;
wire [32:0] \add_33s_33ns_33_2_1_U1.din0 ;
wire [32:0] \add_33s_33ns_33_2_1_U1.din1 ;
wire [32:0] \add_33s_33ns_33_2_1_U1.dout ;
wire \add_33s_33ns_33_2_1_U1.reset ;
wire [32:0] \add_33s_33ns_33_2_1_U1.top_add_33s_33ns_33_2_1_Adder_0_U.a ;
wire [32:0] \add_33s_33ns_33_2_1_U1.top_add_33s_33ns_33_2_1_Adder_0_U.ain_s0 ;
wire [32:0] \add_33s_33ns_33_2_1_U1.top_add_33s_33ns_33_2_1_Adder_0_U.b ;
wire [32:0] \add_33s_33ns_33_2_1_U1.top_add_33s_33ns_33_2_1_Adder_0_U.bin_s0 ;
wire \add_33s_33ns_33_2_1_U1.top_add_33s_33ns_33_2_1_Adder_0_U.ce ;
wire \add_33s_33ns_33_2_1_U1.top_add_33s_33ns_33_2_1_Adder_0_U.clk ;
wire \add_33s_33ns_33_2_1_U1.top_add_33s_33ns_33_2_1_Adder_0_U.facout_s1 ;
wire \add_33s_33ns_33_2_1_U1.top_add_33s_33ns_33_2_1_Adder_0_U.facout_s2 ;
wire [15:0] \add_33s_33ns_33_2_1_U1.top_add_33s_33ns_33_2_1_Adder_0_U.fas_s1 ;
wire [16:0] \add_33s_33ns_33_2_1_U1.top_add_33s_33ns_33_2_1_Adder_0_U.fas_s2 ;
wire \add_33s_33ns_33_2_1_U1.top_add_33s_33ns_33_2_1_Adder_0_U.reset ;
wire [32:0] \add_33s_33ns_33_2_1_U1.top_add_33s_33ns_33_2_1_Adder_0_U.s ;
wire [15:0] \add_33s_33ns_33_2_1_U1.top_add_33s_33ns_33_2_1_Adder_0_U.u1.a ;
wire [15:0] \add_33s_33ns_33_2_1_U1.top_add_33s_33ns_33_2_1_Adder_0_U.u1.b ;
wire \add_33s_33ns_33_2_1_U1.top_add_33s_33ns_33_2_1_Adder_0_U.u1.cin ;
wire \add_33s_33ns_33_2_1_U1.top_add_33s_33ns_33_2_1_Adder_0_U.u1.cout ;
wire [15:0] \add_33s_33ns_33_2_1_U1.top_add_33s_33ns_33_2_1_Adder_0_U.u1.s ;
wire [16:0] \add_33s_33ns_33_2_1_U1.top_add_33s_33ns_33_2_1_Adder_0_U.u2.a ;
wire [16:0] \add_33s_33ns_33_2_1_U1.top_add_33s_33ns_33_2_1_Adder_0_U.u2.b ;
wire \add_33s_33ns_33_2_1_U1.top_add_33s_33ns_33_2_1_Adder_0_U.u2.cin ;
wire \add_33s_33ns_33_2_1_U1.top_add_33s_33ns_33_2_1_Adder_0_U.u2.cout ;
wire [16:0] \add_33s_33ns_33_2_1_U1.top_add_33s_33ns_33_2_1_Adder_0_U.u2.s ;
wire \add_34s_34s_34_2_1_U13.ce ;
wire \add_34s_34s_34_2_1_U13.clk ;
wire [33:0] \add_34s_34s_34_2_1_U13.din0 ;
wire [33:0] \add_34s_34s_34_2_1_U13.din1 ;
wire [33:0] \add_34s_34s_34_2_1_U13.dout ;
wire \add_34s_34s_34_2_1_U13.reset ;
wire [33:0] \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_9_U.a ;
wire [33:0] \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_9_U.ain_s0 ;
wire [33:0] \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_9_U.b ;
wire [33:0] \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_9_U.bin_s0 ;
wire \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_9_U.ce ;
wire \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_9_U.clk ;
wire \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_9_U.facout_s1 ;
wire \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_9_U.facout_s2 ;
wire [16:0] \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_9_U.fas_s1 ;
wire [16:0] \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_9_U.fas_s2 ;
wire \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_9_U.reset ;
wire [33:0] \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_9_U.s ;
wire [16:0] \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_9_U.u1.a ;
wire [16:0] \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_9_U.u1.b ;
wire \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_9_U.u1.cin ;
wire \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_9_U.u1.cout ;
wire [16:0] \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_9_U.u1.s ;
wire [16:0] \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_9_U.u2.a ;
wire [16:0] \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_9_U.u2.b ;
wire \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_9_U.u2.cin ;
wire \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_9_U.u2.cout ;
wire [16:0] \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_9_U.u2.s ;
wire \add_39s_39s_39_2_1_U16.ce ;
wire \add_39s_39s_39_2_1_U16.clk ;
wire [38:0] \add_39s_39s_39_2_1_U16.din0 ;
wire [38:0] \add_39s_39s_39_2_1_U16.din1 ;
wire [38:0] \add_39s_39s_39_2_1_U16.dout ;
wire \add_39s_39s_39_2_1_U16.reset ;
wire [38:0] \add_39s_39s_39_2_1_U16.top_add_39s_39s_39_2_1_Adder_10_U.a ;
wire [38:0] \add_39s_39s_39_2_1_U16.top_add_39s_39s_39_2_1_Adder_10_U.ain_s0 ;
wire [38:0] \add_39s_39s_39_2_1_U16.top_add_39s_39s_39_2_1_Adder_10_U.b ;
wire [38:0] \add_39s_39s_39_2_1_U16.top_add_39s_39s_39_2_1_Adder_10_U.bin_s0 ;
wire \add_39s_39s_39_2_1_U16.top_add_39s_39s_39_2_1_Adder_10_U.ce ;
wire \add_39s_39s_39_2_1_U16.top_add_39s_39s_39_2_1_Adder_10_U.clk ;
wire \add_39s_39s_39_2_1_U16.top_add_39s_39s_39_2_1_Adder_10_U.facout_s1 ;
wire \add_39s_39s_39_2_1_U16.top_add_39s_39s_39_2_1_Adder_10_U.facout_s2 ;
wire [18:0] \add_39s_39s_39_2_1_U16.top_add_39s_39s_39_2_1_Adder_10_U.fas_s1 ;
wire [19:0] \add_39s_39s_39_2_1_U16.top_add_39s_39s_39_2_1_Adder_10_U.fas_s2 ;
wire \add_39s_39s_39_2_1_U16.top_add_39s_39s_39_2_1_Adder_10_U.reset ;
wire [38:0] \add_39s_39s_39_2_1_U16.top_add_39s_39s_39_2_1_Adder_10_U.s ;
wire [18:0] \add_39s_39s_39_2_1_U16.top_add_39s_39s_39_2_1_Adder_10_U.u1.a ;
wire [18:0] \add_39s_39s_39_2_1_U16.top_add_39s_39s_39_2_1_Adder_10_U.u1.b ;
wire \add_39s_39s_39_2_1_U16.top_add_39s_39s_39_2_1_Adder_10_U.u1.cin ;
wire \add_39s_39s_39_2_1_U16.top_add_39s_39s_39_2_1_Adder_10_U.u1.cout ;
wire [18:0] \add_39s_39s_39_2_1_U16.top_add_39s_39s_39_2_1_Adder_10_U.u1.s ;
wire [19:0] \add_39s_39s_39_2_1_U16.top_add_39s_39s_39_2_1_Adder_10_U.u2.a ;
wire [19:0] \add_39s_39s_39_2_1_U16.top_add_39s_39s_39_2_1_Adder_10_U.u2.b ;
wire \add_39s_39s_39_2_1_U16.top_add_39s_39s_39_2_1_Adder_10_U.u2.cin ;
wire \add_39s_39s_39_2_1_U16.top_add_39s_39s_39_2_1_Adder_10_U.u2.cout ;
wire [19:0] \add_39s_39s_39_2_1_U16.top_add_39s_39s_39_2_1_Adder_10_U.u2.s ;
wire \add_56s_56s_56_2_1_U9.ce ;
wire \add_56s_56s_56_2_1_U9.clk ;
wire [55:0] \add_56s_56s_56_2_1_U9.din0 ;
wire [55:0] \add_56s_56s_56_2_1_U9.din1 ;
wire [55:0] \add_56s_56s_56_2_1_U9.dout ;
wire \add_56s_56s_56_2_1_U9.reset ;
wire [55:0] \add_56s_56s_56_2_1_U9.top_add_56s_56s_56_2_1_Adder_6_U.a ;
wire [55:0] \add_56s_56s_56_2_1_U9.top_add_56s_56s_56_2_1_Adder_6_U.ain_s0 ;
wire [55:0] \add_56s_56s_56_2_1_U9.top_add_56s_56s_56_2_1_Adder_6_U.b ;
wire [55:0] \add_56s_56s_56_2_1_U9.top_add_56s_56s_56_2_1_Adder_6_U.bin_s0 ;
wire \add_56s_56s_56_2_1_U9.top_add_56s_56s_56_2_1_Adder_6_U.ce ;
wire \add_56s_56s_56_2_1_U9.top_add_56s_56s_56_2_1_Adder_6_U.clk ;
wire \add_56s_56s_56_2_1_U9.top_add_56s_56s_56_2_1_Adder_6_U.facout_s1 ;
wire \add_56s_56s_56_2_1_U9.top_add_56s_56s_56_2_1_Adder_6_U.facout_s2 ;
wire [27:0] \add_56s_56s_56_2_1_U9.top_add_56s_56s_56_2_1_Adder_6_U.fas_s1 ;
wire [27:0] \add_56s_56s_56_2_1_U9.top_add_56s_56s_56_2_1_Adder_6_U.fas_s2 ;
wire \add_56s_56s_56_2_1_U9.top_add_56s_56s_56_2_1_Adder_6_U.reset ;
wire [55:0] \add_56s_56s_56_2_1_U9.top_add_56s_56s_56_2_1_Adder_6_U.s ;
wire [27:0] \add_56s_56s_56_2_1_U9.top_add_56s_56s_56_2_1_Adder_6_U.u1.a ;
wire [27:0] \add_56s_56s_56_2_1_U9.top_add_56s_56s_56_2_1_Adder_6_U.u1.b ;
wire \add_56s_56s_56_2_1_U9.top_add_56s_56s_56_2_1_Adder_6_U.u1.cin ;
wire \add_56s_56s_56_2_1_U9.top_add_56s_56s_56_2_1_Adder_6_U.u1.cout ;
wire [27:0] \add_56s_56s_56_2_1_U9.top_add_56s_56s_56_2_1_Adder_6_U.u1.s ;
wire [27:0] \add_56s_56s_56_2_1_U9.top_add_56s_56s_56_2_1_Adder_6_U.u2.a ;
wire [27:0] \add_56s_56s_56_2_1_U9.top_add_56s_56s_56_2_1_Adder_6_U.u2.b ;
wire \add_56s_56s_56_2_1_U9.top_add_56s_56s_56_2_1_Adder_6_U.u2.cin ;
wire \add_56s_56s_56_2_1_U9.top_add_56s_56s_56_2_1_Adder_6_U.u2.cout ;
wire [27:0] \add_56s_56s_56_2_1_U9.top_add_56s_56s_56_2_1_Adder_6_U.u2.s ;
wire \add_5s_5ns_5_2_1_U6.ce ;
wire \add_5s_5ns_5_2_1_U6.clk ;
wire [4:0] \add_5s_5ns_5_2_1_U6.din0 ;
wire [4:0] \add_5s_5ns_5_2_1_U6.din1 ;
wire [4:0] \add_5s_5ns_5_2_1_U6.dout ;
wire \add_5s_5ns_5_2_1_U6.reset ;
wire [4:0] \add_5s_5ns_5_2_1_U6.top_add_5s_5ns_5_2_1_Adder_4_U.a ;
wire [4:0] \add_5s_5ns_5_2_1_U6.top_add_5s_5ns_5_2_1_Adder_4_U.ain_s0 ;
wire [4:0] \add_5s_5ns_5_2_1_U6.top_add_5s_5ns_5_2_1_Adder_4_U.b ;
wire [4:0] \add_5s_5ns_5_2_1_U6.top_add_5s_5ns_5_2_1_Adder_4_U.bin_s0 ;
wire \add_5s_5ns_5_2_1_U6.top_add_5s_5ns_5_2_1_Adder_4_U.ce ;
wire \add_5s_5ns_5_2_1_U6.top_add_5s_5ns_5_2_1_Adder_4_U.clk ;
wire \add_5s_5ns_5_2_1_U6.top_add_5s_5ns_5_2_1_Adder_4_U.facout_s1 ;
wire \add_5s_5ns_5_2_1_U6.top_add_5s_5ns_5_2_1_Adder_4_U.facout_s2 ;
wire [1:0] \add_5s_5ns_5_2_1_U6.top_add_5s_5ns_5_2_1_Adder_4_U.fas_s1 ;
wire [2:0] \add_5s_5ns_5_2_1_U6.top_add_5s_5ns_5_2_1_Adder_4_U.fas_s2 ;
wire \add_5s_5ns_5_2_1_U6.top_add_5s_5ns_5_2_1_Adder_4_U.reset ;
wire [4:0] \add_5s_5ns_5_2_1_U6.top_add_5s_5ns_5_2_1_Adder_4_U.s ;
wire [1:0] \add_5s_5ns_5_2_1_U6.top_add_5s_5ns_5_2_1_Adder_4_U.u1.a ;
wire [1:0] \add_5s_5ns_5_2_1_U6.top_add_5s_5ns_5_2_1_Adder_4_U.u1.b ;
wire \add_5s_5ns_5_2_1_U6.top_add_5s_5ns_5_2_1_Adder_4_U.u1.cin ;
wire \add_5s_5ns_5_2_1_U6.top_add_5s_5ns_5_2_1_Adder_4_U.u1.cout ;
wire [1:0] \add_5s_5ns_5_2_1_U6.top_add_5s_5ns_5_2_1_Adder_4_U.u1.s ;
wire [2:0] \add_5s_5ns_5_2_1_U6.top_add_5s_5ns_5_2_1_Adder_4_U.u2.a ;
wire [2:0] \add_5s_5ns_5_2_1_U6.top_add_5s_5ns_5_2_1_Adder_4_U.u2.b ;
wire \add_5s_5ns_5_2_1_U6.top_add_5s_5ns_5_2_1_Adder_4_U.u2.cin ;
wire \add_5s_5ns_5_2_1_U6.top_add_5s_5ns_5_2_1_Adder_4_U.u2.cout ;
wire [2:0] \add_5s_5ns_5_2_1_U6.top_add_5s_5ns_5_2_1_Adder_4_U.u2.s ;
wire ap_CS_fsm_state1;
wire ap_CS_fsm_state10;
wire ap_CS_fsm_state11;
wire ap_CS_fsm_state12;
wire ap_CS_fsm_state13;
wire ap_CS_fsm_state14;
wire ap_CS_fsm_state15;
wire ap_CS_fsm_state16;
wire ap_CS_fsm_state17;
wire ap_CS_fsm_state18;
wire ap_CS_fsm_state19;
wire ap_CS_fsm_state2;
wire ap_CS_fsm_state20;
wire ap_CS_fsm_state21;
wire ap_CS_fsm_state22;
wire ap_CS_fsm_state23;
wire ap_CS_fsm_state24;
wire ap_CS_fsm_state25;
wire ap_CS_fsm_state26;
wire ap_CS_fsm_state27;
wire ap_CS_fsm_state28;
wire ap_CS_fsm_state29;
wire ap_CS_fsm_state3;
wire ap_CS_fsm_state30;
wire ap_CS_fsm_state31;
wire ap_CS_fsm_state32;
wire ap_CS_fsm_state4;
wire ap_CS_fsm_state5;
wire ap_CS_fsm_state6;
wire ap_CS_fsm_state7;
wire ap_CS_fsm_state8;
wire ap_CS_fsm_state9;
wire [31:0] ap_NS_fsm;
wire ap_clk;
wire ap_done;
wire ap_idle;
wire ap_ready;
wire ap_rst;
wire ap_start;
wire [15:0] empty_16_fu_361_p0;
wire [9:0] empty_16_fu_361_p1;
wire [2:0] empty_fu_247_p1;
wire [32:0] grp_fu_227_p0;
wire [32:0] grp_fu_227_p2;
wire [1:0] grp_fu_267_p0;
wire [1:0] grp_fu_267_p2;
wire [24:0] grp_fu_281_p0;
wire [24:0] grp_fu_281_p2;
wire [24:0] grp_fu_350_p1;
wire [24:0] grp_fu_350_p2;
wire [4:0] grp_fu_355_p0;
wire [4:0] grp_fu_355_p2;
wire [17:0] grp_fu_398_p0;
wire [17:0] grp_fu_398_p1;
wire [17:0] grp_fu_398_p2;
wire [24:0] grp_fu_450_p0;
wire [24:0] grp_fu_450_p2;
wire [55:0] grp_fu_514_p0;
wire [55:0] grp_fu_514_p1;
wire [55:0] grp_fu_514_p2;
wire [31:0] grp_fu_535_p2;
wire [31:0] grp_fu_563_p1;
wire [31:0] grp_fu_563_p2;
wire [31:0] grp_fu_571_p1;
wire [31:0] grp_fu_571_p2;
wire [33:0] grp_fu_591_p0;
wire [33:0] grp_fu_591_p1;
wire [33:0] grp_fu_591_p2;
wire [31:0] grp_fu_607_p2;
wire [31:0] grp_fu_647_p1;
wire [31:0] grp_fu_647_p2;
wire [38:0] grp_fu_667_p0;
wire [38:0] grp_fu_667_p1;
wire [38:0] grp_fu_667_p2;
wire [31:0] grp_fu_693_p2;
wire [31:0] grp_fu_725_p2;
wire icmp_ln851_1_fu_520_p2;
wire icmp_ln851_2_fu_677_p2;
wire icmp_ln851_fu_276_p2;
wire [20:0] lhs_V_fu_407_p3;
wire [1:0] \mul_2s_2s_4_1_1_U4.din0 ;
wire [1:0] \mul_2s_2s_4_1_1_U4.din1 ;
wire [3:0] \mul_2s_2s_4_1_1_U4.dout ;
wire [1:0] \mul_2s_2s_4_1_1_U4.top_mul_2s_2s_4_1_1_Multiplier_0_U.a ;
wire [1:0] \mul_2s_2s_4_1_1_U4.top_mul_2s_2s_4_1_1_Multiplier_0_U.b ;
wire [3:0] \mul_2s_2s_4_1_1_U4.top_mul_2s_2s_4_1_1_Multiplier_0_U.p ;
wire [3:0] op_0;
wire [7:0] op_10;
wire [7:0] op_11;
wire [20:0] op_12_V_fu_371_p3;
wire [31:0] op_13_V_fu_488_p3;
wire [3:0] op_14;
wire [7:0] op_16;
wire op_17_V_fu_616_p2;
wire [31:0] op_18;
wire op_19;
wire [3:0] op_2;
wire [31:0] op_3;
wire [31:0] op_30;
wire op_30_ap_vld;
wire [15:0] op_5;
wire [3:0] op_8;
wire overflow_fu_471_p2;
wire p_Result_1_fu_310_p3;
wire p_Result_4_fu_540_p3;
wire p_Result_5_fu_621_p3;
wire p_Result_6_fu_698_p3;
wire p_Result_s_fu_287_p3;
wire [31:0] p_Val2_3_fu_458_p3;
wire [9:0] r_fu_365_p2;
wire [2:0] ret_V_14_fu_251_p2;
wire [1:0] ret_V_15_fu_303_p3;
wire [24:0] ret_V_17_fu_322_p3;
wire [31:0] ret_V_20_fu_552_p3;
wire [31:0] ret_V_24_fu_637_p3;
wire [31:0] ret_V_26_fu_710_p3;
wire [20:0] ret_V_fu_415_p2;
wire [1:0] ret_fu_332_p0;
wire [1:0] ret_fu_332_p1;
wire [3:0] ret_fu_332_p2;
wire [11:0] rhs_1_fu_383_p3;
wire [32:0] rhs_7_fu_580_p3;
wire [37:0] rhs_9_fu_656_p3;
wire [31:0] select_ln384_fu_480_p3;
wire [31:0] select_ln69_fu_717_p3;
wire [24:0] select_ln850_1_fu_317_p3;
wire [31:0] select_ln850_2_fu_547_p3;
wire [31:0] select_ln850_3_fu_631_p3;
wire [31:0] select_ln850_4_fu_705_p3;
wire [1:0] select_ln850_fu_297_p3;
wire [15:0] sext_ln1192_6_fu_390_p1;
wire [3:0] sext_ln1345_fu_329_p1;
wire [7:0] sext_ln703_2_fu_576_p0;
wire [31:0] sext_ln703_3_fu_652_p0;
wire [15:0] sext_ln703_fu_379_p0;
wire [24:0] sext_ln850_fu_273_p1;
wire [47:0] tmp_fu_503_p3;
wire trunc_ln213_1_fu_612_p1;
wire trunc_ln213_fu_338_p1;
wire [1:0] trunc_ln728_1_fu_404_p1;
wire [16:0] trunc_ln728_fu_455_p1;
wire [8:0] trunc_ln851_1_fu_243_p1;
wire [22:0] trunc_ln851_2_fu_496_p1;
wire [7:0] trunc_ln851_3_fu_628_p0;
wire trunc_ln851_3_fu_628_p1;
wire [31:0] trunc_ln851_4_fu_673_p0;
wire [5:0] trunc_ln851_4_fu_673_p1;
wire trunc_ln851_fu_294_p1;
wire xor_ln340_fu_476_p2;
wire xor_ln785_fu_466_p2;


assign _042_ = ap_CS_fsm[12] & icmp_ln851_1_reg_888;
assign _043_ = icmp_ln851_2_reg_997 & ap_CS_fsm[28];
assign _044_ = _046_ & ap_CS_fsm[0];
assign _045_ = ap_start & ap_CS_fsm[0];
assign overflow_fu_471_p2 = xor_ln785_fu_466_p2 & p_Result_8_reg_852;
assign ret_V_fu_415_p2 = { op_12_V_fu_371_p3[20:19], op_5[7:0], 11'h000 } & { ret_reg_795[1:0], 19'h00000 };
assign xor_ln785_fu_466_p2 = ~ p_Result_7_reg_846;
assign op_12_V_fu_371_p3[20:19] = ~ op_5[9:8];
assign _046_ = ~ ap_start;
always @(posedge \add_18ns_18s_18_2_1_U7.top_add_18ns_18s_18_2_1_Adder_5_U.clk )
\add_18ns_18s_18_2_1_U7.top_add_18ns_18s_18_2_1_Adder_5_U.bin_s1  <= _048_;
always @(posedge \add_18ns_18s_18_2_1_U7.top_add_18ns_18s_18_2_1_Adder_5_U.clk )
\add_18ns_18s_18_2_1_U7.top_add_18ns_18s_18_2_1_Adder_5_U.ain_s1  <= _047_;
always @(posedge \add_18ns_18s_18_2_1_U7.top_add_18ns_18s_18_2_1_Adder_5_U.clk )
\add_18ns_18s_18_2_1_U7.top_add_18ns_18s_18_2_1_Adder_5_U.sum_s1  <= _050_;
always @(posedge \add_18ns_18s_18_2_1_U7.top_add_18ns_18s_18_2_1_Adder_5_U.clk )
\add_18ns_18s_18_2_1_U7.top_add_18ns_18s_18_2_1_Adder_5_U.carry_s1  <= _049_;
assign _048_ = \add_18ns_18s_18_2_1_U7.top_add_18ns_18s_18_2_1_Adder_5_U.ce  ? \add_18ns_18s_18_2_1_U7.top_add_18ns_18s_18_2_1_Adder_5_U.b [17:9] : \add_18ns_18s_18_2_1_U7.top_add_18ns_18s_18_2_1_Adder_5_U.bin_s1 ;
assign _047_ = \add_18ns_18s_18_2_1_U7.top_add_18ns_18s_18_2_1_Adder_5_U.ce  ? \add_18ns_18s_18_2_1_U7.top_add_18ns_18s_18_2_1_Adder_5_U.a [17:9] : \add_18ns_18s_18_2_1_U7.top_add_18ns_18s_18_2_1_Adder_5_U.ain_s1 ;
assign _049_ = \add_18ns_18s_18_2_1_U7.top_add_18ns_18s_18_2_1_Adder_5_U.ce  ? \add_18ns_18s_18_2_1_U7.top_add_18ns_18s_18_2_1_Adder_5_U.facout_s1  : \add_18ns_18s_18_2_1_U7.top_add_18ns_18s_18_2_1_Adder_5_U.carry_s1 ;
assign _050_ = \add_18ns_18s_18_2_1_U7.top_add_18ns_18s_18_2_1_Adder_5_U.ce  ? \add_18ns_18s_18_2_1_U7.top_add_18ns_18s_18_2_1_Adder_5_U.fas_s1  : \add_18ns_18s_18_2_1_U7.top_add_18ns_18s_18_2_1_Adder_5_U.sum_s1 ;
assign _051_ = \add_18ns_18s_18_2_1_U7.top_add_18ns_18s_18_2_1_Adder_5_U.u1.a  + \add_18ns_18s_18_2_1_U7.top_add_18ns_18s_18_2_1_Adder_5_U.u1.b ;
assign { \add_18ns_18s_18_2_1_U7.top_add_18ns_18s_18_2_1_Adder_5_U.u1.cout , \add_18ns_18s_18_2_1_U7.top_add_18ns_18s_18_2_1_Adder_5_U.u1.s  } = _051_ + \add_18ns_18s_18_2_1_U7.top_add_18ns_18s_18_2_1_Adder_5_U.u1.cin ;
assign _052_ = \add_18ns_18s_18_2_1_U7.top_add_18ns_18s_18_2_1_Adder_5_U.u2.a  + \add_18ns_18s_18_2_1_U7.top_add_18ns_18s_18_2_1_Adder_5_U.u2.b ;
assign { \add_18ns_18s_18_2_1_U7.top_add_18ns_18s_18_2_1_Adder_5_U.u2.cout , \add_18ns_18s_18_2_1_U7.top_add_18ns_18s_18_2_1_Adder_5_U.u2.s  } = _052_ + \add_18ns_18s_18_2_1_U7.top_add_18ns_18s_18_2_1_Adder_5_U.u2.cin ;
always @(posedge \add_25ns_25s_25_2_1_U5.top_add_25ns_25s_25_2_1_Adder_3_U.clk )
\add_25ns_25s_25_2_1_U5.top_add_25ns_25s_25_2_1_Adder_3_U.bin_s1  <= _054_;
always @(posedge \add_25ns_25s_25_2_1_U5.top_add_25ns_25s_25_2_1_Adder_3_U.clk )
\add_25ns_25s_25_2_1_U5.top_add_25ns_25s_25_2_1_Adder_3_U.ain_s1  <= _053_;
always @(posedge \add_25ns_25s_25_2_1_U5.top_add_25ns_25s_25_2_1_Adder_3_U.clk )
\add_25ns_25s_25_2_1_U5.top_add_25ns_25s_25_2_1_Adder_3_U.sum_s1  <= _056_;
always @(posedge \add_25ns_25s_25_2_1_U5.top_add_25ns_25s_25_2_1_Adder_3_U.clk )
\add_25ns_25s_25_2_1_U5.top_add_25ns_25s_25_2_1_Adder_3_U.carry_s1  <= _055_;
assign _054_ = \add_25ns_25s_25_2_1_U5.top_add_25ns_25s_25_2_1_Adder_3_U.ce  ? \add_25ns_25s_25_2_1_U5.top_add_25ns_25s_25_2_1_Adder_3_U.b [24:12] : \add_25ns_25s_25_2_1_U5.top_add_25ns_25s_25_2_1_Adder_3_U.bin_s1 ;
assign _053_ = \add_25ns_25s_25_2_1_U5.top_add_25ns_25s_25_2_1_Adder_3_U.ce  ? \add_25ns_25s_25_2_1_U5.top_add_25ns_25s_25_2_1_Adder_3_U.a [24:12] : \add_25ns_25s_25_2_1_U5.top_add_25ns_25s_25_2_1_Adder_3_U.ain_s1 ;
assign _055_ = \add_25ns_25s_25_2_1_U5.top_add_25ns_25s_25_2_1_Adder_3_U.ce  ? \add_25ns_25s_25_2_1_U5.top_add_25ns_25s_25_2_1_Adder_3_U.facout_s1  : \add_25ns_25s_25_2_1_U5.top_add_25ns_25s_25_2_1_Adder_3_U.carry_s1 ;
assign _056_ = \add_25ns_25s_25_2_1_U5.top_add_25ns_25s_25_2_1_Adder_3_U.ce  ? \add_25ns_25s_25_2_1_U5.top_add_25ns_25s_25_2_1_Adder_3_U.fas_s1  : \add_25ns_25s_25_2_1_U5.top_add_25ns_25s_25_2_1_Adder_3_U.sum_s1 ;
assign _057_ = \add_25ns_25s_25_2_1_U5.top_add_25ns_25s_25_2_1_Adder_3_U.u1.a  + \add_25ns_25s_25_2_1_U5.top_add_25ns_25s_25_2_1_Adder_3_U.u1.b ;
assign { \add_25ns_25s_25_2_1_U5.top_add_25ns_25s_25_2_1_Adder_3_U.u1.cout , \add_25ns_25s_25_2_1_U5.top_add_25ns_25s_25_2_1_Adder_3_U.u1.s  } = _057_ + \add_25ns_25s_25_2_1_U5.top_add_25ns_25s_25_2_1_Adder_3_U.u1.cin ;
assign _058_ = \add_25ns_25s_25_2_1_U5.top_add_25ns_25s_25_2_1_Adder_3_U.u2.a  + \add_25ns_25s_25_2_1_U5.top_add_25ns_25s_25_2_1_Adder_3_U.u2.b ;
assign { \add_25ns_25s_25_2_1_U5.top_add_25ns_25s_25_2_1_Adder_3_U.u2.cout , \add_25ns_25s_25_2_1_U5.top_add_25ns_25s_25_2_1_Adder_3_U.u2.s  } = _058_ + \add_25ns_25s_25_2_1_U5.top_add_25ns_25s_25_2_1_Adder_3_U.u2.cin ;
always @(posedge \add_25s_25ns_25_2_1_U3.top_add_25s_25ns_25_2_1_Adder_2_U.clk )
\add_25s_25ns_25_2_1_U3.top_add_25s_25ns_25_2_1_Adder_2_U.bin_s1  <= _060_;
always @(posedge \add_25s_25ns_25_2_1_U3.top_add_25s_25ns_25_2_1_Adder_2_U.clk )
\add_25s_25ns_25_2_1_U3.top_add_25s_25ns_25_2_1_Adder_2_U.ain_s1  <= _059_;
always @(posedge \add_25s_25ns_25_2_1_U3.top_add_25s_25ns_25_2_1_Adder_2_U.clk )
\add_25s_25ns_25_2_1_U3.top_add_25s_25ns_25_2_1_Adder_2_U.sum_s1  <= _062_;
always @(posedge \add_25s_25ns_25_2_1_U3.top_add_25s_25ns_25_2_1_Adder_2_U.clk )
\add_25s_25ns_25_2_1_U3.top_add_25s_25ns_25_2_1_Adder_2_U.carry_s1  <= _061_;
assign _060_ = \add_25s_25ns_25_2_1_U3.top_add_25s_25ns_25_2_1_Adder_2_U.ce  ? \add_25s_25ns_25_2_1_U3.top_add_25s_25ns_25_2_1_Adder_2_U.b [24:12] : \add_25s_25ns_25_2_1_U3.top_add_25s_25ns_25_2_1_Adder_2_U.bin_s1 ;
assign _059_ = \add_25s_25ns_25_2_1_U3.top_add_25s_25ns_25_2_1_Adder_2_U.ce  ? \add_25s_25ns_25_2_1_U3.top_add_25s_25ns_25_2_1_Adder_2_U.a [24:12] : \add_25s_25ns_25_2_1_U3.top_add_25s_25ns_25_2_1_Adder_2_U.ain_s1 ;
assign _061_ = \add_25s_25ns_25_2_1_U3.top_add_25s_25ns_25_2_1_Adder_2_U.ce  ? \add_25s_25ns_25_2_1_U3.top_add_25s_25ns_25_2_1_Adder_2_U.facout_s1  : \add_25s_25ns_25_2_1_U3.top_add_25s_25ns_25_2_1_Adder_2_U.carry_s1 ;
assign _062_ = \add_25s_25ns_25_2_1_U3.top_add_25s_25ns_25_2_1_Adder_2_U.ce  ? \add_25s_25ns_25_2_1_U3.top_add_25s_25ns_25_2_1_Adder_2_U.fas_s1  : \add_25s_25ns_25_2_1_U3.top_add_25s_25ns_25_2_1_Adder_2_U.sum_s1 ;
assign _063_ = \add_25s_25ns_25_2_1_U3.top_add_25s_25ns_25_2_1_Adder_2_U.u1.a  + \add_25s_25ns_25_2_1_U3.top_add_25s_25ns_25_2_1_Adder_2_U.u1.b ;
assign { \add_25s_25ns_25_2_1_U3.top_add_25s_25ns_25_2_1_Adder_2_U.u1.cout , \add_25s_25ns_25_2_1_U3.top_add_25s_25ns_25_2_1_Adder_2_U.u1.s  } = _063_ + \add_25s_25ns_25_2_1_U3.top_add_25s_25ns_25_2_1_Adder_2_U.u1.cin ;
assign _064_ = \add_25s_25ns_25_2_1_U3.top_add_25s_25ns_25_2_1_Adder_2_U.u2.a  + \add_25s_25ns_25_2_1_U3.top_add_25s_25ns_25_2_1_Adder_2_U.u2.b ;
assign { \add_25s_25ns_25_2_1_U3.top_add_25s_25ns_25_2_1_Adder_2_U.u2.cout , \add_25s_25ns_25_2_1_U3.top_add_25s_25ns_25_2_1_Adder_2_U.u2.s  } = _064_ + \add_25s_25ns_25_2_1_U3.top_add_25s_25ns_25_2_1_Adder_2_U.u2.cin ;
always @(posedge \add_25s_25ns_25_2_1_U8.top_add_25s_25ns_25_2_1_Adder_2_U.clk )
\add_25s_25ns_25_2_1_U8.top_add_25s_25ns_25_2_1_Adder_2_U.bin_s1  <= _066_;
always @(posedge \add_25s_25ns_25_2_1_U8.top_add_25s_25ns_25_2_1_Adder_2_U.clk )
\add_25s_25ns_25_2_1_U8.top_add_25s_25ns_25_2_1_Adder_2_U.ain_s1  <= _065_;
always @(posedge \add_25s_25ns_25_2_1_U8.top_add_25s_25ns_25_2_1_Adder_2_U.clk )
\add_25s_25ns_25_2_1_U8.top_add_25s_25ns_25_2_1_Adder_2_U.sum_s1  <= _068_;
always @(posedge \add_25s_25ns_25_2_1_U8.top_add_25s_25ns_25_2_1_Adder_2_U.clk )
\add_25s_25ns_25_2_1_U8.top_add_25s_25ns_25_2_1_Adder_2_U.carry_s1  <= _067_;
assign _066_ = \add_25s_25ns_25_2_1_U8.top_add_25s_25ns_25_2_1_Adder_2_U.ce  ? \add_25s_25ns_25_2_1_U8.top_add_25s_25ns_25_2_1_Adder_2_U.b [24:12] : \add_25s_25ns_25_2_1_U8.top_add_25s_25ns_25_2_1_Adder_2_U.bin_s1 ;
assign _065_ = \add_25s_25ns_25_2_1_U8.top_add_25s_25ns_25_2_1_Adder_2_U.ce  ? \add_25s_25ns_25_2_1_U8.top_add_25s_25ns_25_2_1_Adder_2_U.a [24:12] : \add_25s_25ns_25_2_1_U8.top_add_25s_25ns_25_2_1_Adder_2_U.ain_s1 ;
assign _067_ = \add_25s_25ns_25_2_1_U8.top_add_25s_25ns_25_2_1_Adder_2_U.ce  ? \add_25s_25ns_25_2_1_U8.top_add_25s_25ns_25_2_1_Adder_2_U.facout_s1  : \add_25s_25ns_25_2_1_U8.top_add_25s_25ns_25_2_1_Adder_2_U.carry_s1 ;
assign _068_ = \add_25s_25ns_25_2_1_U8.top_add_25s_25ns_25_2_1_Adder_2_U.ce  ? \add_25s_25ns_25_2_1_U8.top_add_25s_25ns_25_2_1_Adder_2_U.fas_s1  : \add_25s_25ns_25_2_1_U8.top_add_25s_25ns_25_2_1_Adder_2_U.sum_s1 ;
assign _069_ = \add_25s_25ns_25_2_1_U8.top_add_25s_25ns_25_2_1_Adder_2_U.u1.a  + \add_25s_25ns_25_2_1_U8.top_add_25s_25ns_25_2_1_Adder_2_U.u1.b ;
assign { \add_25s_25ns_25_2_1_U8.top_add_25s_25ns_25_2_1_Adder_2_U.u1.cout , \add_25s_25ns_25_2_1_U8.top_add_25s_25ns_25_2_1_Adder_2_U.u1.s  } = _069_ + \add_25s_25ns_25_2_1_U8.top_add_25s_25ns_25_2_1_Adder_2_U.u1.cin ;
assign _070_ = \add_25s_25ns_25_2_1_U8.top_add_25s_25ns_25_2_1_Adder_2_U.u2.a  + \add_25s_25ns_25_2_1_U8.top_add_25s_25ns_25_2_1_Adder_2_U.u2.b ;
assign { \add_25s_25ns_25_2_1_U8.top_add_25s_25ns_25_2_1_Adder_2_U.u2.cout , \add_25s_25ns_25_2_1_U8.top_add_25s_25ns_25_2_1_Adder_2_U.u2.s  } = _070_ + \add_25s_25ns_25_2_1_U8.top_add_25s_25ns_25_2_1_Adder_2_U.u2.cin ;
always @(posedge \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.clk )
\add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.bin_s1  <= _072_;
always @(posedge \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.clk )
\add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.ain_s1  <= _071_;
always @(posedge \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.clk )
\add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.sum_s1  <= _074_;
always @(posedge \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.clk )
\add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.carry_s1  <= _073_;
assign _072_ = \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.ce  ? \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.b [1] : \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.bin_s1 ;
assign _071_ = \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.ce  ? \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.a [1] : \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.ain_s1 ;
assign _073_ = \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.ce  ? \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.facout_s1  : \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.carry_s1 ;
assign _074_ = \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.ce  ? \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.fas_s1  : \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.sum_s1 ;
assign _075_ = \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.a  + \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.b ;
assign { \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.cout , \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.s  } = _075_ + \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.cin ;
assign _076_ = \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.a  + \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.b ;
assign { \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.cout , \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.s  } = _076_ + \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.cin ;
always @(posedge \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.clk )
\add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s1  <= _078_;
always @(posedge \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.clk )
\add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s1  <= _077_;
always @(posedge \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.clk )
\add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.sum_s1  <= _080_;
always @(posedge \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.clk )
\add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.carry_s1  <= _079_;
assign _078_ = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.ce  ? \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.b [31:16] : \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s1 ;
assign _077_ = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.ce  ? \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.a [31:16] : \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s1 ;
assign _079_ = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.ce  ? \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.facout_s1  : \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.carry_s1 ;
assign _080_ = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.ce  ? \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s1  : \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.sum_s1 ;
assign _081_ = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.a  + \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.b ;
assign { \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cout , \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.s  } = _081_ + \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cin ;
assign _082_ = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.a  + \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.b ;
assign { \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cout , \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.s  } = _082_ + \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cin ;
always @(posedge \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.clk )
\add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s1  <= _084_;
always @(posedge \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.clk )
\add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s1  <= _083_;
always @(posedge \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.clk )
\add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.sum_s1  <= _086_;
always @(posedge \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.clk )
\add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.carry_s1  <= _085_;
assign _084_ = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.ce  ? \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.b [31:16] : \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s1 ;
assign _083_ = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.ce  ? \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.a [31:16] : \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s1 ;
assign _085_ = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.ce  ? \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.facout_s1  : \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.carry_s1 ;
assign _086_ = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.ce  ? \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s1  : \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.sum_s1 ;
assign _087_ = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.a  + \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.b ;
assign { \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cout , \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.s  } = _087_ + \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cin ;
assign _088_ = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.a  + \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.b ;
assign { \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cout , \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.s  } = _088_ + \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cin ;
always @(posedge \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.clk )
\add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s1  <= _090_;
always @(posedge \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.clk )
\add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s1  <= _089_;
always @(posedge \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.clk )
\add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.sum_s1  <= _092_;
always @(posedge \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.clk )
\add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.carry_s1  <= _091_;
assign _090_ = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.ce  ? \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.b [31:16] : \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s1 ;
assign _089_ = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.ce  ? \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.a [31:16] : \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s1 ;
assign _091_ = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.ce  ? \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.facout_s1  : \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.carry_s1 ;
assign _092_ = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.ce  ? \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s1  : \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.sum_s1 ;
assign _093_ = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.a  + \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.b ;
assign { \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cout , \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.s  } = _093_ + \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cin ;
assign _094_ = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.a  + \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.b ;
assign { \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cout , \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.s  } = _094_ + \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cin ;
always @(posedge \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_7_U.clk )
\add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s1  <= _096_;
always @(posedge \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_7_U.clk )
\add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s1  <= _095_;
always @(posedge \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_7_U.clk )
\add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_7_U.sum_s1  <= _098_;
always @(posedge \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_7_U.clk )
\add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_7_U.carry_s1  <= _097_;
assign _096_ = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_7_U.ce  ? \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_7_U.b [31:16] : \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s1 ;
assign _095_ = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_7_U.ce  ? \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_7_U.a [31:16] : \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s1 ;
assign _097_ = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_7_U.ce  ? \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_7_U.facout_s1  : \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_7_U.carry_s1 ;
assign _098_ = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_7_U.ce  ? \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s1  : \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_7_U.sum_s1 ;
assign _099_ = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.a  + \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.b ;
assign { \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cout , \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.s  } = _099_ + \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cin ;
assign _100_ = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.a  + \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.b ;
assign { \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cout , \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.s  } = _100_ + \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cin ;
always @(posedge \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.clk )
\add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s1  <= _102_;
always @(posedge \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.clk )
\add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s1  <= _101_;
always @(posedge \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.clk )
\add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.sum_s1  <= _104_;
always @(posedge \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.clk )
\add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.carry_s1  <= _103_;
assign _102_ = \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.ce  ? \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.b [31:16] : \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s1 ;
assign _101_ = \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.ce  ? \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.a [31:16] : \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s1 ;
assign _103_ = \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.ce  ? \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.facout_s1  : \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.carry_s1 ;
assign _104_ = \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.ce  ? \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s1  : \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.sum_s1 ;
assign _105_ = \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.a  + \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.b ;
assign { \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cout , \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.s  } = _105_ + \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cin ;
assign _106_ = \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.a  + \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.b ;
assign { \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cout , \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.s  } = _106_ + \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cin ;
always @(posedge \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.clk )
\add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.bin_s1  <= _108_;
always @(posedge \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.clk )
\add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.ain_s1  <= _107_;
always @(posedge \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.clk )
\add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.sum_s1  <= _110_;
always @(posedge \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.clk )
\add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.carry_s1  <= _109_;
assign _108_ = \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.ce  ? \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.b [31:16] : \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.bin_s1 ;
assign _107_ = \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.ce  ? \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.a [31:16] : \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.ain_s1 ;
assign _109_ = \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.ce  ? \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.facout_s1  : \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.carry_s1 ;
assign _110_ = \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.ce  ? \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.fas_s1  : \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.sum_s1 ;
assign _111_ = \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.u1.a  + \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.u1.b ;
assign { \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.u1.cout , \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.u1.s  } = _111_ + \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.u1.cin ;
assign _112_ = \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.u2.a  + \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.u2.b ;
assign { \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.u2.cout , \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.u2.s  } = _112_ + \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.u2.cin ;
always @(posedge \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.clk )
\add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.bin_s1  <= _114_;
always @(posedge \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.clk )
\add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.ain_s1  <= _113_;
always @(posedge \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.clk )
\add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.sum_s1  <= _116_;
always @(posedge \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.clk )
\add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.carry_s1  <= _115_;
assign _114_ = \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.ce  ? \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.b [31:16] : \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.bin_s1 ;
assign _113_ = \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.ce  ? \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.a [31:16] : \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.ain_s1 ;
assign _115_ = \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.ce  ? \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.facout_s1  : \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.carry_s1 ;
assign _116_ = \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.ce  ? \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.fas_s1  : \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.sum_s1 ;
assign _117_ = \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.u1.a  + \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.u1.b ;
assign { \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.u1.cout , \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.u1.s  } = _117_ + \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.u1.cin ;
assign _118_ = \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.u2.a  + \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.u2.b ;
assign { \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.u2.cout , \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.u2.s  } = _118_ + \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.u2.cin ;
always @(posedge \add_33s_33ns_33_2_1_U1.top_add_33s_33ns_33_2_1_Adder_0_U.clk )
\add_33s_33ns_33_2_1_U1.top_add_33s_33ns_33_2_1_Adder_0_U.bin_s1  <= _120_;
always @(posedge \add_33s_33ns_33_2_1_U1.top_add_33s_33ns_33_2_1_Adder_0_U.clk )
\add_33s_33ns_33_2_1_U1.top_add_33s_33ns_33_2_1_Adder_0_U.ain_s1  <= _119_;
always @(posedge \add_33s_33ns_33_2_1_U1.top_add_33s_33ns_33_2_1_Adder_0_U.clk )
\add_33s_33ns_33_2_1_U1.top_add_33s_33ns_33_2_1_Adder_0_U.sum_s1  <= _122_;
always @(posedge \add_33s_33ns_33_2_1_U1.top_add_33s_33ns_33_2_1_Adder_0_U.clk )
\add_33s_33ns_33_2_1_U1.top_add_33s_33ns_33_2_1_Adder_0_U.carry_s1  <= _121_;
assign _120_ = \add_33s_33ns_33_2_1_U1.top_add_33s_33ns_33_2_1_Adder_0_U.ce  ? \add_33s_33ns_33_2_1_U1.top_add_33s_33ns_33_2_1_Adder_0_U.b [32:16] : \add_33s_33ns_33_2_1_U1.top_add_33s_33ns_33_2_1_Adder_0_U.bin_s1 ;
assign _119_ = \add_33s_33ns_33_2_1_U1.top_add_33s_33ns_33_2_1_Adder_0_U.ce  ? \add_33s_33ns_33_2_1_U1.top_add_33s_33ns_33_2_1_Adder_0_U.a [32:16] : \add_33s_33ns_33_2_1_U1.top_add_33s_33ns_33_2_1_Adder_0_U.ain_s1 ;
assign _121_ = \add_33s_33ns_33_2_1_U1.top_add_33s_33ns_33_2_1_Adder_0_U.ce  ? \add_33s_33ns_33_2_1_U1.top_add_33s_33ns_33_2_1_Adder_0_U.facout_s1  : \add_33s_33ns_33_2_1_U1.top_add_33s_33ns_33_2_1_Adder_0_U.carry_s1 ;
assign _122_ = \add_33s_33ns_33_2_1_U1.top_add_33s_33ns_33_2_1_Adder_0_U.ce  ? \add_33s_33ns_33_2_1_U1.top_add_33s_33ns_33_2_1_Adder_0_U.fas_s1  : \add_33s_33ns_33_2_1_U1.top_add_33s_33ns_33_2_1_Adder_0_U.sum_s1 ;
assign _123_ = \add_33s_33ns_33_2_1_U1.top_add_33s_33ns_33_2_1_Adder_0_U.u1.a  + \add_33s_33ns_33_2_1_U1.top_add_33s_33ns_33_2_1_Adder_0_U.u1.b ;
assign { \add_33s_33ns_33_2_1_U1.top_add_33s_33ns_33_2_1_Adder_0_U.u1.cout , \add_33s_33ns_33_2_1_U1.top_add_33s_33ns_33_2_1_Adder_0_U.u1.s  } = _123_ + \add_33s_33ns_33_2_1_U1.top_add_33s_33ns_33_2_1_Adder_0_U.u1.cin ;
assign _124_ = \add_33s_33ns_33_2_1_U1.top_add_33s_33ns_33_2_1_Adder_0_U.u2.a  + \add_33s_33ns_33_2_1_U1.top_add_33s_33ns_33_2_1_Adder_0_U.u2.b ;
assign { \add_33s_33ns_33_2_1_U1.top_add_33s_33ns_33_2_1_Adder_0_U.u2.cout , \add_33s_33ns_33_2_1_U1.top_add_33s_33ns_33_2_1_Adder_0_U.u2.s  } = _124_ + \add_33s_33ns_33_2_1_U1.top_add_33s_33ns_33_2_1_Adder_0_U.u2.cin ;
always @(posedge \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_9_U.clk )
\add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_9_U.bin_s1  <= _126_;
always @(posedge \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_9_U.clk )
\add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_9_U.ain_s1  <= _125_;
always @(posedge \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_9_U.clk )
\add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_9_U.sum_s1  <= _128_;
always @(posedge \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_9_U.clk )
\add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_9_U.carry_s1  <= _127_;
assign _126_ = \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_9_U.ce  ? \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_9_U.b [33:17] : \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_9_U.bin_s1 ;
assign _125_ = \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_9_U.ce  ? \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_9_U.a [33:17] : \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_9_U.ain_s1 ;
assign _127_ = \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_9_U.ce  ? \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_9_U.facout_s1  : \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_9_U.carry_s1 ;
assign _128_ = \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_9_U.ce  ? \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_9_U.fas_s1  : \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_9_U.sum_s1 ;
assign _129_ = \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_9_U.u1.a  + \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_9_U.u1.b ;
assign { \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_9_U.u1.cout , \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_9_U.u1.s  } = _129_ + \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_9_U.u1.cin ;
assign _130_ = \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_9_U.u2.a  + \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_9_U.u2.b ;
assign { \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_9_U.u2.cout , \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_9_U.u2.s  } = _130_ + \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_9_U.u2.cin ;
always @(posedge \add_39s_39s_39_2_1_U16.top_add_39s_39s_39_2_1_Adder_10_U.clk )
\add_39s_39s_39_2_1_U16.top_add_39s_39s_39_2_1_Adder_10_U.bin_s1  <= _132_;
always @(posedge \add_39s_39s_39_2_1_U16.top_add_39s_39s_39_2_1_Adder_10_U.clk )
\add_39s_39s_39_2_1_U16.top_add_39s_39s_39_2_1_Adder_10_U.ain_s1  <= _131_;
always @(posedge \add_39s_39s_39_2_1_U16.top_add_39s_39s_39_2_1_Adder_10_U.clk )
\add_39s_39s_39_2_1_U16.top_add_39s_39s_39_2_1_Adder_10_U.sum_s1  <= _134_;
always @(posedge \add_39s_39s_39_2_1_U16.top_add_39s_39s_39_2_1_Adder_10_U.clk )
\add_39s_39s_39_2_1_U16.top_add_39s_39s_39_2_1_Adder_10_U.carry_s1  <= _133_;
assign _132_ = \add_39s_39s_39_2_1_U16.top_add_39s_39s_39_2_1_Adder_10_U.ce  ? \add_39s_39s_39_2_1_U16.top_add_39s_39s_39_2_1_Adder_10_U.b [38:19] : \add_39s_39s_39_2_1_U16.top_add_39s_39s_39_2_1_Adder_10_U.bin_s1 ;
assign _131_ = \add_39s_39s_39_2_1_U16.top_add_39s_39s_39_2_1_Adder_10_U.ce  ? \add_39s_39s_39_2_1_U16.top_add_39s_39s_39_2_1_Adder_10_U.a [38:19] : \add_39s_39s_39_2_1_U16.top_add_39s_39s_39_2_1_Adder_10_U.ain_s1 ;
assign _133_ = \add_39s_39s_39_2_1_U16.top_add_39s_39s_39_2_1_Adder_10_U.ce  ? \add_39s_39s_39_2_1_U16.top_add_39s_39s_39_2_1_Adder_10_U.facout_s1  : \add_39s_39s_39_2_1_U16.top_add_39s_39s_39_2_1_Adder_10_U.carry_s1 ;
assign _134_ = \add_39s_39s_39_2_1_U16.top_add_39s_39s_39_2_1_Adder_10_U.ce  ? \add_39s_39s_39_2_1_U16.top_add_39s_39s_39_2_1_Adder_10_U.fas_s1  : \add_39s_39s_39_2_1_U16.top_add_39s_39s_39_2_1_Adder_10_U.sum_s1 ;
assign _135_ = \add_39s_39s_39_2_1_U16.top_add_39s_39s_39_2_1_Adder_10_U.u1.a  + \add_39s_39s_39_2_1_U16.top_add_39s_39s_39_2_1_Adder_10_U.u1.b ;
assign { \add_39s_39s_39_2_1_U16.top_add_39s_39s_39_2_1_Adder_10_U.u1.cout , \add_39s_39s_39_2_1_U16.top_add_39s_39s_39_2_1_Adder_10_U.u1.s  } = _135_ + \add_39s_39s_39_2_1_U16.top_add_39s_39s_39_2_1_Adder_10_U.u1.cin ;
assign _136_ = \add_39s_39s_39_2_1_U16.top_add_39s_39s_39_2_1_Adder_10_U.u2.a  + \add_39s_39s_39_2_1_U16.top_add_39s_39s_39_2_1_Adder_10_U.u2.b ;
assign { \add_39s_39s_39_2_1_U16.top_add_39s_39s_39_2_1_Adder_10_U.u2.cout , \add_39s_39s_39_2_1_U16.top_add_39s_39s_39_2_1_Adder_10_U.u2.s  } = _136_ + \add_39s_39s_39_2_1_U16.top_add_39s_39s_39_2_1_Adder_10_U.u2.cin ;
always @(posedge \add_56s_56s_56_2_1_U9.top_add_56s_56s_56_2_1_Adder_6_U.clk )
\add_56s_56s_56_2_1_U9.top_add_56s_56s_56_2_1_Adder_6_U.bin_s1  <= _138_;
always @(posedge \add_56s_56s_56_2_1_U9.top_add_56s_56s_56_2_1_Adder_6_U.clk )
\add_56s_56s_56_2_1_U9.top_add_56s_56s_56_2_1_Adder_6_U.ain_s1  <= _137_;
always @(posedge \add_56s_56s_56_2_1_U9.top_add_56s_56s_56_2_1_Adder_6_U.clk )
\add_56s_56s_56_2_1_U9.top_add_56s_56s_56_2_1_Adder_6_U.sum_s1  <= _140_;
always @(posedge \add_56s_56s_56_2_1_U9.top_add_56s_56s_56_2_1_Adder_6_U.clk )
\add_56s_56s_56_2_1_U9.top_add_56s_56s_56_2_1_Adder_6_U.carry_s1  <= _139_;
assign _138_ = \add_56s_56s_56_2_1_U9.top_add_56s_56s_56_2_1_Adder_6_U.ce  ? \add_56s_56s_56_2_1_U9.top_add_56s_56s_56_2_1_Adder_6_U.b [55:28] : \add_56s_56s_56_2_1_U9.top_add_56s_56s_56_2_1_Adder_6_U.bin_s1 ;
assign _137_ = \add_56s_56s_56_2_1_U9.top_add_56s_56s_56_2_1_Adder_6_U.ce  ? \add_56s_56s_56_2_1_U9.top_add_56s_56s_56_2_1_Adder_6_U.a [55:28] : \add_56s_56s_56_2_1_U9.top_add_56s_56s_56_2_1_Adder_6_U.ain_s1 ;
assign _139_ = \add_56s_56s_56_2_1_U9.top_add_56s_56s_56_2_1_Adder_6_U.ce  ? \add_56s_56s_56_2_1_U9.top_add_56s_56s_56_2_1_Adder_6_U.facout_s1  : \add_56s_56s_56_2_1_U9.top_add_56s_56s_56_2_1_Adder_6_U.carry_s1 ;
assign _140_ = \add_56s_56s_56_2_1_U9.top_add_56s_56s_56_2_1_Adder_6_U.ce  ? \add_56s_56s_56_2_1_U9.top_add_56s_56s_56_2_1_Adder_6_U.fas_s1  : \add_56s_56s_56_2_1_U9.top_add_56s_56s_56_2_1_Adder_6_U.sum_s1 ;
assign _141_ = \add_56s_56s_56_2_1_U9.top_add_56s_56s_56_2_1_Adder_6_U.u1.a  + \add_56s_56s_56_2_1_U9.top_add_56s_56s_56_2_1_Adder_6_U.u1.b ;
assign { \add_56s_56s_56_2_1_U9.top_add_56s_56s_56_2_1_Adder_6_U.u1.cout , \add_56s_56s_56_2_1_U9.top_add_56s_56s_56_2_1_Adder_6_U.u1.s  } = _141_ + \add_56s_56s_56_2_1_U9.top_add_56s_56s_56_2_1_Adder_6_U.u1.cin ;
assign _142_ = \add_56s_56s_56_2_1_U9.top_add_56s_56s_56_2_1_Adder_6_U.u2.a  + \add_56s_56s_56_2_1_U9.top_add_56s_56s_56_2_1_Adder_6_U.u2.b ;
assign { \add_56s_56s_56_2_1_U9.top_add_56s_56s_56_2_1_Adder_6_U.u2.cout , \add_56s_56s_56_2_1_U9.top_add_56s_56s_56_2_1_Adder_6_U.u2.s  } = _142_ + \add_56s_56s_56_2_1_U9.top_add_56s_56s_56_2_1_Adder_6_U.u2.cin ;
always @(posedge \add_5s_5ns_5_2_1_U6.top_add_5s_5ns_5_2_1_Adder_4_U.clk )
\add_5s_5ns_5_2_1_U6.top_add_5s_5ns_5_2_1_Adder_4_U.bin_s1  <= _144_;
always @(posedge \add_5s_5ns_5_2_1_U6.top_add_5s_5ns_5_2_1_Adder_4_U.clk )
\add_5s_5ns_5_2_1_U6.top_add_5s_5ns_5_2_1_Adder_4_U.ain_s1  <= _143_;
always @(posedge \add_5s_5ns_5_2_1_U6.top_add_5s_5ns_5_2_1_Adder_4_U.clk )
\add_5s_5ns_5_2_1_U6.top_add_5s_5ns_5_2_1_Adder_4_U.sum_s1  <= _146_;
always @(posedge \add_5s_5ns_5_2_1_U6.top_add_5s_5ns_5_2_1_Adder_4_U.clk )
\add_5s_5ns_5_2_1_U6.top_add_5s_5ns_5_2_1_Adder_4_U.carry_s1  <= _145_;
assign _144_ = \add_5s_5ns_5_2_1_U6.top_add_5s_5ns_5_2_1_Adder_4_U.ce  ? \add_5s_5ns_5_2_1_U6.top_add_5s_5ns_5_2_1_Adder_4_U.b [4:2] : \add_5s_5ns_5_2_1_U6.top_add_5s_5ns_5_2_1_Adder_4_U.bin_s1 ;
assign _143_ = \add_5s_5ns_5_2_1_U6.top_add_5s_5ns_5_2_1_Adder_4_U.ce  ? \add_5s_5ns_5_2_1_U6.top_add_5s_5ns_5_2_1_Adder_4_U.a [4:2] : \add_5s_5ns_5_2_1_U6.top_add_5s_5ns_5_2_1_Adder_4_U.ain_s1 ;
assign _145_ = \add_5s_5ns_5_2_1_U6.top_add_5s_5ns_5_2_1_Adder_4_U.ce  ? \add_5s_5ns_5_2_1_U6.top_add_5s_5ns_5_2_1_Adder_4_U.facout_s1  : \add_5s_5ns_5_2_1_U6.top_add_5s_5ns_5_2_1_Adder_4_U.carry_s1 ;
assign _146_ = \add_5s_5ns_5_2_1_U6.top_add_5s_5ns_5_2_1_Adder_4_U.ce  ? \add_5s_5ns_5_2_1_U6.top_add_5s_5ns_5_2_1_Adder_4_U.fas_s1  : \add_5s_5ns_5_2_1_U6.top_add_5s_5ns_5_2_1_Adder_4_U.sum_s1 ;
assign _147_ = \add_5s_5ns_5_2_1_U6.top_add_5s_5ns_5_2_1_Adder_4_U.u1.a  + \add_5s_5ns_5_2_1_U6.top_add_5s_5ns_5_2_1_Adder_4_U.u1.b ;
assign { \add_5s_5ns_5_2_1_U6.top_add_5s_5ns_5_2_1_Adder_4_U.u1.cout , \add_5s_5ns_5_2_1_U6.top_add_5s_5ns_5_2_1_Adder_4_U.u1.s  } = _147_ + \add_5s_5ns_5_2_1_U6.top_add_5s_5ns_5_2_1_Adder_4_U.u1.cin ;
assign _148_ = \add_5s_5ns_5_2_1_U6.top_add_5s_5ns_5_2_1_Adder_4_U.u2.a  + \add_5s_5ns_5_2_1_U6.top_add_5s_5ns_5_2_1_Adder_4_U.u2.b ;
assign { \add_5s_5ns_5_2_1_U6.top_add_5s_5ns_5_2_1_Adder_4_U.u2.cout , \add_5s_5ns_5_2_1_U6.top_add_5s_5ns_5_2_1_Adder_4_U.u2.s  } = _148_ + \add_5s_5ns_5_2_1_U6.top_add_5s_5ns_5_2_1_Adder_4_U.u2.cin ;
assign \mul_2s_2s_4_1_1_U4.top_mul_2s_2s_4_1_1_Multiplier_0_U.p  = $signed(\mul_2s_2s_4_1_1_U4.top_mul_2s_2s_4_1_1_Multiplier_0_U.a ) * $signed(\mul_2s_2s_4_1_1_U4.top_mul_2s_2s_4_1_1_Multiplier_0_U.b );
assign _149_ = | trunc_ln851_2_reg_873;
assign _150_ = | op_18[5:0];
assign _151_ = | trunc_ln851_1_reg_745;
always @(posedge ap_clk)
ret_reg_795 <= _034_;
always @(posedge ap_clk)
trunc_ln213_reg_801 <= _038_;
always @(posedge ap_clk)
ret_V_26_reg_1019 <= _031_;
always @(posedge ap_clk)
select_ln69_reg_1024 <= _035_;
always @(posedge ap_clk)
ret_V_22_reg_930 <= _027_;
always @(posedge ap_clk)
ret_V_21_reg_920 <= _026_;
always @(posedge ap_clk)
ret_V_25_reg_1002 <= _030_;
always @(posedge ap_clk)
ret_V_21_cast_reg_1007 <= _025_;
always @(posedge ap_clk)
ret_V_20_reg_910 <= _024_;
always @(posedge ap_clk)
ret_V_19_reg_893 <= _023_;
always @(posedge ap_clk)
ret_V_8_cast_reg_898 <= _032_;
always @(posedge ap_clk)
ret_V_23_reg_950 <= _028_;
always @(posedge ap_clk)
ret_V_19_cast_reg_955 <= _022_;
always @(posedge ap_clk)
ret_V_16_reg_735 <= _019_;
always @(posedge ap_clk)
tmp_1_reg_740 <= _037_;
always @(posedge ap_clk)
trunc_ln851_1_reg_745 <= _039_;
always @(posedge ap_clk)
ret_V_15_reg_785 <= _018_;
always @(posedge ap_clk)
ret_V_17_reg_790 <= _020_;
always @(posedge ap_clk)
ret_V_18_reg_841 <= _021_;
always @(posedge ap_clk)
p_Result_7_reg_846 <= _016_;
always @(posedge ap_clk)
p_Result_8_reg_852 <= _017_;
always @(posedge ap_clk)
op_28_V_reg_982 <= _015_;
always @(posedge ap_clk)
op_17_V_reg_967 <= _013_;
always @(posedge ap_clk)
ret_V_24_reg_972 <= _029_;
always @(posedge ap_clk)
op_13_V_reg_863 <= _011_;
always @(posedge ap_clk)
op_23_V_reg_868 <= _014_;
always @(posedge ap_clk)
trunc_ln851_2_reg_873 <= _040_;
always @(posedge ap_clk)
ret_V_cast_reg_756 <= _033_;
always @(posedge ap_clk)
sext_ln850_reg_763 <= _036_;
always @(posedge ap_clk)
icmp_ln851_reg_770 <= _010_;
always @(posedge ap_clk)
icmp_ln851_2_reg_997 <= _009_;
always @(posedge ap_clk)
icmp_ln851_1_reg_888 <= _008_;
always @(posedge ap_clk)
op_15_V_reg_826 <= _012_;
always @(posedge ap_clk)
add_ln69_reg_831 <= _006_;
always @(posedge ap_clk)
add_ln69_1_reg_836 <= _005_;
always @(posedge ap_clk)
add_ln691_4_reg_1014 <= _003_;
always @(posedge ap_clk)
add_ln691_3_reg_962 <= _002_;
always @(posedge ap_clk)
add_ln691_2_reg_905 <= _001_;
always @(posedge ap_clk)
add_ln691_reg_775 <= _004_;
always @(posedge ap_clk)
add_ln691_1_reg_780 <= _000_;
always @(posedge ap_clk)
ap_CS_fsm <= _007_;
assign _041_ = _045_ ? 2'h2 : 2'h1;
assign _152_ = ap_CS_fsm == 1'h1;
function [31:0] _444_;
input [31:0] a;
input [1023:0] b;
input [31:0] s;
case (s)
32'b00000000000000000000000000000001:
_444_ = b[31:0];
32'b00000000000000000000000000000010:
_444_ = b[63:32];
32'b00000000000000000000000000000100:
_444_ = b[95:64];
32'b00000000000000000000000000001000:
_444_ = b[127:96];
32'b00000000000000000000000000010000:
_444_ = b[159:128];
32'b00000000000000000000000000100000:
_444_ = b[191:160];
32'b00000000000000000000000001000000:
_444_ = b[223:192];
32'b00000000000000000000000010000000:
_444_ = b[255:224];
32'b00000000000000000000000100000000:
_444_ = b[287:256];
32'b00000000000000000000001000000000:
_444_ = b[319:288];
32'b00000000000000000000010000000000:
_444_ = b[351:320];
32'b00000000000000000000100000000000:
_444_ = b[383:352];
32'b00000000000000000001000000000000:
_444_ = b[415:384];
32'b00000000000000000010000000000000:
_444_ = b[447:416];
32'b00000000000000000100000000000000:
_444_ = b[479:448];
32'b00000000000000001000000000000000:
_444_ = b[511:480];
32'b00000000000000010000000000000000:
_444_ = b[543:512];
32'b00000000000000100000000000000000:
_444_ = b[575:544];
32'b00000000000001000000000000000000:
_444_ = b[607:576];
32'b00000000000010000000000000000000:
_444_ = b[639:608];
32'b00000000000100000000000000000000:
_444_ = b[671:640];
32'b00000000001000000000000000000000:
_444_ = b[703:672];
32'b00000000010000000000000000000000:
_444_ = b[735:704];
32'b00000000100000000000000000000000:
_444_ = b[767:736];
32'b00000001000000000000000000000000:
_444_ = b[799:768];
32'b00000010000000000000000000000000:
_444_ = b[831:800];
32'b00000100000000000000000000000000:
_444_ = b[863:832];
32'b00001000000000000000000000000000:
_444_ = b[895:864];
32'b00010000000000000000000000000000:
_444_ = b[927:896];
32'b00100000000000000000000000000000:
_444_ = b[959:928];
32'b01000000000000000000000000000000:
_444_ = b[991:960];
32'b10000000000000000000000000000000:
_444_ = b[1023:992];
32'b00000000000000000000000000000000:
_444_ = a;
default:
_444_ = 32'bx;
endcase
endfunction
assign ap_NS_fsm = _444_(32'hxxxxxxxx, { 30'h00000000, _041_, 992'h00000004000000080000001000000020000000400000008000000100000002000000040000000800000010000000200000004000000080000001000000020000000400000008000000100000002000000040000000800000010000000200000004000000080000001000000020000000400000008000000000000001 }, { _152_, _183_, _182_, _181_, _180_, _179_, _178_, _177_, _176_, _175_, _174_, _173_, _172_, _171_, _170_, _169_, _168_, _167_, _166_, _165_, _164_, _163_, _162_, _161_, _160_, _159_, _158_, _157_, _156_, _155_, _154_, _153_ });
assign _153_ = ap_CS_fsm == 32'd2147483648;
assign _154_ = ap_CS_fsm == 31'h40000000;
assign _155_ = ap_CS_fsm == 30'h20000000;
assign _156_ = ap_CS_fsm == 29'h10000000;
assign _157_ = ap_CS_fsm == 28'h8000000;
assign _158_ = ap_CS_fsm == 27'h4000000;
assign _159_ = ap_CS_fsm == 26'h2000000;
assign _160_ = ap_CS_fsm == 25'h1000000;
assign _161_ = ap_CS_fsm == 24'h800000;
assign _162_ = ap_CS_fsm == 23'h400000;
assign _163_ = ap_CS_fsm == 22'h200000;
assign _164_ = ap_CS_fsm == 21'h100000;
assign _165_ = ap_CS_fsm == 20'h80000;
assign _166_ = ap_CS_fsm == 19'h40000;
assign _167_ = ap_CS_fsm == 18'h20000;
assign _168_ = ap_CS_fsm == 17'h10000;
assign _169_ = ap_CS_fsm == 16'h8000;
assign _170_ = ap_CS_fsm == 15'h4000;
assign _171_ = ap_CS_fsm == 14'h2000;
assign _172_ = ap_CS_fsm == 13'h1000;
assign _173_ = ap_CS_fsm == 12'h800;
assign _174_ = ap_CS_fsm == 11'h400;
assign _175_ = ap_CS_fsm == 10'h200;
assign _176_ = ap_CS_fsm == 9'h100;
assign _177_ = ap_CS_fsm == 8'h80;
assign _178_ = ap_CS_fsm == 7'h40;
assign _179_ = ap_CS_fsm == 6'h20;
assign _180_ = ap_CS_fsm == 5'h10;
assign _181_ = ap_CS_fsm == 4'h8;
assign _182_ = ap_CS_fsm == 3'h4;
assign _183_ = ap_CS_fsm == 2'h2;
assign op_30_ap_vld = ap_CS_fsm[31] ? 1'h1 : 1'h0;
assign ap_idle = _044_ ? 1'h1 : 1'h0;
assign _038_ = ap_CS_fsm[5] ? ret_fu_332_p2[0] : trunc_ln213_reg_801;
assign _034_ = ap_CS_fsm[5] ? ret_fu_332_p2 : ret_reg_795;
assign _035_ = ap_CS_fsm[29] ? select_ln69_fu_717_p3 : select_ln69_reg_1024;
assign _031_ = ap_CS_fsm[29] ? ret_V_26_fu_710_p3 : ret_V_26_reg_1019;
assign _027_ = ap_CS_fsm[17] ? grp_fu_571_p2 : ret_V_22_reg_930;
assign _026_ = ap_CS_fsm[15] ? grp_fu_563_p2 : ret_V_21_reg_920;
assign _025_ = ap_CS_fsm[26] ? grp_fu_667_p2[37:6] : ret_V_21_cast_reg_1007;
assign _030_ = ap_CS_fsm[26] ? grp_fu_667_p2 : ret_V_25_reg_1002;
assign _024_ = ap_CS_fsm[13] ? ret_V_20_fu_552_p3 : ret_V_20_reg_910;
assign _032_ = ap_CS_fsm[10] ? grp_fu_514_p2[54:23] : ret_V_8_cast_reg_898;
assign _023_ = ap_CS_fsm[10] ? grp_fu_514_p2 : ret_V_19_reg_893;
assign _022_ = ap_CS_fsm[19] ? grp_fu_591_p2[32:1] : ret_V_19_cast_reg_955;
assign _028_ = ap_CS_fsm[19] ? grp_fu_591_p2 : ret_V_23_reg_950;
assign _039_ = ap_CS_fsm[1] ? grp_fu_227_p2[8:0] : trunc_ln851_1_reg_745;
assign _037_ = ap_CS_fsm[1] ? grp_fu_227_p2[32:9] : tmp_1_reg_740;
assign _019_ = ap_CS_fsm[1] ? grp_fu_227_p2 : ret_V_16_reg_735;
assign _020_ = ap_CS_fsm[4] ? ret_V_17_fu_322_p3 : ret_V_17_reg_790;
assign _018_ = ap_CS_fsm[4] ? ret_V_15_fu_303_p3 : ret_V_15_reg_785;
assign _017_ = ap_CS_fsm[7] ? grp_fu_398_p2[16] : p_Result_8_reg_852;
assign _016_ = ap_CS_fsm[7] ? grp_fu_398_p2[17] : p_Result_7_reg_846;
assign _021_ = ap_CS_fsm[7] ? grp_fu_398_p2 : ret_V_18_reg_841;
assign _015_ = ap_CS_fsm[24] ? grp_fu_647_p2 : op_28_V_reg_982;
assign _029_ = ap_CS_fsm[22] ? ret_V_24_fu_637_p3 : ret_V_24_reg_972;
assign _013_ = ap_CS_fsm[22] ? op_17_V_fu_616_p2 : op_17_V_reg_967;
assign _040_ = ap_CS_fsm[8] ? op_13_V_fu_488_p3[22:0] : trunc_ln851_2_reg_873;
assign _014_ = ap_CS_fsm[8] ? grp_fu_450_p2 : op_23_V_reg_868;
assign _011_ = ap_CS_fsm[8] ? op_13_V_fu_488_p3 : op_13_V_reg_863;
assign _010_ = ap_CS_fsm[2] ? icmp_ln851_fu_276_p2 : icmp_ln851_reg_770;
assign _036_ = ap_CS_fsm[2] ? { tmp_1_reg_740[23], tmp_1_reg_740 } : sext_ln850_reg_763;
assign _033_ = ap_CS_fsm[2] ? { op_2[2], 1'h1 } : ret_V_cast_reg_756;
assign _009_ = ap_CS_fsm[25] ? icmp_ln851_2_fu_677_p2 : icmp_ln851_2_reg_997;
assign _008_ = ap_CS_fsm[9] ? icmp_ln851_1_fu_520_p2 : icmp_ln851_1_reg_888;
assign _005_ = ap_CS_fsm[6] ? grp_fu_355_p2 : add_ln69_1_reg_836;
assign _006_ = ap_CS_fsm[6] ? grp_fu_350_p2 : add_ln69_reg_831;
assign _012_ = ap_CS_fsm[6] ? ret_V_fu_415_p2[20:19] : op_15_V_reg_826;
assign _003_ = _043_ ? grp_fu_693_p2 : add_ln691_4_reg_1014;
assign _002_ = ap_CS_fsm[21] ? grp_fu_607_p2 : add_ln691_3_reg_962;
assign _001_ = _042_ ? grp_fu_535_p2 : add_ln691_2_reg_905;
assign _000_ = ap_CS_fsm[3] ? grp_fu_281_p2 : add_ln691_1_reg_780;
assign _004_ = ap_CS_fsm[3] ? grp_fu_267_p2 : add_ln691_reg_775;
assign _007_ = ap_rst ? 32'd1 : ap_NS_fsm;
assign icmp_ln851_1_fu_520_p2 = _149_ ? 1'h1 : 1'h0;
assign icmp_ln851_2_fu_677_p2 = _150_ ? 1'h1 : 1'h0;
assign icmp_ln851_fu_276_p2 = _151_ ? 1'h1 : 1'h0;
assign op_13_V_fu_488_p3 = xor_ln340_fu_476_p2 ? select_ln384_fu_480_p3 : { ret_V_18_reg_841[16:0], 15'h0000 };
assign ret_V_15_fu_303_p3 = op_2[3] ? select_ln850_fu_297_p3 : ret_V_cast_reg_756;
assign ret_V_17_fu_322_p3 = ret_V_16_reg_735[32] ? select_ln850_1_fu_317_p3 : sext_ln850_reg_763;
assign ret_V_20_fu_552_p3 = ret_V_19_reg_893[55] ? select_ln850_2_fu_547_p3 : ret_V_8_cast_reg_898;
assign ret_V_24_fu_637_p3 = ret_V_23_reg_950[33] ? select_ln850_3_fu_631_p3 : ret_V_19_cast_reg_955;
assign ret_V_26_fu_710_p3 = ret_V_25_reg_1002[38] ? select_ln850_4_fu_705_p3 : ret_V_21_cast_reg_1007;
assign select_ln384_fu_480_p3 = overflow_fu_471_p2 ? 32'd2147483647 : 32'd2147483648;
assign select_ln69_fu_717_p3 = op_19 ? 32'd4294967295 : 32'd0;
assign select_ln850_1_fu_317_p3 = icmp_ln851_reg_770 ? add_ln691_1_reg_780 : sext_ln850_reg_763;
assign select_ln850_2_fu_547_p3 = icmp_ln851_1_reg_888 ? add_ln691_2_reg_905 : ret_V_8_cast_reg_898;
assign select_ln850_3_fu_631_p3 = op_16[0] ? add_ln691_3_reg_962 : ret_V_19_cast_reg_955;
assign select_ln850_4_fu_705_p3 = icmp_ln851_2_reg_997 ? add_ln691_4_reg_1014 : ret_V_21_cast_reg_1007;
assign select_ln850_fu_297_p3 = op_2[0] ? add_ln691_reg_775 : ret_V_cast_reg_756;
assign op_17_V_fu_616_p2 = trunc_ln213_reg_801 ^ op_10[0];
assign xor_ln340_fu_476_p2 = p_Result_8_reg_852 ^ p_Result_7_reg_846;
assign ap_CS_fsm_state1 = ap_CS_fsm[0];
assign ap_CS_fsm_state10 = ap_CS_fsm[9];
assign ap_CS_fsm_state11 = ap_CS_fsm[10];
assign ap_CS_fsm_state12 = ap_CS_fsm[11];
assign ap_CS_fsm_state13 = ap_CS_fsm[12];
assign ap_CS_fsm_state14 = ap_CS_fsm[13];
assign ap_CS_fsm_state15 = ap_CS_fsm[14];
assign ap_CS_fsm_state16 = ap_CS_fsm[15];
assign ap_CS_fsm_state17 = ap_CS_fsm[16];
assign ap_CS_fsm_state18 = ap_CS_fsm[17];
assign ap_CS_fsm_state19 = ap_CS_fsm[18];
assign ap_CS_fsm_state2 = ap_CS_fsm[1];
assign ap_CS_fsm_state20 = ap_CS_fsm[19];
assign ap_CS_fsm_state21 = ap_CS_fsm[20];
assign ap_CS_fsm_state22 = ap_CS_fsm[21];
assign ap_CS_fsm_state23 = ap_CS_fsm[22];
assign ap_CS_fsm_state24 = ap_CS_fsm[23];
assign ap_CS_fsm_state25 = ap_CS_fsm[24];
assign ap_CS_fsm_state26 = ap_CS_fsm[25];
assign ap_CS_fsm_state27 = ap_CS_fsm[26];
assign ap_CS_fsm_state28 = ap_CS_fsm[27];
assign ap_CS_fsm_state29 = ap_CS_fsm[28];
assign ap_CS_fsm_state3 = ap_CS_fsm[2];
assign ap_CS_fsm_state30 = ap_CS_fsm[29];
assign ap_CS_fsm_state31 = ap_CS_fsm[30];
assign ap_CS_fsm_state32 = ap_CS_fsm[31];
assign ap_CS_fsm_state4 = ap_CS_fsm[3];
assign ap_CS_fsm_state5 = ap_CS_fsm[4];
assign ap_CS_fsm_state6 = ap_CS_fsm[5];
assign ap_CS_fsm_state7 = ap_CS_fsm[6];
assign ap_CS_fsm_state8 = ap_CS_fsm[7];
assign ap_CS_fsm_state9 = ap_CS_fsm[8];
assign ap_done = op_30_ap_vld;
assign ap_ready = op_30_ap_vld;
assign empty_16_fu_361_p0 = op_5;
assign empty_16_fu_361_p1 = op_5[9:0];
assign empty_fu_247_p1 = op_2[2:0];
assign grp_fu_227_p0 = { op_3[31], op_3 };
assign grp_fu_267_p0 = { op_2[2], 1'h1 };
assign grp_fu_281_p0 = { tmp_1_reg_740[23], tmp_1_reg_740 };
assign grp_fu_350_p1 = { op_11[7], op_11[7], op_11[7], op_11[7], op_11[7], op_11[7], op_11[7], op_11[7], op_11[7], op_11[7], op_11[7], op_11[7], op_11[7], op_11[7], op_11[7], op_11[7], op_11[7], op_11 };
assign grp_fu_355_p0 = { op_8[3], op_8 };
assign grp_fu_398_p0 = { 2'h0, ret_reg_795[3], ret_reg_795[3], ret_reg_795[3], ret_reg_795[3], ret_reg_795, 8'h00 };
assign grp_fu_398_p1 = { op_5[15], op_5[15], op_5 };
assign grp_fu_450_p0 = { add_ln69_1_reg_836[4], add_ln69_1_reg_836[4], add_ln69_1_reg_836[4], add_ln69_1_reg_836[4], add_ln69_1_reg_836[4], add_ln69_1_reg_836[4], add_ln69_1_reg_836[4], add_ln69_1_reg_836[4], add_ln69_1_reg_836[4], add_ln69_1_reg_836[4], add_ln69_1_reg_836[4], add_ln69_1_reg_836[4], add_ln69_1_reg_836[4], add_ln69_1_reg_836[4], add_ln69_1_reg_836[4], add_ln69_1_reg_836[4], add_ln69_1_reg_836[4], add_ln69_1_reg_836[4], add_ln69_1_reg_836[4], add_ln69_1_reg_836[4], add_ln69_1_reg_836 };
assign grp_fu_514_p0 = { op_23_V_reg_868[24], op_23_V_reg_868[24], op_23_V_reg_868[24], op_23_V_reg_868[24], op_23_V_reg_868[24], op_23_V_reg_868[24], op_23_V_reg_868[24], op_23_V_reg_868[24], op_23_V_reg_868, 23'h000000 };
assign grp_fu_514_p1 = { op_13_V_reg_863[31], op_13_V_reg_863[31], op_13_V_reg_863[31], op_13_V_reg_863[31], op_13_V_reg_863[31], op_13_V_reg_863[31], op_13_V_reg_863[31], op_13_V_reg_863[31], op_13_V_reg_863[31], op_13_V_reg_863[31], op_13_V_reg_863[31], op_13_V_reg_863[31], op_13_V_reg_863[31], op_13_V_reg_863[31], op_13_V_reg_863[31], op_13_V_reg_863[31], op_13_V_reg_863[31], op_13_V_reg_863[31], op_13_V_reg_863[31], op_13_V_reg_863[31], op_13_V_reg_863[31], op_13_V_reg_863[31], op_13_V_reg_863[31], op_13_V_reg_863[31], op_13_V_reg_863 };
assign grp_fu_563_p1 = { op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14 };
assign grp_fu_571_p1 = { op_15_V_reg_826[1], op_15_V_reg_826[1], op_15_V_reg_826[1], op_15_V_reg_826[1], op_15_V_reg_826[1], op_15_V_reg_826[1], op_15_V_reg_826[1], op_15_V_reg_826[1], op_15_V_reg_826[1], op_15_V_reg_826[1], op_15_V_reg_826[1], op_15_V_reg_826[1], op_15_V_reg_826[1], op_15_V_reg_826[1], op_15_V_reg_826[1], op_15_V_reg_826[1], op_15_V_reg_826[1], op_15_V_reg_826[1], op_15_V_reg_826[1], op_15_V_reg_826[1], op_15_V_reg_826[1], op_15_V_reg_826[1], op_15_V_reg_826[1], op_15_V_reg_826[1], op_15_V_reg_826[1], op_15_V_reg_826[1], op_15_V_reg_826[1], op_15_V_reg_826[1], op_15_V_reg_826[1], op_15_V_reg_826[1], op_15_V_reg_826 };
assign grp_fu_591_p0 = { ret_V_22_reg_930[31], ret_V_22_reg_930, 1'h0 };
assign grp_fu_591_p1 = { op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16 };
assign grp_fu_647_p1 = { 31'h00000000, op_17_V_reg_967 };
assign grp_fu_667_p0 = { op_28_V_reg_982[31], op_28_V_reg_982, 6'h00 };
assign grp_fu_667_p1 = { op_18[31], op_18[31], op_18[31], op_18[31], op_18[31], op_18[31], op_18[31], op_18 };
assign lhs_V_fu_407_p3 = { ret_reg_795[1:0], 19'h00000 };
assign op_12_V_fu_371_p3[18:0] = { op_5[7:0], 11'h000 };
assign op_30 = grp_fu_725_p2;
assign p_Result_1_fu_310_p3 = ret_V_16_reg_735[32];
assign p_Result_4_fu_540_p3 = ret_V_19_reg_893[55];
assign p_Result_5_fu_621_p3 = ret_V_23_reg_950[33];
assign p_Result_6_fu_698_p3 = ret_V_25_reg_1002[38];
assign p_Result_s_fu_287_p3 = op_2[3];
assign p_Val2_3_fu_458_p3 = { ret_V_18_reg_841[16:0], 15'h0000 };
assign r_fu_365_p2 = { op_12_V_fu_371_p3[20:19], op_5[7:0] };
assign ret_V_14_fu_251_p2 = { op_2[2], 1'h1, op_2[0] };
assign ret_fu_332_p0 = ret_V_15_reg_785;
assign ret_fu_332_p1 = ret_V_15_reg_785;
assign rhs_1_fu_383_p3 = { ret_reg_795, 8'h00 };
assign rhs_7_fu_580_p3 = { ret_V_22_reg_930, 1'h0 };
assign rhs_9_fu_656_p3 = { op_28_V_reg_982, 6'h00 };
assign sext_ln1192_6_fu_390_p1 = { ret_reg_795[3], ret_reg_795[3], ret_reg_795[3], ret_reg_795[3], ret_reg_795, 8'h00 };
assign sext_ln1345_fu_329_p1 = { ret_V_15_reg_785[1], ret_V_15_reg_785[1], ret_V_15_reg_785 };
assign sext_ln703_2_fu_576_p0 = op_16;
assign sext_ln703_3_fu_652_p0 = op_18;
assign sext_ln703_fu_379_p0 = op_5;
assign sext_ln850_fu_273_p1 = { tmp_1_reg_740[23], tmp_1_reg_740 };
assign tmp_fu_503_p3 = { op_23_V_reg_868, 23'h000000 };
assign trunc_ln213_1_fu_612_p1 = op_10[0];
assign trunc_ln213_fu_338_p1 = ret_fu_332_p2[0];
assign trunc_ln728_1_fu_404_p1 = ret_reg_795[1:0];
assign trunc_ln728_fu_455_p1 = ret_V_18_reg_841[16:0];
assign trunc_ln851_1_fu_243_p1 = grp_fu_227_p2[8:0];
assign trunc_ln851_2_fu_496_p1 = op_13_V_fu_488_p3[22:0];
assign trunc_ln851_3_fu_628_p0 = op_16;
assign trunc_ln851_3_fu_628_p1 = op_16[0];
assign trunc_ln851_4_fu_673_p0 = op_18;
assign trunc_ln851_4_fu_673_p1 = op_18[5:0];
assign trunc_ln851_fu_294_p1 = op_2[0];
assign \mul_2s_2s_4_1_1_U4.top_mul_2s_2s_4_1_1_Multiplier_0_U.a  = \mul_2s_2s_4_1_1_U4.din0 ;
assign \mul_2s_2s_4_1_1_U4.top_mul_2s_2s_4_1_1_Multiplier_0_U.b  = \mul_2s_2s_4_1_1_U4.din1 ;
assign \mul_2s_2s_4_1_1_U4.dout  = \mul_2s_2s_4_1_1_U4.top_mul_2s_2s_4_1_1_Multiplier_0_U.p ;
assign \mul_2s_2s_4_1_1_U4.din0  = ret_V_15_reg_785;
assign \mul_2s_2s_4_1_1_U4.din1  = ret_V_15_reg_785;
assign ret_fu_332_p2 = \mul_2s_2s_4_1_1_U4.dout ;
assign \add_5s_5ns_5_2_1_U6.top_add_5s_5ns_5_2_1_Adder_4_U.ain_s0  = \add_5s_5ns_5_2_1_U6.top_add_5s_5ns_5_2_1_Adder_4_U.a ;
assign \add_5s_5ns_5_2_1_U6.top_add_5s_5ns_5_2_1_Adder_4_U.bin_s0  = \add_5s_5ns_5_2_1_U6.top_add_5s_5ns_5_2_1_Adder_4_U.b ;
assign \add_5s_5ns_5_2_1_U6.top_add_5s_5ns_5_2_1_Adder_4_U.s  = { \add_5s_5ns_5_2_1_U6.top_add_5s_5ns_5_2_1_Adder_4_U.fas_s2 , \add_5s_5ns_5_2_1_U6.top_add_5s_5ns_5_2_1_Adder_4_U.sum_s1  };
assign \add_5s_5ns_5_2_1_U6.top_add_5s_5ns_5_2_1_Adder_4_U.u2.a  = \add_5s_5ns_5_2_1_U6.top_add_5s_5ns_5_2_1_Adder_4_U.ain_s1 ;
assign \add_5s_5ns_5_2_1_U6.top_add_5s_5ns_5_2_1_Adder_4_U.u2.b  = \add_5s_5ns_5_2_1_U6.top_add_5s_5ns_5_2_1_Adder_4_U.bin_s1 ;
assign \add_5s_5ns_5_2_1_U6.top_add_5s_5ns_5_2_1_Adder_4_U.u2.cin  = \add_5s_5ns_5_2_1_U6.top_add_5s_5ns_5_2_1_Adder_4_U.carry_s1 ;
assign \add_5s_5ns_5_2_1_U6.top_add_5s_5ns_5_2_1_Adder_4_U.facout_s2  = \add_5s_5ns_5_2_1_U6.top_add_5s_5ns_5_2_1_Adder_4_U.u2.cout ;
assign \add_5s_5ns_5_2_1_U6.top_add_5s_5ns_5_2_1_Adder_4_U.fas_s2  = \add_5s_5ns_5_2_1_U6.top_add_5s_5ns_5_2_1_Adder_4_U.u2.s ;
assign \add_5s_5ns_5_2_1_U6.top_add_5s_5ns_5_2_1_Adder_4_U.u1.a  = \add_5s_5ns_5_2_1_U6.top_add_5s_5ns_5_2_1_Adder_4_U.a [1:0];
assign \add_5s_5ns_5_2_1_U6.top_add_5s_5ns_5_2_1_Adder_4_U.u1.b  = \add_5s_5ns_5_2_1_U6.top_add_5s_5ns_5_2_1_Adder_4_U.b [1:0];
assign \add_5s_5ns_5_2_1_U6.top_add_5s_5ns_5_2_1_Adder_4_U.u1.cin  = 1'h0;
assign \add_5s_5ns_5_2_1_U6.top_add_5s_5ns_5_2_1_Adder_4_U.facout_s1  = \add_5s_5ns_5_2_1_U6.top_add_5s_5ns_5_2_1_Adder_4_U.u1.cout ;
assign \add_5s_5ns_5_2_1_U6.top_add_5s_5ns_5_2_1_Adder_4_U.fas_s1  = \add_5s_5ns_5_2_1_U6.top_add_5s_5ns_5_2_1_Adder_4_U.u1.s ;
assign \add_5s_5ns_5_2_1_U6.top_add_5s_5ns_5_2_1_Adder_4_U.a  = \add_5s_5ns_5_2_1_U6.din0 ;
assign \add_5s_5ns_5_2_1_U6.top_add_5s_5ns_5_2_1_Adder_4_U.b  = \add_5s_5ns_5_2_1_U6.din1 ;
assign \add_5s_5ns_5_2_1_U6.top_add_5s_5ns_5_2_1_Adder_4_U.ce  = \add_5s_5ns_5_2_1_U6.ce ;
assign \add_5s_5ns_5_2_1_U6.top_add_5s_5ns_5_2_1_Adder_4_U.clk  = \add_5s_5ns_5_2_1_U6.clk ;
assign \add_5s_5ns_5_2_1_U6.top_add_5s_5ns_5_2_1_Adder_4_U.reset  = \add_5s_5ns_5_2_1_U6.reset ;
assign \add_5s_5ns_5_2_1_U6.dout  = \add_5s_5ns_5_2_1_U6.top_add_5s_5ns_5_2_1_Adder_4_U.s ;
assign \add_5s_5ns_5_2_1_U6.ce  = 1'h1;
assign \add_5s_5ns_5_2_1_U6.clk  = ap_clk;
assign \add_5s_5ns_5_2_1_U6.din0  = { op_8[3], op_8 };
assign \add_5s_5ns_5_2_1_U6.din1  = 5'h01;
assign grp_fu_355_p2 = \add_5s_5ns_5_2_1_U6.dout ;
assign \add_5s_5ns_5_2_1_U6.reset  = ap_rst;
assign \add_56s_56s_56_2_1_U9.top_add_56s_56s_56_2_1_Adder_6_U.ain_s0  = \add_56s_56s_56_2_1_U9.top_add_56s_56s_56_2_1_Adder_6_U.a ;
assign \add_56s_56s_56_2_1_U9.top_add_56s_56s_56_2_1_Adder_6_U.bin_s0  = \add_56s_56s_56_2_1_U9.top_add_56s_56s_56_2_1_Adder_6_U.b ;
assign \add_56s_56s_56_2_1_U9.top_add_56s_56s_56_2_1_Adder_6_U.s  = { \add_56s_56s_56_2_1_U9.top_add_56s_56s_56_2_1_Adder_6_U.fas_s2 , \add_56s_56s_56_2_1_U9.top_add_56s_56s_56_2_1_Adder_6_U.sum_s1  };
assign \add_56s_56s_56_2_1_U9.top_add_56s_56s_56_2_1_Adder_6_U.u2.a  = \add_56s_56s_56_2_1_U9.top_add_56s_56s_56_2_1_Adder_6_U.ain_s1 ;
assign \add_56s_56s_56_2_1_U9.top_add_56s_56s_56_2_1_Adder_6_U.u2.b  = \add_56s_56s_56_2_1_U9.top_add_56s_56s_56_2_1_Adder_6_U.bin_s1 ;
assign \add_56s_56s_56_2_1_U9.top_add_56s_56s_56_2_1_Adder_6_U.u2.cin  = \add_56s_56s_56_2_1_U9.top_add_56s_56s_56_2_1_Adder_6_U.carry_s1 ;
assign \add_56s_56s_56_2_1_U9.top_add_56s_56s_56_2_1_Adder_6_U.facout_s2  = \add_56s_56s_56_2_1_U9.top_add_56s_56s_56_2_1_Adder_6_U.u2.cout ;
assign \add_56s_56s_56_2_1_U9.top_add_56s_56s_56_2_1_Adder_6_U.fas_s2  = \add_56s_56s_56_2_1_U9.top_add_56s_56s_56_2_1_Adder_6_U.u2.s ;
assign \add_56s_56s_56_2_1_U9.top_add_56s_56s_56_2_1_Adder_6_U.u1.a  = \add_56s_56s_56_2_1_U9.top_add_56s_56s_56_2_1_Adder_6_U.a [27:0];
assign \add_56s_56s_56_2_1_U9.top_add_56s_56s_56_2_1_Adder_6_U.u1.b  = \add_56s_56s_56_2_1_U9.top_add_56s_56s_56_2_1_Adder_6_U.b [27:0];
assign \add_56s_56s_56_2_1_U9.top_add_56s_56s_56_2_1_Adder_6_U.u1.cin  = 1'h0;
assign \add_56s_56s_56_2_1_U9.top_add_56s_56s_56_2_1_Adder_6_U.facout_s1  = \add_56s_56s_56_2_1_U9.top_add_56s_56s_56_2_1_Adder_6_U.u1.cout ;
assign \add_56s_56s_56_2_1_U9.top_add_56s_56s_56_2_1_Adder_6_U.fas_s1  = \add_56s_56s_56_2_1_U9.top_add_56s_56s_56_2_1_Adder_6_U.u1.s ;
assign \add_56s_56s_56_2_1_U9.top_add_56s_56s_56_2_1_Adder_6_U.a  = \add_56s_56s_56_2_1_U9.din0 ;
assign \add_56s_56s_56_2_1_U9.top_add_56s_56s_56_2_1_Adder_6_U.b  = \add_56s_56s_56_2_1_U9.din1 ;
assign \add_56s_56s_56_2_1_U9.top_add_56s_56s_56_2_1_Adder_6_U.ce  = \add_56s_56s_56_2_1_U9.ce ;
assign \add_56s_56s_56_2_1_U9.top_add_56s_56s_56_2_1_Adder_6_U.clk  = \add_56s_56s_56_2_1_U9.clk ;
assign \add_56s_56s_56_2_1_U9.top_add_56s_56s_56_2_1_Adder_6_U.reset  = \add_56s_56s_56_2_1_U9.reset ;
assign \add_56s_56s_56_2_1_U9.dout  = \add_56s_56s_56_2_1_U9.top_add_56s_56s_56_2_1_Adder_6_U.s ;
assign \add_56s_56s_56_2_1_U9.ce  = 1'h1;
assign \add_56s_56s_56_2_1_U9.clk  = ap_clk;
assign \add_56s_56s_56_2_1_U9.din0  = { op_23_V_reg_868[24], op_23_V_reg_868[24], op_23_V_reg_868[24], op_23_V_reg_868[24], op_23_V_reg_868[24], op_23_V_reg_868[24], op_23_V_reg_868[24], op_23_V_reg_868[24], op_23_V_reg_868, 23'h000000 };
assign \add_56s_56s_56_2_1_U9.din1  = { op_13_V_reg_863[31], op_13_V_reg_863[31], op_13_V_reg_863[31], op_13_V_reg_863[31], op_13_V_reg_863[31], op_13_V_reg_863[31], op_13_V_reg_863[31], op_13_V_reg_863[31], op_13_V_reg_863[31], op_13_V_reg_863[31], op_13_V_reg_863[31], op_13_V_reg_863[31], op_13_V_reg_863[31], op_13_V_reg_863[31], op_13_V_reg_863[31], op_13_V_reg_863[31], op_13_V_reg_863[31], op_13_V_reg_863[31], op_13_V_reg_863[31], op_13_V_reg_863[31], op_13_V_reg_863[31], op_13_V_reg_863[31], op_13_V_reg_863[31], op_13_V_reg_863[31], op_13_V_reg_863 };
assign grp_fu_514_p2 = \add_56s_56s_56_2_1_U9.dout ;
assign \add_56s_56s_56_2_1_U9.reset  = ap_rst;
assign \add_39s_39s_39_2_1_U16.top_add_39s_39s_39_2_1_Adder_10_U.ain_s0  = \add_39s_39s_39_2_1_U16.top_add_39s_39s_39_2_1_Adder_10_U.a ;
assign \add_39s_39s_39_2_1_U16.top_add_39s_39s_39_2_1_Adder_10_U.bin_s0  = \add_39s_39s_39_2_1_U16.top_add_39s_39s_39_2_1_Adder_10_U.b ;
assign \add_39s_39s_39_2_1_U16.top_add_39s_39s_39_2_1_Adder_10_U.s  = { \add_39s_39s_39_2_1_U16.top_add_39s_39s_39_2_1_Adder_10_U.fas_s2 , \add_39s_39s_39_2_1_U16.top_add_39s_39s_39_2_1_Adder_10_U.sum_s1  };
assign \add_39s_39s_39_2_1_U16.top_add_39s_39s_39_2_1_Adder_10_U.u2.a  = \add_39s_39s_39_2_1_U16.top_add_39s_39s_39_2_1_Adder_10_U.ain_s1 ;
assign \add_39s_39s_39_2_1_U16.top_add_39s_39s_39_2_1_Adder_10_U.u2.b  = \add_39s_39s_39_2_1_U16.top_add_39s_39s_39_2_1_Adder_10_U.bin_s1 ;
assign \add_39s_39s_39_2_1_U16.top_add_39s_39s_39_2_1_Adder_10_U.u2.cin  = \add_39s_39s_39_2_1_U16.top_add_39s_39s_39_2_1_Adder_10_U.carry_s1 ;
assign \add_39s_39s_39_2_1_U16.top_add_39s_39s_39_2_1_Adder_10_U.facout_s2  = \add_39s_39s_39_2_1_U16.top_add_39s_39s_39_2_1_Adder_10_U.u2.cout ;
assign \add_39s_39s_39_2_1_U16.top_add_39s_39s_39_2_1_Adder_10_U.fas_s2  = \add_39s_39s_39_2_1_U16.top_add_39s_39s_39_2_1_Adder_10_U.u2.s ;
assign \add_39s_39s_39_2_1_U16.top_add_39s_39s_39_2_1_Adder_10_U.u1.a  = \add_39s_39s_39_2_1_U16.top_add_39s_39s_39_2_1_Adder_10_U.a [18:0];
assign \add_39s_39s_39_2_1_U16.top_add_39s_39s_39_2_1_Adder_10_U.u1.b  = \add_39s_39s_39_2_1_U16.top_add_39s_39s_39_2_1_Adder_10_U.b [18:0];
assign \add_39s_39s_39_2_1_U16.top_add_39s_39s_39_2_1_Adder_10_U.u1.cin  = 1'h0;
assign \add_39s_39s_39_2_1_U16.top_add_39s_39s_39_2_1_Adder_10_U.facout_s1  = \add_39s_39s_39_2_1_U16.top_add_39s_39s_39_2_1_Adder_10_U.u1.cout ;
assign \add_39s_39s_39_2_1_U16.top_add_39s_39s_39_2_1_Adder_10_U.fas_s1  = \add_39s_39s_39_2_1_U16.top_add_39s_39s_39_2_1_Adder_10_U.u1.s ;
assign \add_39s_39s_39_2_1_U16.top_add_39s_39s_39_2_1_Adder_10_U.a  = \add_39s_39s_39_2_1_U16.din0 ;
assign \add_39s_39s_39_2_1_U16.top_add_39s_39s_39_2_1_Adder_10_U.b  = \add_39s_39s_39_2_1_U16.din1 ;
assign \add_39s_39s_39_2_1_U16.top_add_39s_39s_39_2_1_Adder_10_U.ce  = \add_39s_39s_39_2_1_U16.ce ;
assign \add_39s_39s_39_2_1_U16.top_add_39s_39s_39_2_1_Adder_10_U.clk  = \add_39s_39s_39_2_1_U16.clk ;
assign \add_39s_39s_39_2_1_U16.top_add_39s_39s_39_2_1_Adder_10_U.reset  = \add_39s_39s_39_2_1_U16.reset ;
assign \add_39s_39s_39_2_1_U16.dout  = \add_39s_39s_39_2_1_U16.top_add_39s_39s_39_2_1_Adder_10_U.s ;
assign \add_39s_39s_39_2_1_U16.ce  = 1'h1;
assign \add_39s_39s_39_2_1_U16.clk  = ap_clk;
assign \add_39s_39s_39_2_1_U16.din0  = { op_28_V_reg_982[31], op_28_V_reg_982, 6'h00 };
assign \add_39s_39s_39_2_1_U16.din1  = { op_18[31], op_18[31], op_18[31], op_18[31], op_18[31], op_18[31], op_18[31], op_18 };
assign grp_fu_667_p2 = \add_39s_39s_39_2_1_U16.dout ;
assign \add_39s_39s_39_2_1_U16.reset  = ap_rst;
assign \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_9_U.ain_s0  = \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_9_U.a ;
assign \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_9_U.bin_s0  = \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_9_U.b ;
assign \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_9_U.s  = { \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_9_U.fas_s2 , \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_9_U.sum_s1  };
assign \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_9_U.u2.a  = \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_9_U.ain_s1 ;
assign \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_9_U.u2.b  = \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_9_U.bin_s1 ;
assign \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_9_U.u2.cin  = \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_9_U.carry_s1 ;
assign \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_9_U.facout_s2  = \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_9_U.u2.cout ;
assign \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_9_U.fas_s2  = \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_9_U.u2.s ;
assign \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_9_U.u1.a  = \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_9_U.a [16:0];
assign \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_9_U.u1.b  = \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_9_U.b [16:0];
assign \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_9_U.u1.cin  = 1'h0;
assign \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_9_U.facout_s1  = \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_9_U.u1.cout ;
assign \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_9_U.fas_s1  = \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_9_U.u1.s ;
assign \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_9_U.a  = \add_34s_34s_34_2_1_U13.din0 ;
assign \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_9_U.b  = \add_34s_34s_34_2_1_U13.din1 ;
assign \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_9_U.ce  = \add_34s_34s_34_2_1_U13.ce ;
assign \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_9_U.clk  = \add_34s_34s_34_2_1_U13.clk ;
assign \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_9_U.reset  = \add_34s_34s_34_2_1_U13.reset ;
assign \add_34s_34s_34_2_1_U13.dout  = \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_9_U.s ;
assign \add_34s_34s_34_2_1_U13.ce  = 1'h1;
assign \add_34s_34s_34_2_1_U13.clk  = ap_clk;
assign \add_34s_34s_34_2_1_U13.din0  = { ret_V_22_reg_930[31], ret_V_22_reg_930, 1'h0 };
assign \add_34s_34s_34_2_1_U13.din1  = { op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16 };
assign grp_fu_591_p2 = \add_34s_34s_34_2_1_U13.dout ;
assign \add_34s_34s_34_2_1_U13.reset  = ap_rst;
assign \add_33s_33ns_33_2_1_U1.top_add_33s_33ns_33_2_1_Adder_0_U.ain_s0  = \add_33s_33ns_33_2_1_U1.top_add_33s_33ns_33_2_1_Adder_0_U.a ;
assign \add_33s_33ns_33_2_1_U1.top_add_33s_33ns_33_2_1_Adder_0_U.bin_s0  = \add_33s_33ns_33_2_1_U1.top_add_33s_33ns_33_2_1_Adder_0_U.b ;
assign \add_33s_33ns_33_2_1_U1.top_add_33s_33ns_33_2_1_Adder_0_U.s  = { \add_33s_33ns_33_2_1_U1.top_add_33s_33ns_33_2_1_Adder_0_U.fas_s2 , \add_33s_33ns_33_2_1_U1.top_add_33s_33ns_33_2_1_Adder_0_U.sum_s1  };
assign \add_33s_33ns_33_2_1_U1.top_add_33s_33ns_33_2_1_Adder_0_U.u2.a  = \add_33s_33ns_33_2_1_U1.top_add_33s_33ns_33_2_1_Adder_0_U.ain_s1 ;
assign \add_33s_33ns_33_2_1_U1.top_add_33s_33ns_33_2_1_Adder_0_U.u2.b  = \add_33s_33ns_33_2_1_U1.top_add_33s_33ns_33_2_1_Adder_0_U.bin_s1 ;
assign \add_33s_33ns_33_2_1_U1.top_add_33s_33ns_33_2_1_Adder_0_U.u2.cin  = \add_33s_33ns_33_2_1_U1.top_add_33s_33ns_33_2_1_Adder_0_U.carry_s1 ;
assign \add_33s_33ns_33_2_1_U1.top_add_33s_33ns_33_2_1_Adder_0_U.facout_s2  = \add_33s_33ns_33_2_1_U1.top_add_33s_33ns_33_2_1_Adder_0_U.u2.cout ;
assign \add_33s_33ns_33_2_1_U1.top_add_33s_33ns_33_2_1_Adder_0_U.fas_s2  = \add_33s_33ns_33_2_1_U1.top_add_33s_33ns_33_2_1_Adder_0_U.u2.s ;
assign \add_33s_33ns_33_2_1_U1.top_add_33s_33ns_33_2_1_Adder_0_U.u1.a  = \add_33s_33ns_33_2_1_U1.top_add_33s_33ns_33_2_1_Adder_0_U.a [15:0];
assign \add_33s_33ns_33_2_1_U1.top_add_33s_33ns_33_2_1_Adder_0_U.u1.b  = \add_33s_33ns_33_2_1_U1.top_add_33s_33ns_33_2_1_Adder_0_U.b [15:0];
assign \add_33s_33ns_33_2_1_U1.top_add_33s_33ns_33_2_1_Adder_0_U.u1.cin  = 1'h0;
assign \add_33s_33ns_33_2_1_U1.top_add_33s_33ns_33_2_1_Adder_0_U.facout_s1  = \add_33s_33ns_33_2_1_U1.top_add_33s_33ns_33_2_1_Adder_0_U.u1.cout ;
assign \add_33s_33ns_33_2_1_U1.top_add_33s_33ns_33_2_1_Adder_0_U.fas_s1  = \add_33s_33ns_33_2_1_U1.top_add_33s_33ns_33_2_1_Adder_0_U.u1.s ;
assign \add_33s_33ns_33_2_1_U1.top_add_33s_33ns_33_2_1_Adder_0_U.a  = \add_33s_33ns_33_2_1_U1.din0 ;
assign \add_33s_33ns_33_2_1_U1.top_add_33s_33ns_33_2_1_Adder_0_U.b  = \add_33s_33ns_33_2_1_U1.din1 ;
assign \add_33s_33ns_33_2_1_U1.top_add_33s_33ns_33_2_1_Adder_0_U.ce  = \add_33s_33ns_33_2_1_U1.ce ;
assign \add_33s_33ns_33_2_1_U1.top_add_33s_33ns_33_2_1_Adder_0_U.clk  = \add_33s_33ns_33_2_1_U1.clk ;
assign \add_33s_33ns_33_2_1_U1.top_add_33s_33ns_33_2_1_Adder_0_U.reset  = \add_33s_33ns_33_2_1_U1.reset ;
assign \add_33s_33ns_33_2_1_U1.dout  = \add_33s_33ns_33_2_1_U1.top_add_33s_33ns_33_2_1_Adder_0_U.s ;
assign \add_33s_33ns_33_2_1_U1.ce  = 1'h1;
assign \add_33s_33ns_33_2_1_U1.clk  = ap_clk;
assign \add_33s_33ns_33_2_1_U1.din0  = { op_3[31], op_3 };
assign \add_33s_33ns_33_2_1_U1.din1  = 33'h000000200;
assign grp_fu_227_p2 = \add_33s_33ns_33_2_1_U1.dout ;
assign \add_33s_33ns_33_2_1_U1.reset  = ap_rst;
assign \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.ain_s0  = \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.a ;
assign \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.bin_s0  = \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.b ;
assign \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.s  = { \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.fas_s2 , \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.sum_s1  };
assign \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.u2.a  = \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.ain_s1 ;
assign \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.u2.b  = \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.bin_s1 ;
assign \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.u2.cin  = \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.carry_s1 ;
assign \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.facout_s2  = \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.u2.cout ;
assign \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.fas_s2  = \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.u2.s ;
assign \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.u1.a  = \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.a [15:0];
assign \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.u1.b  = \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.b [15:0];
assign \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.u1.cin  = 1'h0;
assign \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.facout_s1  = \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.u1.cout ;
assign \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.fas_s1  = \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.u1.s ;
assign \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.a  = \add_32ns_32s_32_2_1_U12.din0 ;
assign \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.b  = \add_32ns_32s_32_2_1_U12.din1 ;
assign \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.ce  = \add_32ns_32s_32_2_1_U12.ce ;
assign \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.clk  = \add_32ns_32s_32_2_1_U12.clk ;
assign \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.reset  = \add_32ns_32s_32_2_1_U12.reset ;
assign \add_32ns_32s_32_2_1_U12.dout  = \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.s ;
assign \add_32ns_32s_32_2_1_U12.ce  = 1'h1;
assign \add_32ns_32s_32_2_1_U12.clk  = ap_clk;
assign \add_32ns_32s_32_2_1_U12.din0  = ret_V_21_reg_920;
assign \add_32ns_32s_32_2_1_U12.din1  = { op_15_V_reg_826[1], op_15_V_reg_826[1], op_15_V_reg_826[1], op_15_V_reg_826[1], op_15_V_reg_826[1], op_15_V_reg_826[1], op_15_V_reg_826[1], op_15_V_reg_826[1], op_15_V_reg_826[1], op_15_V_reg_826[1], op_15_V_reg_826[1], op_15_V_reg_826[1], op_15_V_reg_826[1], op_15_V_reg_826[1], op_15_V_reg_826[1], op_15_V_reg_826[1], op_15_V_reg_826[1], op_15_V_reg_826[1], op_15_V_reg_826[1], op_15_V_reg_826[1], op_15_V_reg_826[1], op_15_V_reg_826[1], op_15_V_reg_826[1], op_15_V_reg_826[1], op_15_V_reg_826[1], op_15_V_reg_826[1], op_15_V_reg_826[1], op_15_V_reg_826[1], op_15_V_reg_826[1], op_15_V_reg_826[1], op_15_V_reg_826 };
assign grp_fu_571_p2 = \add_32ns_32s_32_2_1_U12.dout ;
assign \add_32ns_32s_32_2_1_U12.reset  = ap_rst;
assign \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.ain_s0  = \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.a ;
assign \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.bin_s0  = \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.b ;
assign \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.s  = { \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.fas_s2 , \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.sum_s1  };
assign \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.u2.a  = \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.ain_s1 ;
assign \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.u2.b  = \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.bin_s1 ;
assign \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.u2.cin  = \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.carry_s1 ;
assign \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.facout_s2  = \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.u2.cout ;
assign \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.fas_s2  = \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.u2.s ;
assign \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.u1.a  = \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.a [15:0];
assign \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.u1.b  = \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.b [15:0];
assign \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.u1.cin  = 1'h0;
assign \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.facout_s1  = \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.u1.cout ;
assign \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.fas_s1  = \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.u1.s ;
assign \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.a  = \add_32ns_32s_32_2_1_U11.din0 ;
assign \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.b  = \add_32ns_32s_32_2_1_U11.din1 ;
assign \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.ce  = \add_32ns_32s_32_2_1_U11.ce ;
assign \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.clk  = \add_32ns_32s_32_2_1_U11.clk ;
assign \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.reset  = \add_32ns_32s_32_2_1_U11.reset ;
assign \add_32ns_32s_32_2_1_U11.dout  = \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.s ;
assign \add_32ns_32s_32_2_1_U11.ce  = 1'h1;
assign \add_32ns_32s_32_2_1_U11.clk  = ap_clk;
assign \add_32ns_32s_32_2_1_U11.din0  = ret_V_20_reg_910;
assign \add_32ns_32s_32_2_1_U11.din1  = { op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14 };
assign grp_fu_563_p2 = \add_32ns_32s_32_2_1_U11.dout ;
assign \add_32ns_32s_32_2_1_U11.reset  = ap_rst;
assign \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s0  = \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.a ;
assign \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s0  = \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.b ;
assign \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.s  = { \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s2 , \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.sum_s1  };
assign \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.a  = \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s1 ;
assign \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.b  = \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s1 ;
assign \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cin  = \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.carry_s1 ;
assign \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.facout_s2  = \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cout ;
assign \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s2  = \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.s ;
assign \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.a  = \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.a [15:0];
assign \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.b  = \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.b [15:0];
assign \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cin  = 1'h0;
assign \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.facout_s1  = \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cout ;
assign \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s1  = \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.s ;
assign \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.a  = \add_32ns_32ns_32_2_1_U18.din0 ;
assign \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.b  = \add_32ns_32ns_32_2_1_U18.din1 ;
assign \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.ce  = \add_32ns_32ns_32_2_1_U18.ce ;
assign \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.clk  = \add_32ns_32ns_32_2_1_U18.clk ;
assign \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.reset  = \add_32ns_32ns_32_2_1_U18.reset ;
assign \add_32ns_32ns_32_2_1_U18.dout  = \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.s ;
assign \add_32ns_32ns_32_2_1_U18.ce  = 1'h1;
assign \add_32ns_32ns_32_2_1_U18.clk  = ap_clk;
assign \add_32ns_32ns_32_2_1_U18.din0  = ret_V_26_reg_1019;
assign \add_32ns_32ns_32_2_1_U18.din1  = select_ln69_reg_1024;
assign grp_fu_725_p2 = \add_32ns_32ns_32_2_1_U18.dout ;
assign \add_32ns_32ns_32_2_1_U18.reset  = ap_rst;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s0  = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_7_U.a ;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s0  = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_7_U.b ;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_7_U.s  = { \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s2 , \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_7_U.sum_s1  };
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.a  = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s1 ;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.b  = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s1 ;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cin  = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_7_U.carry_s1 ;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_7_U.facout_s2  = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cout ;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s2  = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.s ;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.a  = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_7_U.a [15:0];
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.b  = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_7_U.b [15:0];
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cin  = 1'h0;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_7_U.facout_s1  = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cout ;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s1  = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.s ;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_7_U.a  = \add_32ns_32ns_32_2_1_U17.din0 ;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_7_U.b  = \add_32ns_32ns_32_2_1_U17.din1 ;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_7_U.ce  = \add_32ns_32ns_32_2_1_U17.ce ;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_7_U.clk  = \add_32ns_32ns_32_2_1_U17.clk ;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_7_U.reset  = \add_32ns_32ns_32_2_1_U17.reset ;
assign \add_32ns_32ns_32_2_1_U17.dout  = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_7_U.s ;
assign \add_32ns_32ns_32_2_1_U17.ce  = 1'h1;
assign \add_32ns_32ns_32_2_1_U17.clk  = ap_clk;
assign \add_32ns_32ns_32_2_1_U17.din0  = ret_V_21_cast_reg_1007;
assign \add_32ns_32ns_32_2_1_U17.din1  = 32'd1;
assign grp_fu_693_p2 = \add_32ns_32ns_32_2_1_U17.dout ;
assign \add_32ns_32ns_32_2_1_U17.reset  = ap_rst;
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s0  = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.a ;
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s0  = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.b ;
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.s  = { \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s2 , \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.sum_s1  };
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.a  = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s1 ;
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.b  = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s1 ;
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cin  = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.carry_s1 ;
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.facout_s2  = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cout ;
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s2  = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.s ;
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.a  = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.a [15:0];
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.b  = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.b [15:0];
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cin  = 1'h0;
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.facout_s1  = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cout ;
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s1  = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.s ;
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.a  = \add_32ns_32ns_32_2_1_U15.din0 ;
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.b  = \add_32ns_32ns_32_2_1_U15.din1 ;
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.ce  = \add_32ns_32ns_32_2_1_U15.ce ;
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.clk  = \add_32ns_32ns_32_2_1_U15.clk ;
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.reset  = \add_32ns_32ns_32_2_1_U15.reset ;
assign \add_32ns_32ns_32_2_1_U15.dout  = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.s ;
assign \add_32ns_32ns_32_2_1_U15.ce  = 1'h1;
assign \add_32ns_32ns_32_2_1_U15.clk  = ap_clk;
assign \add_32ns_32ns_32_2_1_U15.din0  = ret_V_24_reg_972;
assign \add_32ns_32ns_32_2_1_U15.din1  = { 31'h00000000, op_17_V_reg_967 };
assign grp_fu_647_p2 = \add_32ns_32ns_32_2_1_U15.dout ;
assign \add_32ns_32ns_32_2_1_U15.reset  = ap_rst;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s0  = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.a ;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s0  = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.b ;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.s  = { \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s2 , \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.sum_s1  };
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.a  = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s1 ;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.b  = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s1 ;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cin  = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.carry_s1 ;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.facout_s2  = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cout ;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s2  = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.s ;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.a  = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.a [15:0];
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.b  = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.b [15:0];
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cin  = 1'h0;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.facout_s1  = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cout ;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s1  = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.s ;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.a  = \add_32ns_32ns_32_2_1_U14.din0 ;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.b  = \add_32ns_32ns_32_2_1_U14.din1 ;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.ce  = \add_32ns_32ns_32_2_1_U14.ce ;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.clk  = \add_32ns_32ns_32_2_1_U14.clk ;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.reset  = \add_32ns_32ns_32_2_1_U14.reset ;
assign \add_32ns_32ns_32_2_1_U14.dout  = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.s ;
assign \add_32ns_32ns_32_2_1_U14.ce  = 1'h1;
assign \add_32ns_32ns_32_2_1_U14.clk  = ap_clk;
assign \add_32ns_32ns_32_2_1_U14.din0  = ret_V_19_cast_reg_955;
assign \add_32ns_32ns_32_2_1_U14.din1  = 32'd1;
assign grp_fu_607_p2 = \add_32ns_32ns_32_2_1_U14.dout ;
assign \add_32ns_32ns_32_2_1_U14.reset  = ap_rst;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s0  = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.a ;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s0  = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.b ;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.s  = { \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s2 , \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.sum_s1  };
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.a  = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s1 ;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.b  = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s1 ;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cin  = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.carry_s1 ;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.facout_s2  = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cout ;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s2  = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.s ;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.a  = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.a [15:0];
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.b  = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.b [15:0];
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cin  = 1'h0;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.facout_s1  = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cout ;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s1  = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.s ;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.a  = \add_32ns_32ns_32_2_1_U10.din0 ;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.b  = \add_32ns_32ns_32_2_1_U10.din1 ;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.ce  = \add_32ns_32ns_32_2_1_U10.ce ;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.clk  = \add_32ns_32ns_32_2_1_U10.clk ;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.reset  = \add_32ns_32ns_32_2_1_U10.reset ;
assign \add_32ns_32ns_32_2_1_U10.dout  = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.s ;
assign \add_32ns_32ns_32_2_1_U10.ce  = 1'h1;
assign \add_32ns_32ns_32_2_1_U10.clk  = ap_clk;
assign \add_32ns_32ns_32_2_1_U10.din0  = ret_V_8_cast_reg_898;
assign \add_32ns_32ns_32_2_1_U10.din1  = 32'd1;
assign grp_fu_535_p2 = \add_32ns_32ns_32_2_1_U10.dout ;
assign \add_32ns_32ns_32_2_1_U10.reset  = ap_rst;
assign \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.ain_s0  = \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.a ;
assign \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.bin_s0  = \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.b ;
assign \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.s  = { \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.fas_s2 , \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.sum_s1  };
assign \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.a  = \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.ain_s1 ;
assign \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.b  = \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.bin_s1 ;
assign \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.cin  = \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.carry_s1 ;
assign \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.facout_s2  = \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.cout ;
assign \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.fas_s2  = \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.s ;
assign \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.a  = \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.a [0];
assign \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.b  = \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.b [0];
assign \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.cin  = 1'h0;
assign \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.facout_s1  = \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.cout ;
assign \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.fas_s1  = \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.s ;
assign \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.a  = \add_2ns_2ns_2_2_1_U2.din0 ;
assign \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.b  = \add_2ns_2ns_2_2_1_U2.din1 ;
assign \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.ce  = \add_2ns_2ns_2_2_1_U2.ce ;
assign \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.clk  = \add_2ns_2ns_2_2_1_U2.clk ;
assign \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.reset  = \add_2ns_2ns_2_2_1_U2.reset ;
assign \add_2ns_2ns_2_2_1_U2.dout  = \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.s ;
assign \add_2ns_2ns_2_2_1_U2.ce  = 1'h1;
assign \add_2ns_2ns_2_2_1_U2.clk  = ap_clk;
assign \add_2ns_2ns_2_2_1_U2.din0  = { op_2[2], 1'h1 };
assign \add_2ns_2ns_2_2_1_U2.din1  = 2'h1;
assign grp_fu_267_p2 = \add_2ns_2ns_2_2_1_U2.dout ;
assign \add_2ns_2ns_2_2_1_U2.reset  = ap_rst;
assign \add_25s_25ns_25_2_1_U8.top_add_25s_25ns_25_2_1_Adder_2_U.ain_s0  = \add_25s_25ns_25_2_1_U8.top_add_25s_25ns_25_2_1_Adder_2_U.a ;
assign \add_25s_25ns_25_2_1_U8.top_add_25s_25ns_25_2_1_Adder_2_U.bin_s0  = \add_25s_25ns_25_2_1_U8.top_add_25s_25ns_25_2_1_Adder_2_U.b ;
assign \add_25s_25ns_25_2_1_U8.top_add_25s_25ns_25_2_1_Adder_2_U.s  = { \add_25s_25ns_25_2_1_U8.top_add_25s_25ns_25_2_1_Adder_2_U.fas_s2 , \add_25s_25ns_25_2_1_U8.top_add_25s_25ns_25_2_1_Adder_2_U.sum_s1  };
assign \add_25s_25ns_25_2_1_U8.top_add_25s_25ns_25_2_1_Adder_2_U.u2.a  = \add_25s_25ns_25_2_1_U8.top_add_25s_25ns_25_2_1_Adder_2_U.ain_s1 ;
assign \add_25s_25ns_25_2_1_U8.top_add_25s_25ns_25_2_1_Adder_2_U.u2.b  = \add_25s_25ns_25_2_1_U8.top_add_25s_25ns_25_2_1_Adder_2_U.bin_s1 ;
assign \add_25s_25ns_25_2_1_U8.top_add_25s_25ns_25_2_1_Adder_2_U.u2.cin  = \add_25s_25ns_25_2_1_U8.top_add_25s_25ns_25_2_1_Adder_2_U.carry_s1 ;
assign \add_25s_25ns_25_2_1_U8.top_add_25s_25ns_25_2_1_Adder_2_U.facout_s2  = \add_25s_25ns_25_2_1_U8.top_add_25s_25ns_25_2_1_Adder_2_U.u2.cout ;
assign \add_25s_25ns_25_2_1_U8.top_add_25s_25ns_25_2_1_Adder_2_U.fas_s2  = \add_25s_25ns_25_2_1_U8.top_add_25s_25ns_25_2_1_Adder_2_U.u2.s ;
assign \add_25s_25ns_25_2_1_U8.top_add_25s_25ns_25_2_1_Adder_2_U.u1.a  = \add_25s_25ns_25_2_1_U8.top_add_25s_25ns_25_2_1_Adder_2_U.a [11:0];
assign \add_25s_25ns_25_2_1_U8.top_add_25s_25ns_25_2_1_Adder_2_U.u1.b  = \add_25s_25ns_25_2_1_U8.top_add_25s_25ns_25_2_1_Adder_2_U.b [11:0];
assign \add_25s_25ns_25_2_1_U8.top_add_25s_25ns_25_2_1_Adder_2_U.u1.cin  = 1'h0;
assign \add_25s_25ns_25_2_1_U8.top_add_25s_25ns_25_2_1_Adder_2_U.facout_s1  = \add_25s_25ns_25_2_1_U8.top_add_25s_25ns_25_2_1_Adder_2_U.u1.cout ;
assign \add_25s_25ns_25_2_1_U8.top_add_25s_25ns_25_2_1_Adder_2_U.fas_s1  = \add_25s_25ns_25_2_1_U8.top_add_25s_25ns_25_2_1_Adder_2_U.u1.s ;
assign \add_25s_25ns_25_2_1_U8.top_add_25s_25ns_25_2_1_Adder_2_U.a  = \add_25s_25ns_25_2_1_U8.din0 ;
assign \add_25s_25ns_25_2_1_U8.top_add_25s_25ns_25_2_1_Adder_2_U.b  = \add_25s_25ns_25_2_1_U8.din1 ;
assign \add_25s_25ns_25_2_1_U8.top_add_25s_25ns_25_2_1_Adder_2_U.ce  = \add_25s_25ns_25_2_1_U8.ce ;
assign \add_25s_25ns_25_2_1_U8.top_add_25s_25ns_25_2_1_Adder_2_U.clk  = \add_25s_25ns_25_2_1_U8.clk ;
assign \add_25s_25ns_25_2_1_U8.top_add_25s_25ns_25_2_1_Adder_2_U.reset  = \add_25s_25ns_25_2_1_U8.reset ;
assign \add_25s_25ns_25_2_1_U8.dout  = \add_25s_25ns_25_2_1_U8.top_add_25s_25ns_25_2_1_Adder_2_U.s ;
assign \add_25s_25ns_25_2_1_U8.ce  = 1'h1;
assign \add_25s_25ns_25_2_1_U8.clk  = ap_clk;
assign \add_25s_25ns_25_2_1_U8.din0  = { add_ln69_1_reg_836[4], add_ln69_1_reg_836[4], add_ln69_1_reg_836[4], add_ln69_1_reg_836[4], add_ln69_1_reg_836[4], add_ln69_1_reg_836[4], add_ln69_1_reg_836[4], add_ln69_1_reg_836[4], add_ln69_1_reg_836[4], add_ln69_1_reg_836[4], add_ln69_1_reg_836[4], add_ln69_1_reg_836[4], add_ln69_1_reg_836[4], add_ln69_1_reg_836[4], add_ln69_1_reg_836[4], add_ln69_1_reg_836[4], add_ln69_1_reg_836[4], add_ln69_1_reg_836[4], add_ln69_1_reg_836[4], add_ln69_1_reg_836[4], add_ln69_1_reg_836 };
assign \add_25s_25ns_25_2_1_U8.din1  = add_ln69_reg_831;
assign grp_fu_450_p2 = \add_25s_25ns_25_2_1_U8.dout ;
assign \add_25s_25ns_25_2_1_U8.reset  = ap_rst;
assign \add_25s_25ns_25_2_1_U3.top_add_25s_25ns_25_2_1_Adder_2_U.ain_s0  = \add_25s_25ns_25_2_1_U3.top_add_25s_25ns_25_2_1_Adder_2_U.a ;
assign \add_25s_25ns_25_2_1_U3.top_add_25s_25ns_25_2_1_Adder_2_U.bin_s0  = \add_25s_25ns_25_2_1_U3.top_add_25s_25ns_25_2_1_Adder_2_U.b ;
assign \add_25s_25ns_25_2_1_U3.top_add_25s_25ns_25_2_1_Adder_2_U.s  = { \add_25s_25ns_25_2_1_U3.top_add_25s_25ns_25_2_1_Adder_2_U.fas_s2 , \add_25s_25ns_25_2_1_U3.top_add_25s_25ns_25_2_1_Adder_2_U.sum_s1  };
assign \add_25s_25ns_25_2_1_U3.top_add_25s_25ns_25_2_1_Adder_2_U.u2.a  = \add_25s_25ns_25_2_1_U3.top_add_25s_25ns_25_2_1_Adder_2_U.ain_s1 ;
assign \add_25s_25ns_25_2_1_U3.top_add_25s_25ns_25_2_1_Adder_2_U.u2.b  = \add_25s_25ns_25_2_1_U3.top_add_25s_25ns_25_2_1_Adder_2_U.bin_s1 ;
assign \add_25s_25ns_25_2_1_U3.top_add_25s_25ns_25_2_1_Adder_2_U.u2.cin  = \add_25s_25ns_25_2_1_U3.top_add_25s_25ns_25_2_1_Adder_2_U.carry_s1 ;
assign \add_25s_25ns_25_2_1_U3.top_add_25s_25ns_25_2_1_Adder_2_U.facout_s2  = \add_25s_25ns_25_2_1_U3.top_add_25s_25ns_25_2_1_Adder_2_U.u2.cout ;
assign \add_25s_25ns_25_2_1_U3.top_add_25s_25ns_25_2_1_Adder_2_U.fas_s2  = \add_25s_25ns_25_2_1_U3.top_add_25s_25ns_25_2_1_Adder_2_U.u2.s ;
assign \add_25s_25ns_25_2_1_U3.top_add_25s_25ns_25_2_1_Adder_2_U.u1.a  = \add_25s_25ns_25_2_1_U3.top_add_25s_25ns_25_2_1_Adder_2_U.a [11:0];
assign \add_25s_25ns_25_2_1_U3.top_add_25s_25ns_25_2_1_Adder_2_U.u1.b  = \add_25s_25ns_25_2_1_U3.top_add_25s_25ns_25_2_1_Adder_2_U.b [11:0];
assign \add_25s_25ns_25_2_1_U3.top_add_25s_25ns_25_2_1_Adder_2_U.u1.cin  = 1'h0;
assign \add_25s_25ns_25_2_1_U3.top_add_25s_25ns_25_2_1_Adder_2_U.facout_s1  = \add_25s_25ns_25_2_1_U3.top_add_25s_25ns_25_2_1_Adder_2_U.u1.cout ;
assign \add_25s_25ns_25_2_1_U3.top_add_25s_25ns_25_2_1_Adder_2_U.fas_s1  = \add_25s_25ns_25_2_1_U3.top_add_25s_25ns_25_2_1_Adder_2_U.u1.s ;
assign \add_25s_25ns_25_2_1_U3.top_add_25s_25ns_25_2_1_Adder_2_U.a  = \add_25s_25ns_25_2_1_U3.din0 ;
assign \add_25s_25ns_25_2_1_U3.top_add_25s_25ns_25_2_1_Adder_2_U.b  = \add_25s_25ns_25_2_1_U3.din1 ;
assign \add_25s_25ns_25_2_1_U3.top_add_25s_25ns_25_2_1_Adder_2_U.ce  = \add_25s_25ns_25_2_1_U3.ce ;
assign \add_25s_25ns_25_2_1_U3.top_add_25s_25ns_25_2_1_Adder_2_U.clk  = \add_25s_25ns_25_2_1_U3.clk ;
assign \add_25s_25ns_25_2_1_U3.top_add_25s_25ns_25_2_1_Adder_2_U.reset  = \add_25s_25ns_25_2_1_U3.reset ;
assign \add_25s_25ns_25_2_1_U3.dout  = \add_25s_25ns_25_2_1_U3.top_add_25s_25ns_25_2_1_Adder_2_U.s ;
assign \add_25s_25ns_25_2_1_U3.ce  = 1'h1;
assign \add_25s_25ns_25_2_1_U3.clk  = ap_clk;
assign \add_25s_25ns_25_2_1_U3.din0  = { tmp_1_reg_740[23], tmp_1_reg_740 };
assign \add_25s_25ns_25_2_1_U3.din1  = 25'h0000001;
assign grp_fu_281_p2 = \add_25s_25ns_25_2_1_U3.dout ;
assign \add_25s_25ns_25_2_1_U3.reset  = ap_rst;
assign \add_25ns_25s_25_2_1_U5.top_add_25ns_25s_25_2_1_Adder_3_U.ain_s0  = \add_25ns_25s_25_2_1_U5.top_add_25ns_25s_25_2_1_Adder_3_U.a ;
assign \add_25ns_25s_25_2_1_U5.top_add_25ns_25s_25_2_1_Adder_3_U.bin_s0  = \add_25ns_25s_25_2_1_U5.top_add_25ns_25s_25_2_1_Adder_3_U.b ;
assign \add_25ns_25s_25_2_1_U5.top_add_25ns_25s_25_2_1_Adder_3_U.s  = { \add_25ns_25s_25_2_1_U5.top_add_25ns_25s_25_2_1_Adder_3_U.fas_s2 , \add_25ns_25s_25_2_1_U5.top_add_25ns_25s_25_2_1_Adder_3_U.sum_s1  };
assign \add_25ns_25s_25_2_1_U5.top_add_25ns_25s_25_2_1_Adder_3_U.u2.a  = \add_25ns_25s_25_2_1_U5.top_add_25ns_25s_25_2_1_Adder_3_U.ain_s1 ;
assign \add_25ns_25s_25_2_1_U5.top_add_25ns_25s_25_2_1_Adder_3_U.u2.b  = \add_25ns_25s_25_2_1_U5.top_add_25ns_25s_25_2_1_Adder_3_U.bin_s1 ;
assign \add_25ns_25s_25_2_1_U5.top_add_25ns_25s_25_2_1_Adder_3_U.u2.cin  = \add_25ns_25s_25_2_1_U5.top_add_25ns_25s_25_2_1_Adder_3_U.carry_s1 ;
assign \add_25ns_25s_25_2_1_U5.top_add_25ns_25s_25_2_1_Adder_3_U.facout_s2  = \add_25ns_25s_25_2_1_U5.top_add_25ns_25s_25_2_1_Adder_3_U.u2.cout ;
assign \add_25ns_25s_25_2_1_U5.top_add_25ns_25s_25_2_1_Adder_3_U.fas_s2  = \add_25ns_25s_25_2_1_U5.top_add_25ns_25s_25_2_1_Adder_3_U.u2.s ;
assign \add_25ns_25s_25_2_1_U5.top_add_25ns_25s_25_2_1_Adder_3_U.u1.a  = \add_25ns_25s_25_2_1_U5.top_add_25ns_25s_25_2_1_Adder_3_U.a [11:0];
assign \add_25ns_25s_25_2_1_U5.top_add_25ns_25s_25_2_1_Adder_3_U.u1.b  = \add_25ns_25s_25_2_1_U5.top_add_25ns_25s_25_2_1_Adder_3_U.b [11:0];
assign \add_25ns_25s_25_2_1_U5.top_add_25ns_25s_25_2_1_Adder_3_U.u1.cin  = 1'h0;
assign \add_25ns_25s_25_2_1_U5.top_add_25ns_25s_25_2_1_Adder_3_U.facout_s1  = \add_25ns_25s_25_2_1_U5.top_add_25ns_25s_25_2_1_Adder_3_U.u1.cout ;
assign \add_25ns_25s_25_2_1_U5.top_add_25ns_25s_25_2_1_Adder_3_U.fas_s1  = \add_25ns_25s_25_2_1_U5.top_add_25ns_25s_25_2_1_Adder_3_U.u1.s ;
assign \add_25ns_25s_25_2_1_U5.top_add_25ns_25s_25_2_1_Adder_3_U.a  = \add_25ns_25s_25_2_1_U5.din0 ;
assign \add_25ns_25s_25_2_1_U5.top_add_25ns_25s_25_2_1_Adder_3_U.b  = \add_25ns_25s_25_2_1_U5.din1 ;
assign \add_25ns_25s_25_2_1_U5.top_add_25ns_25s_25_2_1_Adder_3_U.ce  = \add_25ns_25s_25_2_1_U5.ce ;
assign \add_25ns_25s_25_2_1_U5.top_add_25ns_25s_25_2_1_Adder_3_U.clk  = \add_25ns_25s_25_2_1_U5.clk ;
assign \add_25ns_25s_25_2_1_U5.top_add_25ns_25s_25_2_1_Adder_3_U.reset  = \add_25ns_25s_25_2_1_U5.reset ;
assign \add_25ns_25s_25_2_1_U5.dout  = \add_25ns_25s_25_2_1_U5.top_add_25ns_25s_25_2_1_Adder_3_U.s ;
assign \add_25ns_25s_25_2_1_U5.ce  = 1'h1;
assign \add_25ns_25s_25_2_1_U5.clk  = ap_clk;
assign \add_25ns_25s_25_2_1_U5.din0  = ret_V_17_reg_790;
assign \add_25ns_25s_25_2_1_U5.din1  = { op_11[7], op_11[7], op_11[7], op_11[7], op_11[7], op_11[7], op_11[7], op_11[7], op_11[7], op_11[7], op_11[7], op_11[7], op_11[7], op_11[7], op_11[7], op_11[7], op_11[7], op_11 };
assign grp_fu_350_p2 = \add_25ns_25s_25_2_1_U5.dout ;
assign \add_25ns_25s_25_2_1_U5.reset  = ap_rst;
assign \add_18ns_18s_18_2_1_U7.top_add_18ns_18s_18_2_1_Adder_5_U.ain_s0  = \add_18ns_18s_18_2_1_U7.top_add_18ns_18s_18_2_1_Adder_5_U.a ;
assign \add_18ns_18s_18_2_1_U7.top_add_18ns_18s_18_2_1_Adder_5_U.bin_s0  = \add_18ns_18s_18_2_1_U7.top_add_18ns_18s_18_2_1_Adder_5_U.b ;
assign \add_18ns_18s_18_2_1_U7.top_add_18ns_18s_18_2_1_Adder_5_U.s  = { \add_18ns_18s_18_2_1_U7.top_add_18ns_18s_18_2_1_Adder_5_U.fas_s2 , \add_18ns_18s_18_2_1_U7.top_add_18ns_18s_18_2_1_Adder_5_U.sum_s1  };
assign \add_18ns_18s_18_2_1_U7.top_add_18ns_18s_18_2_1_Adder_5_U.u2.a  = \add_18ns_18s_18_2_1_U7.top_add_18ns_18s_18_2_1_Adder_5_U.ain_s1 ;
assign \add_18ns_18s_18_2_1_U7.top_add_18ns_18s_18_2_1_Adder_5_U.u2.b  = \add_18ns_18s_18_2_1_U7.top_add_18ns_18s_18_2_1_Adder_5_U.bin_s1 ;
assign \add_18ns_18s_18_2_1_U7.top_add_18ns_18s_18_2_1_Adder_5_U.u2.cin  = \add_18ns_18s_18_2_1_U7.top_add_18ns_18s_18_2_1_Adder_5_U.carry_s1 ;
assign \add_18ns_18s_18_2_1_U7.top_add_18ns_18s_18_2_1_Adder_5_U.facout_s2  = \add_18ns_18s_18_2_1_U7.top_add_18ns_18s_18_2_1_Adder_5_U.u2.cout ;
assign \add_18ns_18s_18_2_1_U7.top_add_18ns_18s_18_2_1_Adder_5_U.fas_s2  = \add_18ns_18s_18_2_1_U7.top_add_18ns_18s_18_2_1_Adder_5_U.u2.s ;
assign \add_18ns_18s_18_2_1_U7.top_add_18ns_18s_18_2_1_Adder_5_U.u1.a  = \add_18ns_18s_18_2_1_U7.top_add_18ns_18s_18_2_1_Adder_5_U.a [8:0];
assign \add_18ns_18s_18_2_1_U7.top_add_18ns_18s_18_2_1_Adder_5_U.u1.b  = \add_18ns_18s_18_2_1_U7.top_add_18ns_18s_18_2_1_Adder_5_U.b [8:0];
assign \add_18ns_18s_18_2_1_U7.top_add_18ns_18s_18_2_1_Adder_5_U.u1.cin  = 1'h0;
assign \add_18ns_18s_18_2_1_U7.top_add_18ns_18s_18_2_1_Adder_5_U.facout_s1  = \add_18ns_18s_18_2_1_U7.top_add_18ns_18s_18_2_1_Adder_5_U.u1.cout ;
assign \add_18ns_18s_18_2_1_U7.top_add_18ns_18s_18_2_1_Adder_5_U.fas_s1  = \add_18ns_18s_18_2_1_U7.top_add_18ns_18s_18_2_1_Adder_5_U.u1.s ;
assign \add_18ns_18s_18_2_1_U7.top_add_18ns_18s_18_2_1_Adder_5_U.a  = \add_18ns_18s_18_2_1_U7.din0 ;
assign \add_18ns_18s_18_2_1_U7.top_add_18ns_18s_18_2_1_Adder_5_U.b  = \add_18ns_18s_18_2_1_U7.din1 ;
assign \add_18ns_18s_18_2_1_U7.top_add_18ns_18s_18_2_1_Adder_5_U.ce  = \add_18ns_18s_18_2_1_U7.ce ;
assign \add_18ns_18s_18_2_1_U7.top_add_18ns_18s_18_2_1_Adder_5_U.clk  = \add_18ns_18s_18_2_1_U7.clk ;
assign \add_18ns_18s_18_2_1_U7.top_add_18ns_18s_18_2_1_Adder_5_U.reset  = \add_18ns_18s_18_2_1_U7.reset ;
assign \add_18ns_18s_18_2_1_U7.dout  = \add_18ns_18s_18_2_1_U7.top_add_18ns_18s_18_2_1_Adder_5_U.s ;
assign \add_18ns_18s_18_2_1_U7.ce  = 1'h1;
assign \add_18ns_18s_18_2_1_U7.clk  = ap_clk;
assign \add_18ns_18s_18_2_1_U7.din0  = { 2'h0, ret_reg_795[3], ret_reg_795[3], ret_reg_795[3], ret_reg_795[3], ret_reg_795, 8'h00 };
assign \add_18ns_18s_18_2_1_U7.din1  = { op_5[15], op_5[15], op_5 };
assign grp_fu_398_p2 = \add_18ns_18s_18_2_1_U7.dout ;
assign \add_18ns_18s_18_2_1_U7.reset  = ap_rst;
endmodule


// Product machine:
module top_A_times_top_B (ap_start, op_0, op_10, op_11, op_14, op_16, op_18, op_19, op_2, op_3, op_5, op_8, ap_clk, unsafe_signal);
input ap_start;
input [3:0] op_0;
input [7:0] op_10;
input [7:0] op_11;
input [3:0] op_14;
input [7:0] op_16;
input [31:0] op_18;
input op_19;
input [3:0] op_2;
input [31:0] op_3;
input [15:0] op_5;
input [3:0] op_8;
input ap_clk;
output unsafe_signal;
reg _setup;
initial _setup = 1'b0;
always @ (posedge ap_clk) _setup <= 1'b1;
reg ap_start_internal;
always @ (posedge ap_clk) if (!_setup) ap_start_internal <= ap_start;
reg [3:0] op_0_internal;
always @ (posedge ap_clk) if (!_setup) op_0_internal <= op_0;
reg [7:0] op_10_internal;
always @ (posedge ap_clk) if (!_setup) op_10_internal <= op_10;
reg [7:0] op_11_internal;
always @ (posedge ap_clk) if (!_setup) op_11_internal <= op_11;
reg [3:0] op_14_internal;
always @ (posedge ap_clk) if (!_setup) op_14_internal <= op_14;
reg [7:0] op_16_internal;
always @ (posedge ap_clk) if (!_setup) op_16_internal <= op_16;
reg [31:0] op_18_internal;
always @ (posedge ap_clk) if (!_setup) op_18_internal <= op_18;
reg op_19_internal;
always @ (posedge ap_clk) if (!_setup) op_19_internal <= op_19;
reg [3:0] op_2_internal;
always @ (posedge ap_clk) if (!_setup) op_2_internal <= op_2;
reg [31:0] op_3_internal;
always @ (posedge ap_clk) if (!_setup) op_3_internal <= op_3;
reg [15:0] op_5_internal;
always @ (posedge ap_clk) if (!_setup) op_5_internal <= op_5;
reg [3:0] op_8_internal;
always @ (posedge ap_clk) if (!_setup) op_8_internal <= op_8;
wire ap_done_A;
wire ap_done_B;
wire ap_done_eq;
assign ap_done_eq = ap_done_A == ap_done_B;
wire ap_idle_A;
wire ap_idle_B;
wire ap_idle_eq;
assign ap_idle_eq = ap_idle_A == ap_idle_B;
wire ap_ready_A;
wire ap_ready_B;
wire ap_ready_eq;
assign ap_ready_eq = ap_ready_A == ap_ready_B;
wire [31:0] op_30_A;
wire [31:0] op_30_B;
wire op_30_eq;
assign op_30_eq = op_30_A == op_30_B;
wire op_30_ap_vld_A;
wire op_30_ap_vld_B;
wire clk_enable_A;
wire clk_enable_B;
assign clk_enable_A = _setup & (~op_30_ap_vld_A | op_30_ap_vld_B);
assign clk_enable_B = _setup;
wire divergent;
assign divergent = ~(ap_done_eq & ap_idle_eq & ap_ready_eq & op_30_eq);
assign unsafe_signal = op_30_ap_vld_A & op_30_ap_vld_B & divergent;
top_A instance_A (
    .ap_clk(ap_clk),
    .clk_enable(clk_enable_A),
    .ap_start(ap_start_internal),
    .op_0(op_0_internal),
    .op_10(op_10_internal),
    .op_11(op_11_internal),
    .op_14(op_14_internal),
    .op_16(op_16_internal),
    .op_18(op_18_internal),
    .op_19(op_19_internal),
    .op_2(op_2_internal),
    .op_3(op_3_internal),
    .op_5(op_5_internal),
    .op_8(op_8_internal),
    .ap_done(ap_done_A),
    .ap_idle(ap_idle_A),
    .ap_ready(ap_ready_A),
    .op_30(op_30_A),
    .op_30_ap_vld(op_30_ap_vld_A)
);
top_B instance_B (
    .ap_clk(ap_clk),
    .clk_enable(clk_enable_B),
    .ap_start(ap_start_internal),
    .op_0(op_0_internal),
    .op_10(op_10_internal),
    .op_11(op_11_internal),
    .op_14(op_14_internal),
    .op_16(op_16_internal),
    .op_18(op_18_internal),
    .op_19(op_19_internal),
    .op_2(op_2_internal),
    .op_3(op_3_internal),
    .op_5(op_5_internal),
    .op_8(op_8_internal),
    .ap_done(ap_done_B),
    .ap_idle(ap_idle_B),
    .ap_ready(ap_ready_B),
    .op_30(op_30_B),
    .op_30_ap_vld(op_30_ap_vld_B)
);
endmodule
