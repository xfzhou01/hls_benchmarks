// Processed by function `construct_kairos` in `verilog_tricks.py`.
// Machine A:
// Processed by function `add_clk_enable_signal` in `verilog_tricks.py`.
// Processed by function `remove_reset_signal` in `verilog_tricks.py`.
module top_A (
  ap_clk,
  ap_start,
  ap_done,
  ap_idle,
  ap_ready,
  op_0,
  op_1,
  op_4,
  op_6,
  op_8,
  op_9,
  op_10,
  op_12,
  op_13,
  op_14,
  op_15,
  op_17,
  op_18,
  op_19,
  op_31,
  op_31_ap_vld,
clk_enable
);
input clk_enable;


input ap_clk;
wire ap_rst;
assign ap_rst = op_31_ap_vld;
input ap_start;
input [1:0] op_0;
input [3:0] op_1;
input [3:0] op_10;
input [31:0] op_12;
input [7:0] op_13;
input [1:0] op_14;
input [3:0] op_15;
input op_17;
input op_18;
input [31:0] op_19;
input [31:0] op_4;
input [3:0] op_6;
input [7:0] op_8;
input op_9;
output ap_done;
output ap_idle;
output ap_ready;
output [31:0] op_31;
output op_31_ap_vld;


reg [8:0] \add_18ns_18ns_18_2_1_U5.top_add_18ns_18ns_18_2_1_Adder_2_U.ain_s1 ;
reg [8:0] \add_18ns_18ns_18_2_1_U5.top_add_18ns_18ns_18_2_1_Adder_2_U.bin_s1 ;
reg \add_18ns_18ns_18_2_1_U5.top_add_18ns_18ns_18_2_1_Adder_2_U.carry_s1 ;
reg [8:0] \add_18ns_18ns_18_2_1_U5.top_add_18ns_18ns_18_2_1_Adder_2_U.sum_s1 ;
reg [8:0] \add_18ns_18s_18_2_1_U4.top_add_18ns_18s_18_2_1_Adder_1_U.ain_s1 ;
reg [8:0] \add_18ns_18s_18_2_1_U4.top_add_18ns_18s_18_2_1_Adder_1_U.bin_s1 ;
reg \add_18ns_18s_18_2_1_U4.top_add_18ns_18s_18_2_1_Adder_1_U.carry_s1 ;
reg [8:0] \add_18ns_18s_18_2_1_U4.top_add_18ns_18s_18_2_1_Adder_1_U.sum_s1 ;
reg [10:0] \add_22s_22s_22_2_1_U7.top_add_22s_22s_22_2_1_Adder_4_U.ain_s1 ;
reg [10:0] \add_22s_22s_22_2_1_U7.top_add_22s_22s_22_2_1_Adder_4_U.bin_s1 ;
reg \add_22s_22s_22_2_1_U7.top_add_22s_22s_22_2_1_Adder_4_U.carry_s1 ;
reg [10:0] \add_22s_22s_22_2_1_U7.top_add_22s_22s_22_2_1_Adder_4_U.sum_s1 ;
reg \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_11_U.ain_s1 ;
reg \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_11_U.bin_s1 ;
reg \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_11_U.carry_s1 ;
reg \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_11_U.sum_s1 ;
reg \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_11_U.ain_s1 ;
reg \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_11_U.bin_s1 ;
reg \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_11_U.carry_s1 ;
reg \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_11_U.sum_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s1 ;
reg \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.carry_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.sum_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s1 ;
reg \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.carry_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.sum_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s1 ;
reg \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.carry_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.sum_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s1 ;
reg \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.carry_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.sum_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s1 ;
reg \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.carry_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.sum_s1 ;
reg [15:0] \add_32ns_32s_32_2_1_U13.top_add_32ns_32s_32_2_1_Adder_9_U.ain_s1 ;
reg [15:0] \add_32ns_32s_32_2_1_U13.top_add_32ns_32s_32_2_1_Adder_9_U.bin_s1 ;
reg \add_32ns_32s_32_2_1_U13.top_add_32ns_32s_32_2_1_Adder_9_U.carry_s1 ;
reg [15:0] \add_32ns_32s_32_2_1_U13.top_add_32ns_32s_32_2_1_Adder_9_U.sum_s1 ;
reg [15:0] \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_5_U.ain_s1 ;
reg [15:0] \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_5_U.bin_s1 ;
reg \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_5_U.carry_s1 ;
reg [15:0] \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_5_U.sum_s1 ;
reg [15:0] \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.ain_s1 ;
reg [15:0] \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.bin_s1 ;
reg \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.carry_s1 ;
reg [15:0] \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.sum_s1 ;
reg [17:0] \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_10_U.ain_s1 ;
reg [17:0] \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_10_U.bin_s1 ;
reg \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_10_U.carry_s1 ;
reg [16:0] \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_10_U.sum_s1 ;
reg [17:0] \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_6_U.ain_s1 ;
reg [17:0] \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_6_U.bin_s1 ;
reg \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_6_U.carry_s1 ;
reg [17:0] \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_6_U.sum_s1 ;
reg [23:0] \add_47s_47s_47_2_1_U11.top_add_47s_47s_47_2_1_Adder_8_U.ain_s1 ;
reg [23:0] \add_47s_47s_47_2_1_U11.top_add_47s_47s_47_2_1_Adder_8_U.bin_s1 ;
reg \add_47s_47s_47_2_1_U11.top_add_47s_47s_47_2_1_Adder_8_U.carry_s1 ;
reg [22:0] \add_47s_47s_47_2_1_U11.top_add_47s_47s_47_2_1_Adder_8_U.sum_s1 ;
reg [31:0] add_ln691_1_reg_913;
reg [31:0] add_ln691_2_reg_950;
reg [31:0] add_ln691_3_reg_1012;
reg [31:0] add_ln691_reg_866;
reg [1:0] add_ln69_1_reg_1032;
reg [1:0] add_ln69_2_reg_1047;
reg [31:0] add_ln69_reg_1042;
reg [41:0] ap_CS_fsm = 42'h00000000001;
reg [3:0] \ashr_4ns_4ns_4_7_1_U2.din1_cast_array[0] ;
reg [3:0] \ashr_4ns_4ns_4_7_1_U2.din1_cast_array[1] ;
reg [3:0] \ashr_4ns_4ns_4_7_1_U2.din1_cast_array[2] ;
reg [3:0] \ashr_4ns_4ns_4_7_1_U2.din1_cast_array[3] ;
reg [3:0] \ashr_4ns_4ns_4_7_1_U2.din1_cast_array[4] ;
reg [3:0] \ashr_4ns_4ns_4_7_1_U2.din1_cast_array[5] ;
reg [3:0] \ashr_4ns_4ns_4_7_1_U2.dout_array[0] ;
reg [3:0] \ashr_4ns_4ns_4_7_1_U2.dout_array[1] ;
reg [3:0] \ashr_4ns_4ns_4_7_1_U2.dout_array[2] ;
reg [3:0] \ashr_4ns_4ns_4_7_1_U2.dout_array[3] ;
reg [3:0] \ashr_4ns_4ns_4_7_1_U2.dout_array[4] ;
reg [3:0] \ashr_4ns_4ns_4_7_1_U2.dout_array[5] ;
reg [3:0] ashr_ln799_reg_744;
reg icmp_ln768_reg_843;
reg icmp_ln786_reg_848;
reg icmp_ln851_1_reg_896;
reg icmp_ln851_2_reg_933;
reg icmp_ln851_3_reg_990;
reg icmp_ln851_reg_805;
reg [3:0] op_11_V_reg_871;
reg [31:0] op_26_V_reg_975;
reg overflow_reg_860;
reg p_Result_4_reg_734;
reg p_Result_5_reg_815;
reg p_Result_6_reg_821;
reg [3:0] r_reg_754;
reg [31:0] ret_V_16_cast_reg_1000;
reg [35:0] ret_V_1_reg_810;
reg [17:0] ret_V_2_reg_780;
reg [31:0] ret_V_3_cast_reg_906;
reg [21:0] ret_V_3_reg_833;
reg [35:0] ret_V_4_reg_901;
reg [46:0] ret_V_5_reg_938;
reg [31:0] ret_V_6_cast_reg_943;
reg [31:0] ret_V_6_reg_955;
reg [31:0] ret_V_7_reg_965;
reg [34:0] ret_V_8_reg_995;
reg [31:0] ret_V_9_reg_1022;
reg [17:0] ret_V_reg_770;
reg [17:0] select_ln1192_reg_775;
reg [31:0] select_ln353_1_reg_918;
reg [31:0] select_ln353_reg_876;
reg [1:0] select_ln69_1_reg_1027;
reg [1:0] select_ln69_reg_1007;
reg [31:0] sext_ln831_reg_853;
reg [3:0] sh_reg_739;
reg [3:0] \shl_4ns_4ns_4_7_1_U3.din1_cast_array[0] ;
reg [3:0] \shl_4ns_4ns_4_7_1_U3.din1_cast_array[1] ;
reg [3:0] \shl_4ns_4ns_4_7_1_U3.din1_cast_array[2] ;
reg [3:0] \shl_4ns_4ns_4_7_1_U3.din1_cast_array[3] ;
reg [3:0] \shl_4ns_4ns_4_7_1_U3.din1_cast_array[4] ;
reg [3:0] \shl_4ns_4ns_4_7_1_U3.din1_cast_array[5] ;
reg [3:0] \shl_4ns_4ns_4_7_1_U3.dout_array[0] ;
reg [3:0] \shl_4ns_4ns_4_7_1_U3.dout_array[1] ;
reg [3:0] \shl_4ns_4ns_4_7_1_U3.dout_array[2] ;
reg [3:0] \shl_4ns_4ns_4_7_1_U3.dout_array[3] ;
reg [3:0] \shl_4ns_4ns_4_7_1_U3.dout_array[4] ;
reg [3:0] \shl_4ns_4ns_4_7_1_U3.dout_array[5] ;
reg [3:0] shl_ln781_reg_749;
reg [17:0] \sub_36s_36ns_36_2_1_U6.top_sub_36s_36ns_36_2_1_Adder_3_U.ain_s1 ;
reg [17:0] \sub_36s_36ns_36_2_1_U6.top_sub_36s_36ns_36_2_1_Adder_3_U.bin_s1 ;
reg \sub_36s_36ns_36_2_1_U6.top_sub_36s_36ns_36_2_1_Adder_3_U.carry_s1 ;
reg [17:0] \sub_36s_36ns_36_2_1_U6.top_sub_36s_36ns_36_2_1_Adder_3_U.sum_s1 ;
reg [1:0] \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.ain_s1 ;
reg [1:0] \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.bin_s1 ;
reg \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.carry_s1 ;
reg [1:0] \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.sum_s1 ;
reg [31:0] tmp_2_reg_827;
reg [18:0] tmp_reg_838;
reg [2:0] trunc_ln851_1_reg_881;
wire [31:0] _000_;
wire [31:0] _001_;
wire [31:0] _002_;
wire [31:0] _003_;
wire [1:0] _004_;
wire [1:0] _005_;
wire [31:0] _006_;
wire [41:0] _007_;
wire [3:0] _008_;
wire _009_;
wire _010_;
wire _011_;
wire _012_;
wire _013_;
wire _014_;
wire [3:0] _015_;
wire [31:0] _016_;
wire _017_;
wire _018_;
wire _019_;
wire _020_;
wire [3:0] _021_;
wire [31:0] _022_;
wire [35:0] _023_;
wire [17:0] _024_;
wire [31:0] _025_;
wire [21:0] _026_;
wire [35:0] _027_;
wire [46:0] _028_;
wire [31:0] _029_;
wire [31:0] _030_;
wire [31:0] _031_;
wire [34:0] _032_;
wire [31:0] _033_;
wire [17:0] _034_;
wire [17:0] _035_;
wire [31:0] _036_;
wire [31:0] _037_;
wire [1:0] _038_;
wire [1:0] _039_;
wire [31:0] _040_;
wire [3:0] _041_;
wire [3:0] _042_;
wire [31:0] _043_;
wire [18:0] _044_;
wire [2:0] _045_;
wire [1:0] _046_;
wire _047_;
wire _048_;
wire _049_;
wire _050_;
wire _051_;
wire _052_;
wire _053_;
wire _054_;
wire _055_;
wire _056_;
wire [8:0] _057_;
wire [8:0] _058_;
wire _059_;
wire [8:0] _060_;
wire [9:0] _061_;
wire [9:0] _062_;
wire [8:0] _063_;
wire [8:0] _064_;
wire _065_;
wire [8:0] _066_;
wire [9:0] _067_;
wire [9:0] _068_;
wire [10:0] _069_;
wire [10:0] _070_;
wire _071_;
wire [10:0] _072_;
wire [11:0] _073_;
wire [11:0] _074_;
wire _075_;
wire _076_;
wire _077_;
wire _078_;
wire [1:0] _079_;
wire [1:0] _080_;
wire _081_;
wire _082_;
wire _083_;
wire _084_;
wire [1:0] _085_;
wire [1:0] _086_;
wire [15:0] _087_;
wire [15:0] _088_;
wire _089_;
wire [15:0] _090_;
wire [16:0] _091_;
wire [16:0] _092_;
wire [15:0] _093_;
wire [15:0] _094_;
wire _095_;
wire [15:0] _096_;
wire [16:0] _097_;
wire [16:0] _098_;
wire [15:0] _099_;
wire [15:0] _100_;
wire _101_;
wire [15:0] _102_;
wire [16:0] _103_;
wire [16:0] _104_;
wire [15:0] _105_;
wire [15:0] _106_;
wire _107_;
wire [15:0] _108_;
wire [16:0] _109_;
wire [16:0] _110_;
wire [15:0] _111_;
wire [15:0] _112_;
wire _113_;
wire [15:0] _114_;
wire [16:0] _115_;
wire [16:0] _116_;
wire [15:0] _117_;
wire [15:0] _118_;
wire _119_;
wire [15:0] _120_;
wire [16:0] _121_;
wire [16:0] _122_;
wire [15:0] _123_;
wire [15:0] _124_;
wire _125_;
wire [15:0] _126_;
wire [16:0] _127_;
wire [16:0] _128_;
wire [15:0] _129_;
wire [15:0] _130_;
wire _131_;
wire [15:0] _132_;
wire [16:0] _133_;
wire [16:0] _134_;
wire [17:0] _135_;
wire [17:0] _136_;
wire _137_;
wire [16:0] _138_;
wire [17:0] _139_;
wire [18:0] _140_;
wire [17:0] _141_;
wire [17:0] _142_;
wire _143_;
wire [17:0] _144_;
wire [18:0] _145_;
wire [18:0] _146_;
wire [23:0] _147_;
wire [23:0] _148_;
wire _149_;
wire [22:0] _150_;
wire [23:0] _151_;
wire [24:0] _152_;
wire [3:0] _153_;
wire [3:0] _154_;
wire [3:0] _155_;
wire [3:0] _156_;
wire [3:0] _157_;
wire [3:0] _158_;
wire [3:0] _159_;
wire [3:0] _160_;
wire [3:0] _161_;
wire [3:0] _162_;
wire [3:0] _163_;
wire [3:0] _164_;
wire [3:0] _165_;
wire [3:0] _166_;
wire [3:0] _167_;
wire [3:0] _168_;
wire [3:0] _169_;
wire [3:0] _170_;
wire [3:0] _171_;
wire [3:0] _172_;
wire [3:0] _173_;
wire [3:0] _174_;
wire [3:0] _175_;
wire [3:0] _176_;
wire [3:0] _177_;
wire [3:0] _178_;
wire [3:0] _179_;
wire [3:0] _180_;
wire [3:0] _181_;
wire [3:0] _182_;
wire [3:0] _183_;
wire [3:0] _184_;
wire [3:0] _185_;
wire [3:0] _186_;
wire [3:0] _187_;
wire [3:0] _188_;
wire [3:0] _189_;
wire [3:0] _190_;
wire [3:0] _191_;
wire [3:0] _192_;
wire [3:0] _193_;
wire [3:0] _194_;
wire [3:0] _195_;
wire [3:0] _196_;
wire [3:0] _197_;
wire [3:0] _198_;
wire [3:0] _199_;
wire [3:0] _200_;
wire [3:0] _201_;
wire [3:0] _202_;
wire [3:0] _203_;
wire [3:0] _204_;
wire [3:0] _205_;
wire [3:0] _206_;
wire [17:0] _207_;
wire [17:0] _208_;
wire _209_;
wire [17:0] _210_;
wire [18:0] _211_;
wire [18:0] _212_;
wire [1:0] _213_;
wire [1:0] _214_;
wire _215_;
wire [1:0] _216_;
wire [2:0] _217_;
wire [2:0] _218_;
wire _219_;
wire _220_;
wire _221_;
wire _222_;
wire _223_;
wire _224_;
wire _225_;
wire _226_;
wire _227_;
wire _228_;
wire _229_;
wire _230_;
wire _231_;
wire _232_;
wire _233_;
wire _234_;
wire _235_;
wire _236_;
wire _237_;
wire _238_;
wire _239_;
wire _240_;
wire _241_;
wire _242_;
wire _243_;
wire _244_;
wire _245_;
wire _246_;
wire _247_;
wire _248_;
wire _249_;
wire _250_;
wire _251_;
wire _252_;
wire _253_;
wire _254_;
wire _255_;
wire _256_;
wire _257_;
wire _258_;
wire _259_;
wire _260_;
wire _261_;
wire _262_;
wire _263_;
wire _264_;
wire _265_;
wire _266_;
wire \add_18ns_18ns_18_2_1_U5.ce ;
wire \add_18ns_18ns_18_2_1_U5.clk ;
wire [17:0] \add_18ns_18ns_18_2_1_U5.din0 ;
wire [17:0] \add_18ns_18ns_18_2_1_U5.din1 ;
wire [17:0] \add_18ns_18ns_18_2_1_U5.dout ;
wire \add_18ns_18ns_18_2_1_U5.reset ;
wire [17:0] \add_18ns_18ns_18_2_1_U5.top_add_18ns_18ns_18_2_1_Adder_2_U.a ;
wire [17:0] \add_18ns_18ns_18_2_1_U5.top_add_18ns_18ns_18_2_1_Adder_2_U.ain_s0 ;
wire [17:0] \add_18ns_18ns_18_2_1_U5.top_add_18ns_18ns_18_2_1_Adder_2_U.b ;
wire [17:0] \add_18ns_18ns_18_2_1_U5.top_add_18ns_18ns_18_2_1_Adder_2_U.bin_s0 ;
wire \add_18ns_18ns_18_2_1_U5.top_add_18ns_18ns_18_2_1_Adder_2_U.ce ;
wire \add_18ns_18ns_18_2_1_U5.top_add_18ns_18ns_18_2_1_Adder_2_U.clk ;
wire \add_18ns_18ns_18_2_1_U5.top_add_18ns_18ns_18_2_1_Adder_2_U.facout_s1 ;
wire \add_18ns_18ns_18_2_1_U5.top_add_18ns_18ns_18_2_1_Adder_2_U.facout_s2 ;
wire [8:0] \add_18ns_18ns_18_2_1_U5.top_add_18ns_18ns_18_2_1_Adder_2_U.fas_s1 ;
wire [8:0] \add_18ns_18ns_18_2_1_U5.top_add_18ns_18ns_18_2_1_Adder_2_U.fas_s2 ;
wire \add_18ns_18ns_18_2_1_U5.top_add_18ns_18ns_18_2_1_Adder_2_U.reset ;
wire [17:0] \add_18ns_18ns_18_2_1_U5.top_add_18ns_18ns_18_2_1_Adder_2_U.s ;
wire [8:0] \add_18ns_18ns_18_2_1_U5.top_add_18ns_18ns_18_2_1_Adder_2_U.u1.a ;
wire [8:0] \add_18ns_18ns_18_2_1_U5.top_add_18ns_18ns_18_2_1_Adder_2_U.u1.b ;
wire \add_18ns_18ns_18_2_1_U5.top_add_18ns_18ns_18_2_1_Adder_2_U.u1.cin ;
wire \add_18ns_18ns_18_2_1_U5.top_add_18ns_18ns_18_2_1_Adder_2_U.u1.cout ;
wire [8:0] \add_18ns_18ns_18_2_1_U5.top_add_18ns_18ns_18_2_1_Adder_2_U.u1.s ;
wire [8:0] \add_18ns_18ns_18_2_1_U5.top_add_18ns_18ns_18_2_1_Adder_2_U.u2.a ;
wire [8:0] \add_18ns_18ns_18_2_1_U5.top_add_18ns_18ns_18_2_1_Adder_2_U.u2.b ;
wire \add_18ns_18ns_18_2_1_U5.top_add_18ns_18ns_18_2_1_Adder_2_U.u2.cin ;
wire \add_18ns_18ns_18_2_1_U5.top_add_18ns_18ns_18_2_1_Adder_2_U.u2.cout ;
wire [8:0] \add_18ns_18ns_18_2_1_U5.top_add_18ns_18ns_18_2_1_Adder_2_U.u2.s ;
wire \add_18ns_18s_18_2_1_U4.ce ;
wire \add_18ns_18s_18_2_1_U4.clk ;
wire [17:0] \add_18ns_18s_18_2_1_U4.din0 ;
wire [17:0] \add_18ns_18s_18_2_1_U4.din1 ;
wire [17:0] \add_18ns_18s_18_2_1_U4.dout ;
wire \add_18ns_18s_18_2_1_U4.reset ;
wire [17:0] \add_18ns_18s_18_2_1_U4.top_add_18ns_18s_18_2_1_Adder_1_U.a ;
wire [17:0] \add_18ns_18s_18_2_1_U4.top_add_18ns_18s_18_2_1_Adder_1_U.ain_s0 ;
wire [17:0] \add_18ns_18s_18_2_1_U4.top_add_18ns_18s_18_2_1_Adder_1_U.b ;
wire [17:0] \add_18ns_18s_18_2_1_U4.top_add_18ns_18s_18_2_1_Adder_1_U.bin_s0 ;
wire \add_18ns_18s_18_2_1_U4.top_add_18ns_18s_18_2_1_Adder_1_U.ce ;
wire \add_18ns_18s_18_2_1_U4.top_add_18ns_18s_18_2_1_Adder_1_U.clk ;
wire \add_18ns_18s_18_2_1_U4.top_add_18ns_18s_18_2_1_Adder_1_U.facout_s1 ;
wire \add_18ns_18s_18_2_1_U4.top_add_18ns_18s_18_2_1_Adder_1_U.facout_s2 ;
wire [8:0] \add_18ns_18s_18_2_1_U4.top_add_18ns_18s_18_2_1_Adder_1_U.fas_s1 ;
wire [8:0] \add_18ns_18s_18_2_1_U4.top_add_18ns_18s_18_2_1_Adder_1_U.fas_s2 ;
wire \add_18ns_18s_18_2_1_U4.top_add_18ns_18s_18_2_1_Adder_1_U.reset ;
wire [17:0] \add_18ns_18s_18_2_1_U4.top_add_18ns_18s_18_2_1_Adder_1_U.s ;
wire [8:0] \add_18ns_18s_18_2_1_U4.top_add_18ns_18s_18_2_1_Adder_1_U.u1.a ;
wire [8:0] \add_18ns_18s_18_2_1_U4.top_add_18ns_18s_18_2_1_Adder_1_U.u1.b ;
wire \add_18ns_18s_18_2_1_U4.top_add_18ns_18s_18_2_1_Adder_1_U.u1.cin ;
wire \add_18ns_18s_18_2_1_U4.top_add_18ns_18s_18_2_1_Adder_1_U.u1.cout ;
wire [8:0] \add_18ns_18s_18_2_1_U4.top_add_18ns_18s_18_2_1_Adder_1_U.u1.s ;
wire [8:0] \add_18ns_18s_18_2_1_U4.top_add_18ns_18s_18_2_1_Adder_1_U.u2.a ;
wire [8:0] \add_18ns_18s_18_2_1_U4.top_add_18ns_18s_18_2_1_Adder_1_U.u2.b ;
wire \add_18ns_18s_18_2_1_U4.top_add_18ns_18s_18_2_1_Adder_1_U.u2.cin ;
wire \add_18ns_18s_18_2_1_U4.top_add_18ns_18s_18_2_1_Adder_1_U.u2.cout ;
wire [8:0] \add_18ns_18s_18_2_1_U4.top_add_18ns_18s_18_2_1_Adder_1_U.u2.s ;
wire \add_22s_22s_22_2_1_U7.ce ;
wire \add_22s_22s_22_2_1_U7.clk ;
wire [21:0] \add_22s_22s_22_2_1_U7.din0 ;
wire [21:0] \add_22s_22s_22_2_1_U7.din1 ;
wire [21:0] \add_22s_22s_22_2_1_U7.dout ;
wire \add_22s_22s_22_2_1_U7.reset ;
wire [21:0] \add_22s_22s_22_2_1_U7.top_add_22s_22s_22_2_1_Adder_4_U.a ;
wire [21:0] \add_22s_22s_22_2_1_U7.top_add_22s_22s_22_2_1_Adder_4_U.ain_s0 ;
wire [21:0] \add_22s_22s_22_2_1_U7.top_add_22s_22s_22_2_1_Adder_4_U.b ;
wire [21:0] \add_22s_22s_22_2_1_U7.top_add_22s_22s_22_2_1_Adder_4_U.bin_s0 ;
wire \add_22s_22s_22_2_1_U7.top_add_22s_22s_22_2_1_Adder_4_U.ce ;
wire \add_22s_22s_22_2_1_U7.top_add_22s_22s_22_2_1_Adder_4_U.clk ;
wire \add_22s_22s_22_2_1_U7.top_add_22s_22s_22_2_1_Adder_4_U.facout_s1 ;
wire \add_22s_22s_22_2_1_U7.top_add_22s_22s_22_2_1_Adder_4_U.facout_s2 ;
wire [10:0] \add_22s_22s_22_2_1_U7.top_add_22s_22s_22_2_1_Adder_4_U.fas_s1 ;
wire [10:0] \add_22s_22s_22_2_1_U7.top_add_22s_22s_22_2_1_Adder_4_U.fas_s2 ;
wire \add_22s_22s_22_2_1_U7.top_add_22s_22s_22_2_1_Adder_4_U.reset ;
wire [21:0] \add_22s_22s_22_2_1_U7.top_add_22s_22s_22_2_1_Adder_4_U.s ;
wire [10:0] \add_22s_22s_22_2_1_U7.top_add_22s_22s_22_2_1_Adder_4_U.u1.a ;
wire [10:0] \add_22s_22s_22_2_1_U7.top_add_22s_22s_22_2_1_Adder_4_U.u1.b ;
wire \add_22s_22s_22_2_1_U7.top_add_22s_22s_22_2_1_Adder_4_U.u1.cin ;
wire \add_22s_22s_22_2_1_U7.top_add_22s_22s_22_2_1_Adder_4_U.u1.cout ;
wire [10:0] \add_22s_22s_22_2_1_U7.top_add_22s_22s_22_2_1_Adder_4_U.u1.s ;
wire [10:0] \add_22s_22s_22_2_1_U7.top_add_22s_22s_22_2_1_Adder_4_U.u2.a ;
wire [10:0] \add_22s_22s_22_2_1_U7.top_add_22s_22s_22_2_1_Adder_4_U.u2.b ;
wire \add_22s_22s_22_2_1_U7.top_add_22s_22s_22_2_1_Adder_4_U.u2.cin ;
wire \add_22s_22s_22_2_1_U7.top_add_22s_22s_22_2_1_Adder_4_U.u2.cout ;
wire [10:0] \add_22s_22s_22_2_1_U7.top_add_22s_22s_22_2_1_Adder_4_U.u2.s ;
wire \add_2ns_2ns_2_2_1_U17.ce ;
wire \add_2ns_2ns_2_2_1_U17.clk ;
wire [1:0] \add_2ns_2ns_2_2_1_U17.din0 ;
wire [1:0] \add_2ns_2ns_2_2_1_U17.din1 ;
wire [1:0] \add_2ns_2ns_2_2_1_U17.dout ;
wire \add_2ns_2ns_2_2_1_U17.reset ;
wire [1:0] \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_11_U.a ;
wire [1:0] \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_11_U.ain_s0 ;
wire [1:0] \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_11_U.b ;
wire [1:0] \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_11_U.bin_s0 ;
wire \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_11_U.ce ;
wire \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_11_U.clk ;
wire \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_11_U.facout_s1 ;
wire \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_11_U.facout_s2 ;
wire \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_11_U.fas_s1 ;
wire \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_11_U.fas_s2 ;
wire \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_11_U.reset ;
wire [1:0] \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_11_U.s ;
wire \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_11_U.u1.a ;
wire \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_11_U.u1.b ;
wire \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_11_U.u1.cin ;
wire \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_11_U.u1.cout ;
wire \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_11_U.u1.s ;
wire \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_11_U.u2.a ;
wire \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_11_U.u2.b ;
wire \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_11_U.u2.cin ;
wire \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_11_U.u2.cout ;
wire \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_11_U.u2.s ;
wire \add_2ns_2ns_2_2_1_U19.ce ;
wire \add_2ns_2ns_2_2_1_U19.clk ;
wire [1:0] \add_2ns_2ns_2_2_1_U19.din0 ;
wire [1:0] \add_2ns_2ns_2_2_1_U19.din1 ;
wire [1:0] \add_2ns_2ns_2_2_1_U19.dout ;
wire \add_2ns_2ns_2_2_1_U19.reset ;
wire [1:0] \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_11_U.a ;
wire [1:0] \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_11_U.ain_s0 ;
wire [1:0] \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_11_U.b ;
wire [1:0] \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_11_U.bin_s0 ;
wire \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_11_U.ce ;
wire \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_11_U.clk ;
wire \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_11_U.facout_s1 ;
wire \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_11_U.facout_s2 ;
wire \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_11_U.fas_s1 ;
wire \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_11_U.fas_s2 ;
wire \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_11_U.reset ;
wire [1:0] \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_11_U.s ;
wire \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_11_U.u1.a ;
wire \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_11_U.u1.b ;
wire \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_11_U.u1.cin ;
wire \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_11_U.u1.cout ;
wire \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_11_U.u1.s ;
wire \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_11_U.u2.a ;
wire \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_11_U.u2.b ;
wire \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_11_U.u2.cin ;
wire \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_11_U.u2.cout ;
wire \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_11_U.u2.s ;
wire \add_32ns_32ns_32_2_1_U10.ce ;
wire \add_32ns_32ns_32_2_1_U10.clk ;
wire [31:0] \add_32ns_32ns_32_2_1_U10.din0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U10.din1 ;
wire [31:0] \add_32ns_32ns_32_2_1_U10.dout ;
wire \add_32ns_32ns_32_2_1_U10.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.a ;
wire [31:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.b ;
wire [31:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s0 ;
wire \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.ce ;
wire \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.clk ;
wire \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.facout_s1 ;
wire \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.facout_s2 ;
wire [15:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s1 ;
wire [15:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s2 ;
wire \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.b ;
wire \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cin ;
wire \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.b ;
wire \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cin ;
wire \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.s ;
wire \add_32ns_32ns_32_2_1_U12.ce ;
wire \add_32ns_32ns_32_2_1_U12.clk ;
wire [31:0] \add_32ns_32ns_32_2_1_U12.din0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U12.din1 ;
wire [31:0] \add_32ns_32ns_32_2_1_U12.dout ;
wire \add_32ns_32ns_32_2_1_U12.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.a ;
wire [31:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.b ;
wire [31:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s0 ;
wire \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.ce ;
wire \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.clk ;
wire \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.facout_s1 ;
wire \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.facout_s2 ;
wire [15:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s1 ;
wire [15:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s2 ;
wire \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.b ;
wire \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cin ;
wire \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.b ;
wire \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cin ;
wire \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.s ;
wire \add_32ns_32ns_32_2_1_U14.ce ;
wire \add_32ns_32ns_32_2_1_U14.clk ;
wire [31:0] \add_32ns_32ns_32_2_1_U14.din0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U14.din1 ;
wire [31:0] \add_32ns_32ns_32_2_1_U14.dout ;
wire \add_32ns_32ns_32_2_1_U14.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.a ;
wire [31:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.b ;
wire [31:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s0 ;
wire \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.ce ;
wire \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.clk ;
wire \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.facout_s1 ;
wire \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.facout_s2 ;
wire [15:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s1 ;
wire [15:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s2 ;
wire \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.b ;
wire \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cin ;
wire \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.b ;
wire \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cin ;
wire \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.s ;
wire \add_32ns_32ns_32_2_1_U16.ce ;
wire \add_32ns_32ns_32_2_1_U16.clk ;
wire [31:0] \add_32ns_32ns_32_2_1_U16.din0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U16.din1 ;
wire [31:0] \add_32ns_32ns_32_2_1_U16.dout ;
wire \add_32ns_32ns_32_2_1_U16.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.a ;
wire [31:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.b ;
wire [31:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s0 ;
wire \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.ce ;
wire \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.clk ;
wire \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.facout_s1 ;
wire \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.facout_s2 ;
wire [15:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s1 ;
wire [15:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s2 ;
wire \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.b ;
wire \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cin ;
wire \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.b ;
wire \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cin ;
wire \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.s ;
wire \add_32ns_32ns_32_2_1_U18.ce ;
wire \add_32ns_32ns_32_2_1_U18.clk ;
wire [31:0] \add_32ns_32ns_32_2_1_U18.din0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U18.din1 ;
wire [31:0] \add_32ns_32ns_32_2_1_U18.dout ;
wire \add_32ns_32ns_32_2_1_U18.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.a ;
wire [31:0] \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.b ;
wire [31:0] \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s0 ;
wire \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.ce ;
wire \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.clk ;
wire \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.facout_s1 ;
wire \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.facout_s2 ;
wire [15:0] \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s1 ;
wire [15:0] \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s2 ;
wire \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.b ;
wire \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cin ;
wire \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.b ;
wire \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cin ;
wire \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.s ;
wire \add_32ns_32s_32_2_1_U13.ce ;
wire \add_32ns_32s_32_2_1_U13.clk ;
wire [31:0] \add_32ns_32s_32_2_1_U13.din0 ;
wire [31:0] \add_32ns_32s_32_2_1_U13.din1 ;
wire [31:0] \add_32ns_32s_32_2_1_U13.dout ;
wire \add_32ns_32s_32_2_1_U13.reset ;
wire [31:0] \add_32ns_32s_32_2_1_U13.top_add_32ns_32s_32_2_1_Adder_9_U.a ;
wire [31:0] \add_32ns_32s_32_2_1_U13.top_add_32ns_32s_32_2_1_Adder_9_U.ain_s0 ;
wire [31:0] \add_32ns_32s_32_2_1_U13.top_add_32ns_32s_32_2_1_Adder_9_U.b ;
wire [31:0] \add_32ns_32s_32_2_1_U13.top_add_32ns_32s_32_2_1_Adder_9_U.bin_s0 ;
wire \add_32ns_32s_32_2_1_U13.top_add_32ns_32s_32_2_1_Adder_9_U.ce ;
wire \add_32ns_32s_32_2_1_U13.top_add_32ns_32s_32_2_1_Adder_9_U.clk ;
wire \add_32ns_32s_32_2_1_U13.top_add_32ns_32s_32_2_1_Adder_9_U.facout_s1 ;
wire \add_32ns_32s_32_2_1_U13.top_add_32ns_32s_32_2_1_Adder_9_U.facout_s2 ;
wire [15:0] \add_32ns_32s_32_2_1_U13.top_add_32ns_32s_32_2_1_Adder_9_U.fas_s1 ;
wire [15:0] \add_32ns_32s_32_2_1_U13.top_add_32ns_32s_32_2_1_Adder_9_U.fas_s2 ;
wire \add_32ns_32s_32_2_1_U13.top_add_32ns_32s_32_2_1_Adder_9_U.reset ;
wire [31:0] \add_32ns_32s_32_2_1_U13.top_add_32ns_32s_32_2_1_Adder_9_U.s ;
wire [15:0] \add_32ns_32s_32_2_1_U13.top_add_32ns_32s_32_2_1_Adder_9_U.u1.a ;
wire [15:0] \add_32ns_32s_32_2_1_U13.top_add_32ns_32s_32_2_1_Adder_9_U.u1.b ;
wire \add_32ns_32s_32_2_1_U13.top_add_32ns_32s_32_2_1_Adder_9_U.u1.cin ;
wire \add_32ns_32s_32_2_1_U13.top_add_32ns_32s_32_2_1_Adder_9_U.u1.cout ;
wire [15:0] \add_32ns_32s_32_2_1_U13.top_add_32ns_32s_32_2_1_Adder_9_U.u1.s ;
wire [15:0] \add_32ns_32s_32_2_1_U13.top_add_32ns_32s_32_2_1_Adder_9_U.u2.a ;
wire [15:0] \add_32ns_32s_32_2_1_U13.top_add_32ns_32s_32_2_1_Adder_9_U.u2.b ;
wire \add_32ns_32s_32_2_1_U13.top_add_32ns_32s_32_2_1_Adder_9_U.u2.cin ;
wire \add_32ns_32s_32_2_1_U13.top_add_32ns_32s_32_2_1_Adder_9_U.u2.cout ;
wire [15:0] \add_32ns_32s_32_2_1_U13.top_add_32ns_32s_32_2_1_Adder_9_U.u2.s ;
wire \add_32s_32ns_32_2_1_U20.ce ;
wire \add_32s_32ns_32_2_1_U20.clk ;
wire [31:0] \add_32s_32ns_32_2_1_U20.din0 ;
wire [31:0] \add_32s_32ns_32_2_1_U20.din1 ;
wire [31:0] \add_32s_32ns_32_2_1_U20.dout ;
wire \add_32s_32ns_32_2_1_U20.reset ;
wire [31:0] \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_5_U.a ;
wire [31:0] \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_5_U.ain_s0 ;
wire [31:0] \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_5_U.b ;
wire [31:0] \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_5_U.bin_s0 ;
wire \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_5_U.ce ;
wire \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_5_U.clk ;
wire \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_5_U.facout_s1 ;
wire \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_5_U.facout_s2 ;
wire [15:0] \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_5_U.fas_s1 ;
wire [15:0] \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_5_U.fas_s2 ;
wire \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_5_U.reset ;
wire [31:0] \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_5_U.s ;
wire [15:0] \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_5_U.u1.a ;
wire [15:0] \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_5_U.u1.b ;
wire \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_5_U.u1.cin ;
wire \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_5_U.u1.cout ;
wire [15:0] \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_5_U.u1.s ;
wire [15:0] \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_5_U.u2.a ;
wire [15:0] \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_5_U.u2.b ;
wire \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_5_U.u2.cin ;
wire \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_5_U.u2.cout ;
wire [15:0] \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_5_U.u2.s ;
wire \add_32s_32ns_32_2_1_U8.ce ;
wire \add_32s_32ns_32_2_1_U8.clk ;
wire [31:0] \add_32s_32ns_32_2_1_U8.din0 ;
wire [31:0] \add_32s_32ns_32_2_1_U8.din1 ;
wire [31:0] \add_32s_32ns_32_2_1_U8.dout ;
wire \add_32s_32ns_32_2_1_U8.reset ;
wire [31:0] \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.a ;
wire [31:0] \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.ain_s0 ;
wire [31:0] \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.b ;
wire [31:0] \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.bin_s0 ;
wire \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.ce ;
wire \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.clk ;
wire \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.facout_s1 ;
wire \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.facout_s2 ;
wire [15:0] \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.fas_s1 ;
wire [15:0] \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.fas_s2 ;
wire \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.reset ;
wire [31:0] \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.s ;
wire [15:0] \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.u1.a ;
wire [15:0] \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.u1.b ;
wire \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.u1.cin ;
wire \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.u1.cout ;
wire [15:0] \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.u1.s ;
wire [15:0] \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.u2.a ;
wire [15:0] \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.u2.b ;
wire \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.u2.cin ;
wire \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.u2.cout ;
wire [15:0] \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.u2.s ;
wire \add_35s_35s_35_2_1_U15.ce ;
wire \add_35s_35s_35_2_1_U15.clk ;
wire [34:0] \add_35s_35s_35_2_1_U15.din0 ;
wire [34:0] \add_35s_35s_35_2_1_U15.din1 ;
wire [34:0] \add_35s_35s_35_2_1_U15.dout ;
wire \add_35s_35s_35_2_1_U15.reset ;
wire [34:0] \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_10_U.a ;
wire [34:0] \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_10_U.ain_s0 ;
wire [34:0] \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_10_U.b ;
wire [34:0] \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_10_U.bin_s0 ;
wire \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_10_U.ce ;
wire \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_10_U.clk ;
wire \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_10_U.facout_s1 ;
wire \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_10_U.facout_s2 ;
wire [16:0] \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_10_U.fas_s1 ;
wire [17:0] \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_10_U.fas_s2 ;
wire \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_10_U.reset ;
wire [34:0] \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_10_U.s ;
wire [16:0] \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_10_U.u1.a ;
wire [16:0] \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_10_U.u1.b ;
wire \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_10_U.u1.cin ;
wire \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_10_U.u1.cout ;
wire [16:0] \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_10_U.u1.s ;
wire [17:0] \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_10_U.u2.a ;
wire [17:0] \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_10_U.u2.b ;
wire \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_10_U.u2.cin ;
wire \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_10_U.u2.cout ;
wire [17:0] \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_10_U.u2.s ;
wire \add_36s_36s_36_2_1_U9.ce ;
wire \add_36s_36s_36_2_1_U9.clk ;
wire [35:0] \add_36s_36s_36_2_1_U9.din0 ;
wire [35:0] \add_36s_36s_36_2_1_U9.din1 ;
wire [35:0] \add_36s_36s_36_2_1_U9.dout ;
wire \add_36s_36s_36_2_1_U9.reset ;
wire [35:0] \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_6_U.a ;
wire [35:0] \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_6_U.ain_s0 ;
wire [35:0] \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_6_U.b ;
wire [35:0] \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_6_U.bin_s0 ;
wire \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_6_U.ce ;
wire \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_6_U.clk ;
wire \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_6_U.facout_s1 ;
wire \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_6_U.facout_s2 ;
wire [17:0] \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_6_U.fas_s1 ;
wire [17:0] \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_6_U.fas_s2 ;
wire \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_6_U.reset ;
wire [35:0] \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_6_U.s ;
wire [17:0] \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_6_U.u1.a ;
wire [17:0] \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_6_U.u1.b ;
wire \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_6_U.u1.cin ;
wire \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_6_U.u1.cout ;
wire [17:0] \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_6_U.u1.s ;
wire [17:0] \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_6_U.u2.a ;
wire [17:0] \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_6_U.u2.b ;
wire \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_6_U.u2.cin ;
wire \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_6_U.u2.cout ;
wire [17:0] \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_6_U.u2.s ;
wire \add_47s_47s_47_2_1_U11.ce ;
wire \add_47s_47s_47_2_1_U11.clk ;
wire [46:0] \add_47s_47s_47_2_1_U11.din0 ;
wire [46:0] \add_47s_47s_47_2_1_U11.din1 ;
wire [46:0] \add_47s_47s_47_2_1_U11.dout ;
wire \add_47s_47s_47_2_1_U11.reset ;
wire [46:0] \add_47s_47s_47_2_1_U11.top_add_47s_47s_47_2_1_Adder_8_U.a ;
wire [46:0] \add_47s_47s_47_2_1_U11.top_add_47s_47s_47_2_1_Adder_8_U.ain_s0 ;
wire [46:0] \add_47s_47s_47_2_1_U11.top_add_47s_47s_47_2_1_Adder_8_U.b ;
wire [46:0] \add_47s_47s_47_2_1_U11.top_add_47s_47s_47_2_1_Adder_8_U.bin_s0 ;
wire \add_47s_47s_47_2_1_U11.top_add_47s_47s_47_2_1_Adder_8_U.ce ;
wire \add_47s_47s_47_2_1_U11.top_add_47s_47s_47_2_1_Adder_8_U.clk ;
wire \add_47s_47s_47_2_1_U11.top_add_47s_47s_47_2_1_Adder_8_U.facout_s1 ;
wire \add_47s_47s_47_2_1_U11.top_add_47s_47s_47_2_1_Adder_8_U.facout_s2 ;
wire [22:0] \add_47s_47s_47_2_1_U11.top_add_47s_47s_47_2_1_Adder_8_U.fas_s1 ;
wire [23:0] \add_47s_47s_47_2_1_U11.top_add_47s_47s_47_2_1_Adder_8_U.fas_s2 ;
wire \add_47s_47s_47_2_1_U11.top_add_47s_47s_47_2_1_Adder_8_U.reset ;
wire [46:0] \add_47s_47s_47_2_1_U11.top_add_47s_47s_47_2_1_Adder_8_U.s ;
wire [22:0] \add_47s_47s_47_2_1_U11.top_add_47s_47s_47_2_1_Adder_8_U.u1.a ;
wire [22:0] \add_47s_47s_47_2_1_U11.top_add_47s_47s_47_2_1_Adder_8_U.u1.b ;
wire \add_47s_47s_47_2_1_U11.top_add_47s_47s_47_2_1_Adder_8_U.u1.cin ;
wire \add_47s_47s_47_2_1_U11.top_add_47s_47s_47_2_1_Adder_8_U.u1.cout ;
wire [22:0] \add_47s_47s_47_2_1_U11.top_add_47s_47s_47_2_1_Adder_8_U.u1.s ;
wire [23:0] \add_47s_47s_47_2_1_U11.top_add_47s_47s_47_2_1_Adder_8_U.u2.a ;
wire [23:0] \add_47s_47s_47_2_1_U11.top_add_47s_47s_47_2_1_Adder_8_U.u2.b ;
wire \add_47s_47s_47_2_1_U11.top_add_47s_47s_47_2_1_Adder_8_U.u2.cin ;
wire \add_47s_47s_47_2_1_U11.top_add_47s_47s_47_2_1_Adder_8_U.u2.cout ;
wire [23:0] \add_47s_47s_47_2_1_U11.top_add_47s_47s_47_2_1_Adder_8_U.u2.s ;
wire ap_CS_fsm_state1;
wire ap_CS_fsm_state10;
wire ap_CS_fsm_state11;
wire ap_CS_fsm_state12;
wire ap_CS_fsm_state13;
wire ap_CS_fsm_state14;
wire ap_CS_fsm_state15;
wire ap_CS_fsm_state16;
wire ap_CS_fsm_state17;
wire ap_CS_fsm_state18;
wire ap_CS_fsm_state19;
wire ap_CS_fsm_state2;
wire ap_CS_fsm_state20;
wire ap_CS_fsm_state21;
wire ap_CS_fsm_state22;
wire ap_CS_fsm_state23;
wire ap_CS_fsm_state24;
wire ap_CS_fsm_state25;
wire ap_CS_fsm_state26;
wire ap_CS_fsm_state27;
wire ap_CS_fsm_state28;
wire ap_CS_fsm_state29;
wire ap_CS_fsm_state3;
wire ap_CS_fsm_state30;
wire ap_CS_fsm_state31;
wire ap_CS_fsm_state32;
wire ap_CS_fsm_state33;
wire ap_CS_fsm_state34;
wire ap_CS_fsm_state35;
wire ap_CS_fsm_state36;
wire ap_CS_fsm_state37;
wire ap_CS_fsm_state38;
wire ap_CS_fsm_state39;
wire ap_CS_fsm_state40;
wire ap_CS_fsm_state41;
wire ap_CS_fsm_state42;
wire ap_CS_fsm_state9;
wire [41:0] ap_NS_fsm;
wire ap_clk;
wire ap_done;
wire ap_idle;
wire ap_ready;
wire ap_rst;
wire ap_start;
wire \ashr_4ns_4ns_4_7_1_U2.ce ;
wire \ashr_4ns_4ns_4_7_1_U2.clk ;
wire [3:0] \ashr_4ns_4ns_4_7_1_U2.din0 ;
wire [3:0] \ashr_4ns_4ns_4_7_1_U2.din1 ;
wire [3:0] \ashr_4ns_4ns_4_7_1_U2.din1_cast ;
wire [3:0] \ashr_4ns_4ns_4_7_1_U2.din1_mask ;
wire [3:0] \ashr_4ns_4ns_4_7_1_U2.dout ;
wire \ashr_4ns_4ns_4_7_1_U2.reset ;
wire [3:0] grp_fu_227_p2;
wire [3:0] grp_fu_233_p2;
wire [3:0] grp_fu_237_p2;
wire [17:0] grp_fu_257_p0;
wire [17:0] grp_fu_257_p1;
wire [17:0] grp_fu_257_p2;
wire [17:0] grp_fu_271_p2;
wire [35:0] grp_fu_294_p0;
wire [35:0] grp_fu_294_p1;
wire [35:0] grp_fu_294_p2;
wire [21:0] grp_fu_315_p0;
wire [21:0] grp_fu_315_p1;
wire [21:0] grp_fu_315_p2;
wire [31:0] grp_fu_380_p0;
wire [31:0] grp_fu_380_p2;
wire [35:0] grp_fu_476_p0;
wire [35:0] grp_fu_476_p1;
wire [35:0] grp_fu_476_p2;
wire [31:0] grp_fu_497_p2;
wire [46:0] grp_fu_536_p0;
wire [46:0] grp_fu_536_p1;
wire [46:0] grp_fu_536_p2;
wire [31:0] grp_fu_562_p2;
wire [31:0] grp_fu_590_p1;
wire [31:0] grp_fu_590_p2;
wire [31:0] grp_fu_599_p1;
wire [31:0] grp_fu_599_p2;
wire [34:0] grp_fu_619_p0;
wire [34:0] grp_fu_619_p1;
wire [34:0] grp_fu_619_p2;
wire [31:0] grp_fu_659_p2;
wire [1:0] grp_fu_676_p1;
wire [1:0] grp_fu_676_p2;
wire [31:0] grp_fu_708_p2;
wire [1:0] grp_fu_713_p2;
wire [31:0] grp_fu_720_p0;
wire [31:0] grp_fu_720_p2;
wire icmp_ln768_fu_367_p2;
wire icmp_ln786_fu_372_p2;
wire icmp_ln851_1_fu_482_p2;
wire icmp_ln851_2_fu_546_p2;
wire icmp_ln851_3_fu_629_p2;
wire icmp_ln851_fu_325_p2;
wire [1:0] op_0;
wire [3:0] op_1;
wire [3:0] op_10;
wire [3:0] op_11_V_fu_431_p3;
wire [31:0] op_12;
wire [7:0] op_13;
wire [1:0] op_14;
wire [3:0] op_15;
wire op_16_V_fu_653_p2;
wire op_17;
wire op_18;
wire [31:0] op_19;
wire [31:0] op_31;
wire op_31_ap_vld;
wire [31:0] op_4;
wire [3:0] op_6;
wire [7:0] op_8;
wire op_9;
wire or_ln384_fu_426_p2;
wire or_ln785_fu_386_p2;
wire or_ln786_fu_409_p2;
wire overflow_fu_395_p2;
wire p_Result_1_fu_502_p3;
wire p_Result_2_fu_567_p3;
wire p_Result_3_fu_681_p3;
wire p_Result_s_fu_439_p3;
wire [3:0] p_Val2_1_fu_401_p1;
wire [3:0] r_fu_241_p3;
wire [31:0] ret_V_6_fu_579_p3;
wire [31:0] ret_V_9_fu_693_p3;
wire [6:0] rhs_1_fu_279_p3;
wire [34:0] rhs_3_fu_465_p3;
wire [45:0] rhs_4_fu_525_p3;
wire [33:0] rhs_7_fu_608_p3;
wire [17:0] select_ln1192_fu_263_p3;
wire [31:0] select_ln353_1_fu_514_p3;
wire [31:0] select_ln353_fu_451_p3;
wire [3:0] select_ln384_fu_419_p3;
wire [1:0] select_ln69_1_fu_700_p3;
wire [1:0] select_ln69_fu_664_p3;
wire [31:0] select_ln850_1_fu_509_p3;
wire [31:0] select_ln850_2_fu_574_p3;
wire [31:0] select_ln850_3_fu_688_p3;
wire [31:0] select_ln850_fu_446_p3;
wire [3:0] sext_ln1192_fu_300_p0;
wire [34:0] sext_ln1193_1_fu_286_p1;
wire [15:0] sext_ln703_1_fu_250_p1;
wire [31:0] sext_ln703_3_fu_521_p0;
wire [3:0] sext_ln703_4_fu_604_p0;
wire [31:0] sext_ln831_fu_377_p1;
wire \shl_4ns_4ns_4_7_1_U3.ce ;
wire \shl_4ns_4ns_4_7_1_U3.clk ;
wire [3:0] \shl_4ns_4ns_4_7_1_U3.din0 ;
wire [3:0] \shl_4ns_4ns_4_7_1_U3.din1 ;
wire [3:0] \shl_4ns_4ns_4_7_1_U3.din1_cast ;
wire [3:0] \shl_4ns_4ns_4_7_1_U3.din1_mask ;
wire [3:0] \shl_4ns_4ns_4_7_1_U3.dout ;
wire \shl_4ns_4ns_4_7_1_U3.reset ;
wire \sub_36s_36ns_36_2_1_U6.ce ;
wire \sub_36s_36ns_36_2_1_U6.clk ;
wire [35:0] \sub_36s_36ns_36_2_1_U6.din0 ;
wire [35:0] \sub_36s_36ns_36_2_1_U6.din1 ;
wire [35:0] \sub_36s_36ns_36_2_1_U6.dout ;
wire \sub_36s_36ns_36_2_1_U6.reset ;
wire [35:0] \sub_36s_36ns_36_2_1_U6.top_sub_36s_36ns_36_2_1_Adder_3_U.a ;
wire [35:0] \sub_36s_36ns_36_2_1_U6.top_sub_36s_36ns_36_2_1_Adder_3_U.ain_s0 ;
wire [35:0] \sub_36s_36ns_36_2_1_U6.top_sub_36s_36ns_36_2_1_Adder_3_U.b ;
wire [35:0] \sub_36s_36ns_36_2_1_U6.top_sub_36s_36ns_36_2_1_Adder_3_U.bin_s0 ;
wire \sub_36s_36ns_36_2_1_U6.top_sub_36s_36ns_36_2_1_Adder_3_U.ce ;
wire \sub_36s_36ns_36_2_1_U6.top_sub_36s_36ns_36_2_1_Adder_3_U.clk ;
wire \sub_36s_36ns_36_2_1_U6.top_sub_36s_36ns_36_2_1_Adder_3_U.facout_s1 ;
wire \sub_36s_36ns_36_2_1_U6.top_sub_36s_36ns_36_2_1_Adder_3_U.facout_s2 ;
wire [17:0] \sub_36s_36ns_36_2_1_U6.top_sub_36s_36ns_36_2_1_Adder_3_U.fas_s1 ;
wire [17:0] \sub_36s_36ns_36_2_1_U6.top_sub_36s_36ns_36_2_1_Adder_3_U.fas_s2 ;
wire \sub_36s_36ns_36_2_1_U6.top_sub_36s_36ns_36_2_1_Adder_3_U.reset ;
wire [35:0] \sub_36s_36ns_36_2_1_U6.top_sub_36s_36ns_36_2_1_Adder_3_U.s ;
wire [17:0] \sub_36s_36ns_36_2_1_U6.top_sub_36s_36ns_36_2_1_Adder_3_U.u1.a ;
wire [17:0] \sub_36s_36ns_36_2_1_U6.top_sub_36s_36ns_36_2_1_Adder_3_U.u1.b ;
wire \sub_36s_36ns_36_2_1_U6.top_sub_36s_36ns_36_2_1_Adder_3_U.u1.cin ;
wire \sub_36s_36ns_36_2_1_U6.top_sub_36s_36ns_36_2_1_Adder_3_U.u1.cout ;
wire [17:0] \sub_36s_36ns_36_2_1_U6.top_sub_36s_36ns_36_2_1_Adder_3_U.u1.s ;
wire [17:0] \sub_36s_36ns_36_2_1_U6.top_sub_36s_36ns_36_2_1_Adder_3_U.u2.a ;
wire [17:0] \sub_36s_36ns_36_2_1_U6.top_sub_36s_36ns_36_2_1_Adder_3_U.u2.b ;
wire \sub_36s_36ns_36_2_1_U6.top_sub_36s_36ns_36_2_1_Adder_3_U.u2.cin ;
wire \sub_36s_36ns_36_2_1_U6.top_sub_36s_36ns_36_2_1_Adder_3_U.u2.cout ;
wire [17:0] \sub_36s_36ns_36_2_1_U6.top_sub_36s_36ns_36_2_1_Adder_3_U.u2.s ;
wire \sub_4ns_4ns_4_2_1_U1.ce ;
wire \sub_4ns_4ns_4_2_1_U1.clk ;
wire [3:0] \sub_4ns_4ns_4_2_1_U1.din0 ;
wire [3:0] \sub_4ns_4ns_4_2_1_U1.din1 ;
wire [3:0] \sub_4ns_4ns_4_2_1_U1.dout ;
wire \sub_4ns_4ns_4_2_1_U1.reset ;
wire [3:0] \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.a ;
wire [3:0] \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.ain_s0 ;
wire [3:0] \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.b ;
wire [3:0] \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.bin_s0 ;
wire \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.ce ;
wire \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.clk ;
wire \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.facout_s1 ;
wire \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.facout_s2 ;
wire [1:0] \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.fas_s1 ;
wire [1:0] \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.fas_s2 ;
wire \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.reset ;
wire [3:0] \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.s ;
wire [1:0] \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.u1.a ;
wire [1:0] \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.u1.b ;
wire \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.u1.cin ;
wire \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.u1.cout ;
wire [1:0] \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.u1.s ;
wire [1:0] \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.u2.a ;
wire [1:0] \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.u2.b ;
wire \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.u2.cin ;
wire \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.u2.cout ;
wire [1:0] \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.u2.s ;
wire [20:0] tmp_5_fu_304_p3;
wire trunc_ln69_1_fu_649_p1;
wire trunc_ln69_fu_645_p1;
wire [2:0] trunc_ln851_1_fu_458_p1;
wire [31:0] trunc_ln851_2_fu_542_p0;
wire [13:0] trunc_ln851_2_fu_542_p1;
wire [3:0] trunc_ln851_3_fu_625_p0;
wire [1:0] trunc_ln851_3_fu_625_p1;
wire [3:0] trunc_ln851_fu_321_p0;
wire [2:0] trunc_ln851_fu_321_p1;
wire underflow_fu_414_p2;
wire xor_ln785_fu_390_p2;
wire xor_ln786_fu_404_p2;


assign _047_ = icmp_ln851_1_reg_896 & ap_CS_fsm[22];
assign _048_ = icmp_ln851_2_reg_933 & ap_CS_fsm[27];
assign _049_ = icmp_ln851_3_reg_990 & ap_CS_fsm[36];
assign _050_ = ap_CS_fsm[17] & icmp_ln851_reg_805;
assign _051_ = p_Result_4_reg_734 & ap_CS_fsm[8];
assign _052_ = _055_ & ap_CS_fsm[8];
assign _053_ = _056_ & ap_CS_fsm[0];
assign _054_ = ap_start & ap_CS_fsm[0];
assign op_16_V_fu_653_p2 = op_4[0] & op_8[0];
assign overflow_fu_395_p2 = xor_ln785_fu_390_p2 & or_ln785_fu_386_p2;
assign underflow_fu_414_p2 = p_Result_5_reg_815 & or_ln786_fu_409_p2;
assign xor_ln786_fu_404_p2 = ~ p_Result_6_reg_821;
assign xor_ln785_fu_390_p2 = ~ p_Result_5_reg_815;
assign _055_ = ~ p_Result_4_reg_734;
assign _056_ = ~ ap_start;
always @(posedge \add_18ns_18ns_18_2_1_U5.top_add_18ns_18ns_18_2_1_Adder_2_U.clk )
\add_18ns_18ns_18_2_1_U5.top_add_18ns_18ns_18_2_1_Adder_2_U.bin_s1  <= _058_;
always @(posedge \add_18ns_18ns_18_2_1_U5.top_add_18ns_18ns_18_2_1_Adder_2_U.clk )
\add_18ns_18ns_18_2_1_U5.top_add_18ns_18ns_18_2_1_Adder_2_U.ain_s1  <= _057_;
always @(posedge \add_18ns_18ns_18_2_1_U5.top_add_18ns_18ns_18_2_1_Adder_2_U.clk )
\add_18ns_18ns_18_2_1_U5.top_add_18ns_18ns_18_2_1_Adder_2_U.sum_s1  <= _060_;
always @(posedge \add_18ns_18ns_18_2_1_U5.top_add_18ns_18ns_18_2_1_Adder_2_U.clk )
\add_18ns_18ns_18_2_1_U5.top_add_18ns_18ns_18_2_1_Adder_2_U.carry_s1  <= _059_;
assign _058_ = \add_18ns_18ns_18_2_1_U5.top_add_18ns_18ns_18_2_1_Adder_2_U.ce  ? \add_18ns_18ns_18_2_1_U5.top_add_18ns_18ns_18_2_1_Adder_2_U.b [17:9] : \add_18ns_18ns_18_2_1_U5.top_add_18ns_18ns_18_2_1_Adder_2_U.bin_s1 ;
assign _057_ = \add_18ns_18ns_18_2_1_U5.top_add_18ns_18ns_18_2_1_Adder_2_U.ce  ? \add_18ns_18ns_18_2_1_U5.top_add_18ns_18ns_18_2_1_Adder_2_U.a [17:9] : \add_18ns_18ns_18_2_1_U5.top_add_18ns_18ns_18_2_1_Adder_2_U.ain_s1 ;
assign _059_ = \add_18ns_18ns_18_2_1_U5.top_add_18ns_18ns_18_2_1_Adder_2_U.ce  ? \add_18ns_18ns_18_2_1_U5.top_add_18ns_18ns_18_2_1_Adder_2_U.facout_s1  : \add_18ns_18ns_18_2_1_U5.top_add_18ns_18ns_18_2_1_Adder_2_U.carry_s1 ;
assign _060_ = \add_18ns_18ns_18_2_1_U5.top_add_18ns_18ns_18_2_1_Adder_2_U.ce  ? \add_18ns_18ns_18_2_1_U5.top_add_18ns_18ns_18_2_1_Adder_2_U.fas_s1  : \add_18ns_18ns_18_2_1_U5.top_add_18ns_18ns_18_2_1_Adder_2_U.sum_s1 ;
assign _061_ = \add_18ns_18ns_18_2_1_U5.top_add_18ns_18ns_18_2_1_Adder_2_U.u1.a  + \add_18ns_18ns_18_2_1_U5.top_add_18ns_18ns_18_2_1_Adder_2_U.u1.b ;
assign { \add_18ns_18ns_18_2_1_U5.top_add_18ns_18ns_18_2_1_Adder_2_U.u1.cout , \add_18ns_18ns_18_2_1_U5.top_add_18ns_18ns_18_2_1_Adder_2_U.u1.s  } = _061_ + \add_18ns_18ns_18_2_1_U5.top_add_18ns_18ns_18_2_1_Adder_2_U.u1.cin ;
assign _062_ = \add_18ns_18ns_18_2_1_U5.top_add_18ns_18ns_18_2_1_Adder_2_U.u2.a  + \add_18ns_18ns_18_2_1_U5.top_add_18ns_18ns_18_2_1_Adder_2_U.u2.b ;
assign { \add_18ns_18ns_18_2_1_U5.top_add_18ns_18ns_18_2_1_Adder_2_U.u2.cout , \add_18ns_18ns_18_2_1_U5.top_add_18ns_18ns_18_2_1_Adder_2_U.u2.s  } = _062_ + \add_18ns_18ns_18_2_1_U5.top_add_18ns_18ns_18_2_1_Adder_2_U.u2.cin ;
always @(posedge \add_18ns_18s_18_2_1_U4.top_add_18ns_18s_18_2_1_Adder_1_U.clk )
\add_18ns_18s_18_2_1_U4.top_add_18ns_18s_18_2_1_Adder_1_U.bin_s1  <= _064_;
always @(posedge \add_18ns_18s_18_2_1_U4.top_add_18ns_18s_18_2_1_Adder_1_U.clk )
\add_18ns_18s_18_2_1_U4.top_add_18ns_18s_18_2_1_Adder_1_U.ain_s1  <= _063_;
always @(posedge \add_18ns_18s_18_2_1_U4.top_add_18ns_18s_18_2_1_Adder_1_U.clk )
\add_18ns_18s_18_2_1_U4.top_add_18ns_18s_18_2_1_Adder_1_U.sum_s1  <= _066_;
always @(posedge \add_18ns_18s_18_2_1_U4.top_add_18ns_18s_18_2_1_Adder_1_U.clk )
\add_18ns_18s_18_2_1_U4.top_add_18ns_18s_18_2_1_Adder_1_U.carry_s1  <= _065_;
assign _064_ = \add_18ns_18s_18_2_1_U4.top_add_18ns_18s_18_2_1_Adder_1_U.ce  ? \add_18ns_18s_18_2_1_U4.top_add_18ns_18s_18_2_1_Adder_1_U.b [17:9] : \add_18ns_18s_18_2_1_U4.top_add_18ns_18s_18_2_1_Adder_1_U.bin_s1 ;
assign _063_ = \add_18ns_18s_18_2_1_U4.top_add_18ns_18s_18_2_1_Adder_1_U.ce  ? \add_18ns_18s_18_2_1_U4.top_add_18ns_18s_18_2_1_Adder_1_U.a [17:9] : \add_18ns_18s_18_2_1_U4.top_add_18ns_18s_18_2_1_Adder_1_U.ain_s1 ;
assign _065_ = \add_18ns_18s_18_2_1_U4.top_add_18ns_18s_18_2_1_Adder_1_U.ce  ? \add_18ns_18s_18_2_1_U4.top_add_18ns_18s_18_2_1_Adder_1_U.facout_s1  : \add_18ns_18s_18_2_1_U4.top_add_18ns_18s_18_2_1_Adder_1_U.carry_s1 ;
assign _066_ = \add_18ns_18s_18_2_1_U4.top_add_18ns_18s_18_2_1_Adder_1_U.ce  ? \add_18ns_18s_18_2_1_U4.top_add_18ns_18s_18_2_1_Adder_1_U.fas_s1  : \add_18ns_18s_18_2_1_U4.top_add_18ns_18s_18_2_1_Adder_1_U.sum_s1 ;
assign _067_ = \add_18ns_18s_18_2_1_U4.top_add_18ns_18s_18_2_1_Adder_1_U.u1.a  + \add_18ns_18s_18_2_1_U4.top_add_18ns_18s_18_2_1_Adder_1_U.u1.b ;
assign { \add_18ns_18s_18_2_1_U4.top_add_18ns_18s_18_2_1_Adder_1_U.u1.cout , \add_18ns_18s_18_2_1_U4.top_add_18ns_18s_18_2_1_Adder_1_U.u1.s  } = _067_ + \add_18ns_18s_18_2_1_U4.top_add_18ns_18s_18_2_1_Adder_1_U.u1.cin ;
assign _068_ = \add_18ns_18s_18_2_1_U4.top_add_18ns_18s_18_2_1_Adder_1_U.u2.a  + \add_18ns_18s_18_2_1_U4.top_add_18ns_18s_18_2_1_Adder_1_U.u2.b ;
assign { \add_18ns_18s_18_2_1_U4.top_add_18ns_18s_18_2_1_Adder_1_U.u2.cout , \add_18ns_18s_18_2_1_U4.top_add_18ns_18s_18_2_1_Adder_1_U.u2.s  } = _068_ + \add_18ns_18s_18_2_1_U4.top_add_18ns_18s_18_2_1_Adder_1_U.u2.cin ;
always @(posedge \add_22s_22s_22_2_1_U7.top_add_22s_22s_22_2_1_Adder_4_U.clk )
\add_22s_22s_22_2_1_U7.top_add_22s_22s_22_2_1_Adder_4_U.bin_s1  <= _070_;
always @(posedge \add_22s_22s_22_2_1_U7.top_add_22s_22s_22_2_1_Adder_4_U.clk )
\add_22s_22s_22_2_1_U7.top_add_22s_22s_22_2_1_Adder_4_U.ain_s1  <= _069_;
always @(posedge \add_22s_22s_22_2_1_U7.top_add_22s_22s_22_2_1_Adder_4_U.clk )
\add_22s_22s_22_2_1_U7.top_add_22s_22s_22_2_1_Adder_4_U.sum_s1  <= _072_;
always @(posedge \add_22s_22s_22_2_1_U7.top_add_22s_22s_22_2_1_Adder_4_U.clk )
\add_22s_22s_22_2_1_U7.top_add_22s_22s_22_2_1_Adder_4_U.carry_s1  <= _071_;
assign _070_ = \add_22s_22s_22_2_1_U7.top_add_22s_22s_22_2_1_Adder_4_U.ce  ? \add_22s_22s_22_2_1_U7.top_add_22s_22s_22_2_1_Adder_4_U.b [21:11] : \add_22s_22s_22_2_1_U7.top_add_22s_22s_22_2_1_Adder_4_U.bin_s1 ;
assign _069_ = \add_22s_22s_22_2_1_U7.top_add_22s_22s_22_2_1_Adder_4_U.ce  ? \add_22s_22s_22_2_1_U7.top_add_22s_22s_22_2_1_Adder_4_U.a [21:11] : \add_22s_22s_22_2_1_U7.top_add_22s_22s_22_2_1_Adder_4_U.ain_s1 ;
assign _071_ = \add_22s_22s_22_2_1_U7.top_add_22s_22s_22_2_1_Adder_4_U.ce  ? \add_22s_22s_22_2_1_U7.top_add_22s_22s_22_2_1_Adder_4_U.facout_s1  : \add_22s_22s_22_2_1_U7.top_add_22s_22s_22_2_1_Adder_4_U.carry_s1 ;
assign _072_ = \add_22s_22s_22_2_1_U7.top_add_22s_22s_22_2_1_Adder_4_U.ce  ? \add_22s_22s_22_2_1_U7.top_add_22s_22s_22_2_1_Adder_4_U.fas_s1  : \add_22s_22s_22_2_1_U7.top_add_22s_22s_22_2_1_Adder_4_U.sum_s1 ;
assign _073_ = \add_22s_22s_22_2_1_U7.top_add_22s_22s_22_2_1_Adder_4_U.u1.a  + \add_22s_22s_22_2_1_U7.top_add_22s_22s_22_2_1_Adder_4_U.u1.b ;
assign { \add_22s_22s_22_2_1_U7.top_add_22s_22s_22_2_1_Adder_4_U.u1.cout , \add_22s_22s_22_2_1_U7.top_add_22s_22s_22_2_1_Adder_4_U.u1.s  } = _073_ + \add_22s_22s_22_2_1_U7.top_add_22s_22s_22_2_1_Adder_4_U.u1.cin ;
assign _074_ = \add_22s_22s_22_2_1_U7.top_add_22s_22s_22_2_1_Adder_4_U.u2.a  + \add_22s_22s_22_2_1_U7.top_add_22s_22s_22_2_1_Adder_4_U.u2.b ;
assign { \add_22s_22s_22_2_1_U7.top_add_22s_22s_22_2_1_Adder_4_U.u2.cout , \add_22s_22s_22_2_1_U7.top_add_22s_22s_22_2_1_Adder_4_U.u2.s  } = _074_ + \add_22s_22s_22_2_1_U7.top_add_22s_22s_22_2_1_Adder_4_U.u2.cin ;
always @(posedge \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_11_U.clk )
\add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_11_U.bin_s1  <= _076_;
always @(posedge \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_11_U.clk )
\add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_11_U.ain_s1  <= _075_;
always @(posedge \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_11_U.clk )
\add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_11_U.sum_s1  <= _078_;
always @(posedge \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_11_U.clk )
\add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_11_U.carry_s1  <= _077_;
assign _076_ = \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_11_U.ce  ? \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_11_U.b [1] : \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_11_U.bin_s1 ;
assign _075_ = \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_11_U.ce  ? \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_11_U.a [1] : \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_11_U.ain_s1 ;
assign _077_ = \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_11_U.ce  ? \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_11_U.facout_s1  : \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_11_U.carry_s1 ;
assign _078_ = \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_11_U.ce  ? \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_11_U.fas_s1  : \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_11_U.sum_s1 ;
assign _079_ = \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_11_U.u1.a  + \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_11_U.u1.b ;
assign { \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_11_U.u1.cout , \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_11_U.u1.s  } = _079_ + \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_11_U.u1.cin ;
assign _080_ = \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_11_U.u2.a  + \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_11_U.u2.b ;
assign { \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_11_U.u2.cout , \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_11_U.u2.s  } = _080_ + \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_11_U.u2.cin ;
always @(posedge \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_11_U.clk )
\add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_11_U.bin_s1  <= _082_;
always @(posedge \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_11_U.clk )
\add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_11_U.ain_s1  <= _081_;
always @(posedge \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_11_U.clk )
\add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_11_U.sum_s1  <= _084_;
always @(posedge \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_11_U.clk )
\add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_11_U.carry_s1  <= _083_;
assign _082_ = \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_11_U.ce  ? \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_11_U.b [1] : \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_11_U.bin_s1 ;
assign _081_ = \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_11_U.ce  ? \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_11_U.a [1] : \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_11_U.ain_s1 ;
assign _083_ = \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_11_U.ce  ? \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_11_U.facout_s1  : \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_11_U.carry_s1 ;
assign _084_ = \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_11_U.ce  ? \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_11_U.fas_s1  : \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_11_U.sum_s1 ;
assign _085_ = \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_11_U.u1.a  + \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_11_U.u1.b ;
assign { \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_11_U.u1.cout , \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_11_U.u1.s  } = _085_ + \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_11_U.u1.cin ;
assign _086_ = \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_11_U.u2.a  + \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_11_U.u2.b ;
assign { \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_11_U.u2.cout , \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_11_U.u2.s  } = _086_ + \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_11_U.u2.cin ;
always @(posedge \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.clk )
\add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s1  <= _088_;
always @(posedge \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.clk )
\add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s1  <= _087_;
always @(posedge \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.clk )
\add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.sum_s1  <= _090_;
always @(posedge \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.clk )
\add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.carry_s1  <= _089_;
assign _088_ = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.ce  ? \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.b [31:16] : \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s1 ;
assign _087_ = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.ce  ? \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.a [31:16] : \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s1 ;
assign _089_ = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.ce  ? \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.facout_s1  : \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.carry_s1 ;
assign _090_ = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.ce  ? \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s1  : \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.sum_s1 ;
assign _091_ = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.a  + \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.b ;
assign { \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cout , \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.s  } = _091_ + \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cin ;
assign _092_ = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.a  + \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.b ;
assign { \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cout , \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.s  } = _092_ + \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cin ;
always @(posedge \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.clk )
\add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s1  <= _094_;
always @(posedge \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.clk )
\add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s1  <= _093_;
always @(posedge \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.clk )
\add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.sum_s1  <= _096_;
always @(posedge \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.clk )
\add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.carry_s1  <= _095_;
assign _094_ = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.ce  ? \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.b [31:16] : \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s1 ;
assign _093_ = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.ce  ? \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.a [31:16] : \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s1 ;
assign _095_ = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.ce  ? \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.facout_s1  : \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.carry_s1 ;
assign _096_ = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.ce  ? \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s1  : \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.sum_s1 ;
assign _097_ = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.a  + \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.b ;
assign { \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cout , \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.s  } = _097_ + \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cin ;
assign _098_ = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.a  + \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.b ;
assign { \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cout , \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.s  } = _098_ + \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cin ;
always @(posedge \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.clk )
\add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s1  <= _100_;
always @(posedge \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.clk )
\add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s1  <= _099_;
always @(posedge \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.clk )
\add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.sum_s1  <= _102_;
always @(posedge \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.clk )
\add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.carry_s1  <= _101_;
assign _100_ = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.ce  ? \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.b [31:16] : \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s1 ;
assign _099_ = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.ce  ? \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.a [31:16] : \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s1 ;
assign _101_ = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.ce  ? \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.facout_s1  : \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.carry_s1 ;
assign _102_ = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.ce  ? \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s1  : \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.sum_s1 ;
assign _103_ = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.a  + \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.b ;
assign { \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cout , \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.s  } = _103_ + \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cin ;
assign _104_ = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.a  + \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.b ;
assign { \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cout , \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.s  } = _104_ + \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cin ;
always @(posedge \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.clk )
\add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s1  <= _106_;
always @(posedge \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.clk )
\add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s1  <= _105_;
always @(posedge \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.clk )
\add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.sum_s1  <= _108_;
always @(posedge \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.clk )
\add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.carry_s1  <= _107_;
assign _106_ = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.ce  ? \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.b [31:16] : \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s1 ;
assign _105_ = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.ce  ? \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.a [31:16] : \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s1 ;
assign _107_ = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.ce  ? \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.facout_s1  : \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.carry_s1 ;
assign _108_ = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.ce  ? \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s1  : \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.sum_s1 ;
assign _109_ = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.a  + \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.b ;
assign { \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cout , \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.s  } = _109_ + \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cin ;
assign _110_ = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.a  + \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.b ;
assign { \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cout , \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.s  } = _110_ + \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cin ;
always @(posedge \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.clk )
\add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s1  <= _112_;
always @(posedge \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.clk )
\add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s1  <= _111_;
always @(posedge \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.clk )
\add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.sum_s1  <= _114_;
always @(posedge \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.clk )
\add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.carry_s1  <= _113_;
assign _112_ = \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.ce  ? \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.b [31:16] : \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s1 ;
assign _111_ = \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.ce  ? \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.a [31:16] : \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s1 ;
assign _113_ = \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.ce  ? \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.facout_s1  : \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.carry_s1 ;
assign _114_ = \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.ce  ? \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s1  : \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.sum_s1 ;
assign _115_ = \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.a  + \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.b ;
assign { \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cout , \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.s  } = _115_ + \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cin ;
assign _116_ = \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.a  + \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.b ;
assign { \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cout , \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.s  } = _116_ + \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cin ;
always @(posedge \add_32ns_32s_32_2_1_U13.top_add_32ns_32s_32_2_1_Adder_9_U.clk )
\add_32ns_32s_32_2_1_U13.top_add_32ns_32s_32_2_1_Adder_9_U.bin_s1  <= _118_;
always @(posedge \add_32ns_32s_32_2_1_U13.top_add_32ns_32s_32_2_1_Adder_9_U.clk )
\add_32ns_32s_32_2_1_U13.top_add_32ns_32s_32_2_1_Adder_9_U.ain_s1  <= _117_;
always @(posedge \add_32ns_32s_32_2_1_U13.top_add_32ns_32s_32_2_1_Adder_9_U.clk )
\add_32ns_32s_32_2_1_U13.top_add_32ns_32s_32_2_1_Adder_9_U.sum_s1  <= _120_;
always @(posedge \add_32ns_32s_32_2_1_U13.top_add_32ns_32s_32_2_1_Adder_9_U.clk )
\add_32ns_32s_32_2_1_U13.top_add_32ns_32s_32_2_1_Adder_9_U.carry_s1  <= _119_;
assign _118_ = \add_32ns_32s_32_2_1_U13.top_add_32ns_32s_32_2_1_Adder_9_U.ce  ? \add_32ns_32s_32_2_1_U13.top_add_32ns_32s_32_2_1_Adder_9_U.b [31:16] : \add_32ns_32s_32_2_1_U13.top_add_32ns_32s_32_2_1_Adder_9_U.bin_s1 ;
assign _117_ = \add_32ns_32s_32_2_1_U13.top_add_32ns_32s_32_2_1_Adder_9_U.ce  ? \add_32ns_32s_32_2_1_U13.top_add_32ns_32s_32_2_1_Adder_9_U.a [31:16] : \add_32ns_32s_32_2_1_U13.top_add_32ns_32s_32_2_1_Adder_9_U.ain_s1 ;
assign _119_ = \add_32ns_32s_32_2_1_U13.top_add_32ns_32s_32_2_1_Adder_9_U.ce  ? \add_32ns_32s_32_2_1_U13.top_add_32ns_32s_32_2_1_Adder_9_U.facout_s1  : \add_32ns_32s_32_2_1_U13.top_add_32ns_32s_32_2_1_Adder_9_U.carry_s1 ;
assign _120_ = \add_32ns_32s_32_2_1_U13.top_add_32ns_32s_32_2_1_Adder_9_U.ce  ? \add_32ns_32s_32_2_1_U13.top_add_32ns_32s_32_2_1_Adder_9_U.fas_s1  : \add_32ns_32s_32_2_1_U13.top_add_32ns_32s_32_2_1_Adder_9_U.sum_s1 ;
assign _121_ = \add_32ns_32s_32_2_1_U13.top_add_32ns_32s_32_2_1_Adder_9_U.u1.a  + \add_32ns_32s_32_2_1_U13.top_add_32ns_32s_32_2_1_Adder_9_U.u1.b ;
assign { \add_32ns_32s_32_2_1_U13.top_add_32ns_32s_32_2_1_Adder_9_U.u1.cout , \add_32ns_32s_32_2_1_U13.top_add_32ns_32s_32_2_1_Adder_9_U.u1.s  } = _121_ + \add_32ns_32s_32_2_1_U13.top_add_32ns_32s_32_2_1_Adder_9_U.u1.cin ;
assign _122_ = \add_32ns_32s_32_2_1_U13.top_add_32ns_32s_32_2_1_Adder_9_U.u2.a  + \add_32ns_32s_32_2_1_U13.top_add_32ns_32s_32_2_1_Adder_9_U.u2.b ;
assign { \add_32ns_32s_32_2_1_U13.top_add_32ns_32s_32_2_1_Adder_9_U.u2.cout , \add_32ns_32s_32_2_1_U13.top_add_32ns_32s_32_2_1_Adder_9_U.u2.s  } = _122_ + \add_32ns_32s_32_2_1_U13.top_add_32ns_32s_32_2_1_Adder_9_U.u2.cin ;
always @(posedge \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_5_U.clk )
\add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_5_U.bin_s1  <= _124_;
always @(posedge \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_5_U.clk )
\add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_5_U.ain_s1  <= _123_;
always @(posedge \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_5_U.clk )
\add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_5_U.sum_s1  <= _126_;
always @(posedge \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_5_U.clk )
\add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_5_U.carry_s1  <= _125_;
assign _124_ = \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_5_U.ce  ? \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_5_U.b [31:16] : \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_5_U.bin_s1 ;
assign _123_ = \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_5_U.ce  ? \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_5_U.a [31:16] : \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_5_U.ain_s1 ;
assign _125_ = \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_5_U.ce  ? \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_5_U.facout_s1  : \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_5_U.carry_s1 ;
assign _126_ = \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_5_U.ce  ? \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_5_U.fas_s1  : \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_5_U.sum_s1 ;
assign _127_ = \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_5_U.u1.a  + \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_5_U.u1.b ;
assign { \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_5_U.u1.cout , \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_5_U.u1.s  } = _127_ + \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_5_U.u1.cin ;
assign _128_ = \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_5_U.u2.a  + \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_5_U.u2.b ;
assign { \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_5_U.u2.cout , \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_5_U.u2.s  } = _128_ + \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_5_U.u2.cin ;
always @(posedge \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.clk )
\add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.bin_s1  <= _130_;
always @(posedge \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.clk )
\add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.ain_s1  <= _129_;
always @(posedge \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.clk )
\add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.sum_s1  <= _132_;
always @(posedge \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.clk )
\add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.carry_s1  <= _131_;
assign _130_ = \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.ce  ? \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.b [31:16] : \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.bin_s1 ;
assign _129_ = \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.ce  ? \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.a [31:16] : \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.ain_s1 ;
assign _131_ = \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.ce  ? \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.facout_s1  : \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.carry_s1 ;
assign _132_ = \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.ce  ? \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.fas_s1  : \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.sum_s1 ;
assign _133_ = \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.u1.a  + \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.u1.b ;
assign { \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.u1.cout , \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.u1.s  } = _133_ + \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.u1.cin ;
assign _134_ = \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.u2.a  + \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.u2.b ;
assign { \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.u2.cout , \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.u2.s  } = _134_ + \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.u2.cin ;
always @(posedge \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_10_U.clk )
\add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_10_U.bin_s1  <= _136_;
always @(posedge \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_10_U.clk )
\add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_10_U.ain_s1  <= _135_;
always @(posedge \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_10_U.clk )
\add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_10_U.sum_s1  <= _138_;
always @(posedge \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_10_U.clk )
\add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_10_U.carry_s1  <= _137_;
assign _136_ = \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_10_U.ce  ? \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_10_U.b [34:17] : \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_10_U.bin_s1 ;
assign _135_ = \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_10_U.ce  ? \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_10_U.a [34:17] : \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_10_U.ain_s1 ;
assign _137_ = \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_10_U.ce  ? \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_10_U.facout_s1  : \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_10_U.carry_s1 ;
assign _138_ = \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_10_U.ce  ? \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_10_U.fas_s1  : \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_10_U.sum_s1 ;
assign _139_ = \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_10_U.u1.a  + \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_10_U.u1.b ;
assign { \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_10_U.u1.cout , \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_10_U.u1.s  } = _139_ + \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_10_U.u1.cin ;
assign _140_ = \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_10_U.u2.a  + \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_10_U.u2.b ;
assign { \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_10_U.u2.cout , \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_10_U.u2.s  } = _140_ + \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_10_U.u2.cin ;
always @(posedge \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_6_U.clk )
\add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_6_U.bin_s1  <= _142_;
always @(posedge \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_6_U.clk )
\add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_6_U.ain_s1  <= _141_;
always @(posedge \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_6_U.clk )
\add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_6_U.sum_s1  <= _144_;
always @(posedge \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_6_U.clk )
\add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_6_U.carry_s1  <= _143_;
assign _142_ = \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_6_U.ce  ? \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_6_U.b [35:18] : \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_6_U.bin_s1 ;
assign _141_ = \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_6_U.ce  ? \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_6_U.a [35:18] : \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_6_U.ain_s1 ;
assign _143_ = \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_6_U.ce  ? \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_6_U.facout_s1  : \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_6_U.carry_s1 ;
assign _144_ = \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_6_U.ce  ? \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_6_U.fas_s1  : \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_6_U.sum_s1 ;
assign _145_ = \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_6_U.u1.a  + \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_6_U.u1.b ;
assign { \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_6_U.u1.cout , \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_6_U.u1.s  } = _145_ + \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_6_U.u1.cin ;
assign _146_ = \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_6_U.u2.a  + \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_6_U.u2.b ;
assign { \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_6_U.u2.cout , \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_6_U.u2.s  } = _146_ + \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_6_U.u2.cin ;
always @(posedge \add_47s_47s_47_2_1_U11.top_add_47s_47s_47_2_1_Adder_8_U.clk )
\add_47s_47s_47_2_1_U11.top_add_47s_47s_47_2_1_Adder_8_U.bin_s1  <= _148_;
always @(posedge \add_47s_47s_47_2_1_U11.top_add_47s_47s_47_2_1_Adder_8_U.clk )
\add_47s_47s_47_2_1_U11.top_add_47s_47s_47_2_1_Adder_8_U.ain_s1  <= _147_;
always @(posedge \add_47s_47s_47_2_1_U11.top_add_47s_47s_47_2_1_Adder_8_U.clk )
\add_47s_47s_47_2_1_U11.top_add_47s_47s_47_2_1_Adder_8_U.sum_s1  <= _150_;
always @(posedge \add_47s_47s_47_2_1_U11.top_add_47s_47s_47_2_1_Adder_8_U.clk )
\add_47s_47s_47_2_1_U11.top_add_47s_47s_47_2_1_Adder_8_U.carry_s1  <= _149_;
assign _148_ = \add_47s_47s_47_2_1_U11.top_add_47s_47s_47_2_1_Adder_8_U.ce  ? \add_47s_47s_47_2_1_U11.top_add_47s_47s_47_2_1_Adder_8_U.b [46:23] : \add_47s_47s_47_2_1_U11.top_add_47s_47s_47_2_1_Adder_8_U.bin_s1 ;
assign _147_ = \add_47s_47s_47_2_1_U11.top_add_47s_47s_47_2_1_Adder_8_U.ce  ? \add_47s_47s_47_2_1_U11.top_add_47s_47s_47_2_1_Adder_8_U.a [46:23] : \add_47s_47s_47_2_1_U11.top_add_47s_47s_47_2_1_Adder_8_U.ain_s1 ;
assign _149_ = \add_47s_47s_47_2_1_U11.top_add_47s_47s_47_2_1_Adder_8_U.ce  ? \add_47s_47s_47_2_1_U11.top_add_47s_47s_47_2_1_Adder_8_U.facout_s1  : \add_47s_47s_47_2_1_U11.top_add_47s_47s_47_2_1_Adder_8_U.carry_s1 ;
assign _150_ = \add_47s_47s_47_2_1_U11.top_add_47s_47s_47_2_1_Adder_8_U.ce  ? \add_47s_47s_47_2_1_U11.top_add_47s_47s_47_2_1_Adder_8_U.fas_s1  : \add_47s_47s_47_2_1_U11.top_add_47s_47s_47_2_1_Adder_8_U.sum_s1 ;
assign _151_ = \add_47s_47s_47_2_1_U11.top_add_47s_47s_47_2_1_Adder_8_U.u1.a  + \add_47s_47s_47_2_1_U11.top_add_47s_47s_47_2_1_Adder_8_U.u1.b ;
assign { \add_47s_47s_47_2_1_U11.top_add_47s_47s_47_2_1_Adder_8_U.u1.cout , \add_47s_47s_47_2_1_U11.top_add_47s_47s_47_2_1_Adder_8_U.u1.s  } = _151_ + \add_47s_47s_47_2_1_U11.top_add_47s_47s_47_2_1_Adder_8_U.u1.cin ;
assign _152_ = \add_47s_47s_47_2_1_U11.top_add_47s_47s_47_2_1_Adder_8_U.u2.a  + \add_47s_47s_47_2_1_U11.top_add_47s_47s_47_2_1_Adder_8_U.u2.b ;
assign { \add_47s_47s_47_2_1_U11.top_add_47s_47s_47_2_1_Adder_8_U.u2.cout , \add_47s_47s_47_2_1_U11.top_add_47s_47s_47_2_1_Adder_8_U.u2.s  } = _152_ + \add_47s_47s_47_2_1_U11.top_add_47s_47s_47_2_1_Adder_8_U.u2.cin ;
always @(posedge \ashr_4ns_4ns_4_7_1_U2.clk )
\ashr_4ns_4ns_4_7_1_U2.dout_array[5]  <= _164_;
always @(posedge \ashr_4ns_4ns_4_7_1_U2.clk )
\ashr_4ns_4ns_4_7_1_U2.din1_cast_array[5]  <= _158_;
always @(posedge \ashr_4ns_4ns_4_7_1_U2.clk )
\ashr_4ns_4ns_4_7_1_U2.dout_array[4]  <= _163_;
always @(posedge \ashr_4ns_4ns_4_7_1_U2.clk )
\ashr_4ns_4ns_4_7_1_U2.din1_cast_array[4]  <= _157_;
always @(posedge \ashr_4ns_4ns_4_7_1_U2.clk )
\ashr_4ns_4ns_4_7_1_U2.dout_array[3]  <= _162_;
always @(posedge \ashr_4ns_4ns_4_7_1_U2.clk )
\ashr_4ns_4ns_4_7_1_U2.din1_cast_array[3]  <= _156_;
always @(posedge \ashr_4ns_4ns_4_7_1_U2.clk )
\ashr_4ns_4ns_4_7_1_U2.dout_array[2]  <= _161_;
always @(posedge \ashr_4ns_4ns_4_7_1_U2.clk )
\ashr_4ns_4ns_4_7_1_U2.din1_cast_array[2]  <= _155_;
always @(posedge \ashr_4ns_4ns_4_7_1_U2.clk )
\ashr_4ns_4ns_4_7_1_U2.dout_array[1]  <= _160_;
always @(posedge \ashr_4ns_4ns_4_7_1_U2.clk )
\ashr_4ns_4ns_4_7_1_U2.din1_cast_array[1]  <= _154_;
always @(posedge \ashr_4ns_4ns_4_7_1_U2.clk )
\ashr_4ns_4ns_4_7_1_U2.dout_array[0]  <= _159_;
always @(posedge \ashr_4ns_4ns_4_7_1_U2.clk )
\ashr_4ns_4ns_4_7_1_U2.din1_cast_array[0]  <= _153_;
assign _165_ = \ashr_4ns_4ns_4_7_1_U2.ce  ? \ashr_4ns_4ns_4_7_1_U2.din1_cast_array[4]  : \ashr_4ns_4ns_4_7_1_U2.din1_cast_array[5] ;
assign _158_ = \ashr_4ns_4ns_4_7_1_U2.reset  ? 4'h0 : _165_;
assign _166_ = \ashr_4ns_4ns_4_7_1_U2.ce  ? _179_ : \ashr_4ns_4ns_4_7_1_U2.dout_array[5] ;
assign _164_ = \ashr_4ns_4ns_4_7_1_U2.reset  ? 4'h0 : _166_;
assign _167_ = \ashr_4ns_4ns_4_7_1_U2.ce  ? \ashr_4ns_4ns_4_7_1_U2.din1_cast_array[3]  : \ashr_4ns_4ns_4_7_1_U2.din1_cast_array[4] ;
assign _157_ = \ashr_4ns_4ns_4_7_1_U2.reset  ? 4'h0 : _167_;
assign _168_ = \ashr_4ns_4ns_4_7_1_U2.ce  ? _178_ : \ashr_4ns_4ns_4_7_1_U2.dout_array[4] ;
assign _163_ = \ashr_4ns_4ns_4_7_1_U2.reset  ? 4'h0 : _168_;
assign _169_ = \ashr_4ns_4ns_4_7_1_U2.ce  ? \ashr_4ns_4ns_4_7_1_U2.din1_cast_array[2]  : \ashr_4ns_4ns_4_7_1_U2.din1_cast_array[3] ;
assign _156_ = \ashr_4ns_4ns_4_7_1_U2.reset  ? 4'h0 : _169_;
assign _170_ = \ashr_4ns_4ns_4_7_1_U2.ce  ? _177_ : \ashr_4ns_4ns_4_7_1_U2.dout_array[3] ;
assign _162_ = \ashr_4ns_4ns_4_7_1_U2.reset  ? 4'h0 : _170_;
assign _171_ = \ashr_4ns_4ns_4_7_1_U2.ce  ? \ashr_4ns_4ns_4_7_1_U2.din1_cast_array[1]  : \ashr_4ns_4ns_4_7_1_U2.din1_cast_array[2] ;
assign _155_ = \ashr_4ns_4ns_4_7_1_U2.reset  ? 4'h0 : _171_;
assign _172_ = \ashr_4ns_4ns_4_7_1_U2.ce  ? \ashr_4ns_4ns_4_7_1_U2.dout_array[1]  : \ashr_4ns_4ns_4_7_1_U2.dout_array[2] ;
assign _161_ = \ashr_4ns_4ns_4_7_1_U2.reset  ? 4'h0 : _172_;
assign _173_ = \ashr_4ns_4ns_4_7_1_U2.ce  ? \ashr_4ns_4ns_4_7_1_U2.din1_cast_array[0]  : \ashr_4ns_4ns_4_7_1_U2.din1_cast_array[1] ;
assign _154_ = \ashr_4ns_4ns_4_7_1_U2.reset  ? 4'h0 : _173_;
assign _174_ = \ashr_4ns_4ns_4_7_1_U2.ce  ? \ashr_4ns_4ns_4_7_1_U2.dout_array[0]  : \ashr_4ns_4ns_4_7_1_U2.dout_array[1] ;
assign _160_ = \ashr_4ns_4ns_4_7_1_U2.reset  ? 4'h0 : _174_;
assign _175_ = \ashr_4ns_4ns_4_7_1_U2.ce  ? \ashr_4ns_4ns_4_7_1_U2.din1  : \ashr_4ns_4ns_4_7_1_U2.din1_cast_array[0] ;
assign _153_ = \ashr_4ns_4ns_4_7_1_U2.reset  ? 4'h0 : _175_;
assign _176_ = \ashr_4ns_4ns_4_7_1_U2.ce  ? \ashr_4ns_4ns_4_7_1_U2.din0  : \ashr_4ns_4ns_4_7_1_U2.dout_array[0] ;
assign _159_ = \ashr_4ns_4ns_4_7_1_U2.reset  ? 4'h0 : _176_;
assign _177_ = $signed(\ashr_4ns_4ns_4_7_1_U2.dout_array[2] ) >>> { \ashr_4ns_4ns_4_7_1_U2.din1_cast_array[2] [3], 3'h0 };
assign _178_ = $signed(\ashr_4ns_4ns_4_7_1_U2.dout_array[3] ) >>> { \ashr_4ns_4ns_4_7_1_U2.din1_cast_array[3] [2], 2'h0 };
assign _179_ = $signed(\ashr_4ns_4ns_4_7_1_U2.dout_array[4] ) >>> { \ashr_4ns_4ns_4_7_1_U2.din1_cast_array[4] [1], 1'h0 };
assign \ashr_4ns_4ns_4_7_1_U2.dout  = $signed(\ashr_4ns_4ns_4_7_1_U2.dout_array[5] ) >>> \ashr_4ns_4ns_4_7_1_U2.din1_cast_array[5] [0];
always @(posedge \shl_4ns_4ns_4_7_1_U3.clk )
\shl_4ns_4ns_4_7_1_U3.dout_array[5]  <= _191_;
always @(posedge \shl_4ns_4ns_4_7_1_U3.clk )
\shl_4ns_4ns_4_7_1_U3.din1_cast_array[5]  <= _185_;
always @(posedge \shl_4ns_4ns_4_7_1_U3.clk )
\shl_4ns_4ns_4_7_1_U3.dout_array[4]  <= _190_;
always @(posedge \shl_4ns_4ns_4_7_1_U3.clk )
\shl_4ns_4ns_4_7_1_U3.din1_cast_array[4]  <= _184_;
always @(posedge \shl_4ns_4ns_4_7_1_U3.clk )
\shl_4ns_4ns_4_7_1_U3.dout_array[3]  <= _189_;
always @(posedge \shl_4ns_4ns_4_7_1_U3.clk )
\shl_4ns_4ns_4_7_1_U3.din1_cast_array[3]  <= _183_;
always @(posedge \shl_4ns_4ns_4_7_1_U3.clk )
\shl_4ns_4ns_4_7_1_U3.dout_array[2]  <= _188_;
always @(posedge \shl_4ns_4ns_4_7_1_U3.clk )
\shl_4ns_4ns_4_7_1_U3.din1_cast_array[2]  <= _182_;
always @(posedge \shl_4ns_4ns_4_7_1_U3.clk )
\shl_4ns_4ns_4_7_1_U3.dout_array[1]  <= _187_;
always @(posedge \shl_4ns_4ns_4_7_1_U3.clk )
\shl_4ns_4ns_4_7_1_U3.din1_cast_array[1]  <= _181_;
always @(posedge \shl_4ns_4ns_4_7_1_U3.clk )
\shl_4ns_4ns_4_7_1_U3.dout_array[0]  <= _186_;
always @(posedge \shl_4ns_4ns_4_7_1_U3.clk )
\shl_4ns_4ns_4_7_1_U3.din1_cast_array[0]  <= _180_;
assign _192_ = \shl_4ns_4ns_4_7_1_U3.ce  ? \shl_4ns_4ns_4_7_1_U3.din1_cast_array[4]  : \shl_4ns_4ns_4_7_1_U3.din1_cast_array[5] ;
assign _185_ = \shl_4ns_4ns_4_7_1_U3.reset  ? 4'h0 : _192_;
assign _193_ = \shl_4ns_4ns_4_7_1_U3.ce  ? _206_ : \shl_4ns_4ns_4_7_1_U3.dout_array[5] ;
assign _191_ = \shl_4ns_4ns_4_7_1_U3.reset  ? 4'h0 : _193_;
assign _194_ = \shl_4ns_4ns_4_7_1_U3.ce  ? \shl_4ns_4ns_4_7_1_U3.din1_cast_array[3]  : \shl_4ns_4ns_4_7_1_U3.din1_cast_array[4] ;
assign _184_ = \shl_4ns_4ns_4_7_1_U3.reset  ? 4'h0 : _194_;
assign _195_ = \shl_4ns_4ns_4_7_1_U3.ce  ? _205_ : \shl_4ns_4ns_4_7_1_U3.dout_array[4] ;
assign _190_ = \shl_4ns_4ns_4_7_1_U3.reset  ? 4'h0 : _195_;
assign _196_ = \shl_4ns_4ns_4_7_1_U3.ce  ? \shl_4ns_4ns_4_7_1_U3.din1_cast_array[2]  : \shl_4ns_4ns_4_7_1_U3.din1_cast_array[3] ;
assign _183_ = \shl_4ns_4ns_4_7_1_U3.reset  ? 4'h0 : _196_;
assign _197_ = \shl_4ns_4ns_4_7_1_U3.ce  ? _204_ : \shl_4ns_4ns_4_7_1_U3.dout_array[3] ;
assign _189_ = \shl_4ns_4ns_4_7_1_U3.reset  ? 4'h0 : _197_;
assign _198_ = \shl_4ns_4ns_4_7_1_U3.ce  ? \shl_4ns_4ns_4_7_1_U3.din1_cast_array[1]  : \shl_4ns_4ns_4_7_1_U3.din1_cast_array[2] ;
assign _182_ = \shl_4ns_4ns_4_7_1_U3.reset  ? 4'h0 : _198_;
assign _199_ = \shl_4ns_4ns_4_7_1_U3.ce  ? \shl_4ns_4ns_4_7_1_U3.dout_array[1]  : \shl_4ns_4ns_4_7_1_U3.dout_array[2] ;
assign _188_ = \shl_4ns_4ns_4_7_1_U3.reset  ? 4'h0 : _199_;
assign _200_ = \shl_4ns_4ns_4_7_1_U3.ce  ? \shl_4ns_4ns_4_7_1_U3.din1_cast_array[0]  : \shl_4ns_4ns_4_7_1_U3.din1_cast_array[1] ;
assign _181_ = \shl_4ns_4ns_4_7_1_U3.reset  ? 4'h0 : _200_;
assign _201_ = \shl_4ns_4ns_4_7_1_U3.ce  ? \shl_4ns_4ns_4_7_1_U3.dout_array[0]  : \shl_4ns_4ns_4_7_1_U3.dout_array[1] ;
assign _187_ = \shl_4ns_4ns_4_7_1_U3.reset  ? 4'h0 : _201_;
assign _202_ = \shl_4ns_4ns_4_7_1_U3.ce  ? \shl_4ns_4ns_4_7_1_U3.din1  : \shl_4ns_4ns_4_7_1_U3.din1_cast_array[0] ;
assign _180_ = \shl_4ns_4ns_4_7_1_U3.reset  ? 4'h0 : _202_;
assign _203_ = \shl_4ns_4ns_4_7_1_U3.ce  ? \shl_4ns_4ns_4_7_1_U3.din0  : \shl_4ns_4ns_4_7_1_U3.dout_array[0] ;
assign _186_ = \shl_4ns_4ns_4_7_1_U3.reset  ? 4'h0 : _203_;
assign _204_ = \shl_4ns_4ns_4_7_1_U3.dout_array[2]  << { \shl_4ns_4ns_4_7_1_U3.din1_cast_array[2] [3], 3'h0 };
assign _205_ = \shl_4ns_4ns_4_7_1_U3.dout_array[3]  << { \shl_4ns_4ns_4_7_1_U3.din1_cast_array[3] [2], 2'h0 };
assign _206_ = \shl_4ns_4ns_4_7_1_U3.dout_array[4]  << { \shl_4ns_4ns_4_7_1_U3.din1_cast_array[4] [1], 1'h0 };
assign \shl_4ns_4ns_4_7_1_U3.dout  = \shl_4ns_4ns_4_7_1_U3.dout_array[5]  << \shl_4ns_4ns_4_7_1_U3.din1_cast_array[5] [0];
assign \sub_36s_36ns_36_2_1_U6.top_sub_36s_36ns_36_2_1_Adder_3_U.bin_s0  = ~ \sub_36s_36ns_36_2_1_U6.top_sub_36s_36ns_36_2_1_Adder_3_U.b ;
always @(posedge \sub_36s_36ns_36_2_1_U6.top_sub_36s_36ns_36_2_1_Adder_3_U.clk )
\sub_36s_36ns_36_2_1_U6.top_sub_36s_36ns_36_2_1_Adder_3_U.bin_s1  <= _208_;
always @(posedge \sub_36s_36ns_36_2_1_U6.top_sub_36s_36ns_36_2_1_Adder_3_U.clk )
\sub_36s_36ns_36_2_1_U6.top_sub_36s_36ns_36_2_1_Adder_3_U.ain_s1  <= _207_;
always @(posedge \sub_36s_36ns_36_2_1_U6.top_sub_36s_36ns_36_2_1_Adder_3_U.clk )
\sub_36s_36ns_36_2_1_U6.top_sub_36s_36ns_36_2_1_Adder_3_U.sum_s1  <= _210_;
always @(posedge \sub_36s_36ns_36_2_1_U6.top_sub_36s_36ns_36_2_1_Adder_3_U.clk )
\sub_36s_36ns_36_2_1_U6.top_sub_36s_36ns_36_2_1_Adder_3_U.carry_s1  <= _209_;
assign _208_ = \sub_36s_36ns_36_2_1_U6.top_sub_36s_36ns_36_2_1_Adder_3_U.ce  ? \sub_36s_36ns_36_2_1_U6.top_sub_36s_36ns_36_2_1_Adder_3_U.bin_s0 [35:18] : \sub_36s_36ns_36_2_1_U6.top_sub_36s_36ns_36_2_1_Adder_3_U.bin_s1 ;
assign _207_ = \sub_36s_36ns_36_2_1_U6.top_sub_36s_36ns_36_2_1_Adder_3_U.ce  ? \sub_36s_36ns_36_2_1_U6.top_sub_36s_36ns_36_2_1_Adder_3_U.a [35:18] : \sub_36s_36ns_36_2_1_U6.top_sub_36s_36ns_36_2_1_Adder_3_U.ain_s1 ;
assign _209_ = \sub_36s_36ns_36_2_1_U6.top_sub_36s_36ns_36_2_1_Adder_3_U.ce  ? \sub_36s_36ns_36_2_1_U6.top_sub_36s_36ns_36_2_1_Adder_3_U.facout_s1  : \sub_36s_36ns_36_2_1_U6.top_sub_36s_36ns_36_2_1_Adder_3_U.carry_s1 ;
assign _210_ = \sub_36s_36ns_36_2_1_U6.top_sub_36s_36ns_36_2_1_Adder_3_U.ce  ? \sub_36s_36ns_36_2_1_U6.top_sub_36s_36ns_36_2_1_Adder_3_U.fas_s1  : \sub_36s_36ns_36_2_1_U6.top_sub_36s_36ns_36_2_1_Adder_3_U.sum_s1 ;
assign _211_ = \sub_36s_36ns_36_2_1_U6.top_sub_36s_36ns_36_2_1_Adder_3_U.u1.a  + \sub_36s_36ns_36_2_1_U6.top_sub_36s_36ns_36_2_1_Adder_3_U.u1.b ;
assign { \sub_36s_36ns_36_2_1_U6.top_sub_36s_36ns_36_2_1_Adder_3_U.u1.cout , \sub_36s_36ns_36_2_1_U6.top_sub_36s_36ns_36_2_1_Adder_3_U.u1.s  } = _211_ + \sub_36s_36ns_36_2_1_U6.top_sub_36s_36ns_36_2_1_Adder_3_U.u1.cin ;
assign _212_ = \sub_36s_36ns_36_2_1_U6.top_sub_36s_36ns_36_2_1_Adder_3_U.u2.a  + \sub_36s_36ns_36_2_1_U6.top_sub_36s_36ns_36_2_1_Adder_3_U.u2.b ;
assign { \sub_36s_36ns_36_2_1_U6.top_sub_36s_36ns_36_2_1_Adder_3_U.u2.cout , \sub_36s_36ns_36_2_1_U6.top_sub_36s_36ns_36_2_1_Adder_3_U.u2.s  } = _212_ + \sub_36s_36ns_36_2_1_U6.top_sub_36s_36ns_36_2_1_Adder_3_U.u2.cin ;
assign \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.bin_s0  = ~ \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.b ;
always @(posedge \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.clk )
\sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.bin_s1  <= _214_;
always @(posedge \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.clk )
\sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.ain_s1  <= _213_;
always @(posedge \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.clk )
\sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.sum_s1  <= _216_;
always @(posedge \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.clk )
\sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.carry_s1  <= _215_;
assign _214_ = \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.ce  ? \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.bin_s0 [3:2] : \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.bin_s1 ;
assign _213_ = \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.ce  ? \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.a [3:2] : \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.ain_s1 ;
assign _215_ = \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.ce  ? \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.facout_s1  : \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.carry_s1 ;
assign _216_ = \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.ce  ? \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.fas_s1  : \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.sum_s1 ;
assign _217_ = \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.u1.a  + \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.u1.b ;
assign { \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.u1.cout , \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.u1.s  } = _217_ + \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.u1.cin ;
assign _218_ = \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.u2.a  + \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.u2.b ;
assign { \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.u2.cout , \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.u2.s  } = _218_ + \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.u2.cin ;
assign _219_ = | tmp_2_reg_827;
assign _220_ = tmp_2_reg_827 != 32'd4294967295;
assign _221_ = | trunc_ln851_1_reg_881;
assign _222_ = | op_12[13:0];
assign _223_ = | op_15[1:0];
assign _224_ = | op_10[2:0];
assign or_ln384_fu_426_p2 = underflow_fu_414_p2 | overflow_reg_860;
assign or_ln785_fu_386_p2 = p_Result_6_reg_821 | icmp_ln768_reg_843;
assign or_ln786_fu_409_p2 = xor_ln786_fu_404_p2 | icmp_ln786_reg_848;
always @(posedge ap_clk)
shl_ln781_reg_749 <= _042_;
always @(posedge ap_clk)
sh_reg_739 <= _041_;
always @(posedge ap_clk)
select_ln69_reg_1007 <= _039_;
always @(posedge ap_clk)
select_ln353_1_reg_918 <= _036_;
always @(posedge ap_clk)
ret_V_reg_770 <= _034_;
always @(posedge ap_clk)
select_ln1192_reg_775 <= _035_;
always @(posedge ap_clk)
ret_V_7_reg_965 <= _031_;
always @(posedge ap_clk)
ret_V_6_reg_955 <= _030_;
always @(posedge ap_clk)
ret_V_5_reg_938 <= _028_;
always @(posedge ap_clk)
ret_V_6_cast_reg_943 <= _029_;
always @(posedge ap_clk)
ret_V_4_reg_901 <= _027_;
always @(posedge ap_clk)
ret_V_3_cast_reg_906 <= _025_;
always @(posedge ap_clk)
ret_V_2_reg_780 <= _024_;
always @(posedge ap_clk)
ret_V_8_reg_995 <= _032_;
always @(posedge ap_clk)
ret_V_16_cast_reg_1000 <= _022_;
always @(posedge ap_clk)
r_reg_754 <= _021_;
always @(posedge ap_clk)
ret_V_1_reg_810 <= _023_;
always @(posedge ap_clk)
p_Result_5_reg_815 <= _019_;
always @(posedge ap_clk)
p_Result_6_reg_821 <= _020_;
always @(posedge ap_clk)
tmp_2_reg_827 <= _043_;
always @(posedge ap_clk)
ret_V_3_reg_833 <= _026_;
always @(posedge ap_clk)
tmp_reg_838 <= _044_;
always @(posedge ap_clk)
p_Result_4_reg_734 <= _018_;
always @(posedge ap_clk)
overflow_reg_860 <= _017_;
always @(posedge ap_clk)
op_26_V_reg_975 <= _016_;
always @(posedge ap_clk)
op_11_V_reg_871 <= _015_;
always @(posedge ap_clk)
select_ln353_reg_876 <= _037_;
always @(posedge ap_clk)
trunc_ln851_1_reg_881 <= _045_;
always @(posedge ap_clk)
icmp_ln851_reg_805 <= _014_;
always @(posedge ap_clk)
icmp_ln851_3_reg_990 <= _013_;
always @(posedge ap_clk)
icmp_ln851_2_reg_933 <= _012_;
always @(posedge ap_clk)
icmp_ln851_1_reg_896 <= _011_;
always @(posedge ap_clk)
icmp_ln768_reg_843 <= _009_;
always @(posedge ap_clk)
icmp_ln786_reg_848 <= _010_;
always @(posedge ap_clk)
sext_ln831_reg_853 <= _040_;
always @(posedge ap_clk)
ashr_ln799_reg_744 <= _008_;
always @(posedge ap_clk)
add_ln69_reg_1042 <= _006_;
always @(posedge ap_clk)
add_ln69_2_reg_1047 <= _005_;
always @(posedge ap_clk)
ret_V_9_reg_1022 <= _033_;
always @(posedge ap_clk)
select_ln69_1_reg_1027 <= _038_;
always @(posedge ap_clk)
add_ln69_1_reg_1032 <= _004_;
always @(posedge ap_clk)
add_ln691_reg_866 <= _003_;
always @(posedge ap_clk)
add_ln691_3_reg_1012 <= _002_;
always @(posedge ap_clk)
add_ln691_2_reg_950 <= _001_;
always @(posedge ap_clk)
add_ln691_1_reg_913 <= _000_;
always @(posedge ap_clk)
ap_CS_fsm <= _007_;
assign _046_ = _054_ ? 2'h2 : 2'h1;
assign _225_ = ap_CS_fsm == 1'h1;
function [41:0] _637_;
input [41:0] a;
input [1763:0] b;
input [41:0] s;
case (s)
42'b000000000000000000000000000000000000000001:
_637_ = b[41:0];
42'b000000000000000000000000000000000000000010:
_637_ = b[83:42];
42'b000000000000000000000000000000000000000100:
_637_ = b[125:84];
42'b000000000000000000000000000000000000001000:
_637_ = b[167:126];
42'b000000000000000000000000000000000000010000:
_637_ = b[209:168];
42'b000000000000000000000000000000000000100000:
_637_ = b[251:210];
42'b000000000000000000000000000000000001000000:
_637_ = b[293:252];
42'b000000000000000000000000000000000010000000:
_637_ = b[335:294];
42'b000000000000000000000000000000000100000000:
_637_ = b[377:336];
42'b000000000000000000000000000000001000000000:
_637_ = b[419:378];
42'b000000000000000000000000000000010000000000:
_637_ = b[461:420];
42'b000000000000000000000000000000100000000000:
_637_ = b[503:462];
42'b000000000000000000000000000001000000000000:
_637_ = b[545:504];
42'b000000000000000000000000000010000000000000:
_637_ = b[587:546];
42'b000000000000000000000000000100000000000000:
_637_ = b[629:588];
42'b000000000000000000000000001000000000000000:
_637_ = b[671:630];
42'b000000000000000000000000010000000000000000:
_637_ = b[713:672];
42'b000000000000000000000000100000000000000000:
_637_ = b[755:714];
42'b000000000000000000000001000000000000000000:
_637_ = b[797:756];
42'b000000000000000000000010000000000000000000:
_637_ = b[839:798];
42'b000000000000000000000100000000000000000000:
_637_ = b[881:840];
42'b000000000000000000001000000000000000000000:
_637_ = b[923:882];
42'b000000000000000000010000000000000000000000:
_637_ = b[965:924];
42'b000000000000000000100000000000000000000000:
_637_ = b[1007:966];
42'b000000000000000001000000000000000000000000:
_637_ = b[1049:1008];
42'b000000000000000010000000000000000000000000:
_637_ = b[1091:1050];
42'b000000000000000100000000000000000000000000:
_637_ = b[1133:1092];
42'b000000000000001000000000000000000000000000:
_637_ = b[1175:1134];
42'b000000000000010000000000000000000000000000:
_637_ = b[1217:1176];
42'b000000000000100000000000000000000000000000:
_637_ = b[1259:1218];
42'b000000000001000000000000000000000000000000:
_637_ = b[1301:1260];
42'b000000000010000000000000000000000000000000:
_637_ = b[1343:1302];
42'b000000000100000000000000000000000000000000:
_637_ = b[1385:1344];
42'b000000001000000000000000000000000000000000:
_637_ = b[1427:1386];
42'b000000010000000000000000000000000000000000:
_637_ = b[1469:1428];
42'b000000100000000000000000000000000000000000:
_637_ = b[1511:1470];
42'b000001000000000000000000000000000000000000:
_637_ = b[1553:1512];
42'b000010000000000000000000000000000000000000:
_637_ = b[1595:1554];
42'b000100000000000000000000000000000000000000:
_637_ = b[1637:1596];
42'b001000000000000000000000000000000000000000:
_637_ = b[1679:1638];
42'b010000000000000000000000000000000000000000:
_637_ = b[1721:1680];
42'b100000000000000000000000000000000000000000:
_637_ = b[1763:1722];
42'b000000000000000000000000000000000000000000:
_637_ = a;
default:
_637_ = 42'bx;
endcase
endfunction
assign ap_NS_fsm = _637_(42'hxxxxxxxxxxx, { 40'h0000000000, _046_, 1722'h00000000004000000000200000000010000000000800000000040000000002000000000100000000008000000000400000000020000000001000000000080000000004000000000200000000010000000000800000000040000000002000000000100000000008000000000400000000020000000001000000000080000000004000000000200000000010000000000800000000040000000002000000000100000000008000000000400000000020000000001000000000080000000004000000000200000000010000000000800000000000000000001 }, { _225_, _266_, _265_, _264_, _263_, _262_, _261_, _260_, _259_, _258_, _257_, _256_, _255_, _254_, _253_, _252_, _251_, _250_, _249_, _248_, _247_, _246_, _245_, _244_, _243_, _242_, _241_, _240_, _239_, _238_, _237_, _236_, _235_, _234_, _233_, _232_, _231_, _230_, _229_, _228_, _227_, _226_ });
assign _226_ = ap_CS_fsm == 42'h20000000000;
assign _227_ = ap_CS_fsm == 41'h10000000000;
assign _228_ = ap_CS_fsm == 40'h8000000000;
assign _229_ = ap_CS_fsm == 39'h4000000000;
assign _230_ = ap_CS_fsm == 38'h2000000000;
assign _231_ = ap_CS_fsm == 37'h1000000000;
assign _232_ = ap_CS_fsm == 36'h800000000;
assign _233_ = ap_CS_fsm == 35'h400000000;
assign _234_ = ap_CS_fsm == 34'h200000000;
assign _235_ = ap_CS_fsm == 33'h100000000;
assign _236_ = ap_CS_fsm == 32'd2147483648;
assign _237_ = ap_CS_fsm == 31'h40000000;
assign _238_ = ap_CS_fsm == 30'h20000000;
assign _239_ = ap_CS_fsm == 29'h10000000;
assign _240_ = ap_CS_fsm == 28'h8000000;
assign _241_ = ap_CS_fsm == 27'h4000000;
assign _242_ = ap_CS_fsm == 26'h2000000;
assign _243_ = ap_CS_fsm == 25'h1000000;
assign _244_ = ap_CS_fsm == 24'h800000;
assign _245_ = ap_CS_fsm == 23'h400000;
assign _246_ = ap_CS_fsm == 22'h200000;
assign _247_ = ap_CS_fsm == 21'h100000;
assign _248_ = ap_CS_fsm == 20'h80000;
assign _249_ = ap_CS_fsm == 19'h40000;
assign _250_ = ap_CS_fsm == 18'h20000;
assign _251_ = ap_CS_fsm == 17'h10000;
assign _252_ = ap_CS_fsm == 16'h8000;
assign _253_ = ap_CS_fsm == 15'h4000;
assign _254_ = ap_CS_fsm == 14'h2000;
assign _255_ = ap_CS_fsm == 13'h1000;
assign _256_ = ap_CS_fsm == 12'h800;
assign _257_ = ap_CS_fsm == 11'h400;
assign _258_ = ap_CS_fsm == 10'h200;
assign _259_ = ap_CS_fsm == 9'h100;
assign _260_ = ap_CS_fsm == 8'h80;
assign _261_ = ap_CS_fsm == 7'h40;
assign _262_ = ap_CS_fsm == 6'h20;
assign _263_ = ap_CS_fsm == 5'h10;
assign _264_ = ap_CS_fsm == 4'h8;
assign _265_ = ap_CS_fsm == 3'h4;
assign _266_ = ap_CS_fsm == 2'h2;
assign op_31_ap_vld = ap_CS_fsm[41] ? 1'h1 : 1'h0;
assign ap_idle = _053_ ? 1'h1 : 1'h0;
assign _042_ = _052_ ? grp_fu_237_p2 : shl_ln781_reg_749;
assign _041_ = ap_CS_fsm[1] ? grp_fu_227_p2 : sh_reg_739;
assign _039_ = ap_CS_fsm[35] ? select_ln69_fu_664_p3 : select_ln69_reg_1007;
assign _036_ = ap_CS_fsm[23] ? select_ln353_1_fu_514_p3 : select_ln353_1_reg_918;
assign _035_ = ap_CS_fsm[11] ? select_ln1192_fu_263_p3 : select_ln1192_reg_775;
assign _034_ = ap_CS_fsm[11] ? grp_fu_257_p2 : ret_V_reg_770;
assign _031_ = ap_CS_fsm[30] ? grp_fu_590_p2 : ret_V_7_reg_965;
assign _030_ = ap_CS_fsm[28] ? ret_V_6_fu_579_p3 : ret_V_6_reg_955;
assign _029_ = ap_CS_fsm[25] ? grp_fu_536_p2[45:14] : ret_V_6_cast_reg_943;
assign _028_ = ap_CS_fsm[25] ? grp_fu_536_p2 : ret_V_5_reg_938;
assign _025_ = ap_CS_fsm[20] ? grp_fu_476_p2[34:3] : ret_V_3_cast_reg_906;
assign _027_ = ap_CS_fsm[20] ? grp_fu_476_p2 : ret_V_4_reg_901;
assign _024_ = ap_CS_fsm[13] ? grp_fu_271_p2 : ret_V_2_reg_780;
assign _022_ = ap_CS_fsm[34] ? grp_fu_619_p2[33:2] : ret_V_16_cast_reg_1000;
assign _032_ = ap_CS_fsm[34] ? grp_fu_619_p2 : ret_V_8_reg_995;
assign _021_ = ap_CS_fsm[9] ? r_fu_241_p3 : r_reg_754;
assign _044_ = ap_CS_fsm[15] ? grp_fu_315_p2[21:3] : tmp_reg_838;
assign _026_ = ap_CS_fsm[15] ? grp_fu_315_p2 : ret_V_3_reg_833;
assign _043_ = ap_CS_fsm[15] ? grp_fu_294_p2[35:4] : tmp_2_reg_827;
assign _020_ = ap_CS_fsm[15] ? grp_fu_294_p2[3] : p_Result_6_reg_821;
assign _019_ = ap_CS_fsm[15] ? grp_fu_294_p2[35] : p_Result_5_reg_815;
assign _023_ = ap_CS_fsm[15] ? grp_fu_294_p2 : ret_V_1_reg_810;
assign _018_ = ap_CS_fsm[0] ? op_1[3] : p_Result_4_reg_734;
assign _017_ = ap_CS_fsm[17] ? overflow_fu_395_p2 : overflow_reg_860;
assign _016_ = ap_CS_fsm[32] ? grp_fu_599_p2 : op_26_V_reg_975;
assign _045_ = ap_CS_fsm[18] ? op_11_V_fu_431_p3[2:0] : trunc_ln851_1_reg_881;
assign _037_ = ap_CS_fsm[18] ? select_ln353_fu_451_p3 : select_ln353_reg_876;
assign _015_ = ap_CS_fsm[18] ? op_11_V_fu_431_p3 : op_11_V_reg_871;
assign _014_ = ap_CS_fsm[14] ? icmp_ln851_fu_325_p2 : icmp_ln851_reg_805;
assign _013_ = ap_CS_fsm[33] ? icmp_ln851_3_fu_629_p2 : icmp_ln851_3_reg_990;
assign _012_ = ap_CS_fsm[24] ? icmp_ln851_2_fu_546_p2 : icmp_ln851_2_reg_933;
assign _011_ = ap_CS_fsm[19] ? icmp_ln851_1_fu_482_p2 : icmp_ln851_1_reg_896;
assign _040_ = ap_CS_fsm[16] ? { tmp_reg_838[18], tmp_reg_838[18], tmp_reg_838[18], tmp_reg_838[18], tmp_reg_838[18], tmp_reg_838[18], tmp_reg_838[18], tmp_reg_838[18], tmp_reg_838[18], tmp_reg_838[18], tmp_reg_838[18], tmp_reg_838[18], tmp_reg_838[18], tmp_reg_838 } : sext_ln831_reg_853;
assign _010_ = ap_CS_fsm[16] ? icmp_ln786_fu_372_p2 : icmp_ln786_reg_848;
assign _009_ = ap_CS_fsm[16] ? icmp_ln768_fu_367_p2 : icmp_ln768_reg_843;
assign _008_ = _051_ ? grp_fu_233_p2 : ashr_ln799_reg_744;
assign _005_ = ap_CS_fsm[39] ? grp_fu_713_p2 : add_ln69_2_reg_1047;
assign _006_ = ap_CS_fsm[39] ? grp_fu_708_p2 : add_ln69_reg_1042;
assign _004_ = ap_CS_fsm[37] ? grp_fu_676_p2 : add_ln69_1_reg_1032;
assign _038_ = ap_CS_fsm[37] ? select_ln69_1_fu_700_p3 : select_ln69_1_reg_1027;
assign _033_ = ap_CS_fsm[37] ? ret_V_9_fu_693_p3 : ret_V_9_reg_1022;
assign _003_ = _050_ ? grp_fu_380_p2 : add_ln691_reg_866;
assign _002_ = _049_ ? grp_fu_659_p2 : add_ln691_3_reg_1012;
assign _001_ = _048_ ? grp_fu_562_p2 : add_ln691_2_reg_950;
assign _000_ = _047_ ? grp_fu_497_p2 : add_ln691_1_reg_913;
assign _007_ = ap_rst ? 42'h00000000001 : ap_NS_fsm;
assign icmp_ln768_fu_367_p2 = _219_ ? 1'h1 : 1'h0;
assign icmp_ln786_fu_372_p2 = _220_ ? 1'h1 : 1'h0;
assign icmp_ln851_1_fu_482_p2 = _221_ ? 1'h1 : 1'h0;
assign icmp_ln851_2_fu_546_p2 = _222_ ? 1'h1 : 1'h0;
assign icmp_ln851_3_fu_629_p2 = _223_ ? 1'h1 : 1'h0;
assign icmp_ln851_fu_325_p2 = _224_ ? 1'h1 : 1'h0;
assign op_11_V_fu_431_p3 = or_ln384_fu_426_p2 ? select_ln384_fu_419_p3 : ret_V_1_reg_810[3:0];
assign r_fu_241_p3 = p_Result_4_reg_734 ? ashr_ln799_reg_744 : shl_ln781_reg_749;
assign ret_V_6_fu_579_p3 = ret_V_5_reg_938[46] ? select_ln850_2_fu_574_p3 : ret_V_6_cast_reg_943;
assign ret_V_9_fu_693_p3 = ret_V_8_reg_995[34] ? select_ln850_3_fu_688_p3 : ret_V_16_cast_reg_1000;
assign select_ln1192_fu_263_p3 = op_9 ? 18'h3ffff : 18'h00000;
assign select_ln353_1_fu_514_p3 = ret_V_4_reg_901[35] ? select_ln850_1_fu_509_p3 : ret_V_3_cast_reg_906;
assign select_ln353_fu_451_p3 = ret_V_3_reg_833[21] ? select_ln850_fu_446_p3 : sext_ln831_reg_853;
assign select_ln384_fu_419_p3 = overflow_reg_860 ? 4'h7 : 4'h8;
assign select_ln69_1_fu_700_p3 = op_17 ? 2'h3 : 2'h0;
assign select_ln69_fu_664_p3 = op_16_V_fu_653_p2 ? 2'h3 : 2'h0;
assign select_ln850_1_fu_509_p3 = icmp_ln851_1_reg_896 ? add_ln691_1_reg_913 : ret_V_3_cast_reg_906;
assign select_ln850_2_fu_574_p3 = icmp_ln851_2_reg_933 ? add_ln691_2_reg_950 : ret_V_6_cast_reg_943;
assign select_ln850_3_fu_688_p3 = icmp_ln851_3_reg_990 ? add_ln691_3_reg_1012 : ret_V_16_cast_reg_1000;
assign select_ln850_fu_446_p3 = icmp_ln851_reg_805 ? add_ln691_reg_866 : sext_ln831_reg_853;
assign ap_CS_fsm_state1 = ap_CS_fsm[0];
assign ap_CS_fsm_state10 = ap_CS_fsm[9];
assign ap_CS_fsm_state11 = ap_CS_fsm[10];
assign ap_CS_fsm_state12 = ap_CS_fsm[11];
assign ap_CS_fsm_state13 = ap_CS_fsm[12];
assign ap_CS_fsm_state14 = ap_CS_fsm[13];
assign ap_CS_fsm_state15 = ap_CS_fsm[14];
assign ap_CS_fsm_state16 = ap_CS_fsm[15];
assign ap_CS_fsm_state17 = ap_CS_fsm[16];
assign ap_CS_fsm_state18 = ap_CS_fsm[17];
assign ap_CS_fsm_state19 = ap_CS_fsm[18];
assign ap_CS_fsm_state2 = ap_CS_fsm[1];
assign ap_CS_fsm_state20 = ap_CS_fsm[19];
assign ap_CS_fsm_state21 = ap_CS_fsm[20];
assign ap_CS_fsm_state22 = ap_CS_fsm[21];
assign ap_CS_fsm_state23 = ap_CS_fsm[22];
assign ap_CS_fsm_state24 = ap_CS_fsm[23];
assign ap_CS_fsm_state25 = ap_CS_fsm[24];
assign ap_CS_fsm_state26 = ap_CS_fsm[25];
assign ap_CS_fsm_state27 = ap_CS_fsm[26];
assign ap_CS_fsm_state28 = ap_CS_fsm[27];
assign ap_CS_fsm_state29 = ap_CS_fsm[28];
assign ap_CS_fsm_state3 = ap_CS_fsm[2];
assign ap_CS_fsm_state30 = ap_CS_fsm[29];
assign ap_CS_fsm_state31 = ap_CS_fsm[30];
assign ap_CS_fsm_state32 = ap_CS_fsm[31];
assign ap_CS_fsm_state33 = ap_CS_fsm[32];
assign ap_CS_fsm_state34 = ap_CS_fsm[33];
assign ap_CS_fsm_state35 = ap_CS_fsm[34];
assign ap_CS_fsm_state36 = ap_CS_fsm[35];
assign ap_CS_fsm_state37 = ap_CS_fsm[36];
assign ap_CS_fsm_state38 = ap_CS_fsm[37];
assign ap_CS_fsm_state39 = ap_CS_fsm[38];
assign ap_CS_fsm_state40 = ap_CS_fsm[39];
assign ap_CS_fsm_state41 = ap_CS_fsm[40];
assign ap_CS_fsm_state42 = ap_CS_fsm[41];
assign ap_CS_fsm_state9 = ap_CS_fsm[8];
assign ap_done = op_31_ap_vld;
assign ap_ready = op_31_ap_vld;
assign grp_fu_257_p0 = { 2'h0, r_reg_754[3], r_reg_754[3], r_reg_754[3], r_reg_754[3], r_reg_754[3], r_reg_754[3], r_reg_754[3], r_reg_754[3], r_reg_754[3], r_reg_754[3], r_reg_754[3], r_reg_754[3], r_reg_754 };
assign grp_fu_257_p1 = { op_0[1], op_0[1], op_0[1], op_0[1], op_0[1], op_0[1], op_0[1], op_0[1], op_0[1], op_0[1], op_0[1], op_0[1], op_0[1], op_0[1], op_0[1], op_0[1], op_0 };
assign grp_fu_294_p0 = { op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6 };
assign grp_fu_294_p1 = { 1'h0, r_reg_754[3], r_reg_754[3], r_reg_754[3], r_reg_754[3], r_reg_754[3], r_reg_754[3], r_reg_754[3], r_reg_754[3], r_reg_754[3], r_reg_754[3], r_reg_754[3], r_reg_754[3], r_reg_754[3], r_reg_754[3], r_reg_754[3], r_reg_754[3], r_reg_754[3], r_reg_754[3], r_reg_754[3], r_reg_754[3], r_reg_754[3], r_reg_754[3], r_reg_754[3], r_reg_754[3], r_reg_754[3], r_reg_754[3], r_reg_754[3], r_reg_754[3], r_reg_754, 3'h0 };
assign grp_fu_315_p0 = { ret_V_2_reg_780[17], ret_V_2_reg_780, 3'h0 };
assign grp_fu_315_p1 = { op_10[3], op_10[3], op_10[3], op_10[3], op_10[3], op_10[3], op_10[3], op_10[3], op_10[3], op_10[3], op_10[3], op_10[3], op_10[3], op_10[3], op_10[3], op_10[3], op_10[3], op_10[3], op_10 };
assign grp_fu_380_p0 = { tmp_reg_838[18], tmp_reg_838[18], tmp_reg_838[18], tmp_reg_838[18], tmp_reg_838[18], tmp_reg_838[18], tmp_reg_838[18], tmp_reg_838[18], tmp_reg_838[18], tmp_reg_838[18], tmp_reg_838[18], tmp_reg_838[18], tmp_reg_838[18], tmp_reg_838 };
assign grp_fu_476_p0 = { select_ln353_reg_876[31], select_ln353_reg_876, 3'h0 };
assign grp_fu_476_p1 = { op_11_V_reg_871[3], op_11_V_reg_871[3], op_11_V_reg_871[3], op_11_V_reg_871[3], op_11_V_reg_871[3], op_11_V_reg_871[3], op_11_V_reg_871[3], op_11_V_reg_871[3], op_11_V_reg_871[3], op_11_V_reg_871[3], op_11_V_reg_871[3], op_11_V_reg_871[3], op_11_V_reg_871[3], op_11_V_reg_871[3], op_11_V_reg_871[3], op_11_V_reg_871[3], op_11_V_reg_871[3], op_11_V_reg_871[3], op_11_V_reg_871[3], op_11_V_reg_871[3], op_11_V_reg_871[3], op_11_V_reg_871[3], op_11_V_reg_871[3], op_11_V_reg_871[3], op_11_V_reg_871[3], op_11_V_reg_871[3], op_11_V_reg_871[3], op_11_V_reg_871[3], op_11_V_reg_871[3], op_11_V_reg_871[3], op_11_V_reg_871[3], op_11_V_reg_871[3], op_11_V_reg_871 };
assign grp_fu_536_p0 = { select_ln353_1_reg_918[31], select_ln353_1_reg_918, 14'h0000 };
assign grp_fu_536_p1 = { op_12[31], op_12[31], op_12[31], op_12[31], op_12[31], op_12[31], op_12[31], op_12[31], op_12[31], op_12[31], op_12[31], op_12[31], op_12[31], op_12[31], op_12[31], op_12 };
assign grp_fu_590_p1 = { op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13 };
assign grp_fu_599_p1 = { 30'h00000000, op_14 };
assign grp_fu_619_p0 = { op_26_V_reg_975[31], op_26_V_reg_975, 2'h0 };
assign grp_fu_619_p1 = { op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15 };
assign grp_fu_676_p1 = { 1'h0, op_18 };
assign grp_fu_720_p0 = { add_ln69_2_reg_1047[1], add_ln69_2_reg_1047[1], add_ln69_2_reg_1047[1], add_ln69_2_reg_1047[1], add_ln69_2_reg_1047[1], add_ln69_2_reg_1047[1], add_ln69_2_reg_1047[1], add_ln69_2_reg_1047[1], add_ln69_2_reg_1047[1], add_ln69_2_reg_1047[1], add_ln69_2_reg_1047[1], add_ln69_2_reg_1047[1], add_ln69_2_reg_1047[1], add_ln69_2_reg_1047[1], add_ln69_2_reg_1047[1], add_ln69_2_reg_1047[1], add_ln69_2_reg_1047[1], add_ln69_2_reg_1047[1], add_ln69_2_reg_1047[1], add_ln69_2_reg_1047[1], add_ln69_2_reg_1047[1], add_ln69_2_reg_1047[1], add_ln69_2_reg_1047[1], add_ln69_2_reg_1047[1], add_ln69_2_reg_1047[1], add_ln69_2_reg_1047[1], add_ln69_2_reg_1047[1], add_ln69_2_reg_1047[1], add_ln69_2_reg_1047[1], add_ln69_2_reg_1047[1], add_ln69_2_reg_1047 };
assign op_31 = grp_fu_720_p2;
assign p_Result_1_fu_502_p3 = ret_V_4_reg_901[35];
assign p_Result_2_fu_567_p3 = ret_V_5_reg_938[46];
assign p_Result_3_fu_681_p3 = ret_V_8_reg_995[34];
assign p_Result_s_fu_439_p3 = ret_V_3_reg_833[21];
assign p_Val2_1_fu_401_p1 = ret_V_1_reg_810[3:0];
assign rhs_1_fu_279_p3 = { r_reg_754, 3'h0 };
assign rhs_3_fu_465_p3 = { select_ln353_reg_876, 3'h0 };
assign rhs_4_fu_525_p3 = { select_ln353_1_reg_918, 14'h0000 };
assign rhs_7_fu_608_p3 = { op_26_V_reg_975, 2'h0 };
assign sext_ln1192_fu_300_p0 = op_10;
assign sext_ln1193_1_fu_286_p1 = { r_reg_754[3], r_reg_754[3], r_reg_754[3], r_reg_754[3], r_reg_754[3], r_reg_754[3], r_reg_754[3], r_reg_754[3], r_reg_754[3], r_reg_754[3], r_reg_754[3], r_reg_754[3], r_reg_754[3], r_reg_754[3], r_reg_754[3], r_reg_754[3], r_reg_754[3], r_reg_754[3], r_reg_754[3], r_reg_754[3], r_reg_754[3], r_reg_754[3], r_reg_754[3], r_reg_754[3], r_reg_754[3], r_reg_754[3], r_reg_754[3], r_reg_754[3], r_reg_754, 3'h0 };
assign sext_ln703_1_fu_250_p1 = { r_reg_754[3], r_reg_754[3], r_reg_754[3], r_reg_754[3], r_reg_754[3], r_reg_754[3], r_reg_754[3], r_reg_754[3], r_reg_754[3], r_reg_754[3], r_reg_754[3], r_reg_754[3], r_reg_754 };
assign sext_ln703_3_fu_521_p0 = op_12;
assign sext_ln703_4_fu_604_p0 = op_15;
assign sext_ln831_fu_377_p1 = { tmp_reg_838[18], tmp_reg_838[18], tmp_reg_838[18], tmp_reg_838[18], tmp_reg_838[18], tmp_reg_838[18], tmp_reg_838[18], tmp_reg_838[18], tmp_reg_838[18], tmp_reg_838[18], tmp_reg_838[18], tmp_reg_838[18], tmp_reg_838[18], tmp_reg_838 };
assign tmp_5_fu_304_p3 = { ret_V_2_reg_780, 3'h0 };
assign trunc_ln69_1_fu_649_p1 = op_8[0];
assign trunc_ln69_fu_645_p1 = op_4[0];
assign trunc_ln851_1_fu_458_p1 = op_11_V_fu_431_p3[2:0];
assign trunc_ln851_2_fu_542_p0 = op_12;
assign trunc_ln851_2_fu_542_p1 = op_12[13:0];
assign trunc_ln851_3_fu_625_p0 = op_15;
assign trunc_ln851_3_fu_625_p1 = op_15[1:0];
assign trunc_ln851_fu_321_p0 = op_10;
assign trunc_ln851_fu_321_p1 = op_10[2:0];
assign \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.ain_s0  = \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.a ;
assign \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.s  = { \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.fas_s2 , \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.sum_s1  };
assign \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.u2.a  = \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.ain_s1 ;
assign \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.u2.b  = \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.bin_s1 ;
assign \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.u2.cin  = \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.carry_s1 ;
assign \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.facout_s2  = \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.u2.cout ;
assign \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.fas_s2  = \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.u2.s ;
assign \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.u1.a  = \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.a [1:0];
assign \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.u1.b  = \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.bin_s0 [1:0];
assign \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.u1.cin  = 1'h1;
assign \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.facout_s1  = \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.u1.cout ;
assign \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.fas_s1  = \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.u1.s ;
assign \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.a  = \sub_4ns_4ns_4_2_1_U1.din0 ;
assign \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.b  = \sub_4ns_4ns_4_2_1_U1.din1 ;
assign \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.ce  = \sub_4ns_4ns_4_2_1_U1.ce ;
assign \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.clk  = \sub_4ns_4ns_4_2_1_U1.clk ;
assign \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.reset  = \sub_4ns_4ns_4_2_1_U1.reset ;
assign \sub_4ns_4ns_4_2_1_U1.dout  = \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.s ;
assign \sub_4ns_4ns_4_2_1_U1.ce  = 1'h1;
assign \sub_4ns_4ns_4_2_1_U1.clk  = ap_clk;
assign \sub_4ns_4ns_4_2_1_U1.din0  = 4'h0;
assign \sub_4ns_4ns_4_2_1_U1.din1  = op_1;
assign grp_fu_227_p2 = \sub_4ns_4ns_4_2_1_U1.dout ;
assign \sub_4ns_4ns_4_2_1_U1.reset  = ap_rst;
assign \sub_36s_36ns_36_2_1_U6.top_sub_36s_36ns_36_2_1_Adder_3_U.ain_s0  = \sub_36s_36ns_36_2_1_U6.top_sub_36s_36ns_36_2_1_Adder_3_U.a ;
assign \sub_36s_36ns_36_2_1_U6.top_sub_36s_36ns_36_2_1_Adder_3_U.s  = { \sub_36s_36ns_36_2_1_U6.top_sub_36s_36ns_36_2_1_Adder_3_U.fas_s2 , \sub_36s_36ns_36_2_1_U6.top_sub_36s_36ns_36_2_1_Adder_3_U.sum_s1  };
assign \sub_36s_36ns_36_2_1_U6.top_sub_36s_36ns_36_2_1_Adder_3_U.u2.a  = \sub_36s_36ns_36_2_1_U6.top_sub_36s_36ns_36_2_1_Adder_3_U.ain_s1 ;
assign \sub_36s_36ns_36_2_1_U6.top_sub_36s_36ns_36_2_1_Adder_3_U.u2.b  = \sub_36s_36ns_36_2_1_U6.top_sub_36s_36ns_36_2_1_Adder_3_U.bin_s1 ;
assign \sub_36s_36ns_36_2_1_U6.top_sub_36s_36ns_36_2_1_Adder_3_U.u2.cin  = \sub_36s_36ns_36_2_1_U6.top_sub_36s_36ns_36_2_1_Adder_3_U.carry_s1 ;
assign \sub_36s_36ns_36_2_1_U6.top_sub_36s_36ns_36_2_1_Adder_3_U.facout_s2  = \sub_36s_36ns_36_2_1_U6.top_sub_36s_36ns_36_2_1_Adder_3_U.u2.cout ;
assign \sub_36s_36ns_36_2_1_U6.top_sub_36s_36ns_36_2_1_Adder_3_U.fas_s2  = \sub_36s_36ns_36_2_1_U6.top_sub_36s_36ns_36_2_1_Adder_3_U.u2.s ;
assign \sub_36s_36ns_36_2_1_U6.top_sub_36s_36ns_36_2_1_Adder_3_U.u1.a  = \sub_36s_36ns_36_2_1_U6.top_sub_36s_36ns_36_2_1_Adder_3_U.a [17:0];
assign \sub_36s_36ns_36_2_1_U6.top_sub_36s_36ns_36_2_1_Adder_3_U.u1.b  = \sub_36s_36ns_36_2_1_U6.top_sub_36s_36ns_36_2_1_Adder_3_U.bin_s0 [17:0];
assign \sub_36s_36ns_36_2_1_U6.top_sub_36s_36ns_36_2_1_Adder_3_U.u1.cin  = 1'h1;
assign \sub_36s_36ns_36_2_1_U6.top_sub_36s_36ns_36_2_1_Adder_3_U.facout_s1  = \sub_36s_36ns_36_2_1_U6.top_sub_36s_36ns_36_2_1_Adder_3_U.u1.cout ;
assign \sub_36s_36ns_36_2_1_U6.top_sub_36s_36ns_36_2_1_Adder_3_U.fas_s1  = \sub_36s_36ns_36_2_1_U6.top_sub_36s_36ns_36_2_1_Adder_3_U.u1.s ;
assign \sub_36s_36ns_36_2_1_U6.top_sub_36s_36ns_36_2_1_Adder_3_U.a  = \sub_36s_36ns_36_2_1_U6.din0 ;
assign \sub_36s_36ns_36_2_1_U6.top_sub_36s_36ns_36_2_1_Adder_3_U.b  = \sub_36s_36ns_36_2_1_U6.din1 ;
assign \sub_36s_36ns_36_2_1_U6.top_sub_36s_36ns_36_2_1_Adder_3_U.ce  = \sub_36s_36ns_36_2_1_U6.ce ;
assign \sub_36s_36ns_36_2_1_U6.top_sub_36s_36ns_36_2_1_Adder_3_U.clk  = \sub_36s_36ns_36_2_1_U6.clk ;
assign \sub_36s_36ns_36_2_1_U6.top_sub_36s_36ns_36_2_1_Adder_3_U.reset  = \sub_36s_36ns_36_2_1_U6.reset ;
assign \sub_36s_36ns_36_2_1_U6.dout  = \sub_36s_36ns_36_2_1_U6.top_sub_36s_36ns_36_2_1_Adder_3_U.s ;
assign \sub_36s_36ns_36_2_1_U6.ce  = 1'h1;
assign \sub_36s_36ns_36_2_1_U6.clk  = ap_clk;
assign \sub_36s_36ns_36_2_1_U6.din0  = { op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6 };
assign \sub_36s_36ns_36_2_1_U6.din1  = { 1'h0, r_reg_754[3], r_reg_754[3], r_reg_754[3], r_reg_754[3], r_reg_754[3], r_reg_754[3], r_reg_754[3], r_reg_754[3], r_reg_754[3], r_reg_754[3], r_reg_754[3], r_reg_754[3], r_reg_754[3], r_reg_754[3], r_reg_754[3], r_reg_754[3], r_reg_754[3], r_reg_754[3], r_reg_754[3], r_reg_754[3], r_reg_754[3], r_reg_754[3], r_reg_754[3], r_reg_754[3], r_reg_754[3], r_reg_754[3], r_reg_754[3], r_reg_754[3], r_reg_754, 3'h0 };
assign grp_fu_294_p2 = \sub_36s_36ns_36_2_1_U6.dout ;
assign \sub_36s_36ns_36_2_1_U6.reset  = ap_rst;
assign \shl_4ns_4ns_4_7_1_U3.din1_cast  = \shl_4ns_4ns_4_7_1_U3.din1 ;
assign \shl_4ns_4ns_4_7_1_U3.din1_mask  = 4'h1;
assign \shl_4ns_4ns_4_7_1_U3.ce  = 1'h1;
assign \shl_4ns_4ns_4_7_1_U3.clk  = ap_clk;
assign \shl_4ns_4ns_4_7_1_U3.din0  = op_1;
assign \shl_4ns_4ns_4_7_1_U3.din1  = op_1;
assign grp_fu_237_p2 = \shl_4ns_4ns_4_7_1_U3.dout ;
assign \shl_4ns_4ns_4_7_1_U3.reset  = ap_rst;
assign \ashr_4ns_4ns_4_7_1_U2.din1_cast  = \ashr_4ns_4ns_4_7_1_U2.din1 ;
assign \ashr_4ns_4ns_4_7_1_U2.din1_mask  = 4'h1;
assign \ashr_4ns_4ns_4_7_1_U2.ce  = 1'h1;
assign \ashr_4ns_4ns_4_7_1_U2.clk  = ap_clk;
assign \ashr_4ns_4ns_4_7_1_U2.din0  = op_1;
assign \ashr_4ns_4ns_4_7_1_U2.din1  = sh_reg_739;
assign grp_fu_233_p2 = \ashr_4ns_4ns_4_7_1_U2.dout ;
assign \ashr_4ns_4ns_4_7_1_U2.reset  = ap_rst;
assign \add_47s_47s_47_2_1_U11.top_add_47s_47s_47_2_1_Adder_8_U.ain_s0  = \add_47s_47s_47_2_1_U11.top_add_47s_47s_47_2_1_Adder_8_U.a ;
assign \add_47s_47s_47_2_1_U11.top_add_47s_47s_47_2_1_Adder_8_U.bin_s0  = \add_47s_47s_47_2_1_U11.top_add_47s_47s_47_2_1_Adder_8_U.b ;
assign \add_47s_47s_47_2_1_U11.top_add_47s_47s_47_2_1_Adder_8_U.s  = { \add_47s_47s_47_2_1_U11.top_add_47s_47s_47_2_1_Adder_8_U.fas_s2 , \add_47s_47s_47_2_1_U11.top_add_47s_47s_47_2_1_Adder_8_U.sum_s1  };
assign \add_47s_47s_47_2_1_U11.top_add_47s_47s_47_2_1_Adder_8_U.u2.a  = \add_47s_47s_47_2_1_U11.top_add_47s_47s_47_2_1_Adder_8_U.ain_s1 ;
assign \add_47s_47s_47_2_1_U11.top_add_47s_47s_47_2_1_Adder_8_U.u2.b  = \add_47s_47s_47_2_1_U11.top_add_47s_47s_47_2_1_Adder_8_U.bin_s1 ;
assign \add_47s_47s_47_2_1_U11.top_add_47s_47s_47_2_1_Adder_8_U.u2.cin  = \add_47s_47s_47_2_1_U11.top_add_47s_47s_47_2_1_Adder_8_U.carry_s1 ;
assign \add_47s_47s_47_2_1_U11.top_add_47s_47s_47_2_1_Adder_8_U.facout_s2  = \add_47s_47s_47_2_1_U11.top_add_47s_47s_47_2_1_Adder_8_U.u2.cout ;
assign \add_47s_47s_47_2_1_U11.top_add_47s_47s_47_2_1_Adder_8_U.fas_s2  = \add_47s_47s_47_2_1_U11.top_add_47s_47s_47_2_1_Adder_8_U.u2.s ;
assign \add_47s_47s_47_2_1_U11.top_add_47s_47s_47_2_1_Adder_8_U.u1.a  = \add_47s_47s_47_2_1_U11.top_add_47s_47s_47_2_1_Adder_8_U.a [22:0];
assign \add_47s_47s_47_2_1_U11.top_add_47s_47s_47_2_1_Adder_8_U.u1.b  = \add_47s_47s_47_2_1_U11.top_add_47s_47s_47_2_1_Adder_8_U.b [22:0];
assign \add_47s_47s_47_2_1_U11.top_add_47s_47s_47_2_1_Adder_8_U.u1.cin  = 1'h0;
assign \add_47s_47s_47_2_1_U11.top_add_47s_47s_47_2_1_Adder_8_U.facout_s1  = \add_47s_47s_47_2_1_U11.top_add_47s_47s_47_2_1_Adder_8_U.u1.cout ;
assign \add_47s_47s_47_2_1_U11.top_add_47s_47s_47_2_1_Adder_8_U.fas_s1  = \add_47s_47s_47_2_1_U11.top_add_47s_47s_47_2_1_Adder_8_U.u1.s ;
assign \add_47s_47s_47_2_1_U11.top_add_47s_47s_47_2_1_Adder_8_U.a  = \add_47s_47s_47_2_1_U11.din0 ;
assign \add_47s_47s_47_2_1_U11.top_add_47s_47s_47_2_1_Adder_8_U.b  = \add_47s_47s_47_2_1_U11.din1 ;
assign \add_47s_47s_47_2_1_U11.top_add_47s_47s_47_2_1_Adder_8_U.ce  = \add_47s_47s_47_2_1_U11.ce ;
assign \add_47s_47s_47_2_1_U11.top_add_47s_47s_47_2_1_Adder_8_U.clk  = \add_47s_47s_47_2_1_U11.clk ;
assign \add_47s_47s_47_2_1_U11.top_add_47s_47s_47_2_1_Adder_8_U.reset  = \add_47s_47s_47_2_1_U11.reset ;
assign \add_47s_47s_47_2_1_U11.dout  = \add_47s_47s_47_2_1_U11.top_add_47s_47s_47_2_1_Adder_8_U.s ;
assign \add_47s_47s_47_2_1_U11.ce  = 1'h1;
assign \add_47s_47s_47_2_1_U11.clk  = ap_clk;
assign \add_47s_47s_47_2_1_U11.din0  = { select_ln353_1_reg_918[31], select_ln353_1_reg_918, 14'h0000 };
assign \add_47s_47s_47_2_1_U11.din1  = { op_12[31], op_12[31], op_12[31], op_12[31], op_12[31], op_12[31], op_12[31], op_12[31], op_12[31], op_12[31], op_12[31], op_12[31], op_12[31], op_12[31], op_12[31], op_12 };
assign grp_fu_536_p2 = \add_47s_47s_47_2_1_U11.dout ;
assign \add_47s_47s_47_2_1_U11.reset  = ap_rst;
assign \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_6_U.ain_s0  = \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_6_U.a ;
assign \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_6_U.bin_s0  = \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_6_U.b ;
assign \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_6_U.s  = { \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_6_U.fas_s2 , \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_6_U.sum_s1  };
assign \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_6_U.u2.a  = \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_6_U.ain_s1 ;
assign \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_6_U.u2.b  = \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_6_U.bin_s1 ;
assign \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_6_U.u2.cin  = \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_6_U.carry_s1 ;
assign \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_6_U.facout_s2  = \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_6_U.u2.cout ;
assign \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_6_U.fas_s2  = \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_6_U.u2.s ;
assign \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_6_U.u1.a  = \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_6_U.a [17:0];
assign \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_6_U.u1.b  = \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_6_U.b [17:0];
assign \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_6_U.u1.cin  = 1'h0;
assign \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_6_U.facout_s1  = \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_6_U.u1.cout ;
assign \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_6_U.fas_s1  = \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_6_U.u1.s ;
assign \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_6_U.a  = \add_36s_36s_36_2_1_U9.din0 ;
assign \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_6_U.b  = \add_36s_36s_36_2_1_U9.din1 ;
assign \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_6_U.ce  = \add_36s_36s_36_2_1_U9.ce ;
assign \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_6_U.clk  = \add_36s_36s_36_2_1_U9.clk ;
assign \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_6_U.reset  = \add_36s_36s_36_2_1_U9.reset ;
assign \add_36s_36s_36_2_1_U9.dout  = \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_6_U.s ;
assign \add_36s_36s_36_2_1_U9.ce  = 1'h1;
assign \add_36s_36s_36_2_1_U9.clk  = ap_clk;
assign \add_36s_36s_36_2_1_U9.din0  = { select_ln353_reg_876[31], select_ln353_reg_876, 3'h0 };
assign \add_36s_36s_36_2_1_U9.din1  = { op_11_V_reg_871[3], op_11_V_reg_871[3], op_11_V_reg_871[3], op_11_V_reg_871[3], op_11_V_reg_871[3], op_11_V_reg_871[3], op_11_V_reg_871[3], op_11_V_reg_871[3], op_11_V_reg_871[3], op_11_V_reg_871[3], op_11_V_reg_871[3], op_11_V_reg_871[3], op_11_V_reg_871[3], op_11_V_reg_871[3], op_11_V_reg_871[3], op_11_V_reg_871[3], op_11_V_reg_871[3], op_11_V_reg_871[3], op_11_V_reg_871[3], op_11_V_reg_871[3], op_11_V_reg_871[3], op_11_V_reg_871[3], op_11_V_reg_871[3], op_11_V_reg_871[3], op_11_V_reg_871[3], op_11_V_reg_871[3], op_11_V_reg_871[3], op_11_V_reg_871[3], op_11_V_reg_871[3], op_11_V_reg_871[3], op_11_V_reg_871[3], op_11_V_reg_871[3], op_11_V_reg_871 };
assign grp_fu_476_p2 = \add_36s_36s_36_2_1_U9.dout ;
assign \add_36s_36s_36_2_1_U9.reset  = ap_rst;
assign \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_10_U.ain_s0  = \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_10_U.a ;
assign \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_10_U.bin_s0  = \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_10_U.b ;
assign \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_10_U.s  = { \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_10_U.fas_s2 , \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_10_U.sum_s1  };
assign \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_10_U.u2.a  = \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_10_U.ain_s1 ;
assign \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_10_U.u2.b  = \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_10_U.bin_s1 ;
assign \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_10_U.u2.cin  = \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_10_U.carry_s1 ;
assign \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_10_U.facout_s2  = \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_10_U.u2.cout ;
assign \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_10_U.fas_s2  = \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_10_U.u2.s ;
assign \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_10_U.u1.a  = \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_10_U.a [16:0];
assign \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_10_U.u1.b  = \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_10_U.b [16:0];
assign \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_10_U.u1.cin  = 1'h0;
assign \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_10_U.facout_s1  = \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_10_U.u1.cout ;
assign \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_10_U.fas_s1  = \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_10_U.u1.s ;
assign \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_10_U.a  = \add_35s_35s_35_2_1_U15.din0 ;
assign \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_10_U.b  = \add_35s_35s_35_2_1_U15.din1 ;
assign \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_10_U.ce  = \add_35s_35s_35_2_1_U15.ce ;
assign \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_10_U.clk  = \add_35s_35s_35_2_1_U15.clk ;
assign \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_10_U.reset  = \add_35s_35s_35_2_1_U15.reset ;
assign \add_35s_35s_35_2_1_U15.dout  = \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_10_U.s ;
assign \add_35s_35s_35_2_1_U15.ce  = 1'h1;
assign \add_35s_35s_35_2_1_U15.clk  = ap_clk;
assign \add_35s_35s_35_2_1_U15.din0  = { op_26_V_reg_975[31], op_26_V_reg_975, 2'h0 };
assign \add_35s_35s_35_2_1_U15.din1  = { op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15 };
assign grp_fu_619_p2 = \add_35s_35s_35_2_1_U15.dout ;
assign \add_35s_35s_35_2_1_U15.reset  = ap_rst;
assign \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.ain_s0  = \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.a ;
assign \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.bin_s0  = \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.b ;
assign \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.s  = { \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.fas_s2 , \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.sum_s1  };
assign \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.u2.a  = \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.ain_s1 ;
assign \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.u2.b  = \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.bin_s1 ;
assign \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.u2.cin  = \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.carry_s1 ;
assign \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.facout_s2  = \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.u2.cout ;
assign \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.fas_s2  = \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.u2.s ;
assign \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.u1.a  = \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.a [15:0];
assign \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.u1.b  = \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.b [15:0];
assign \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.u1.cin  = 1'h0;
assign \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.facout_s1  = \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.u1.cout ;
assign \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.fas_s1  = \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.u1.s ;
assign \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.a  = \add_32s_32ns_32_2_1_U8.din0 ;
assign \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.b  = \add_32s_32ns_32_2_1_U8.din1 ;
assign \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.ce  = \add_32s_32ns_32_2_1_U8.ce ;
assign \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.clk  = \add_32s_32ns_32_2_1_U8.clk ;
assign \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.reset  = \add_32s_32ns_32_2_1_U8.reset ;
assign \add_32s_32ns_32_2_1_U8.dout  = \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.s ;
assign \add_32s_32ns_32_2_1_U8.ce  = 1'h1;
assign \add_32s_32ns_32_2_1_U8.clk  = ap_clk;
assign \add_32s_32ns_32_2_1_U8.din0  = { tmp_reg_838[18], tmp_reg_838[18], tmp_reg_838[18], tmp_reg_838[18], tmp_reg_838[18], tmp_reg_838[18], tmp_reg_838[18], tmp_reg_838[18], tmp_reg_838[18], tmp_reg_838[18], tmp_reg_838[18], tmp_reg_838[18], tmp_reg_838[18], tmp_reg_838 };
assign \add_32s_32ns_32_2_1_U8.din1  = 32'd1;
assign grp_fu_380_p2 = \add_32s_32ns_32_2_1_U8.dout ;
assign \add_32s_32ns_32_2_1_U8.reset  = ap_rst;
assign \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_5_U.ain_s0  = \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_5_U.a ;
assign \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_5_U.bin_s0  = \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_5_U.b ;
assign \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_5_U.s  = { \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_5_U.fas_s2 , \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_5_U.sum_s1  };
assign \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_5_U.u2.a  = \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_5_U.ain_s1 ;
assign \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_5_U.u2.b  = \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_5_U.bin_s1 ;
assign \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_5_U.u2.cin  = \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_5_U.carry_s1 ;
assign \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_5_U.facout_s2  = \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_5_U.u2.cout ;
assign \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_5_U.fas_s2  = \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_5_U.u2.s ;
assign \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_5_U.u1.a  = \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_5_U.a [15:0];
assign \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_5_U.u1.b  = \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_5_U.b [15:0];
assign \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_5_U.u1.cin  = 1'h0;
assign \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_5_U.facout_s1  = \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_5_U.u1.cout ;
assign \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_5_U.fas_s1  = \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_5_U.u1.s ;
assign \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_5_U.a  = \add_32s_32ns_32_2_1_U20.din0 ;
assign \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_5_U.b  = \add_32s_32ns_32_2_1_U20.din1 ;
assign \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_5_U.ce  = \add_32s_32ns_32_2_1_U20.ce ;
assign \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_5_U.clk  = \add_32s_32ns_32_2_1_U20.clk ;
assign \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_5_U.reset  = \add_32s_32ns_32_2_1_U20.reset ;
assign \add_32s_32ns_32_2_1_U20.dout  = \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_5_U.s ;
assign \add_32s_32ns_32_2_1_U20.ce  = 1'h1;
assign \add_32s_32ns_32_2_1_U20.clk  = ap_clk;
assign \add_32s_32ns_32_2_1_U20.din0  = { add_ln69_2_reg_1047[1], add_ln69_2_reg_1047[1], add_ln69_2_reg_1047[1], add_ln69_2_reg_1047[1], add_ln69_2_reg_1047[1], add_ln69_2_reg_1047[1], add_ln69_2_reg_1047[1], add_ln69_2_reg_1047[1], add_ln69_2_reg_1047[1], add_ln69_2_reg_1047[1], add_ln69_2_reg_1047[1], add_ln69_2_reg_1047[1], add_ln69_2_reg_1047[1], add_ln69_2_reg_1047[1], add_ln69_2_reg_1047[1], add_ln69_2_reg_1047[1], add_ln69_2_reg_1047[1], add_ln69_2_reg_1047[1], add_ln69_2_reg_1047[1], add_ln69_2_reg_1047[1], add_ln69_2_reg_1047[1], add_ln69_2_reg_1047[1], add_ln69_2_reg_1047[1], add_ln69_2_reg_1047[1], add_ln69_2_reg_1047[1], add_ln69_2_reg_1047[1], add_ln69_2_reg_1047[1], add_ln69_2_reg_1047[1], add_ln69_2_reg_1047[1], add_ln69_2_reg_1047[1], add_ln69_2_reg_1047 };
assign \add_32s_32ns_32_2_1_U20.din1  = add_ln69_reg_1042;
assign grp_fu_720_p2 = \add_32s_32ns_32_2_1_U20.dout ;
assign \add_32s_32ns_32_2_1_U20.reset  = ap_rst;
assign \add_32ns_32s_32_2_1_U13.top_add_32ns_32s_32_2_1_Adder_9_U.ain_s0  = \add_32ns_32s_32_2_1_U13.top_add_32ns_32s_32_2_1_Adder_9_U.a ;
assign \add_32ns_32s_32_2_1_U13.top_add_32ns_32s_32_2_1_Adder_9_U.bin_s0  = \add_32ns_32s_32_2_1_U13.top_add_32ns_32s_32_2_1_Adder_9_U.b ;
assign \add_32ns_32s_32_2_1_U13.top_add_32ns_32s_32_2_1_Adder_9_U.s  = { \add_32ns_32s_32_2_1_U13.top_add_32ns_32s_32_2_1_Adder_9_U.fas_s2 , \add_32ns_32s_32_2_1_U13.top_add_32ns_32s_32_2_1_Adder_9_U.sum_s1  };
assign \add_32ns_32s_32_2_1_U13.top_add_32ns_32s_32_2_1_Adder_9_U.u2.a  = \add_32ns_32s_32_2_1_U13.top_add_32ns_32s_32_2_1_Adder_9_U.ain_s1 ;
assign \add_32ns_32s_32_2_1_U13.top_add_32ns_32s_32_2_1_Adder_9_U.u2.b  = \add_32ns_32s_32_2_1_U13.top_add_32ns_32s_32_2_1_Adder_9_U.bin_s1 ;
assign \add_32ns_32s_32_2_1_U13.top_add_32ns_32s_32_2_1_Adder_9_U.u2.cin  = \add_32ns_32s_32_2_1_U13.top_add_32ns_32s_32_2_1_Adder_9_U.carry_s1 ;
assign \add_32ns_32s_32_2_1_U13.top_add_32ns_32s_32_2_1_Adder_9_U.facout_s2  = \add_32ns_32s_32_2_1_U13.top_add_32ns_32s_32_2_1_Adder_9_U.u2.cout ;
assign \add_32ns_32s_32_2_1_U13.top_add_32ns_32s_32_2_1_Adder_9_U.fas_s2  = \add_32ns_32s_32_2_1_U13.top_add_32ns_32s_32_2_1_Adder_9_U.u2.s ;
assign \add_32ns_32s_32_2_1_U13.top_add_32ns_32s_32_2_1_Adder_9_U.u1.a  = \add_32ns_32s_32_2_1_U13.top_add_32ns_32s_32_2_1_Adder_9_U.a [15:0];
assign \add_32ns_32s_32_2_1_U13.top_add_32ns_32s_32_2_1_Adder_9_U.u1.b  = \add_32ns_32s_32_2_1_U13.top_add_32ns_32s_32_2_1_Adder_9_U.b [15:0];
assign \add_32ns_32s_32_2_1_U13.top_add_32ns_32s_32_2_1_Adder_9_U.u1.cin  = 1'h0;
assign \add_32ns_32s_32_2_1_U13.top_add_32ns_32s_32_2_1_Adder_9_U.facout_s1  = \add_32ns_32s_32_2_1_U13.top_add_32ns_32s_32_2_1_Adder_9_U.u1.cout ;
assign \add_32ns_32s_32_2_1_U13.top_add_32ns_32s_32_2_1_Adder_9_U.fas_s1  = \add_32ns_32s_32_2_1_U13.top_add_32ns_32s_32_2_1_Adder_9_U.u1.s ;
assign \add_32ns_32s_32_2_1_U13.top_add_32ns_32s_32_2_1_Adder_9_U.a  = \add_32ns_32s_32_2_1_U13.din0 ;
assign \add_32ns_32s_32_2_1_U13.top_add_32ns_32s_32_2_1_Adder_9_U.b  = \add_32ns_32s_32_2_1_U13.din1 ;
assign \add_32ns_32s_32_2_1_U13.top_add_32ns_32s_32_2_1_Adder_9_U.ce  = \add_32ns_32s_32_2_1_U13.ce ;
assign \add_32ns_32s_32_2_1_U13.top_add_32ns_32s_32_2_1_Adder_9_U.clk  = \add_32ns_32s_32_2_1_U13.clk ;
assign \add_32ns_32s_32_2_1_U13.top_add_32ns_32s_32_2_1_Adder_9_U.reset  = \add_32ns_32s_32_2_1_U13.reset ;
assign \add_32ns_32s_32_2_1_U13.dout  = \add_32ns_32s_32_2_1_U13.top_add_32ns_32s_32_2_1_Adder_9_U.s ;
assign \add_32ns_32s_32_2_1_U13.ce  = 1'h1;
assign \add_32ns_32s_32_2_1_U13.clk  = ap_clk;
assign \add_32ns_32s_32_2_1_U13.din0  = ret_V_6_reg_955;
assign \add_32ns_32s_32_2_1_U13.din1  = { op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13 };
assign grp_fu_590_p2 = \add_32ns_32s_32_2_1_U13.dout ;
assign \add_32ns_32s_32_2_1_U13.reset  = ap_rst;
assign \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s0  = \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.a ;
assign \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s0  = \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.b ;
assign \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.s  = { \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s2 , \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.sum_s1  };
assign \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.a  = \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s1 ;
assign \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.b  = \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s1 ;
assign \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cin  = \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.carry_s1 ;
assign \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.facout_s2  = \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cout ;
assign \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s2  = \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.s ;
assign \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.a  = \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.a [15:0];
assign \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.b  = \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.b [15:0];
assign \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cin  = 1'h0;
assign \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.facout_s1  = \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cout ;
assign \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s1  = \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.s ;
assign \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.a  = \add_32ns_32ns_32_2_1_U18.din0 ;
assign \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.b  = \add_32ns_32ns_32_2_1_U18.din1 ;
assign \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.ce  = \add_32ns_32ns_32_2_1_U18.ce ;
assign \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.clk  = \add_32ns_32ns_32_2_1_U18.clk ;
assign \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.reset  = \add_32ns_32ns_32_2_1_U18.reset ;
assign \add_32ns_32ns_32_2_1_U18.dout  = \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.s ;
assign \add_32ns_32ns_32_2_1_U18.ce  = 1'h1;
assign \add_32ns_32ns_32_2_1_U18.clk  = ap_clk;
assign \add_32ns_32ns_32_2_1_U18.din0  = ret_V_9_reg_1022;
assign \add_32ns_32ns_32_2_1_U18.din1  = op_19;
assign grp_fu_708_p2 = \add_32ns_32ns_32_2_1_U18.dout ;
assign \add_32ns_32ns_32_2_1_U18.reset  = ap_rst;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s0  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.a ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s0  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.b ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.s  = { \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s2 , \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.sum_s1  };
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.a  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s1 ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.b  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s1 ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cin  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.carry_s1 ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.facout_s2  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cout ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s2  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.s ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.a  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.a [15:0];
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.b  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.b [15:0];
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cin  = 1'h0;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.facout_s1  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cout ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s1  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.s ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.a  = \add_32ns_32ns_32_2_1_U16.din0 ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.b  = \add_32ns_32ns_32_2_1_U16.din1 ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.ce  = \add_32ns_32ns_32_2_1_U16.ce ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.clk  = \add_32ns_32ns_32_2_1_U16.clk ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.reset  = \add_32ns_32ns_32_2_1_U16.reset ;
assign \add_32ns_32ns_32_2_1_U16.dout  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.s ;
assign \add_32ns_32ns_32_2_1_U16.ce  = 1'h1;
assign \add_32ns_32ns_32_2_1_U16.clk  = ap_clk;
assign \add_32ns_32ns_32_2_1_U16.din0  = ret_V_16_cast_reg_1000;
assign \add_32ns_32ns_32_2_1_U16.din1  = 32'd1;
assign grp_fu_659_p2 = \add_32ns_32ns_32_2_1_U16.dout ;
assign \add_32ns_32ns_32_2_1_U16.reset  = ap_rst;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s0  = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.a ;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s0  = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.b ;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.s  = { \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s2 , \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.sum_s1  };
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.a  = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s1 ;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.b  = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s1 ;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cin  = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.carry_s1 ;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.facout_s2  = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cout ;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s2  = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.s ;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.a  = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.a [15:0];
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.b  = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.b [15:0];
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cin  = 1'h0;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.facout_s1  = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cout ;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s1  = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.s ;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.a  = \add_32ns_32ns_32_2_1_U14.din0 ;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.b  = \add_32ns_32ns_32_2_1_U14.din1 ;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.ce  = \add_32ns_32ns_32_2_1_U14.ce ;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.clk  = \add_32ns_32ns_32_2_1_U14.clk ;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.reset  = \add_32ns_32ns_32_2_1_U14.reset ;
assign \add_32ns_32ns_32_2_1_U14.dout  = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.s ;
assign \add_32ns_32ns_32_2_1_U14.ce  = 1'h1;
assign \add_32ns_32ns_32_2_1_U14.clk  = ap_clk;
assign \add_32ns_32ns_32_2_1_U14.din0  = ret_V_7_reg_965;
assign \add_32ns_32ns_32_2_1_U14.din1  = { 30'h00000000, op_14 };
assign grp_fu_599_p2 = \add_32ns_32ns_32_2_1_U14.dout ;
assign \add_32ns_32ns_32_2_1_U14.reset  = ap_rst;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s0  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.a ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s0  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.b ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.s  = { \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s2 , \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.sum_s1  };
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.a  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s1 ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.b  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s1 ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cin  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.carry_s1 ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.facout_s2  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cout ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s2  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.s ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.a  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.a [15:0];
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.b  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.b [15:0];
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cin  = 1'h0;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.facout_s1  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cout ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s1  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.s ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.a  = \add_32ns_32ns_32_2_1_U12.din0 ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.b  = \add_32ns_32ns_32_2_1_U12.din1 ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.ce  = \add_32ns_32ns_32_2_1_U12.ce ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.clk  = \add_32ns_32ns_32_2_1_U12.clk ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.reset  = \add_32ns_32ns_32_2_1_U12.reset ;
assign \add_32ns_32ns_32_2_1_U12.dout  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.s ;
assign \add_32ns_32ns_32_2_1_U12.ce  = 1'h1;
assign \add_32ns_32ns_32_2_1_U12.clk  = ap_clk;
assign \add_32ns_32ns_32_2_1_U12.din0  = ret_V_6_cast_reg_943;
assign \add_32ns_32ns_32_2_1_U12.din1  = 32'd1;
assign grp_fu_562_p2 = \add_32ns_32ns_32_2_1_U12.dout ;
assign \add_32ns_32ns_32_2_1_U12.reset  = ap_rst;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s0  = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.a ;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s0  = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.b ;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.s  = { \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s2 , \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.sum_s1  };
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.a  = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s1 ;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.b  = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s1 ;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cin  = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.carry_s1 ;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.facout_s2  = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cout ;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s2  = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.s ;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.a  = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.a [15:0];
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.b  = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.b [15:0];
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cin  = 1'h0;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.facout_s1  = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cout ;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s1  = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.s ;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.a  = \add_32ns_32ns_32_2_1_U10.din0 ;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.b  = \add_32ns_32ns_32_2_1_U10.din1 ;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.ce  = \add_32ns_32ns_32_2_1_U10.ce ;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.clk  = \add_32ns_32ns_32_2_1_U10.clk ;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.reset  = \add_32ns_32ns_32_2_1_U10.reset ;
assign \add_32ns_32ns_32_2_1_U10.dout  = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_7_U.s ;
assign \add_32ns_32ns_32_2_1_U10.ce  = 1'h1;
assign \add_32ns_32ns_32_2_1_U10.clk  = ap_clk;
assign \add_32ns_32ns_32_2_1_U10.din0  = ret_V_3_cast_reg_906;
assign \add_32ns_32ns_32_2_1_U10.din1  = 32'd1;
assign grp_fu_497_p2 = \add_32ns_32ns_32_2_1_U10.dout ;
assign \add_32ns_32ns_32_2_1_U10.reset  = ap_rst;
assign \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_11_U.ain_s0  = \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_11_U.a ;
assign \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_11_U.bin_s0  = \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_11_U.b ;
assign \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_11_U.s  = { \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_11_U.fas_s2 , \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_11_U.sum_s1  };
assign \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_11_U.u2.a  = \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_11_U.ain_s1 ;
assign \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_11_U.u2.b  = \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_11_U.bin_s1 ;
assign \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_11_U.u2.cin  = \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_11_U.carry_s1 ;
assign \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_11_U.facout_s2  = \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_11_U.u2.cout ;
assign \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_11_U.fas_s2  = \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_11_U.u2.s ;
assign \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_11_U.u1.a  = \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_11_U.a [0];
assign \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_11_U.u1.b  = \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_11_U.b [0];
assign \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_11_U.u1.cin  = 1'h0;
assign \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_11_U.facout_s1  = \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_11_U.u1.cout ;
assign \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_11_U.fas_s1  = \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_11_U.u1.s ;
assign \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_11_U.a  = \add_2ns_2ns_2_2_1_U19.din0 ;
assign \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_11_U.b  = \add_2ns_2ns_2_2_1_U19.din1 ;
assign \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_11_U.ce  = \add_2ns_2ns_2_2_1_U19.ce ;
assign \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_11_U.clk  = \add_2ns_2ns_2_2_1_U19.clk ;
assign \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_11_U.reset  = \add_2ns_2ns_2_2_1_U19.reset ;
assign \add_2ns_2ns_2_2_1_U19.dout  = \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_11_U.s ;
assign \add_2ns_2ns_2_2_1_U19.ce  = 1'h1;
assign \add_2ns_2ns_2_2_1_U19.clk  = ap_clk;
assign \add_2ns_2ns_2_2_1_U19.din0  = add_ln69_1_reg_1032;
assign \add_2ns_2ns_2_2_1_U19.din1  = select_ln69_1_reg_1027;
assign grp_fu_713_p2 = \add_2ns_2ns_2_2_1_U19.dout ;
assign \add_2ns_2ns_2_2_1_U19.reset  = ap_rst;
assign \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_11_U.ain_s0  = \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_11_U.a ;
assign \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_11_U.bin_s0  = \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_11_U.b ;
assign \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_11_U.s  = { \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_11_U.fas_s2 , \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_11_U.sum_s1  };
assign \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_11_U.u2.a  = \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_11_U.ain_s1 ;
assign \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_11_U.u2.b  = \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_11_U.bin_s1 ;
assign \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_11_U.u2.cin  = \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_11_U.carry_s1 ;
assign \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_11_U.facout_s2  = \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_11_U.u2.cout ;
assign \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_11_U.fas_s2  = \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_11_U.u2.s ;
assign \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_11_U.u1.a  = \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_11_U.a [0];
assign \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_11_U.u1.b  = \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_11_U.b [0];
assign \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_11_U.u1.cin  = 1'h0;
assign \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_11_U.facout_s1  = \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_11_U.u1.cout ;
assign \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_11_U.fas_s1  = \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_11_U.u1.s ;
assign \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_11_U.a  = \add_2ns_2ns_2_2_1_U17.din0 ;
assign \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_11_U.b  = \add_2ns_2ns_2_2_1_U17.din1 ;
assign \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_11_U.ce  = \add_2ns_2ns_2_2_1_U17.ce ;
assign \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_11_U.clk  = \add_2ns_2ns_2_2_1_U17.clk ;
assign \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_11_U.reset  = \add_2ns_2ns_2_2_1_U17.reset ;
assign \add_2ns_2ns_2_2_1_U17.dout  = \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_11_U.s ;
assign \add_2ns_2ns_2_2_1_U17.ce  = 1'h1;
assign \add_2ns_2ns_2_2_1_U17.clk  = ap_clk;
assign \add_2ns_2ns_2_2_1_U17.din0  = select_ln69_reg_1007;
assign \add_2ns_2ns_2_2_1_U17.din1  = { 1'h0, op_18 };
assign grp_fu_676_p2 = \add_2ns_2ns_2_2_1_U17.dout ;
assign \add_2ns_2ns_2_2_1_U17.reset  = ap_rst;
assign \add_22s_22s_22_2_1_U7.top_add_22s_22s_22_2_1_Adder_4_U.ain_s0  = \add_22s_22s_22_2_1_U7.top_add_22s_22s_22_2_1_Adder_4_U.a ;
assign \add_22s_22s_22_2_1_U7.top_add_22s_22s_22_2_1_Adder_4_U.bin_s0  = \add_22s_22s_22_2_1_U7.top_add_22s_22s_22_2_1_Adder_4_U.b ;
assign \add_22s_22s_22_2_1_U7.top_add_22s_22s_22_2_1_Adder_4_U.s  = { \add_22s_22s_22_2_1_U7.top_add_22s_22s_22_2_1_Adder_4_U.fas_s2 , \add_22s_22s_22_2_1_U7.top_add_22s_22s_22_2_1_Adder_4_U.sum_s1  };
assign \add_22s_22s_22_2_1_U7.top_add_22s_22s_22_2_1_Adder_4_U.u2.a  = \add_22s_22s_22_2_1_U7.top_add_22s_22s_22_2_1_Adder_4_U.ain_s1 ;
assign \add_22s_22s_22_2_1_U7.top_add_22s_22s_22_2_1_Adder_4_U.u2.b  = \add_22s_22s_22_2_1_U7.top_add_22s_22s_22_2_1_Adder_4_U.bin_s1 ;
assign \add_22s_22s_22_2_1_U7.top_add_22s_22s_22_2_1_Adder_4_U.u2.cin  = \add_22s_22s_22_2_1_U7.top_add_22s_22s_22_2_1_Adder_4_U.carry_s1 ;
assign \add_22s_22s_22_2_1_U7.top_add_22s_22s_22_2_1_Adder_4_U.facout_s2  = \add_22s_22s_22_2_1_U7.top_add_22s_22s_22_2_1_Adder_4_U.u2.cout ;
assign \add_22s_22s_22_2_1_U7.top_add_22s_22s_22_2_1_Adder_4_U.fas_s2  = \add_22s_22s_22_2_1_U7.top_add_22s_22s_22_2_1_Adder_4_U.u2.s ;
assign \add_22s_22s_22_2_1_U7.top_add_22s_22s_22_2_1_Adder_4_U.u1.a  = \add_22s_22s_22_2_1_U7.top_add_22s_22s_22_2_1_Adder_4_U.a [10:0];
assign \add_22s_22s_22_2_1_U7.top_add_22s_22s_22_2_1_Adder_4_U.u1.b  = \add_22s_22s_22_2_1_U7.top_add_22s_22s_22_2_1_Adder_4_U.b [10:0];
assign \add_22s_22s_22_2_1_U7.top_add_22s_22s_22_2_1_Adder_4_U.u1.cin  = 1'h0;
assign \add_22s_22s_22_2_1_U7.top_add_22s_22s_22_2_1_Adder_4_U.facout_s1  = \add_22s_22s_22_2_1_U7.top_add_22s_22s_22_2_1_Adder_4_U.u1.cout ;
assign \add_22s_22s_22_2_1_U7.top_add_22s_22s_22_2_1_Adder_4_U.fas_s1  = \add_22s_22s_22_2_1_U7.top_add_22s_22s_22_2_1_Adder_4_U.u1.s ;
assign \add_22s_22s_22_2_1_U7.top_add_22s_22s_22_2_1_Adder_4_U.a  = \add_22s_22s_22_2_1_U7.din0 ;
assign \add_22s_22s_22_2_1_U7.top_add_22s_22s_22_2_1_Adder_4_U.b  = \add_22s_22s_22_2_1_U7.din1 ;
assign \add_22s_22s_22_2_1_U7.top_add_22s_22s_22_2_1_Adder_4_U.ce  = \add_22s_22s_22_2_1_U7.ce ;
assign \add_22s_22s_22_2_1_U7.top_add_22s_22s_22_2_1_Adder_4_U.clk  = \add_22s_22s_22_2_1_U7.clk ;
assign \add_22s_22s_22_2_1_U7.top_add_22s_22s_22_2_1_Adder_4_U.reset  = \add_22s_22s_22_2_1_U7.reset ;
assign \add_22s_22s_22_2_1_U7.dout  = \add_22s_22s_22_2_1_U7.top_add_22s_22s_22_2_1_Adder_4_U.s ;
assign \add_22s_22s_22_2_1_U7.ce  = 1'h1;
assign \add_22s_22s_22_2_1_U7.clk  = ap_clk;
assign \add_22s_22s_22_2_1_U7.din0  = { ret_V_2_reg_780[17], ret_V_2_reg_780, 3'h0 };
assign \add_22s_22s_22_2_1_U7.din1  = { op_10[3], op_10[3], op_10[3], op_10[3], op_10[3], op_10[3], op_10[3], op_10[3], op_10[3], op_10[3], op_10[3], op_10[3], op_10[3], op_10[3], op_10[3], op_10[3], op_10[3], op_10[3], op_10 };
assign grp_fu_315_p2 = \add_22s_22s_22_2_1_U7.dout ;
assign \add_22s_22s_22_2_1_U7.reset  = ap_rst;
assign \add_18ns_18s_18_2_1_U4.top_add_18ns_18s_18_2_1_Adder_1_U.ain_s0  = \add_18ns_18s_18_2_1_U4.top_add_18ns_18s_18_2_1_Adder_1_U.a ;
assign \add_18ns_18s_18_2_1_U4.top_add_18ns_18s_18_2_1_Adder_1_U.bin_s0  = \add_18ns_18s_18_2_1_U4.top_add_18ns_18s_18_2_1_Adder_1_U.b ;
assign \add_18ns_18s_18_2_1_U4.top_add_18ns_18s_18_2_1_Adder_1_U.s  = { \add_18ns_18s_18_2_1_U4.top_add_18ns_18s_18_2_1_Adder_1_U.fas_s2 , \add_18ns_18s_18_2_1_U4.top_add_18ns_18s_18_2_1_Adder_1_U.sum_s1  };
assign \add_18ns_18s_18_2_1_U4.top_add_18ns_18s_18_2_1_Adder_1_U.u2.a  = \add_18ns_18s_18_2_1_U4.top_add_18ns_18s_18_2_1_Adder_1_U.ain_s1 ;
assign \add_18ns_18s_18_2_1_U4.top_add_18ns_18s_18_2_1_Adder_1_U.u2.b  = \add_18ns_18s_18_2_1_U4.top_add_18ns_18s_18_2_1_Adder_1_U.bin_s1 ;
assign \add_18ns_18s_18_2_1_U4.top_add_18ns_18s_18_2_1_Adder_1_U.u2.cin  = \add_18ns_18s_18_2_1_U4.top_add_18ns_18s_18_2_1_Adder_1_U.carry_s1 ;
assign \add_18ns_18s_18_2_1_U4.top_add_18ns_18s_18_2_1_Adder_1_U.facout_s2  = \add_18ns_18s_18_2_1_U4.top_add_18ns_18s_18_2_1_Adder_1_U.u2.cout ;
assign \add_18ns_18s_18_2_1_U4.top_add_18ns_18s_18_2_1_Adder_1_U.fas_s2  = \add_18ns_18s_18_2_1_U4.top_add_18ns_18s_18_2_1_Adder_1_U.u2.s ;
assign \add_18ns_18s_18_2_1_U4.top_add_18ns_18s_18_2_1_Adder_1_U.u1.a  = \add_18ns_18s_18_2_1_U4.top_add_18ns_18s_18_2_1_Adder_1_U.a [8:0];
assign \add_18ns_18s_18_2_1_U4.top_add_18ns_18s_18_2_1_Adder_1_U.u1.b  = \add_18ns_18s_18_2_1_U4.top_add_18ns_18s_18_2_1_Adder_1_U.b [8:0];
assign \add_18ns_18s_18_2_1_U4.top_add_18ns_18s_18_2_1_Adder_1_U.u1.cin  = 1'h0;
assign \add_18ns_18s_18_2_1_U4.top_add_18ns_18s_18_2_1_Adder_1_U.facout_s1  = \add_18ns_18s_18_2_1_U4.top_add_18ns_18s_18_2_1_Adder_1_U.u1.cout ;
assign \add_18ns_18s_18_2_1_U4.top_add_18ns_18s_18_2_1_Adder_1_U.fas_s1  = \add_18ns_18s_18_2_1_U4.top_add_18ns_18s_18_2_1_Adder_1_U.u1.s ;
assign \add_18ns_18s_18_2_1_U4.top_add_18ns_18s_18_2_1_Adder_1_U.a  = \add_18ns_18s_18_2_1_U4.din0 ;
assign \add_18ns_18s_18_2_1_U4.top_add_18ns_18s_18_2_1_Adder_1_U.b  = \add_18ns_18s_18_2_1_U4.din1 ;
assign \add_18ns_18s_18_2_1_U4.top_add_18ns_18s_18_2_1_Adder_1_U.ce  = \add_18ns_18s_18_2_1_U4.ce ;
assign \add_18ns_18s_18_2_1_U4.top_add_18ns_18s_18_2_1_Adder_1_U.clk  = \add_18ns_18s_18_2_1_U4.clk ;
assign \add_18ns_18s_18_2_1_U4.top_add_18ns_18s_18_2_1_Adder_1_U.reset  = \add_18ns_18s_18_2_1_U4.reset ;
assign \add_18ns_18s_18_2_1_U4.dout  = \add_18ns_18s_18_2_1_U4.top_add_18ns_18s_18_2_1_Adder_1_U.s ;
assign \add_18ns_18s_18_2_1_U4.ce  = 1'h1;
assign \add_18ns_18s_18_2_1_U4.clk  = ap_clk;
assign \add_18ns_18s_18_2_1_U4.din0  = { 2'h0, r_reg_754[3], r_reg_754[3], r_reg_754[3], r_reg_754[3], r_reg_754[3], r_reg_754[3], r_reg_754[3], r_reg_754[3], r_reg_754[3], r_reg_754[3], r_reg_754[3], r_reg_754[3], r_reg_754 };
assign \add_18ns_18s_18_2_1_U4.din1  = { op_0[1], op_0[1], op_0[1], op_0[1], op_0[1], op_0[1], op_0[1], op_0[1], op_0[1], op_0[1], op_0[1], op_0[1], op_0[1], op_0[1], op_0[1], op_0[1], op_0 };
assign grp_fu_257_p2 = \add_18ns_18s_18_2_1_U4.dout ;
assign \add_18ns_18s_18_2_1_U4.reset  = ap_rst;
assign \add_18ns_18ns_18_2_1_U5.top_add_18ns_18ns_18_2_1_Adder_2_U.ain_s0  = \add_18ns_18ns_18_2_1_U5.top_add_18ns_18ns_18_2_1_Adder_2_U.a ;
assign \add_18ns_18ns_18_2_1_U5.top_add_18ns_18ns_18_2_1_Adder_2_U.bin_s0  = \add_18ns_18ns_18_2_1_U5.top_add_18ns_18ns_18_2_1_Adder_2_U.b ;
assign \add_18ns_18ns_18_2_1_U5.top_add_18ns_18ns_18_2_1_Adder_2_U.s  = { \add_18ns_18ns_18_2_1_U5.top_add_18ns_18ns_18_2_1_Adder_2_U.fas_s2 , \add_18ns_18ns_18_2_1_U5.top_add_18ns_18ns_18_2_1_Adder_2_U.sum_s1  };
assign \add_18ns_18ns_18_2_1_U5.top_add_18ns_18ns_18_2_1_Adder_2_U.u2.a  = \add_18ns_18ns_18_2_1_U5.top_add_18ns_18ns_18_2_1_Adder_2_U.ain_s1 ;
assign \add_18ns_18ns_18_2_1_U5.top_add_18ns_18ns_18_2_1_Adder_2_U.u2.b  = \add_18ns_18ns_18_2_1_U5.top_add_18ns_18ns_18_2_1_Adder_2_U.bin_s1 ;
assign \add_18ns_18ns_18_2_1_U5.top_add_18ns_18ns_18_2_1_Adder_2_U.u2.cin  = \add_18ns_18ns_18_2_1_U5.top_add_18ns_18ns_18_2_1_Adder_2_U.carry_s1 ;
assign \add_18ns_18ns_18_2_1_U5.top_add_18ns_18ns_18_2_1_Adder_2_U.facout_s2  = \add_18ns_18ns_18_2_1_U5.top_add_18ns_18ns_18_2_1_Adder_2_U.u2.cout ;
assign \add_18ns_18ns_18_2_1_U5.top_add_18ns_18ns_18_2_1_Adder_2_U.fas_s2  = \add_18ns_18ns_18_2_1_U5.top_add_18ns_18ns_18_2_1_Adder_2_U.u2.s ;
assign \add_18ns_18ns_18_2_1_U5.top_add_18ns_18ns_18_2_1_Adder_2_U.u1.a  = \add_18ns_18ns_18_2_1_U5.top_add_18ns_18ns_18_2_1_Adder_2_U.a [8:0];
assign \add_18ns_18ns_18_2_1_U5.top_add_18ns_18ns_18_2_1_Adder_2_U.u1.b  = \add_18ns_18ns_18_2_1_U5.top_add_18ns_18ns_18_2_1_Adder_2_U.b [8:0];
assign \add_18ns_18ns_18_2_1_U5.top_add_18ns_18ns_18_2_1_Adder_2_U.u1.cin  = 1'h0;
assign \add_18ns_18ns_18_2_1_U5.top_add_18ns_18ns_18_2_1_Adder_2_U.facout_s1  = \add_18ns_18ns_18_2_1_U5.top_add_18ns_18ns_18_2_1_Adder_2_U.u1.cout ;
assign \add_18ns_18ns_18_2_1_U5.top_add_18ns_18ns_18_2_1_Adder_2_U.fas_s1  = \add_18ns_18ns_18_2_1_U5.top_add_18ns_18ns_18_2_1_Adder_2_U.u1.s ;
assign \add_18ns_18ns_18_2_1_U5.top_add_18ns_18ns_18_2_1_Adder_2_U.a  = \add_18ns_18ns_18_2_1_U5.din0 ;
assign \add_18ns_18ns_18_2_1_U5.top_add_18ns_18ns_18_2_1_Adder_2_U.b  = \add_18ns_18ns_18_2_1_U5.din1 ;
assign \add_18ns_18ns_18_2_1_U5.top_add_18ns_18ns_18_2_1_Adder_2_U.ce  = \add_18ns_18ns_18_2_1_U5.ce ;
assign \add_18ns_18ns_18_2_1_U5.top_add_18ns_18ns_18_2_1_Adder_2_U.clk  = \add_18ns_18ns_18_2_1_U5.clk ;
assign \add_18ns_18ns_18_2_1_U5.top_add_18ns_18ns_18_2_1_Adder_2_U.reset  = \add_18ns_18ns_18_2_1_U5.reset ;
assign \add_18ns_18ns_18_2_1_U5.dout  = \add_18ns_18ns_18_2_1_U5.top_add_18ns_18ns_18_2_1_Adder_2_U.s ;
assign \add_18ns_18ns_18_2_1_U5.ce  = 1'h1;
assign \add_18ns_18ns_18_2_1_U5.clk  = ap_clk;
assign \add_18ns_18ns_18_2_1_U5.din0  = ret_V_reg_770;
assign \add_18ns_18ns_18_2_1_U5.din1  = select_ln1192_reg_775;
assign grp_fu_271_p2 = \add_18ns_18ns_18_2_1_U5.dout ;
assign \add_18ns_18ns_18_2_1_U5.reset  = ap_rst;
endmodule


// Machine B:
// Processed by function `add_clk_enable_signal` in `verilog_tricks.py`.
// Processed by function `remove_reset_signal` in `verilog_tricks.py`.
module top_B (
  ap_clk,
  ap_start,
  ap_done,
  ap_idle,
  ap_ready,
  op_0,
  op_1,
  op_4,
  op_6,
  op_8,
  op_9,
  op_10,
  op_12,
  op_13,
  op_14,
  op_15,
  op_17,
  op_18,
  op_19,
  op_31,
  op_31_ap_vld,
clk_enable
);
input clk_enable;


input ap_clk;
wire ap_rst;
assign ap_rst = op_31_ap_vld;
input ap_start;
input [1:0] op_0;
input [3:0] op_1;
input [3:0] op_10;
input [31:0] op_12;
input [7:0] op_13;
input [1:0] op_14;
input [3:0] op_15;
input op_17;
input op_18;
input [31:0] op_19;
input [31:0] op_4;
input [3:0] op_6;
input [7:0] op_8;
input op_9;
output ap_done;
output ap_idle;
output ap_ready;
output [31:0] op_31;
output op_31_ap_vld;


reg [31:0] add_ln691_1_reg_833;
reg [31:0] add_ln691_2_reg_854;
reg [31:0] add_ln691_3_reg_880;
reg [31:0] add_ln691_reg_812;
reg [1:0] add_ln69_2_reg_885;
reg [7:0] ap_CS_fsm = 8'h01;
reg icmp_ln768_reg_776;
reg icmp_ln786_reg_781;
reg icmp_ln851_1_reg_817;
reg icmp_ln851_2_reg_849;
reg icmp_ln851_3_reg_875;
reg icmp_ln851_reg_807;
reg [3:0] op_11_V_reg_791;
reg [31:0] op_26_V_reg_859;
reg p_Result_5_reg_764;
reg p_Result_6_reg_770;
reg [3:0] r_reg_753;
reg [31:0] ret_V_16_cast_reg_869;
reg [35:0] ret_V_1_reg_759;
reg [17:0] ret_V_2_reg_786;
reg [31:0] ret_V_3_cast_reg_827;
reg [21:0] ret_V_3_reg_796;
reg [35:0] ret_V_4_reg_822;
reg [46:0] ret_V_5_reg_838;
reg [31:0] ret_V_6_cast_reg_843;
reg [34:0] ret_V_8_reg_864;
reg [31:0] sext_ln831_reg_801;
wire [31:0] _000_;
wire [31:0] _001_;
wire [31:0] _002_;
wire [31:0] _003_;
wire [1:0] _004_;
wire [7:0] _005_;
wire _006_;
wire _007_;
wire _008_;
wire _009_;
wire _010_;
wire _011_;
wire [3:0] _012_;
wire [31:0] _013_;
wire _014_;
wire _015_;
wire [3:0] _016_;
wire [31:0] _017_;
wire [35:0] _018_;
wire [17:0] _019_;
wire [31:0] _020_;
wire [21:0] _021_;
wire [35:0] _022_;
wire [46:0] _023_;
wire [31:0] _024_;
wire [34:0] _025_;
wire [31:0] _026_;
wire [1:0] _027_;
wire _028_;
wire _029_;
wire _030_;
wire _031_;
wire _032_;
wire _033_;
wire _034_;
wire _035_;
wire _036_;
wire _037_;
wire _038_;
wire _039_;
wire _040_;
wire _041_;
wire _042_;
wire _043_;
wire _044_;
wire _045_;
wire [31:0] add_ln691_1_fu_513_p2;
wire [31:0] add_ln691_2_fu_580_p2;
wire [31:0] add_ln691_3_fu_680_p2;
wire [31:0] add_ln691_fu_447_p2;
wire [1:0] add_ln69_1_fu_706_p2;
wire [1:0] add_ln69_2_fu_712_p2;
wire [31:0] add_ln69_fu_737_p2;
wire ap_CS_fsm_state1;
wire ap_CS_fsm_state2;
wire ap_CS_fsm_state3;
wire ap_CS_fsm_state4;
wire ap_CS_fsm_state5;
wire ap_CS_fsm_state6;
wire ap_CS_fsm_state7;
wire ap_CS_fsm_state8;
wire [7:0] ap_NS_fsm;
wire ap_clk;
wire ap_done;
wire ap_idle;
wire ap_ready;
wire ap_rst;
wire ap_start;
wire [3:0] ashr_ln799_fu_233_p2;
wire icmp_ln768_fu_321_p2;
wire icmp_ln786_fu_327_p2;
wire icmp_ln851_1_fu_457_p2;
wire icmp_ln851_2_fu_574_p2;
wire icmp_ln851_3_fu_674_p2;
wire icmp_ln851_fu_441_p2;
wire [1:0] op_0;
wire [3:0] op_1;
wire [3:0] op_10;
wire [3:0] op_11_V_fu_394_p3;
wire [31:0] op_12;
wire [7:0] op_13;
wire [1:0] op_14;
wire [3:0] op_15;
wire op_16_V_fu_633_p2;
wire op_17;
wire op_18;
wire [31:0] op_19;
wire [31:0] op_26_V_fu_619_p2;
wire [31:0] op_31;
wire op_31_ap_vld;
wire [31:0] op_4;
wire [3:0] op_6;
wire [7:0] op_8;
wire op_9;
wire or_ln384_fu_388_p2;
wire or_ln785_fu_350_p2;
wire or_ln786_fu_370_p2;
wire overflow_fu_359_p2;
wire p_Result_1_fu_519_p3;
wire p_Result_2_fu_586_p3;
wire p_Result_3_fu_718_p3;
wire p_Result_4_fu_219_p3;
wire p_Result_s_fu_463_p3;
wire [3:0] p_Val2_1_fu_347_p1;
wire [3:0] r_fu_245_p3;
wire [31:0] ret_V_16_cast_fu_660_p4;
wire [35:0] ret_V_1_fu_289_p2;
wire [17:0] ret_V_2_fu_341_p2;
wire [31:0] ret_V_3_cast_fu_503_p4;
wire [21:0] ret_V_3_fu_417_p2;
wire [35:0] ret_V_4_fu_497_p2;
wire [46:0] ret_V_5_fu_554_p2;
wire [31:0] ret_V_6_cast_fu_560_p4;
wire [31:0] ret_V_6_fu_598_p3;
wire [31:0] ret_V_7_fu_609_p2;
wire [34:0] ret_V_8_fu_654_p2;
wire [31:0] ret_V_9_fu_730_p3;
wire [17:0] ret_V_fu_264_p2;
wire [6:0] rhs_1_fu_274_p3;
wire [34:0] rhs_3_fu_485_p3;
wire [45:0] rhs_4_fu_542_p3;
wire [33:0] rhs_7_fu_643_p3;
wire [17:0] select_ln1192_fu_333_p3;
wire [31:0] select_ln353_1_fu_535_p3;
wire [31:0] select_ln353_fu_478_p3;
wire [3:0] select_ln384_fu_380_p3;
wire [1:0] select_ln69_1_fu_694_p3;
wire [1:0] select_ln69_fu_686_p3;
wire [31:0] select_ln850_1_fu_530_p3;
wire [31:0] select_ln850_2_fu_593_p3;
wire [31:0] select_ln850_3_fu_725_p3;
wire [31:0] select_ln850_fu_473_p3;
wire [21:0] sext_ln1192_1_fu_413_p1;
wire [35:0] sext_ln1192_2_fu_493_p1;
wire [46:0] sext_ln1192_3_fu_550_p1;
wire [31:0] sext_ln1192_4_fu_605_p1;
wire [34:0] sext_ln1192_5_fu_650_p1;
wire [3:0] sext_ln1192_fu_402_p0;
wire [21:0] sext_ln1192_fu_402_p1;
wire [34:0] sext_ln1193_1_fu_281_p1;
wire [35:0] sext_ln1193_fu_270_p1;
wire [31:0] sext_ln69_fu_743_p1;
wire [15:0] sext_ln703_1_fu_257_p1;
wire [35:0] sext_ln703_2_fu_470_p1;
wire [31:0] sext_ln703_3_fu_526_p0;
wire [46:0] sext_ln703_3_fu_526_p1;
wire [3:0] sext_ln703_4_fu_639_p0;
wire [34:0] sext_ln703_4_fu_639_p1;
wire [17:0] sext_ln703_fu_253_p1;
wire [31:0] sext_ln831_fu_433_p1;
wire [3:0] sh_fu_227_p2;
wire [3:0] shl_ln781_fu_239_p2;
wire [31:0] tmp_2_fu_311_p4;
wire [20:0] tmp_5_fu_406_p3;
wire [18:0] tmp_fu_423_p4;
wire trunc_ln69_1_fu_629_p1;
wire trunc_ln69_fu_625_p1;
wire [2:0] trunc_ln851_1_fu_453_p1;
wire [31:0] trunc_ln851_2_fu_570_p0;
wire [13:0] trunc_ln851_2_fu_570_p1;
wire [3:0] trunc_ln851_3_fu_670_p0;
wire [1:0] trunc_ln851_3_fu_670_p1;
wire [3:0] trunc_ln851_fu_437_p0;
wire [2:0] trunc_ln851_fu_437_p1;
wire underflow_fu_375_p2;
wire xor_ln785_fu_354_p2;
wire xor_ln786_fu_365_p2;
wire [35:0] zext_ln1193_fu_285_p1;
wire [1:0] zext_ln69_1_fu_702_p1;
wire [31:0] zext_ln69_fu_615_p1;
wire [17:0] zext_ln703_fu_260_p1;


assign add_ln691_1_fu_513_p2 = ret_V_4_fu_497_p2[34:3] + 1'h1;
assign add_ln691_2_fu_580_p2 = ret_V_5_fu_554_p2[45:14] + 1'h1;
assign add_ln691_3_fu_680_p2 = ret_V_8_fu_654_p2[33:2] + 1'h1;
assign { add_ln691_fu_447_p2[31], add_ln691_fu_447_p2[18:0] } = $signed(ret_V_3_fu_417_p2[21:3]) + $signed(2'h1);
assign add_ln69_1_fu_706_p2 = select_ln69_fu_686_p3 + op_18;
assign add_ln69_2_fu_712_p2 = add_ln69_1_fu_706_p2 + select_ln69_1_fu_694_p3;
assign add_ln69_fu_737_p2 = ret_V_9_fu_730_p3 + op_19;
assign op_26_V_fu_619_p2 = ret_V_7_fu_609_p2 + op_14;
assign op_31 = $signed(add_ln69_2_reg_885) + $signed(add_ln69_fu_737_p2);
assign ret_V_2_fu_341_p2 = ret_V_fu_264_p2 + select_ln1192_fu_333_p3;
assign ret_V_3_fu_417_p2 = $signed({ ret_V_2_reg_786, 3'h0 }) + $signed(op_10);
assign ret_V_4_fu_497_p2 = $signed({ select_ln353_fu_478_p3, 3'h0 }) + $signed(op_11_V_reg_791);
assign ret_V_5_fu_554_p2 = $signed({ select_ln353_1_fu_535_p3, 14'h0000 }) + $signed(op_12);
assign ret_V_7_fu_609_p2 = $signed(ret_V_6_fu_598_p3) + $signed(op_13);
assign ret_V_8_fu_654_p2 = $signed({ op_26_V_reg_859, 2'h0 }) + $signed(op_15);
assign ret_V_fu_264_p2 = $signed({ 1'h0, r_reg_753[3], r_reg_753[3], r_reg_753[3], r_reg_753[3], r_reg_753[3], r_reg_753[3], r_reg_753[3], r_reg_753[3], r_reg_753[3], r_reg_753[3], r_reg_753[3], r_reg_753[3], r_reg_753 }) + $signed(op_0);
assign _028_ = icmp_ln851_1_reg_817 & ap_CS_fsm[3];
assign _029_ = ap_CS_fsm[0] & _031_;
assign _030_ = ap_CS_fsm[0] & ap_start;
assign op_16_V_fu_633_p2 = op_4[0] & op_8[0];
assign overflow_fu_359_p2 = xor_ln785_fu_354_p2 & or_ln785_fu_350_p2;
assign underflow_fu_375_p2 = p_Result_5_reg_764 & or_ln786_fu_370_p2;
assign xor_ln785_fu_354_p2 = ~ p_Result_5_reg_764;
assign xor_ln786_fu_365_p2 = ~ p_Result_6_reg_770;
assign _031_ = ~ ap_start;
assign _032_ = | ret_V_1_fu_289_p2[35:4];
assign _033_ = ret_V_1_fu_289_p2[35:4] != 32'd4294967295;
assign _034_ = | op_11_V_fu_394_p3[2:0];
assign _035_ = | op_12[13:0];
assign _036_ = | op_15[1:0];
assign _037_ = | op_10[2:0];
assign or_ln384_fu_388_p2 = underflow_fu_375_p2 | overflow_fu_359_p2;
assign or_ln785_fu_350_p2 = p_Result_6_reg_770 | icmp_ln768_reg_776;
assign or_ln786_fu_370_p2 = xor_ln786_fu_365_p2 | icmp_ln786_reg_781;
always @(posedge ap_clk)
ret_V_4_reg_822 <= _022_;
always @(posedge ap_clk)
ret_V_3_cast_reg_827 <= _020_;
always @(posedge ap_clk)
r_reg_753 <= _016_;
always @(posedge ap_clk)
op_26_V_reg_859 <= _013_;
always @(posedge ap_clk)
ret_V_1_reg_759 <= _018_;
always @(posedge ap_clk)
p_Result_5_reg_764 <= _014_;
always @(posedge ap_clk)
p_Result_6_reg_770 <= _015_;
always @(posedge ap_clk)
icmp_ln768_reg_776 <= _006_;
always @(posedge ap_clk)
icmp_ln786_reg_781 <= _007_;
always @(posedge ap_clk)
ret_V_2_reg_786 <= _019_;
always @(posedge ap_clk)
op_11_V_reg_791 <= _012_;
always @(posedge ap_clk)
ret_V_3_reg_796 <= _021_;
always @(posedge ap_clk)
sext_ln831_reg_801 <= _026_;
always @(posedge ap_clk)
icmp_ln851_reg_807 <= _011_;
always @(posedge ap_clk)
add_ln691_reg_812 <= _003_;
always @(posedge ap_clk)
icmp_ln851_1_reg_817 <= _008_;
always @(posedge ap_clk)
ret_V_8_reg_864 <= _025_;
always @(posedge ap_clk)
ret_V_16_cast_reg_869 <= _017_;
always @(posedge ap_clk)
icmp_ln851_3_reg_875 <= _010_;
always @(posedge ap_clk)
add_ln691_3_reg_880 <= _002_;
always @(posedge ap_clk)
add_ln69_2_reg_885 <= _004_;
always @(posedge ap_clk)
ret_V_5_reg_838 <= _023_;
always @(posedge ap_clk)
ret_V_6_cast_reg_843 <= _024_;
always @(posedge ap_clk)
icmp_ln851_2_reg_849 <= _009_;
always @(posedge ap_clk)
add_ln691_2_reg_854 <= _001_;
always @(posedge ap_clk)
add_ln691_1_reg_833 <= _000_;
always @(posedge ap_clk)
ap_CS_fsm <= _005_;
assign _027_ = _030_ ? 2'h2 : 2'h1;
assign _038_ = ap_CS_fsm == 1'h1;
function [7:0] _109_;
input [7:0] a;
input [63:0] b;
input [7:0] s;
case (s)
8'b00000001:
_109_ = b[7:0];
8'b00000010:
_109_ = b[15:8];
8'b00000100:
_109_ = b[23:16];
8'b00001000:
_109_ = b[31:24];
8'b00010000:
_109_ = b[39:32];
8'b00100000:
_109_ = b[47:40];
8'b01000000:
_109_ = b[55:48];
8'b10000000:
_109_ = b[63:56];
8'b00000000:
_109_ = a;
default:
_109_ = 8'bx;
endcase
endfunction
assign ap_NS_fsm = _109_(8'hxx, { 6'h00, _027_, 56'h04081020408001 }, { _038_, _045_, _044_, _043_, _042_, _041_, _040_, _039_ });
assign _039_ = ap_CS_fsm == 8'h80;
assign _040_ = ap_CS_fsm == 7'h40;
assign _041_ = ap_CS_fsm == 6'h20;
assign _042_ = ap_CS_fsm == 5'h10;
assign _043_ = ap_CS_fsm == 4'h8;
assign _044_ = ap_CS_fsm == 3'h4;
assign _045_ = ap_CS_fsm == 2'h2;
assign op_31_ap_vld = ap_CS_fsm[7] ? 1'h1 : 1'h0;
assign ap_idle = _029_ ? 1'h1 : 1'h0;
assign _020_ = ap_CS_fsm[3] ? ret_V_4_fu_497_p2[34:3] : ret_V_3_cast_reg_827;
assign _022_ = ap_CS_fsm[3] ? ret_V_4_fu_497_p2 : ret_V_4_reg_822;
assign _016_ = ap_CS_fsm[0] ? r_fu_245_p3 : r_reg_753;
assign _013_ = ap_CS_fsm[5] ? op_26_V_fu_619_p2 : op_26_V_reg_859;
assign _019_ = ap_CS_fsm[1] ? ret_V_2_fu_341_p2 : ret_V_2_reg_786;
assign _007_ = ap_CS_fsm[1] ? icmp_ln786_fu_327_p2 : icmp_ln786_reg_781;
assign _006_ = ap_CS_fsm[1] ? icmp_ln768_fu_321_p2 : icmp_ln768_reg_776;
assign _015_ = ap_CS_fsm[1] ? ret_V_1_fu_289_p2[3] : p_Result_6_reg_770;
assign _014_ = ap_CS_fsm[1] ? ret_V_1_fu_289_p2[35] : p_Result_5_reg_764;
assign _018_ = ap_CS_fsm[1] ? ret_V_1_fu_289_p2 : ret_V_1_reg_759;
assign _008_ = ap_CS_fsm[2] ? icmp_ln851_1_fu_457_p2 : icmp_ln851_1_reg_817;
assign _003_ = ap_CS_fsm[2] ? { add_ln691_fu_447_p2[31], add_ln691_fu_447_p2[31], add_ln691_fu_447_p2[31], add_ln691_fu_447_p2[31], add_ln691_fu_447_p2[31], add_ln691_fu_447_p2[31], add_ln691_fu_447_p2[31], add_ln691_fu_447_p2[31], add_ln691_fu_447_p2[31], add_ln691_fu_447_p2[31], add_ln691_fu_447_p2[31], add_ln691_fu_447_p2[31], add_ln691_fu_447_p2[31], add_ln691_fu_447_p2[18:0] } : add_ln691_reg_812;
assign _011_ = ap_CS_fsm[2] ? icmp_ln851_fu_441_p2 : icmp_ln851_reg_807;
assign _026_ = ap_CS_fsm[2] ? { ret_V_3_fu_417_p2[21], ret_V_3_fu_417_p2[21], ret_V_3_fu_417_p2[21], ret_V_3_fu_417_p2[21], ret_V_3_fu_417_p2[21], ret_V_3_fu_417_p2[21], ret_V_3_fu_417_p2[21], ret_V_3_fu_417_p2[21], ret_V_3_fu_417_p2[21], ret_V_3_fu_417_p2[21], ret_V_3_fu_417_p2[21], ret_V_3_fu_417_p2[21], ret_V_3_fu_417_p2[21], ret_V_3_fu_417_p2[21:3] } : sext_ln831_reg_801;
assign _021_ = ap_CS_fsm[2] ? ret_V_3_fu_417_p2 : ret_V_3_reg_796;
assign _012_ = ap_CS_fsm[2] ? op_11_V_fu_394_p3 : op_11_V_reg_791;
assign _004_ = ap_CS_fsm[6] ? add_ln69_2_fu_712_p2 : add_ln69_2_reg_885;
assign _002_ = ap_CS_fsm[6] ? add_ln691_3_fu_680_p2 : add_ln691_3_reg_880;
assign _010_ = ap_CS_fsm[6] ? icmp_ln851_3_fu_674_p2 : icmp_ln851_3_reg_875;
assign _017_ = ap_CS_fsm[6] ? ret_V_8_fu_654_p2[33:2] : ret_V_16_cast_reg_869;
assign _025_ = ap_CS_fsm[6] ? ret_V_8_fu_654_p2 : ret_V_8_reg_864;
assign _001_ = ap_CS_fsm[4] ? add_ln691_2_fu_580_p2 : add_ln691_2_reg_854;
assign _009_ = ap_CS_fsm[4] ? icmp_ln851_2_fu_574_p2 : icmp_ln851_2_reg_849;
assign _024_ = ap_CS_fsm[4] ? ret_V_5_fu_554_p2[45:14] : ret_V_6_cast_reg_843;
assign _023_ = ap_CS_fsm[4] ? ret_V_5_fu_554_p2 : ret_V_5_reg_838;
assign _000_ = _028_ ? add_ln691_1_fu_513_p2 : add_ln691_1_reg_833;
assign _005_ = ap_rst ? 8'h01 : ap_NS_fsm;
assign shl_ln781_fu_239_p2 = op_1 << op_1;
assign ashr_ln799_fu_233_p2 = $signed(op_1) >>> sh_fu_227_p2;
assign ret_V_1_fu_289_p2 = $signed(op_6) - $signed({ 1'h0, r_reg_753[3], r_reg_753[3], r_reg_753[3], r_reg_753[3], r_reg_753[3], r_reg_753[3], r_reg_753[3], r_reg_753[3], r_reg_753[3], r_reg_753[3], r_reg_753[3], r_reg_753[3], r_reg_753[3], r_reg_753[3], r_reg_753[3], r_reg_753[3], r_reg_753[3], r_reg_753[3], r_reg_753[3], r_reg_753[3], r_reg_753[3], r_reg_753[3], r_reg_753[3], r_reg_753[3], r_reg_753[3], r_reg_753[3], r_reg_753[3], r_reg_753[3], r_reg_753, 3'h0 });
assign sh_fu_227_p2 = 1'h0 - op_1;
assign icmp_ln768_fu_321_p2 = _032_ ? 1'h1 : 1'h0;
assign icmp_ln786_fu_327_p2 = _033_ ? 1'h1 : 1'h0;
assign icmp_ln851_1_fu_457_p2 = _034_ ? 1'h1 : 1'h0;
assign icmp_ln851_2_fu_574_p2 = _035_ ? 1'h1 : 1'h0;
assign icmp_ln851_3_fu_674_p2 = _036_ ? 1'h1 : 1'h0;
assign icmp_ln851_fu_441_p2 = _037_ ? 1'h1 : 1'h0;
assign op_11_V_fu_394_p3 = or_ln384_fu_388_p2 ? select_ln384_fu_380_p3 : ret_V_1_reg_759[3:0];
assign r_fu_245_p3 = op_1[3] ? ashr_ln799_fu_233_p2 : shl_ln781_fu_239_p2;
assign ret_V_6_fu_598_p3 = ret_V_5_reg_838[46] ? select_ln850_2_fu_593_p3 : ret_V_6_cast_reg_843;
assign ret_V_9_fu_730_p3 = ret_V_8_reg_864[34] ? select_ln850_3_fu_725_p3 : ret_V_16_cast_reg_869;
assign select_ln1192_fu_333_p3 = op_9 ? 18'h3ffff : 18'h00000;
assign select_ln353_1_fu_535_p3 = ret_V_4_reg_822[35] ? select_ln850_1_fu_530_p3 : ret_V_3_cast_reg_827;
assign select_ln353_fu_478_p3 = ret_V_3_reg_796[21] ? select_ln850_fu_473_p3 : sext_ln831_reg_801;
assign select_ln384_fu_380_p3 = overflow_fu_359_p2 ? 4'h7 : 4'h8;
assign select_ln69_1_fu_694_p3 = op_17 ? 2'h3 : 2'h0;
assign select_ln69_fu_686_p3 = op_16_V_fu_633_p2 ? 2'h3 : 2'h0;
assign select_ln850_1_fu_530_p3 = icmp_ln851_1_reg_817 ? add_ln691_1_reg_833 : ret_V_3_cast_reg_827;
assign select_ln850_2_fu_593_p3 = icmp_ln851_2_reg_849 ? add_ln691_2_reg_854 : ret_V_6_cast_reg_843;
assign select_ln850_3_fu_725_p3 = icmp_ln851_3_reg_875 ? add_ln691_3_reg_880 : ret_V_16_cast_reg_869;
assign select_ln850_fu_473_p3 = icmp_ln851_reg_807 ? add_ln691_reg_812 : sext_ln831_reg_801;
assign add_ln691_fu_447_p2[30:19] = { add_ln691_fu_447_p2[31], add_ln691_fu_447_p2[31], add_ln691_fu_447_p2[31], add_ln691_fu_447_p2[31], add_ln691_fu_447_p2[31], add_ln691_fu_447_p2[31], add_ln691_fu_447_p2[31], add_ln691_fu_447_p2[31], add_ln691_fu_447_p2[31], add_ln691_fu_447_p2[31], add_ln691_fu_447_p2[31], add_ln691_fu_447_p2[31] };
assign ap_CS_fsm_state1 = ap_CS_fsm[0];
assign ap_CS_fsm_state2 = ap_CS_fsm[1];
assign ap_CS_fsm_state3 = ap_CS_fsm[2];
assign ap_CS_fsm_state4 = ap_CS_fsm[3];
assign ap_CS_fsm_state5 = ap_CS_fsm[4];
assign ap_CS_fsm_state6 = ap_CS_fsm[5];
assign ap_CS_fsm_state7 = ap_CS_fsm[6];
assign ap_CS_fsm_state8 = ap_CS_fsm[7];
assign ap_done = op_31_ap_vld;
assign ap_ready = op_31_ap_vld;
assign p_Result_1_fu_519_p3 = ret_V_4_reg_822[35];
assign p_Result_2_fu_586_p3 = ret_V_5_reg_838[46];
assign p_Result_3_fu_718_p3 = ret_V_8_reg_864[34];
assign p_Result_4_fu_219_p3 = op_1[3];
assign p_Result_s_fu_463_p3 = ret_V_3_reg_796[21];
assign p_Val2_1_fu_347_p1 = ret_V_1_reg_759[3:0];
assign ret_V_16_cast_fu_660_p4 = ret_V_8_fu_654_p2[33:2];
assign ret_V_3_cast_fu_503_p4 = ret_V_4_fu_497_p2[34:3];
assign ret_V_6_cast_fu_560_p4 = ret_V_5_fu_554_p2[45:14];
assign rhs_1_fu_274_p3 = { r_reg_753, 3'h0 };
assign rhs_3_fu_485_p3 = { select_ln353_fu_478_p3, 3'h0 };
assign rhs_4_fu_542_p3 = { select_ln353_1_fu_535_p3, 14'h0000 };
assign rhs_7_fu_643_p3 = { op_26_V_reg_859, 2'h0 };
assign sext_ln1192_1_fu_413_p1 = { ret_V_2_reg_786[17], ret_V_2_reg_786, 3'h0 };
assign sext_ln1192_2_fu_493_p1 = { select_ln353_fu_478_p3[31], select_ln353_fu_478_p3, 3'h0 };
assign sext_ln1192_3_fu_550_p1 = { select_ln353_1_fu_535_p3[31], select_ln353_1_fu_535_p3, 14'h0000 };
assign sext_ln1192_4_fu_605_p1 = { op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13 };
assign sext_ln1192_5_fu_650_p1 = { op_26_V_reg_859[31], op_26_V_reg_859, 2'h0 };
assign sext_ln1192_fu_402_p0 = op_10;
assign sext_ln1192_fu_402_p1 = { op_10[3], op_10[3], op_10[3], op_10[3], op_10[3], op_10[3], op_10[3], op_10[3], op_10[3], op_10[3], op_10[3], op_10[3], op_10[3], op_10[3], op_10[3], op_10[3], op_10[3], op_10[3], op_10 };
assign sext_ln1193_1_fu_281_p1 = { r_reg_753[3], r_reg_753[3], r_reg_753[3], r_reg_753[3], r_reg_753[3], r_reg_753[3], r_reg_753[3], r_reg_753[3], r_reg_753[3], r_reg_753[3], r_reg_753[3], r_reg_753[3], r_reg_753[3], r_reg_753[3], r_reg_753[3], r_reg_753[3], r_reg_753[3], r_reg_753[3], r_reg_753[3], r_reg_753[3], r_reg_753[3], r_reg_753[3], r_reg_753[3], r_reg_753[3], r_reg_753[3], r_reg_753[3], r_reg_753[3], r_reg_753[3], r_reg_753, 3'h0 };
assign sext_ln1193_fu_270_p1 = { op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6 };
assign sext_ln69_fu_743_p1 = { add_ln69_2_reg_885[1], add_ln69_2_reg_885[1], add_ln69_2_reg_885[1], add_ln69_2_reg_885[1], add_ln69_2_reg_885[1], add_ln69_2_reg_885[1], add_ln69_2_reg_885[1], add_ln69_2_reg_885[1], add_ln69_2_reg_885[1], add_ln69_2_reg_885[1], add_ln69_2_reg_885[1], add_ln69_2_reg_885[1], add_ln69_2_reg_885[1], add_ln69_2_reg_885[1], add_ln69_2_reg_885[1], add_ln69_2_reg_885[1], add_ln69_2_reg_885[1], add_ln69_2_reg_885[1], add_ln69_2_reg_885[1], add_ln69_2_reg_885[1], add_ln69_2_reg_885[1], add_ln69_2_reg_885[1], add_ln69_2_reg_885[1], add_ln69_2_reg_885[1], add_ln69_2_reg_885[1], add_ln69_2_reg_885[1], add_ln69_2_reg_885[1], add_ln69_2_reg_885[1], add_ln69_2_reg_885[1], add_ln69_2_reg_885[1], add_ln69_2_reg_885 };
assign sext_ln703_1_fu_257_p1 = { r_reg_753[3], r_reg_753[3], r_reg_753[3], r_reg_753[3], r_reg_753[3], r_reg_753[3], r_reg_753[3], r_reg_753[3], r_reg_753[3], r_reg_753[3], r_reg_753[3], r_reg_753[3], r_reg_753 };
assign sext_ln703_2_fu_470_p1 = { op_11_V_reg_791[3], op_11_V_reg_791[3], op_11_V_reg_791[3], op_11_V_reg_791[3], op_11_V_reg_791[3], op_11_V_reg_791[3], op_11_V_reg_791[3], op_11_V_reg_791[3], op_11_V_reg_791[3], op_11_V_reg_791[3], op_11_V_reg_791[3], op_11_V_reg_791[3], op_11_V_reg_791[3], op_11_V_reg_791[3], op_11_V_reg_791[3], op_11_V_reg_791[3], op_11_V_reg_791[3], op_11_V_reg_791[3], op_11_V_reg_791[3], op_11_V_reg_791[3], op_11_V_reg_791[3], op_11_V_reg_791[3], op_11_V_reg_791[3], op_11_V_reg_791[3], op_11_V_reg_791[3], op_11_V_reg_791[3], op_11_V_reg_791[3], op_11_V_reg_791[3], op_11_V_reg_791[3], op_11_V_reg_791[3], op_11_V_reg_791[3], op_11_V_reg_791[3], op_11_V_reg_791 };
assign sext_ln703_3_fu_526_p0 = op_12;
assign sext_ln703_3_fu_526_p1 = { op_12[31], op_12[31], op_12[31], op_12[31], op_12[31], op_12[31], op_12[31], op_12[31], op_12[31], op_12[31], op_12[31], op_12[31], op_12[31], op_12[31], op_12[31], op_12 };
assign sext_ln703_4_fu_639_p0 = op_15;
assign sext_ln703_4_fu_639_p1 = { op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15 };
assign sext_ln703_fu_253_p1 = { op_0[1], op_0[1], op_0[1], op_0[1], op_0[1], op_0[1], op_0[1], op_0[1], op_0[1], op_0[1], op_0[1], op_0[1], op_0[1], op_0[1], op_0[1], op_0[1], op_0 };
assign sext_ln831_fu_433_p1 = { ret_V_3_fu_417_p2[21], ret_V_3_fu_417_p2[21], ret_V_3_fu_417_p2[21], ret_V_3_fu_417_p2[21], ret_V_3_fu_417_p2[21], ret_V_3_fu_417_p2[21], ret_V_3_fu_417_p2[21], ret_V_3_fu_417_p2[21], ret_V_3_fu_417_p2[21], ret_V_3_fu_417_p2[21], ret_V_3_fu_417_p2[21], ret_V_3_fu_417_p2[21], ret_V_3_fu_417_p2[21], ret_V_3_fu_417_p2[21:3] };
assign tmp_2_fu_311_p4 = ret_V_1_fu_289_p2[35:4];
assign tmp_5_fu_406_p3 = { ret_V_2_reg_786, 3'h0 };
assign tmp_fu_423_p4 = ret_V_3_fu_417_p2[21:3];
assign trunc_ln69_1_fu_629_p1 = op_8[0];
assign trunc_ln69_fu_625_p1 = op_4[0];
assign trunc_ln851_1_fu_453_p1 = op_11_V_fu_394_p3[2:0];
assign trunc_ln851_2_fu_570_p0 = op_12;
assign trunc_ln851_2_fu_570_p1 = op_12[13:0];
assign trunc_ln851_3_fu_670_p0 = op_15;
assign trunc_ln851_3_fu_670_p1 = op_15[1:0];
assign trunc_ln851_fu_437_p0 = op_10;
assign trunc_ln851_fu_437_p1 = op_10[2:0];
assign zext_ln1193_fu_285_p1 = { 1'h0, r_reg_753[3], r_reg_753[3], r_reg_753[3], r_reg_753[3], r_reg_753[3], r_reg_753[3], r_reg_753[3], r_reg_753[3], r_reg_753[3], r_reg_753[3], r_reg_753[3], r_reg_753[3], r_reg_753[3], r_reg_753[3], r_reg_753[3], r_reg_753[3], r_reg_753[3], r_reg_753[3], r_reg_753[3], r_reg_753[3], r_reg_753[3], r_reg_753[3], r_reg_753[3], r_reg_753[3], r_reg_753[3], r_reg_753[3], r_reg_753[3], r_reg_753[3], r_reg_753, 3'h0 };
assign zext_ln69_1_fu_702_p1 = { 1'h0, op_18 };
assign zext_ln69_fu_615_p1 = { 30'h00000000, op_14 };
assign zext_ln703_fu_260_p1 = { 2'h0, r_reg_753[3], r_reg_753[3], r_reg_753[3], r_reg_753[3], r_reg_753[3], r_reg_753[3], r_reg_753[3], r_reg_753[3], r_reg_753[3], r_reg_753[3], r_reg_753[3], r_reg_753[3], r_reg_753 };
endmodule


// Product machine:
module top_A_times_top_B (ap_start, op_0, op_1, op_10, op_12, op_13, op_14, op_15, op_17, op_18, op_19, op_4, op_6, op_8, op_9, ap_clk, unsafe_signal);
input ap_start;
input [1:0] op_0;
input [3:0] op_1;
input [3:0] op_10;
input [31:0] op_12;
input [7:0] op_13;
input [1:0] op_14;
input [3:0] op_15;
input op_17;
input op_18;
input [31:0] op_19;
input [31:0] op_4;
input [3:0] op_6;
input [7:0] op_8;
input op_9;
input ap_clk;
output unsafe_signal;
reg _setup;
initial _setup = 1'b0;
always @ (posedge ap_clk) _setup <= 1'b1;
reg ap_start_internal;
always @ (posedge ap_clk) if (!_setup) ap_start_internal <= ap_start;
reg [1:0] op_0_internal;
always @ (posedge ap_clk) if (!_setup) op_0_internal <= op_0;
reg [3:0] op_1_internal;
always @ (posedge ap_clk) if (!_setup) op_1_internal <= op_1;
reg [3:0] op_10_internal;
always @ (posedge ap_clk) if (!_setup) op_10_internal <= op_10;
reg [31:0] op_12_internal;
always @ (posedge ap_clk) if (!_setup) op_12_internal <= op_12;
reg [7:0] op_13_internal;
always @ (posedge ap_clk) if (!_setup) op_13_internal <= op_13;
reg [1:0] op_14_internal;
always @ (posedge ap_clk) if (!_setup) op_14_internal <= op_14;
reg [3:0] op_15_internal;
always @ (posedge ap_clk) if (!_setup) op_15_internal <= op_15;
reg op_17_internal;
always @ (posedge ap_clk) if (!_setup) op_17_internal <= op_17;
reg op_18_internal;
always @ (posedge ap_clk) if (!_setup) op_18_internal <= op_18;
reg [31:0] op_19_internal;
always @ (posedge ap_clk) if (!_setup) op_19_internal <= op_19;
reg [31:0] op_4_internal;
always @ (posedge ap_clk) if (!_setup) op_4_internal <= op_4;
reg [3:0] op_6_internal;
always @ (posedge ap_clk) if (!_setup) op_6_internal <= op_6;
reg [7:0] op_8_internal;
always @ (posedge ap_clk) if (!_setup) op_8_internal <= op_8;
reg op_9_internal;
always @ (posedge ap_clk) if (!_setup) op_9_internal <= op_9;
wire ap_done_A;
wire ap_done_B;
wire ap_done_eq;
assign ap_done_eq = ap_done_A == ap_done_B;
wire ap_idle_A;
wire ap_idle_B;
wire ap_idle_eq;
assign ap_idle_eq = ap_idle_A == ap_idle_B;
wire ap_ready_A;
wire ap_ready_B;
wire ap_ready_eq;
assign ap_ready_eq = ap_ready_A == ap_ready_B;
wire [31:0] op_31_A;
wire [31:0] op_31_B;
wire op_31_eq;
assign op_31_eq = op_31_A == op_31_B;
wire op_31_ap_vld_A;
wire op_31_ap_vld_B;
wire clk_enable_A;
wire clk_enable_B;
assign clk_enable_A = _setup & (~op_31_ap_vld_A | op_31_ap_vld_B);
assign clk_enable_B = _setup;
wire divergent;
assign divergent = ~(ap_done_eq & ap_idle_eq & ap_ready_eq & op_31_eq);
assign unsafe_signal = op_31_ap_vld_A & op_31_ap_vld_B & divergent;
top_A instance_A (
    .ap_clk(ap_clk),
    .clk_enable(clk_enable_A),
    .ap_start(ap_start_internal),
    .op_0(op_0_internal),
    .op_1(op_1_internal),
    .op_10(op_10_internal),
    .op_12(op_12_internal),
    .op_13(op_13_internal),
    .op_14(op_14_internal),
    .op_15(op_15_internal),
    .op_17(op_17_internal),
    .op_18(op_18_internal),
    .op_19(op_19_internal),
    .op_4(op_4_internal),
    .op_6(op_6_internal),
    .op_8(op_8_internal),
    .op_9(op_9_internal),
    .ap_done(ap_done_A),
    .ap_idle(ap_idle_A),
    .ap_ready(ap_ready_A),
    .op_31(op_31_A),
    .op_31_ap_vld(op_31_ap_vld_A)
);
top_B instance_B (
    .ap_clk(ap_clk),
    .clk_enable(clk_enable_B),
    .ap_start(ap_start_internal),
    .op_0(op_0_internal),
    .op_1(op_1_internal),
    .op_10(op_10_internal),
    .op_12(op_12_internal),
    .op_13(op_13_internal),
    .op_14(op_14_internal),
    .op_15(op_15_internal),
    .op_17(op_17_internal),
    .op_18(op_18_internal),
    .op_19(op_19_internal),
    .op_4(op_4_internal),
    .op_6(op_6_internal),
    .op_8(op_8_internal),
    .op_9(op_9_internal),
    .ap_done(ap_done_B),
    .ap_idle(ap_idle_B),
    .ap_ready(ap_ready_B),
    .op_31(op_31_B),
    .op_31_ap_vld(op_31_ap_vld_B)
);
endmodule
