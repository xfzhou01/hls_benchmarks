// Processed by function `construct_kairos` in `verilog_tricks.py`.
// Machine A:
// Processed by function `add_clk_enable_signal` in `verilog_tricks.py`.
// Processed by function `remove_reset_signal` in `verilog_tricks.py`.
module top_A (
  ap_clk,
  ap_start,
  ap_done,
  ap_idle,
  ap_ready,
  op_0,
  op_1,
  op_2,
  op_3,
  op_4,
  op_8,
  op_10,
  op_11,
  op_14,
  op_15,
  op_16,
  op_17,
  op_31,
  op_31_ap_vld,
clk_enable
);
input clk_enable;


input ap_clk;
wire ap_rst;
assign ap_rst = op_31_ap_vld;
input ap_start;
input [7:0] op_0;
input [15:0] op_1;
input [3:0] op_10;
input op_11;
input op_14;
input [7:0] op_15;
input [3:0] op_16;
input [1:0] op_17;
input op_2;
input [1:0] op_3;
input [1:0] op_4;
input [1:0] op_8;
output ap_done;
output ap_idle;
output ap_ready;
output [31:0] op_31;
output op_31_ap_vld;


reg [31:0] add_ln691_reg_803;
reg [2:0] add_ln69_4_reg_835;
reg [9:0] add_ln69_reg_751;
reg and_ln365_reg_776;
reg [10:0] ap_CS_fsm = 11'h001;
reg icmp_ln851_1_reg_798;
reg icmp_ln851_2_reg_825;
reg icmp_ln851_reg_736;
reg lhs_V_reg_756;
reg [1:0] op_19_V_reg_857;
reg [31:0] op_26_V_reg_808;
reg [31:0] op_30_V_reg_852;
reg or_ln785_reg_771;
reg overflow_reg_846;
reg p_Result_7_reg_766;
reg r_reg_761;
reg [16:0] ret_V_12_reg_724;
reg [10:0] ret_V_14_reg_746;
reg [10:0] ret_V_15_reg_781;
reg [31:0] ret_V_16_cast_reg_867;
reg [39:0] ret_V_16_reg_786;
reg [34:0] ret_V_18_reg_813;
reg [31:0] ret_V_19_reg_830;
reg [33:0] ret_V_20_reg_862;
reg [31:0] ret_V_6_cast_reg_791;
reg [31:0] ret_V_9_cast_reg_818;
reg [9:0] ret_V_reg_729;
wire [31:0] _000_;
wire [2:0] _001_;
wire [9:0] _002_;
wire _003_;
wire [10:0] _004_;
wire _005_;
wire _006_;
wire _007_;
wire _008_;
wire [1:0] _009_;
wire [31:0] _010_;
wire [31:0] _011_;
wire _012_;
wire _013_;
wire _014_;
wire _015_;
wire [16:0] _016_;
wire [10:0] _017_;
wire [10:0] _018_;
wire [31:0] _019_;
wire [39:0] _020_;
wire [34:0] _021_;
wire [31:0] _022_;
wire [33:0] _023_;
wire [31:0] _024_;
wire [31:0] _025_;
wire [9:0] _026_;
wire [1:0] _027_;
wire _028_;
wire _029_;
wire _030_;
wire _031_;
wire _032_;
wire _033_;
wire _034_;
wire _035_;
wire _036_;
wire _037_;
wire _038_;
wire _039_;
wire _040_;
wire _041_;
wire _042_;
wire _043_;
wire _044_;
wire _045_;
wire [31:0] add_ln691_1_fu_558_p2;
wire [31:0] add_ln691_2_fu_704_p2;
wire [31:0] add_ln691_fu_472_p2;
wire [31:0] add_ln69_3_fu_623_p2;
wire [2:0] add_ln69_4_fu_587_p2;
wire [9:0] add_ln69_fu_310_p2;
wire and_ln365_fu_372_p2;
wire ap_CS_fsm_state1;
wire ap_CS_fsm_state10;
wire ap_CS_fsm_state11;
wire ap_CS_fsm_state2;
wire ap_CS_fsm_state3;
wire ap_CS_fsm_state4;
wire ap_CS_fsm_state5;
wire ap_CS_fsm_state6;
wire ap_CS_fsm_state7;
wire ap_CS_fsm_state8;
wire ap_CS_fsm_state9;
wire [10:0] ap_NS_fsm;
wire ap_clk;
wire ap_done;
wire ap_idle;
wire ap_ready;
wire ap_rst;
wire ap_start;
wire empty_fu_322_p1;
wire icmp_ln785_fu_601_p2;
wire icmp_ln851_1_fu_466_p2;
wire icmp_ln851_2_fu_545_p2;
wire icmp_ln851_fu_241_p2;
wire lhs_V_fu_316_p2;
wire [14:0] lhs_fu_205_p3;
wire [7:0] op_0;
wire [15:0] op_1;
wire [3:0] op_10;
wire op_11;
wire [7:0] op_13_V_fu_424_p3;
wire op_14;
wire [7:0] op_15;
wire [3:0] op_16;
wire [1:0] op_17;
wire [1:0] op_19_V_fu_655_p3;
wire op_2;
wire [10:0] op_23_V_fu_381_p2;
wire [31:0] op_26_V_fu_504_p2;
wire [1:0] op_3;
wire [31:0] op_30_V_fu_631_p2;
wire [31:0] op_31;
wire op_31_ap_vld;
wire [1:0] op_4;
wire [1:0] op_8;
wire or_ln384_fu_651_p1;
wire or_ln384_fu_651_p2;
wire or_ln785_1_fu_593_p1;
wire [1:0] or_ln785_1_fu_593_p3;
wire or_ln785_fu_346_p2;
wire overflow_fu_613_p2;
wire [7:0] p_Result_3_fu_408_p4;
wire p_Result_4_fu_477_p3;
wire p_Result_5_fu_551_p3;
wire p_Result_6_fu_694_p3;
wire p_Result_7_fu_340_p2;
wire p_Result_s_fu_247_p3;
wire [7:0] p_Val2_1_fu_395_p3;
wire [6:0] p_Val2_3_fu_402_p2;
wire p_Val2_5_fu_637_p0;
wire [1:0] p_Val2_5_fu_637_p3;
wire r_fu_326_p2;
wire [16:0] ret_V_12_fu_221_p2;
wire [9:0] ret_V_13_fu_265_p3;
wire [10:0] ret_V_14_fu_292_p2;
wire [10:0] ret_V_15_fu_389_p2;
wire [39:0] ret_V_16_fu_446_p2;
wire [31:0] ret_V_17_fu_489_p3;
wire [34:0] ret_V_18_fu_525_p2;
wire [31:0] ret_V_19_fu_569_p3;
wire [33:0] ret_V_20_fu_678_p2;
wire [9:0] ret_V_2_fu_254_p2;
wire [1:0] ret_fu_272_p3;
wire [33:0] rhs_4_fu_514_p3;
wire [32:0] rhs_6_fu_667_p3;
wire [10:0] select_ln1192_fu_280_p3;
wire [1:0] select_ln384_fu_644_p3;
wire [2:0] select_ln69_1_fu_580_p3;
wire [31:0] select_ln69_fu_496_p3;
wire [7:0] select_ln785_fu_417_p3;
wire [31:0] select_ln850_1_fu_484_p3;
wire [31:0] select_ln850_2_fu_563_p3;
wire [31:0] select_ln850_3_fu_709_p3;
wire [9:0] select_ln850_fu_259_p3;
wire [10:0] sext_ln1192_1_fu_288_p1;
wire [39:0] sext_ln1192_2_fu_442_p1;
wire [34:0] sext_ln1192_3_fu_521_p1;
wire [33:0] sext_ln1192_4_fu_674_p1;
wire [16:0] sext_ln1192_fu_213_p1;
wire [31:0] sext_ln69_2_fu_619_p1;
wire [9:0] sext_ln69_3_fu_306_p1;
wire [10:0] sext_ln69_4_fu_378_p1;
wire [2:0] sext_ln69_5_fu_576_p1;
wire [31:0] sext_ln69_6_fu_628_p1;
wire [7:0] sext_ln69_fu_298_p1;
wire [39:0] sext_ln703_1_fu_431_p1;
wire [7:0] sext_ln703_2_fu_510_p0;
wire [34:0] sext_ln703_2_fu_510_p1;
wire [33:0] sext_ln703_3_fu_663_p1;
wire [15:0] sext_ln703_fu_217_p0;
wire [16:0] sext_ln703_fu_217_p1;
wire tmp_1_fu_352_p3;
wire [17:0] tmp_3_fu_435_p3;
wire tmp_fu_332_p3;
wire [6:0] trunc_ln851_1_fu_462_p1;
wire [7:0] trunc_ln851_2_fu_541_p0;
wire [1:0] trunc_ln851_2_fu_541_p1;
wire trunc_ln851_3_fu_701_p1;
wire [15:0] trunc_ln851_fu_237_p0;
wire [6:0] trunc_ln851_fu_237_p1;
wire xor_ln365_1_fu_366_p2;
wire xor_ln365_fu_360_p2;
wire xor_ln785_fu_607_p0;
wire xor_ln785_fu_607_p2;
wire [10:0] zext_ln1192_fu_386_p1;
wire [9:0] zext_ln69_fu_302_p1;


assign add_ln691_1_fu_558_p2 = ret_V_9_cast_reg_818 + 1'h1;
assign add_ln691_2_fu_704_p2 = ret_V_16_cast_reg_867 + 1'h1;
assign add_ln691_fu_472_p2 = ret_V_6_cast_reg_791 + 1'h1;
assign add_ln69_3_fu_623_p2 = $signed(ret_V_19_reg_830) + $signed(op_16);
assign add_ln69_4_fu_587_p2 = $signed(op_17) + $signed(select_ln69_1_fu_580_p3);
assign add_ln69_fu_310_p2 = $signed({ 1'h0, ret_fu_272_p3[1], ret_fu_272_p3[1], ret_fu_272_p3[1], ret_fu_272_p3[1], ret_fu_272_p3[1], ret_fu_272_p3[1], ret_fu_272_p3 }) + $signed(op_10);
assign op_23_V_fu_381_p2 = $signed(add_ln69_reg_751) + $signed(ret_V_14_reg_746);
assign op_26_V_fu_504_p2 = ret_V_17_fu_489_p3 + select_ln69_fu_496_p3;
assign op_30_V_fu_631_p2 = $signed(add_ln69_4_reg_835) + $signed(add_ln69_3_fu_623_p2);
assign ret_V_12_fu_221_p2 = $signed({ op_0, 7'h00 }) + $signed(op_1);
assign ret_V_14_fu_292_p2 = $signed(ret_V_13_fu_265_p3) + $signed(select_ln1192_fu_280_p3);
assign ret_V_15_fu_389_p2 = lhs_V_reg_756 + op_23_V_fu_381_p2;
assign { ret_V_16_fu_446_p2[39], ret_V_16_fu_446_p2[17:0] } = $signed({ ret_V_15_reg_781, 7'h00 }) + $signed(op_13_V_fu_424_p3);
assign ret_V_18_fu_525_p2 = $signed({ op_26_V_reg_808, 2'h0 }) + $signed(op_15);
assign ret_V_20_fu_678_p2 = $signed({ op_30_V_reg_852, 1'h0 }) + $signed(op_19_V_fu_655_p3);
assign ret_V_2_fu_254_p2 = ret_V_reg_729 + 1'h1;
assign _028_ = icmp_ln851_1_reg_798 & ap_CS_fsm[4];
assign _029_ = ap_CS_fsm[0] & _031_;
assign _030_ = ap_CS_fsm[0] & ap_start;
assign and_ln365_fu_372_p2 = xor_ln365_1_fu_366_p2 & or_ln785_fu_346_p2;
assign overflow_fu_613_p2 = xor_ln785_fu_607_p2 & icmp_ln785_fu_601_p2;
assign p_Result_7_fu_340_p2 = ~ op_8[1];
assign r_fu_326_p2 = ~ op_8[0];
assign lhs_V_fu_316_p2 = ~ op_2;
assign xor_ln785_fu_607_p2 = ~ op_11;
assign _031_ = ~ ap_start;
assign _032_ = ! op_1[6:0];
assign _033_ = | op_13_V_fu_424_p3[6:0];
assign _034_ = | op_15[1:0];
assign or_ln384_fu_651_p2 = overflow_reg_846 | op_11;
assign or_ln785_fu_346_p2 = r_fu_326_p2 | p_Result_7_fu_340_p2;
always @(posedge ap_clk)
overflow_reg_846 <= _013_;
always @(posedge ap_clk)
op_30_V_reg_852 <= _011_;
always @(posedge ap_clk)
op_26_V_reg_808 <= _010_;
always @(posedge ap_clk)
op_19_V_reg_857 <= _009_;
always @(posedge ap_clk)
ret_V_20_reg_862 <= _023_;
always @(posedge ap_clk)
ret_V_16_cast_reg_867 <= _019_;
always @(posedge ap_clk)
ret_V_12_reg_724 <= _016_;
always @(posedge ap_clk)
ret_V_reg_729 <= _026_;
always @(posedge ap_clk)
icmp_ln851_reg_736 <= _007_;
always @(posedge ap_clk)
ret_V_18_reg_813 <= _021_;
always @(posedge ap_clk)
ret_V_9_cast_reg_818 <= _025_;
always @(posedge ap_clk)
icmp_ln851_2_reg_825 <= _006_;
always @(posedge ap_clk)
ret_V_16_reg_786 <= _020_;
always @(posedge ap_clk)
ret_V_6_cast_reg_791 <= _024_;
always @(posedge ap_clk)
icmp_ln851_1_reg_798 <= _005_;
always @(posedge ap_clk)
r_reg_761 <= _015_;
always @(posedge ap_clk)
p_Result_7_reg_766 <= _014_;
always @(posedge ap_clk)
or_ln785_reg_771 <= _012_;
always @(posedge ap_clk)
and_ln365_reg_776 <= _003_;
always @(posedge ap_clk)
ret_V_15_reg_781 <= _018_;
always @(posedge ap_clk)
ret_V_14_reg_746 <= _017_;
always @(posedge ap_clk)
add_ln69_reg_751 <= _002_;
always @(posedge ap_clk)
lhs_V_reg_756 <= _008_;
always @(posedge ap_clk)
ret_V_19_reg_830 <= _022_;
always @(posedge ap_clk)
add_ln69_4_reg_835 <= _001_;
always @(posedge ap_clk)
add_ln691_reg_803 <= _000_;
always @(posedge ap_clk)
ap_CS_fsm <= _004_;
assign _027_ = _030_ ? 2'h2 : 2'h1;
assign _035_ = ap_CS_fsm == 1'h1;
function [10:0] _106_;
input [10:0] a;
input [120:0] b;
input [10:0] s;
case (s)
11'b00000000001:
_106_ = b[10:0];
11'b00000000010:
_106_ = b[21:11];
11'b00000000100:
_106_ = b[32:22];
11'b00000001000:
_106_ = b[43:33];
11'b00000010000:
_106_ = b[54:44];
11'b00000100000:
_106_ = b[65:55];
11'b00001000000:
_106_ = b[76:66];
11'b00010000000:
_106_ = b[87:77];
11'b00100000000:
_106_ = b[98:88];
11'b01000000000:
_106_ = b[109:99];
11'b10000000000:
_106_ = b[120:110];
11'b00000000000:
_106_ = a;
default:
_106_ = 11'bx;
endcase
endfunction
assign ap_NS_fsm = _106_(11'hxxx, { 9'h000, _027_, 110'h0020080200802008020080200001 }, { _035_, _045_, _044_, _043_, _042_, _041_, _040_, _039_, _038_, _037_, _036_ });
assign _036_ = ap_CS_fsm == 11'h400;
assign _037_ = ap_CS_fsm == 10'h200;
assign _038_ = ap_CS_fsm == 9'h100;
assign _039_ = ap_CS_fsm == 8'h80;
assign _040_ = ap_CS_fsm == 7'h40;
assign _041_ = ap_CS_fsm == 6'h20;
assign _042_ = ap_CS_fsm == 5'h10;
assign _043_ = ap_CS_fsm == 4'h8;
assign _044_ = ap_CS_fsm == 3'h4;
assign _045_ = ap_CS_fsm == 2'h2;
assign op_31_ap_vld = ap_CS_fsm[10] ? 1'h1 : 1'h0;
assign ap_idle = _029_ ? 1'h1 : 1'h0;
assign _011_ = ap_CS_fsm[8] ? op_30_V_fu_631_p2 : op_30_V_reg_852;
assign _013_ = ap_CS_fsm[8] ? overflow_fu_613_p2 : overflow_reg_846;
assign _010_ = ap_CS_fsm[5] ? op_26_V_fu_504_p2 : op_26_V_reg_808;
assign _019_ = ap_CS_fsm[9] ? ret_V_20_fu_678_p2[32:1] : ret_V_16_cast_reg_867;
assign _023_ = ap_CS_fsm[9] ? ret_V_20_fu_678_p2 : ret_V_20_reg_862;
assign _009_ = ap_CS_fsm[9] ? op_19_V_fu_655_p3 : op_19_V_reg_857;
assign _007_ = ap_CS_fsm[0] ? icmp_ln851_fu_241_p2 : icmp_ln851_reg_736;
assign _026_ = ap_CS_fsm[0] ? ret_V_12_fu_221_p2[16:7] : ret_V_reg_729;
assign _016_ = ap_CS_fsm[0] ? ret_V_12_fu_221_p2 : ret_V_12_reg_724;
assign _006_ = ap_CS_fsm[6] ? icmp_ln851_2_fu_545_p2 : icmp_ln851_2_reg_825;
assign _025_ = ap_CS_fsm[6] ? ret_V_18_fu_525_p2[33:2] : ret_V_9_cast_reg_818;
assign _021_ = ap_CS_fsm[6] ? ret_V_18_fu_525_p2 : ret_V_18_reg_813;
assign _005_ = ap_CS_fsm[3] ? icmp_ln851_1_fu_466_p2 : icmp_ln851_1_reg_798;
assign _024_ = ap_CS_fsm[3] ? { ret_V_16_fu_446_p2[39], ret_V_16_fu_446_p2[39], ret_V_16_fu_446_p2[39], ret_V_16_fu_446_p2[39], ret_V_16_fu_446_p2[39], ret_V_16_fu_446_p2[39], ret_V_16_fu_446_p2[39], ret_V_16_fu_446_p2[39], ret_V_16_fu_446_p2[39], ret_V_16_fu_446_p2[39], ret_V_16_fu_446_p2[39], ret_V_16_fu_446_p2[39], ret_V_16_fu_446_p2[39], ret_V_16_fu_446_p2[39], ret_V_16_fu_446_p2[39], ret_V_16_fu_446_p2[39], ret_V_16_fu_446_p2[39], ret_V_16_fu_446_p2[39], ret_V_16_fu_446_p2[39], ret_V_16_fu_446_p2[39], ret_V_16_fu_446_p2[39], ret_V_16_fu_446_p2[17:7] } : ret_V_6_cast_reg_791;
assign _020_ = ap_CS_fsm[3] ? { ret_V_16_fu_446_p2[39], ret_V_16_fu_446_p2[39], ret_V_16_fu_446_p2[39], ret_V_16_fu_446_p2[39], ret_V_16_fu_446_p2[39], ret_V_16_fu_446_p2[39], ret_V_16_fu_446_p2[39], ret_V_16_fu_446_p2[39], ret_V_16_fu_446_p2[39], ret_V_16_fu_446_p2[39], ret_V_16_fu_446_p2[39], ret_V_16_fu_446_p2[39], ret_V_16_fu_446_p2[39], ret_V_16_fu_446_p2[39], ret_V_16_fu_446_p2[39], ret_V_16_fu_446_p2[39], ret_V_16_fu_446_p2[39], ret_V_16_fu_446_p2[39], ret_V_16_fu_446_p2[39], ret_V_16_fu_446_p2[39], ret_V_16_fu_446_p2[39], ret_V_16_fu_446_p2[39], ret_V_16_fu_446_p2[17:0] } : ret_V_16_reg_786;
assign _018_ = ap_CS_fsm[2] ? ret_V_15_fu_389_p2 : ret_V_15_reg_781;
assign _003_ = ap_CS_fsm[2] ? and_ln365_fu_372_p2 : and_ln365_reg_776;
assign _012_ = ap_CS_fsm[2] ? or_ln785_fu_346_p2 : or_ln785_reg_771;
assign _014_ = ap_CS_fsm[2] ? p_Result_7_fu_340_p2 : p_Result_7_reg_766;
assign _015_ = ap_CS_fsm[2] ? r_fu_326_p2 : r_reg_761;
assign _008_ = ap_CS_fsm[1] ? lhs_V_fu_316_p2 : lhs_V_reg_756;
assign _002_ = ap_CS_fsm[1] ? add_ln69_fu_310_p2 : add_ln69_reg_751;
assign _017_ = ap_CS_fsm[1] ? ret_V_14_fu_292_p2 : ret_V_14_reg_746;
assign _001_ = ap_CS_fsm[7] ? add_ln69_4_fu_587_p2 : add_ln69_4_reg_835;
assign _022_ = ap_CS_fsm[7] ? ret_V_19_fu_569_p3 : ret_V_19_reg_830;
assign _000_ = _028_ ? add_ln691_fu_472_p2 : add_ln691_reg_803;
assign _004_ = ap_rst ? 11'h001 : ap_NS_fsm;
assign icmp_ln785_fu_601_p2 = op_11 ? 1'h1 : 1'h0;
assign icmp_ln851_1_fu_466_p2 = _033_ ? 1'h1 : 1'h0;
assign icmp_ln851_2_fu_545_p2 = _034_ ? 1'h1 : 1'h0;
assign icmp_ln851_fu_241_p2 = _032_ ? 1'h1 : 1'h0;
assign op_13_V_fu_424_p3 = and_ln365_reg_776 ? { r_reg_761, 7'h00 } : select_ln785_fu_417_p3;
assign op_19_V_fu_655_p3 = or_ln384_fu_651_p2 ? select_ln384_fu_644_p3 : p_Val2_5_fu_637_p3;
assign op_31 = ret_V_20_reg_862[33] ? select_ln850_3_fu_709_p3 : ret_V_16_cast_reg_867;
assign p_Val2_5_fu_637_p3 = op_11 ? 2'h2 : 2'h0;
assign ret_V_13_fu_265_p3 = ret_V_12_reg_724[16] ? select_ln850_fu_259_p3 : ret_V_reg_729;
assign ret_V_17_fu_489_p3 = ret_V_16_reg_786[39] ? select_ln850_1_fu_484_p3 : ret_V_6_cast_reg_791;
assign ret_V_19_fu_569_p3 = ret_V_18_reg_813[34] ? select_ln850_2_fu_563_p3 : ret_V_9_cast_reg_818;
assign ret_fu_272_p3 = op_2 ? 2'h3 : op_4;
assign select_ln1192_fu_280_p3 = op_2 ? 11'h7ff : 11'h000;
assign select_ln384_fu_644_p3 = overflow_reg_846 ? 2'h1 : 2'h3;
assign select_ln69_1_fu_580_p3 = op_2 ? 3'h7 : 3'h0;
assign select_ln69_fu_496_p3 = op_14 ? 32'd4294967295 : 32'd0;
assign select_ln785_fu_417_p3 = or_ln785_reg_771 ? { p_Result_7_reg_766, 7'h7f } : 8'h00;
assign select_ln850_1_fu_484_p3 = icmp_ln851_1_reg_798 ? add_ln691_reg_803 : ret_V_6_cast_reg_791;
assign select_ln850_2_fu_563_p3 = icmp_ln851_2_reg_825 ? add_ln691_1_fu_558_p2 : ret_V_9_cast_reg_818;
assign select_ln850_3_fu_709_p3 = op_19_V_reg_857[0] ? add_ln691_2_fu_704_p2 : ret_V_16_cast_reg_867;
assign select_ln850_fu_259_p3 = icmp_ln851_reg_736 ? ret_V_reg_729 : ret_V_2_fu_254_p2;
assign xor_ln365_1_fu_366_p2 = p_Result_7_fu_340_p2 ^ op_8[0];
assign ap_CS_fsm_state1 = ap_CS_fsm[0];
assign ap_CS_fsm_state10 = ap_CS_fsm[9];
assign ap_CS_fsm_state11 = ap_CS_fsm[10];
assign ap_CS_fsm_state2 = ap_CS_fsm[1];
assign ap_CS_fsm_state3 = ap_CS_fsm[2];
assign ap_CS_fsm_state4 = ap_CS_fsm[3];
assign ap_CS_fsm_state5 = ap_CS_fsm[4];
assign ap_CS_fsm_state6 = ap_CS_fsm[5];
assign ap_CS_fsm_state7 = ap_CS_fsm[6];
assign ap_CS_fsm_state8 = ap_CS_fsm[7];
assign ap_CS_fsm_state9 = ap_CS_fsm[8];
assign ap_done = op_31_ap_vld;
assign ap_ready = op_31_ap_vld;
assign empty_fu_322_p1 = op_8[0];
assign lhs_fu_205_p3 = { op_0, 7'h00 };
assign or_ln384_fu_651_p1 = op_11;
assign or_ln785_1_fu_593_p1 = op_11;
assign or_ln785_1_fu_593_p3 = { op_11, 1'h0 };
assign p_Result_3_fu_408_p4 = { p_Result_7_reg_766, 7'h7f };
assign p_Result_4_fu_477_p3 = ret_V_16_reg_786[39];
assign p_Result_5_fu_551_p3 = ret_V_18_reg_813[34];
assign p_Result_6_fu_694_p3 = ret_V_20_reg_862[33];
assign p_Result_s_fu_247_p3 = ret_V_12_reg_724[16];
assign p_Val2_1_fu_395_p3 = { r_reg_761, 7'h00 };
assign p_Val2_3_fu_402_p2 = 7'h7f;
assign p_Val2_5_fu_637_p0 = op_11;
assign ret_V_16_fu_446_p2[38:18] = { ret_V_16_fu_446_p2[39], ret_V_16_fu_446_p2[39], ret_V_16_fu_446_p2[39], ret_V_16_fu_446_p2[39], ret_V_16_fu_446_p2[39], ret_V_16_fu_446_p2[39], ret_V_16_fu_446_p2[39], ret_V_16_fu_446_p2[39], ret_V_16_fu_446_p2[39], ret_V_16_fu_446_p2[39], ret_V_16_fu_446_p2[39], ret_V_16_fu_446_p2[39], ret_V_16_fu_446_p2[39], ret_V_16_fu_446_p2[39], ret_V_16_fu_446_p2[39], ret_V_16_fu_446_p2[39], ret_V_16_fu_446_p2[39], ret_V_16_fu_446_p2[39], ret_V_16_fu_446_p2[39], ret_V_16_fu_446_p2[39], ret_V_16_fu_446_p2[39] };
assign rhs_4_fu_514_p3 = { op_26_V_reg_808, 2'h0 };
assign rhs_6_fu_667_p3 = { op_30_V_reg_852, 1'h0 };
assign sext_ln1192_1_fu_288_p1 = { ret_V_13_fu_265_p3[9], ret_V_13_fu_265_p3 };
assign sext_ln1192_2_fu_442_p1 = { ret_V_15_reg_781[10], ret_V_15_reg_781[10], ret_V_15_reg_781[10], ret_V_15_reg_781[10], ret_V_15_reg_781[10], ret_V_15_reg_781[10], ret_V_15_reg_781[10], ret_V_15_reg_781[10], ret_V_15_reg_781[10], ret_V_15_reg_781[10], ret_V_15_reg_781[10], ret_V_15_reg_781[10], ret_V_15_reg_781[10], ret_V_15_reg_781[10], ret_V_15_reg_781[10], ret_V_15_reg_781[10], ret_V_15_reg_781[10], ret_V_15_reg_781[10], ret_V_15_reg_781[10], ret_V_15_reg_781[10], ret_V_15_reg_781[10], ret_V_15_reg_781[10], ret_V_15_reg_781, 7'h00 };
assign sext_ln1192_3_fu_521_p1 = { op_26_V_reg_808[31], op_26_V_reg_808, 2'h0 };
assign sext_ln1192_4_fu_674_p1 = { op_30_V_reg_852[31], op_30_V_reg_852, 1'h0 };
assign sext_ln1192_fu_213_p1 = { op_0[7], op_0[7], op_0, 7'h00 };
assign sext_ln69_2_fu_619_p1 = { op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16 };
assign sext_ln69_3_fu_306_p1 = { op_10[3], op_10[3], op_10[3], op_10[3], op_10[3], op_10[3], op_10 };
assign sext_ln69_4_fu_378_p1 = { add_ln69_reg_751[9], add_ln69_reg_751 };
assign sext_ln69_5_fu_576_p1 = { op_17[1], op_17 };
assign sext_ln69_6_fu_628_p1 = { add_ln69_4_reg_835[2], add_ln69_4_reg_835[2], add_ln69_4_reg_835[2], add_ln69_4_reg_835[2], add_ln69_4_reg_835[2], add_ln69_4_reg_835[2], add_ln69_4_reg_835[2], add_ln69_4_reg_835[2], add_ln69_4_reg_835[2], add_ln69_4_reg_835[2], add_ln69_4_reg_835[2], add_ln69_4_reg_835[2], add_ln69_4_reg_835[2], add_ln69_4_reg_835[2], add_ln69_4_reg_835[2], add_ln69_4_reg_835[2], add_ln69_4_reg_835[2], add_ln69_4_reg_835[2], add_ln69_4_reg_835[2], add_ln69_4_reg_835[2], add_ln69_4_reg_835[2], add_ln69_4_reg_835[2], add_ln69_4_reg_835[2], add_ln69_4_reg_835[2], add_ln69_4_reg_835[2], add_ln69_4_reg_835[2], add_ln69_4_reg_835[2], add_ln69_4_reg_835[2], add_ln69_4_reg_835[2], add_ln69_4_reg_835 };
assign sext_ln69_fu_298_p1 = { ret_fu_272_p3[1], ret_fu_272_p3[1], ret_fu_272_p3[1], ret_fu_272_p3[1], ret_fu_272_p3[1], ret_fu_272_p3[1], ret_fu_272_p3 };
assign sext_ln703_1_fu_431_p1 = { op_13_V_fu_424_p3[7], op_13_V_fu_424_p3[7], op_13_V_fu_424_p3[7], op_13_V_fu_424_p3[7], op_13_V_fu_424_p3[7], op_13_V_fu_424_p3[7], op_13_V_fu_424_p3[7], op_13_V_fu_424_p3[7], op_13_V_fu_424_p3[7], op_13_V_fu_424_p3[7], op_13_V_fu_424_p3[7], op_13_V_fu_424_p3[7], op_13_V_fu_424_p3[7], op_13_V_fu_424_p3[7], op_13_V_fu_424_p3[7], op_13_V_fu_424_p3[7], op_13_V_fu_424_p3[7], op_13_V_fu_424_p3[7], op_13_V_fu_424_p3[7], op_13_V_fu_424_p3[7], op_13_V_fu_424_p3[7], op_13_V_fu_424_p3[7], op_13_V_fu_424_p3[7], op_13_V_fu_424_p3[7], op_13_V_fu_424_p3[7], op_13_V_fu_424_p3[7], op_13_V_fu_424_p3[7], op_13_V_fu_424_p3[7], op_13_V_fu_424_p3[7], op_13_V_fu_424_p3[7], op_13_V_fu_424_p3[7], op_13_V_fu_424_p3[7], op_13_V_fu_424_p3 };
assign sext_ln703_2_fu_510_p0 = op_15;
assign sext_ln703_2_fu_510_p1 = { op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15 };
assign sext_ln703_3_fu_663_p1 = { op_19_V_fu_655_p3[1], op_19_V_fu_655_p3[1], op_19_V_fu_655_p3[1], op_19_V_fu_655_p3[1], op_19_V_fu_655_p3[1], op_19_V_fu_655_p3[1], op_19_V_fu_655_p3[1], op_19_V_fu_655_p3[1], op_19_V_fu_655_p3[1], op_19_V_fu_655_p3[1], op_19_V_fu_655_p3[1], op_19_V_fu_655_p3[1], op_19_V_fu_655_p3[1], op_19_V_fu_655_p3[1], op_19_V_fu_655_p3[1], op_19_V_fu_655_p3[1], op_19_V_fu_655_p3[1], op_19_V_fu_655_p3[1], op_19_V_fu_655_p3[1], op_19_V_fu_655_p3[1], op_19_V_fu_655_p3[1], op_19_V_fu_655_p3[1], op_19_V_fu_655_p3[1], op_19_V_fu_655_p3[1], op_19_V_fu_655_p3[1], op_19_V_fu_655_p3[1], op_19_V_fu_655_p3[1], op_19_V_fu_655_p3[1], op_19_V_fu_655_p3[1], op_19_V_fu_655_p3[1], op_19_V_fu_655_p3[1], op_19_V_fu_655_p3[1], op_19_V_fu_655_p3 };
assign sext_ln703_fu_217_p0 = op_1;
assign sext_ln703_fu_217_p1 = { op_1[15], op_1 };
assign tmp_1_fu_352_p3 = op_8[1];
assign tmp_3_fu_435_p3 = { ret_V_15_reg_781, 7'h00 };
assign tmp_fu_332_p3 = op_8[1];
assign trunc_ln851_1_fu_462_p1 = op_13_V_fu_424_p3[6:0];
assign trunc_ln851_2_fu_541_p0 = op_15;
assign trunc_ln851_2_fu_541_p1 = op_15[1:0];
assign trunc_ln851_3_fu_701_p1 = op_19_V_reg_857[0];
assign trunc_ln851_fu_237_p0 = op_1;
assign trunc_ln851_fu_237_p1 = op_1[6:0];
assign xor_ln365_fu_360_p2 = p_Result_7_fu_340_p2;
assign xor_ln785_fu_607_p0 = op_11;
assign zext_ln1192_fu_386_p1 = { 10'h000, lhs_V_reg_756 };
assign zext_ln69_fu_302_p1 = { 2'h0, ret_fu_272_p3[1], ret_fu_272_p3[1], ret_fu_272_p3[1], ret_fu_272_p3[1], ret_fu_272_p3[1], ret_fu_272_p3[1], ret_fu_272_p3 };
endmodule


// Machine B:
// Processed by function `add_clk_enable_signal` in `verilog_tricks.py`.
// Processed by function `remove_reset_signal` in `verilog_tricks.py`.
module top_B (
  ap_clk,
  ap_start,
  ap_done,
  ap_idle,
  ap_ready,
  op_0,
  op_1,
  op_2,
  op_3,
  op_4,
  op_8,
  op_10,
  op_11,
  op_14,
  op_15,
  op_16,
  op_17,
  op_31,
  op_31_ap_vld,
clk_enable
);
input clk_enable;


input ap_clk;
wire ap_rst;
assign ap_rst = op_31_ap_vld;
input ap_start;
input [7:0] op_0;
input [15:0] op_1;
input [3:0] op_10;
input op_11;
input op_14;
input [7:0] op_15;
input [3:0] op_16;
input [1:0] op_17;
input op_2;
input [1:0] op_3;
input [1:0] op_4;
input [1:0] op_8;
output ap_done;
output ap_idle;
output ap_ready;
output [31:0] op_31;
output op_31_ap_vld;


reg [4:0] \add_10ns_10ns_10_2_1_U2.top_add_10ns_10ns_10_2_1_Adder_1_U.ain_s1 ;
reg [4:0] \add_10ns_10ns_10_2_1_U2.top_add_10ns_10ns_10_2_1_Adder_1_U.bin_s1 ;
reg \add_10ns_10ns_10_2_1_U2.top_add_10ns_10ns_10_2_1_Adder_1_U.carry_s1 ;
reg [4:0] \add_10ns_10ns_10_2_1_U2.top_add_10ns_10ns_10_2_1_Adder_1_U.sum_s1 ;
reg [4:0] \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.ain_s1 ;
reg [4:0] \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.bin_s1 ;
reg \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.carry_s1 ;
reg [4:0] \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.sum_s1 ;
reg [5:0] \add_11ns_11ns_11_2_1_U6.top_add_11ns_11ns_11_2_1_Adder_4_U.ain_s1 ;
reg [5:0] \add_11ns_11ns_11_2_1_U6.top_add_11ns_11ns_11_2_1_Adder_4_U.bin_s1 ;
reg \add_11ns_11ns_11_2_1_U6.top_add_11ns_11ns_11_2_1_Adder_4_U.carry_s1 ;
reg [4:0] \add_11ns_11ns_11_2_1_U6.top_add_11ns_11ns_11_2_1_Adder_4_U.sum_s1 ;
reg [5:0] \add_11s_11ns_11_2_1_U3.top_add_11s_11ns_11_2_1_Adder_2_U.ain_s1 ;
reg [5:0] \add_11s_11ns_11_2_1_U3.top_add_11s_11ns_11_2_1_Adder_2_U.bin_s1 ;
reg \add_11s_11ns_11_2_1_U3.top_add_11s_11ns_11_2_1_Adder_2_U.carry_s1 ;
reg [4:0] \add_11s_11ns_11_2_1_U3.top_add_11s_11ns_11_2_1_Adder_2_U.sum_s1 ;
reg [5:0] \add_11s_11ns_11_2_1_U5.top_add_11s_11ns_11_2_1_Adder_2_U.ain_s1 ;
reg [5:0] \add_11s_11ns_11_2_1_U5.top_add_11s_11ns_11_2_1_Adder_2_U.bin_s1 ;
reg \add_11s_11ns_11_2_1_U5.top_add_11s_11ns_11_2_1_Adder_2_U.carry_s1 ;
reg [4:0] \add_11s_11ns_11_2_1_U5.top_add_11s_11ns_11_2_1_Adder_2_U.sum_s1 ;
reg [8:0] \add_17s_17s_17_2_1_U1.top_add_17s_17s_17_2_1_Adder_0_U.ain_s1 ;
reg [8:0] \add_17s_17s_17_2_1_U1.top_add_17s_17s_17_2_1_Adder_0_U.bin_s1 ;
reg \add_17s_17s_17_2_1_U1.top_add_17s_17s_17_2_1_Adder_0_U.carry_s1 ;
reg [7:0] \add_17s_17s_17_2_1_U1.top_add_17s_17s_17_2_1_Adder_0_U.sum_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s1 ;
reg \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_6_U.carry_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_6_U.sum_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s1 ;
reg \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.carry_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.sum_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s1 ;
reg \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.carry_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.sum_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s1 ;
reg \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.carry_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.sum_s1 ;
reg [15:0] \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.ain_s1 ;
reg [15:0] \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.bin_s1 ;
reg \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.carry_s1 ;
reg [15:0] \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.sum_s1 ;
reg [15:0] \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_10_U.ain_s1 ;
reg [15:0] \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_10_U.bin_s1 ;
reg \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_10_U.carry_s1 ;
reg [15:0] \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_10_U.sum_s1 ;
reg [16:0] \add_34s_34s_34_2_1_U15.top_add_34s_34s_34_2_1_Adder_11_U.ain_s1 ;
reg [16:0] \add_34s_34s_34_2_1_U15.top_add_34s_34s_34_2_1_Adder_11_U.bin_s1 ;
reg \add_34s_34s_34_2_1_U15.top_add_34s_34s_34_2_1_Adder_11_U.carry_s1 ;
reg [16:0] \add_34s_34s_34_2_1_U15.top_add_34s_34s_34_2_1_Adder_11_U.sum_s1 ;
reg [17:0] \add_35s_35s_35_2_1_U10.top_add_35s_35s_35_2_1_Adder_7_U.ain_s1 ;
reg [17:0] \add_35s_35s_35_2_1_U10.top_add_35s_35s_35_2_1_Adder_7_U.bin_s1 ;
reg \add_35s_35s_35_2_1_U10.top_add_35s_35s_35_2_1_Adder_7_U.carry_s1 ;
reg [16:0] \add_35s_35s_35_2_1_U10.top_add_35s_35s_35_2_1_Adder_7_U.sum_s1 ;
reg [1:0] \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_9_U.ain_s1 ;
reg [1:0] \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_9_U.bin_s1 ;
reg \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_9_U.carry_s1 ;
reg \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_9_U.sum_s1 ;
reg [19:0] \add_40s_40s_40_2_1_U7.top_add_40s_40s_40_2_1_Adder_5_U.ain_s1 ;
reg [19:0] \add_40s_40s_40_2_1_U7.top_add_40s_40s_40_2_1_Adder_5_U.bin_s1 ;
reg \add_40s_40s_40_2_1_U7.top_add_40s_40s_40_2_1_Adder_5_U.carry_s1 ;
reg [19:0] \add_40s_40s_40_2_1_U7.top_add_40s_40s_40_2_1_Adder_5_U.sum_s1 ;
reg [31:0] add_ln691_1_reg_922;
reg [31:0] add_ln691_2_reg_1013;
reg [31:0] add_ln691_reg_875;
reg [31:0] add_ln69_3_reg_959;
reg [2:0] add_ln69_4_reg_964;
reg [9:0] add_ln69_reg_775;
reg and_ln365_reg_823;
reg [31:0] ap_CS_fsm = 32'd1;
reg empty_reg_785;
reg icmp_ln785_reg_954;
reg icmp_ln851_1_reg_858;
reg icmp_ln851_2_reg_905;
reg icmp_ln851_reg_712;
reg lhs_V_reg_818;
reg [7:0] op_13_V_reg_833;
reg [1:0] op_19_V_reg_980;
reg [10:0] op_23_V_reg_813;
reg [31:0] op_26_V_reg_890;
reg [31:0] op_30_V_reg_986;
reg or_ln785_reg_807;
reg overflow_reg_969;
reg p_Result_7_reg_796;
reg r_reg_790;
reg [16:0] ret_V_12_reg_717;
reg [9:0] ret_V_13_reg_740;
reg [10:0] ret_V_14_reg_770;
reg [10:0] ret_V_15_reg_838;
reg [31:0] ret_V_16_cast_reg_1006;
reg [39:0] ret_V_16_reg_863;
reg [31:0] ret_V_17_reg_880;
reg [34:0] ret_V_18_reg_910;
reg [31:0] ret_V_19_reg_927;
reg [33:0] ret_V_20_reg_1001;
reg [9:0] ret_V_2_reg_729;
reg [31:0] ret_V_6_cast_reg_868;
reg [31:0] ret_V_9_cast_reg_915;
reg [9:0] ret_V_reg_722;
reg [1:0] ret_reg_745;
reg [10:0] select_ln1192_reg_750;
reg [2:0] select_ln69_1_reg_932;
reg [31:0] select_ln69_reg_885;
reg [6:0] trunc_ln851_1_reg_843;
wire [31:0] _000_;
wire [31:0] _001_;
wire [31:0] _002_;
wire [31:0] _003_;
wire [2:0] _004_;
wire [9:0] _005_;
wire _006_;
wire [31:0] _007_;
wire _008_;
wire _009_;
wire _010_;
wire _011_;
wire _012_;
wire _013_;
wire [7:0] _014_;
wire [1:0] _015_;
wire [10:0] _016_;
wire [31:0] _017_;
wire [31:0] _018_;
wire _019_;
wire _020_;
wire _021_;
wire _022_;
wire [16:0] _023_;
wire [9:0] _024_;
wire [10:0] _025_;
wire [10:0] _026_;
wire [31:0] _027_;
wire [39:0] _028_;
wire [31:0] _029_;
wire [34:0] _030_;
wire [31:0] _031_;
wire [33:0] _032_;
wire [9:0] _033_;
wire [31:0] _034_;
wire [31:0] _035_;
wire [9:0] _036_;
wire [1:0] _037_;
wire [10:0] _038_;
wire [2:0] _039_;
wire [31:0] _040_;
wire [6:0] _041_;
wire [1:0] _042_;
wire _043_;
wire _044_;
wire _045_;
wire _046_;
wire _047_;
wire _048_;
wire _049_;
wire _050_;
wire [4:0] _051_;
wire [4:0] _052_;
wire _053_;
wire [4:0] _054_;
wire [5:0] _055_;
wire [5:0] _056_;
wire [4:0] _057_;
wire [4:0] _058_;
wire _059_;
wire [4:0] _060_;
wire [5:0] _061_;
wire [5:0] _062_;
wire [5:0] _063_;
wire [5:0] _064_;
wire _065_;
wire [4:0] _066_;
wire [5:0] _067_;
wire [6:0] _068_;
wire [5:0] _069_;
wire [5:0] _070_;
wire _071_;
wire [4:0] _072_;
wire [5:0] _073_;
wire [6:0] _074_;
wire [5:0] _075_;
wire [5:0] _076_;
wire _077_;
wire [4:0] _078_;
wire [5:0] _079_;
wire [6:0] _080_;
wire [8:0] _081_;
wire [8:0] _082_;
wire _083_;
wire [7:0] _084_;
wire [8:0] _085_;
wire [9:0] _086_;
wire [15:0] _087_;
wire [15:0] _088_;
wire _089_;
wire [15:0] _090_;
wire [16:0] _091_;
wire [16:0] _092_;
wire [15:0] _093_;
wire [15:0] _094_;
wire _095_;
wire [15:0] _096_;
wire [16:0] _097_;
wire [16:0] _098_;
wire [15:0] _099_;
wire [15:0] _100_;
wire _101_;
wire [15:0] _102_;
wire [16:0] _103_;
wire [16:0] _104_;
wire [15:0] _105_;
wire [15:0] _106_;
wire _107_;
wire [15:0] _108_;
wire [16:0] _109_;
wire [16:0] _110_;
wire [15:0] _111_;
wire [15:0] _112_;
wire _113_;
wire [15:0] _114_;
wire [16:0] _115_;
wire [16:0] _116_;
wire [15:0] _117_;
wire [15:0] _118_;
wire _119_;
wire [15:0] _120_;
wire [16:0] _121_;
wire [16:0] _122_;
wire [16:0] _123_;
wire [16:0] _124_;
wire _125_;
wire [16:0] _126_;
wire [17:0] _127_;
wire [17:0] _128_;
wire [17:0] _129_;
wire [17:0] _130_;
wire _131_;
wire [16:0] _132_;
wire [17:0] _133_;
wire [18:0] _134_;
wire [1:0] _135_;
wire [1:0] _136_;
wire _137_;
wire _138_;
wire [1:0] _139_;
wire [2:0] _140_;
wire [19:0] _141_;
wire [19:0] _142_;
wire _143_;
wire [19:0] _144_;
wire [20:0] _145_;
wire [20:0] _146_;
wire _147_;
wire _148_;
wire _149_;
wire _150_;
wire _151_;
wire _152_;
wire _153_;
wire _154_;
wire _155_;
wire _156_;
wire _157_;
wire _158_;
wire _159_;
wire _160_;
wire _161_;
wire _162_;
wire _163_;
wire _164_;
wire _165_;
wire _166_;
wire _167_;
wire _168_;
wire _169_;
wire _170_;
wire _171_;
wire _172_;
wire _173_;
wire _174_;
wire _175_;
wire _176_;
wire _177_;
wire _178_;
wire _179_;
wire _180_;
wire \add_10ns_10ns_10_2_1_U2.ce ;
wire \add_10ns_10ns_10_2_1_U2.clk ;
wire [9:0] \add_10ns_10ns_10_2_1_U2.din0 ;
wire [9:0] \add_10ns_10ns_10_2_1_U2.din1 ;
wire [9:0] \add_10ns_10ns_10_2_1_U2.dout ;
wire \add_10ns_10ns_10_2_1_U2.reset ;
wire [9:0] \add_10ns_10ns_10_2_1_U2.top_add_10ns_10ns_10_2_1_Adder_1_U.a ;
wire [9:0] \add_10ns_10ns_10_2_1_U2.top_add_10ns_10ns_10_2_1_Adder_1_U.ain_s0 ;
wire [9:0] \add_10ns_10ns_10_2_1_U2.top_add_10ns_10ns_10_2_1_Adder_1_U.b ;
wire [9:0] \add_10ns_10ns_10_2_1_U2.top_add_10ns_10ns_10_2_1_Adder_1_U.bin_s0 ;
wire \add_10ns_10ns_10_2_1_U2.top_add_10ns_10ns_10_2_1_Adder_1_U.ce ;
wire \add_10ns_10ns_10_2_1_U2.top_add_10ns_10ns_10_2_1_Adder_1_U.clk ;
wire \add_10ns_10ns_10_2_1_U2.top_add_10ns_10ns_10_2_1_Adder_1_U.facout_s1 ;
wire \add_10ns_10ns_10_2_1_U2.top_add_10ns_10ns_10_2_1_Adder_1_U.facout_s2 ;
wire [4:0] \add_10ns_10ns_10_2_1_U2.top_add_10ns_10ns_10_2_1_Adder_1_U.fas_s1 ;
wire [4:0] \add_10ns_10ns_10_2_1_U2.top_add_10ns_10ns_10_2_1_Adder_1_U.fas_s2 ;
wire \add_10ns_10ns_10_2_1_U2.top_add_10ns_10ns_10_2_1_Adder_1_U.reset ;
wire [9:0] \add_10ns_10ns_10_2_1_U2.top_add_10ns_10ns_10_2_1_Adder_1_U.s ;
wire [4:0] \add_10ns_10ns_10_2_1_U2.top_add_10ns_10ns_10_2_1_Adder_1_U.u1.a ;
wire [4:0] \add_10ns_10ns_10_2_1_U2.top_add_10ns_10ns_10_2_1_Adder_1_U.u1.b ;
wire \add_10ns_10ns_10_2_1_U2.top_add_10ns_10ns_10_2_1_Adder_1_U.u1.cin ;
wire \add_10ns_10ns_10_2_1_U2.top_add_10ns_10ns_10_2_1_Adder_1_U.u1.cout ;
wire [4:0] \add_10ns_10ns_10_2_1_U2.top_add_10ns_10ns_10_2_1_Adder_1_U.u1.s ;
wire [4:0] \add_10ns_10ns_10_2_1_U2.top_add_10ns_10ns_10_2_1_Adder_1_U.u2.a ;
wire [4:0] \add_10ns_10ns_10_2_1_U2.top_add_10ns_10ns_10_2_1_Adder_1_U.u2.b ;
wire \add_10ns_10ns_10_2_1_U2.top_add_10ns_10ns_10_2_1_Adder_1_U.u2.cin ;
wire \add_10ns_10ns_10_2_1_U2.top_add_10ns_10ns_10_2_1_Adder_1_U.u2.cout ;
wire [4:0] \add_10ns_10ns_10_2_1_U2.top_add_10ns_10ns_10_2_1_Adder_1_U.u2.s ;
wire \add_10ns_10s_10_2_1_U4.ce ;
wire \add_10ns_10s_10_2_1_U4.clk ;
wire [9:0] \add_10ns_10s_10_2_1_U4.din0 ;
wire [9:0] \add_10ns_10s_10_2_1_U4.din1 ;
wire [9:0] \add_10ns_10s_10_2_1_U4.dout ;
wire \add_10ns_10s_10_2_1_U4.reset ;
wire [9:0] \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.a ;
wire [9:0] \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.ain_s0 ;
wire [9:0] \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.b ;
wire [9:0] \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.bin_s0 ;
wire \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.ce ;
wire \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.clk ;
wire \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.facout_s1 ;
wire \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.facout_s2 ;
wire [4:0] \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.fas_s1 ;
wire [4:0] \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.fas_s2 ;
wire \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.reset ;
wire [9:0] \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.s ;
wire [4:0] \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.u1.a ;
wire [4:0] \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.u1.b ;
wire \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.u1.cin ;
wire \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.u1.cout ;
wire [4:0] \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.u1.s ;
wire [4:0] \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.u2.a ;
wire [4:0] \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.u2.b ;
wire \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.u2.cin ;
wire \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.u2.cout ;
wire [4:0] \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.u2.s ;
wire \add_11ns_11ns_11_2_1_U6.ce ;
wire \add_11ns_11ns_11_2_1_U6.clk ;
wire [10:0] \add_11ns_11ns_11_2_1_U6.din0 ;
wire [10:0] \add_11ns_11ns_11_2_1_U6.din1 ;
wire [10:0] \add_11ns_11ns_11_2_1_U6.dout ;
wire \add_11ns_11ns_11_2_1_U6.reset ;
wire [10:0] \add_11ns_11ns_11_2_1_U6.top_add_11ns_11ns_11_2_1_Adder_4_U.a ;
wire [10:0] \add_11ns_11ns_11_2_1_U6.top_add_11ns_11ns_11_2_1_Adder_4_U.ain_s0 ;
wire [10:0] \add_11ns_11ns_11_2_1_U6.top_add_11ns_11ns_11_2_1_Adder_4_U.b ;
wire [10:0] \add_11ns_11ns_11_2_1_U6.top_add_11ns_11ns_11_2_1_Adder_4_U.bin_s0 ;
wire \add_11ns_11ns_11_2_1_U6.top_add_11ns_11ns_11_2_1_Adder_4_U.ce ;
wire \add_11ns_11ns_11_2_1_U6.top_add_11ns_11ns_11_2_1_Adder_4_U.clk ;
wire \add_11ns_11ns_11_2_1_U6.top_add_11ns_11ns_11_2_1_Adder_4_U.facout_s1 ;
wire \add_11ns_11ns_11_2_1_U6.top_add_11ns_11ns_11_2_1_Adder_4_U.facout_s2 ;
wire [4:0] \add_11ns_11ns_11_2_1_U6.top_add_11ns_11ns_11_2_1_Adder_4_U.fas_s1 ;
wire [5:0] \add_11ns_11ns_11_2_1_U6.top_add_11ns_11ns_11_2_1_Adder_4_U.fas_s2 ;
wire \add_11ns_11ns_11_2_1_U6.top_add_11ns_11ns_11_2_1_Adder_4_U.reset ;
wire [10:0] \add_11ns_11ns_11_2_1_U6.top_add_11ns_11ns_11_2_1_Adder_4_U.s ;
wire [4:0] \add_11ns_11ns_11_2_1_U6.top_add_11ns_11ns_11_2_1_Adder_4_U.u1.a ;
wire [4:0] \add_11ns_11ns_11_2_1_U6.top_add_11ns_11ns_11_2_1_Adder_4_U.u1.b ;
wire \add_11ns_11ns_11_2_1_U6.top_add_11ns_11ns_11_2_1_Adder_4_U.u1.cin ;
wire \add_11ns_11ns_11_2_1_U6.top_add_11ns_11ns_11_2_1_Adder_4_U.u1.cout ;
wire [4:0] \add_11ns_11ns_11_2_1_U6.top_add_11ns_11ns_11_2_1_Adder_4_U.u1.s ;
wire [5:0] \add_11ns_11ns_11_2_1_U6.top_add_11ns_11ns_11_2_1_Adder_4_U.u2.a ;
wire [5:0] \add_11ns_11ns_11_2_1_U6.top_add_11ns_11ns_11_2_1_Adder_4_U.u2.b ;
wire \add_11ns_11ns_11_2_1_U6.top_add_11ns_11ns_11_2_1_Adder_4_U.u2.cin ;
wire \add_11ns_11ns_11_2_1_U6.top_add_11ns_11ns_11_2_1_Adder_4_U.u2.cout ;
wire [5:0] \add_11ns_11ns_11_2_1_U6.top_add_11ns_11ns_11_2_1_Adder_4_U.u2.s ;
wire \add_11s_11ns_11_2_1_U3.ce ;
wire \add_11s_11ns_11_2_1_U3.clk ;
wire [10:0] \add_11s_11ns_11_2_1_U3.din0 ;
wire [10:0] \add_11s_11ns_11_2_1_U3.din1 ;
wire [10:0] \add_11s_11ns_11_2_1_U3.dout ;
wire \add_11s_11ns_11_2_1_U3.reset ;
wire [10:0] \add_11s_11ns_11_2_1_U3.top_add_11s_11ns_11_2_1_Adder_2_U.a ;
wire [10:0] \add_11s_11ns_11_2_1_U3.top_add_11s_11ns_11_2_1_Adder_2_U.ain_s0 ;
wire [10:0] \add_11s_11ns_11_2_1_U3.top_add_11s_11ns_11_2_1_Adder_2_U.b ;
wire [10:0] \add_11s_11ns_11_2_1_U3.top_add_11s_11ns_11_2_1_Adder_2_U.bin_s0 ;
wire \add_11s_11ns_11_2_1_U3.top_add_11s_11ns_11_2_1_Adder_2_U.ce ;
wire \add_11s_11ns_11_2_1_U3.top_add_11s_11ns_11_2_1_Adder_2_U.clk ;
wire \add_11s_11ns_11_2_1_U3.top_add_11s_11ns_11_2_1_Adder_2_U.facout_s1 ;
wire \add_11s_11ns_11_2_1_U3.top_add_11s_11ns_11_2_1_Adder_2_U.facout_s2 ;
wire [4:0] \add_11s_11ns_11_2_1_U3.top_add_11s_11ns_11_2_1_Adder_2_U.fas_s1 ;
wire [5:0] \add_11s_11ns_11_2_1_U3.top_add_11s_11ns_11_2_1_Adder_2_U.fas_s2 ;
wire \add_11s_11ns_11_2_1_U3.top_add_11s_11ns_11_2_1_Adder_2_U.reset ;
wire [10:0] \add_11s_11ns_11_2_1_U3.top_add_11s_11ns_11_2_1_Adder_2_U.s ;
wire [4:0] \add_11s_11ns_11_2_1_U3.top_add_11s_11ns_11_2_1_Adder_2_U.u1.a ;
wire [4:0] \add_11s_11ns_11_2_1_U3.top_add_11s_11ns_11_2_1_Adder_2_U.u1.b ;
wire \add_11s_11ns_11_2_1_U3.top_add_11s_11ns_11_2_1_Adder_2_U.u1.cin ;
wire \add_11s_11ns_11_2_1_U3.top_add_11s_11ns_11_2_1_Adder_2_U.u1.cout ;
wire [4:0] \add_11s_11ns_11_2_1_U3.top_add_11s_11ns_11_2_1_Adder_2_U.u1.s ;
wire [5:0] \add_11s_11ns_11_2_1_U3.top_add_11s_11ns_11_2_1_Adder_2_U.u2.a ;
wire [5:0] \add_11s_11ns_11_2_1_U3.top_add_11s_11ns_11_2_1_Adder_2_U.u2.b ;
wire \add_11s_11ns_11_2_1_U3.top_add_11s_11ns_11_2_1_Adder_2_U.u2.cin ;
wire \add_11s_11ns_11_2_1_U3.top_add_11s_11ns_11_2_1_Adder_2_U.u2.cout ;
wire [5:0] \add_11s_11ns_11_2_1_U3.top_add_11s_11ns_11_2_1_Adder_2_U.u2.s ;
wire \add_11s_11ns_11_2_1_U5.ce ;
wire \add_11s_11ns_11_2_1_U5.clk ;
wire [10:0] \add_11s_11ns_11_2_1_U5.din0 ;
wire [10:0] \add_11s_11ns_11_2_1_U5.din1 ;
wire [10:0] \add_11s_11ns_11_2_1_U5.dout ;
wire \add_11s_11ns_11_2_1_U5.reset ;
wire [10:0] \add_11s_11ns_11_2_1_U5.top_add_11s_11ns_11_2_1_Adder_2_U.a ;
wire [10:0] \add_11s_11ns_11_2_1_U5.top_add_11s_11ns_11_2_1_Adder_2_U.ain_s0 ;
wire [10:0] \add_11s_11ns_11_2_1_U5.top_add_11s_11ns_11_2_1_Adder_2_U.b ;
wire [10:0] \add_11s_11ns_11_2_1_U5.top_add_11s_11ns_11_2_1_Adder_2_U.bin_s0 ;
wire \add_11s_11ns_11_2_1_U5.top_add_11s_11ns_11_2_1_Adder_2_U.ce ;
wire \add_11s_11ns_11_2_1_U5.top_add_11s_11ns_11_2_1_Adder_2_U.clk ;
wire \add_11s_11ns_11_2_1_U5.top_add_11s_11ns_11_2_1_Adder_2_U.facout_s1 ;
wire \add_11s_11ns_11_2_1_U5.top_add_11s_11ns_11_2_1_Adder_2_U.facout_s2 ;
wire [4:0] \add_11s_11ns_11_2_1_U5.top_add_11s_11ns_11_2_1_Adder_2_U.fas_s1 ;
wire [5:0] \add_11s_11ns_11_2_1_U5.top_add_11s_11ns_11_2_1_Adder_2_U.fas_s2 ;
wire \add_11s_11ns_11_2_1_U5.top_add_11s_11ns_11_2_1_Adder_2_U.reset ;
wire [10:0] \add_11s_11ns_11_2_1_U5.top_add_11s_11ns_11_2_1_Adder_2_U.s ;
wire [4:0] \add_11s_11ns_11_2_1_U5.top_add_11s_11ns_11_2_1_Adder_2_U.u1.a ;
wire [4:0] \add_11s_11ns_11_2_1_U5.top_add_11s_11ns_11_2_1_Adder_2_U.u1.b ;
wire \add_11s_11ns_11_2_1_U5.top_add_11s_11ns_11_2_1_Adder_2_U.u1.cin ;
wire \add_11s_11ns_11_2_1_U5.top_add_11s_11ns_11_2_1_Adder_2_U.u1.cout ;
wire [4:0] \add_11s_11ns_11_2_1_U5.top_add_11s_11ns_11_2_1_Adder_2_U.u1.s ;
wire [5:0] \add_11s_11ns_11_2_1_U5.top_add_11s_11ns_11_2_1_Adder_2_U.u2.a ;
wire [5:0] \add_11s_11ns_11_2_1_U5.top_add_11s_11ns_11_2_1_Adder_2_U.u2.b ;
wire \add_11s_11ns_11_2_1_U5.top_add_11s_11ns_11_2_1_Adder_2_U.u2.cin ;
wire \add_11s_11ns_11_2_1_U5.top_add_11s_11ns_11_2_1_Adder_2_U.u2.cout ;
wire [5:0] \add_11s_11ns_11_2_1_U5.top_add_11s_11ns_11_2_1_Adder_2_U.u2.s ;
wire \add_17s_17s_17_2_1_U1.ce ;
wire \add_17s_17s_17_2_1_U1.clk ;
wire [16:0] \add_17s_17s_17_2_1_U1.din0 ;
wire [16:0] \add_17s_17s_17_2_1_U1.din1 ;
wire [16:0] \add_17s_17s_17_2_1_U1.dout ;
wire \add_17s_17s_17_2_1_U1.reset ;
wire [16:0] \add_17s_17s_17_2_1_U1.top_add_17s_17s_17_2_1_Adder_0_U.a ;
wire [16:0] \add_17s_17s_17_2_1_U1.top_add_17s_17s_17_2_1_Adder_0_U.ain_s0 ;
wire [16:0] \add_17s_17s_17_2_1_U1.top_add_17s_17s_17_2_1_Adder_0_U.b ;
wire [16:0] \add_17s_17s_17_2_1_U1.top_add_17s_17s_17_2_1_Adder_0_U.bin_s0 ;
wire \add_17s_17s_17_2_1_U1.top_add_17s_17s_17_2_1_Adder_0_U.ce ;
wire \add_17s_17s_17_2_1_U1.top_add_17s_17s_17_2_1_Adder_0_U.clk ;
wire \add_17s_17s_17_2_1_U1.top_add_17s_17s_17_2_1_Adder_0_U.facout_s1 ;
wire \add_17s_17s_17_2_1_U1.top_add_17s_17s_17_2_1_Adder_0_U.facout_s2 ;
wire [7:0] \add_17s_17s_17_2_1_U1.top_add_17s_17s_17_2_1_Adder_0_U.fas_s1 ;
wire [8:0] \add_17s_17s_17_2_1_U1.top_add_17s_17s_17_2_1_Adder_0_U.fas_s2 ;
wire \add_17s_17s_17_2_1_U1.top_add_17s_17s_17_2_1_Adder_0_U.reset ;
wire [16:0] \add_17s_17s_17_2_1_U1.top_add_17s_17s_17_2_1_Adder_0_U.s ;
wire [7:0] \add_17s_17s_17_2_1_U1.top_add_17s_17s_17_2_1_Adder_0_U.u1.a ;
wire [7:0] \add_17s_17s_17_2_1_U1.top_add_17s_17s_17_2_1_Adder_0_U.u1.b ;
wire \add_17s_17s_17_2_1_U1.top_add_17s_17s_17_2_1_Adder_0_U.u1.cin ;
wire \add_17s_17s_17_2_1_U1.top_add_17s_17s_17_2_1_Adder_0_U.u1.cout ;
wire [7:0] \add_17s_17s_17_2_1_U1.top_add_17s_17s_17_2_1_Adder_0_U.u1.s ;
wire [8:0] \add_17s_17s_17_2_1_U1.top_add_17s_17s_17_2_1_Adder_0_U.u2.a ;
wire [8:0] \add_17s_17s_17_2_1_U1.top_add_17s_17s_17_2_1_Adder_0_U.u2.b ;
wire \add_17s_17s_17_2_1_U1.top_add_17s_17s_17_2_1_Adder_0_U.u2.cin ;
wire \add_17s_17s_17_2_1_U1.top_add_17s_17s_17_2_1_Adder_0_U.u2.cout ;
wire [8:0] \add_17s_17s_17_2_1_U1.top_add_17s_17s_17_2_1_Adder_0_U.u2.s ;
wire \add_32ns_32ns_32_2_1_U11.ce ;
wire \add_32ns_32ns_32_2_1_U11.clk ;
wire [31:0] \add_32ns_32ns_32_2_1_U11.din0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U11.din1 ;
wire [31:0] \add_32ns_32ns_32_2_1_U11.dout ;
wire \add_32ns_32ns_32_2_1_U11.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_6_U.a ;
wire [31:0] \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_6_U.b ;
wire [31:0] \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s0 ;
wire \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_6_U.ce ;
wire \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_6_U.clk ;
wire \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s1 ;
wire \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s2 ;
wire [15:0] \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s1 ;
wire [15:0] \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s2 ;
wire \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_6_U.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_6_U.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.b ;
wire \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cin ;
wire \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.b ;
wire \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cin ;
wire \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.s ;
wire \add_32ns_32ns_32_2_1_U16.ce ;
wire \add_32ns_32ns_32_2_1_U16.clk ;
wire [31:0] \add_32ns_32ns_32_2_1_U16.din0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U16.din1 ;
wire [31:0] \add_32ns_32ns_32_2_1_U16.dout ;
wire \add_32ns_32ns_32_2_1_U16.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.a ;
wire [31:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.b ;
wire [31:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s0 ;
wire \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.ce ;
wire \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.clk ;
wire \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s1 ;
wire \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s2 ;
wire [15:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s1 ;
wire [15:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s2 ;
wire \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.b ;
wire \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cin ;
wire \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.b ;
wire \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cin ;
wire \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.s ;
wire \add_32ns_32ns_32_2_1_U8.ce ;
wire \add_32ns_32ns_32_2_1_U8.clk ;
wire [31:0] \add_32ns_32ns_32_2_1_U8.din0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U8.din1 ;
wire [31:0] \add_32ns_32ns_32_2_1_U8.dout ;
wire \add_32ns_32ns_32_2_1_U8.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.a ;
wire [31:0] \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.b ;
wire [31:0] \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s0 ;
wire \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.ce ;
wire \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.clk ;
wire \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s1 ;
wire \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s2 ;
wire [15:0] \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s1 ;
wire [15:0] \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s2 ;
wire \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.b ;
wire \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cin ;
wire \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.b ;
wire \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cin ;
wire \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.s ;
wire \add_32ns_32ns_32_2_1_U9.ce ;
wire \add_32ns_32ns_32_2_1_U9.clk ;
wire [31:0] \add_32ns_32ns_32_2_1_U9.din0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U9.din1 ;
wire [31:0] \add_32ns_32ns_32_2_1_U9.dout ;
wire \add_32ns_32ns_32_2_1_U9.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.a ;
wire [31:0] \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.b ;
wire [31:0] \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s0 ;
wire \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.ce ;
wire \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.clk ;
wire \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s1 ;
wire \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s2 ;
wire [15:0] \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s1 ;
wire [15:0] \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s2 ;
wire \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.b ;
wire \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cin ;
wire \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.b ;
wire \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cin ;
wire \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.s ;
wire \add_32ns_32s_32_2_1_U12.ce ;
wire \add_32ns_32s_32_2_1_U12.clk ;
wire [31:0] \add_32ns_32s_32_2_1_U12.din0 ;
wire [31:0] \add_32ns_32s_32_2_1_U12.din1 ;
wire [31:0] \add_32ns_32s_32_2_1_U12.dout ;
wire \add_32ns_32s_32_2_1_U12.reset ;
wire [31:0] \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.a ;
wire [31:0] \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.ain_s0 ;
wire [31:0] \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.b ;
wire [31:0] \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.bin_s0 ;
wire \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.ce ;
wire \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.clk ;
wire \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.facout_s1 ;
wire \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.facout_s2 ;
wire [15:0] \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.fas_s1 ;
wire [15:0] \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.fas_s2 ;
wire \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.reset ;
wire [31:0] \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.s ;
wire [15:0] \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.u1.a ;
wire [15:0] \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.u1.b ;
wire \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.u1.cin ;
wire \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.u1.cout ;
wire [15:0] \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.u1.s ;
wire [15:0] \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.u2.a ;
wire [15:0] \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.u2.b ;
wire \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.u2.cin ;
wire \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.u2.cout ;
wire [15:0] \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.u2.s ;
wire \add_32s_32ns_32_2_1_U14.ce ;
wire \add_32s_32ns_32_2_1_U14.clk ;
wire [31:0] \add_32s_32ns_32_2_1_U14.din0 ;
wire [31:0] \add_32s_32ns_32_2_1_U14.din1 ;
wire [31:0] \add_32s_32ns_32_2_1_U14.dout ;
wire \add_32s_32ns_32_2_1_U14.reset ;
wire [31:0] \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_10_U.a ;
wire [31:0] \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_10_U.ain_s0 ;
wire [31:0] \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_10_U.b ;
wire [31:0] \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_10_U.bin_s0 ;
wire \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_10_U.ce ;
wire \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_10_U.clk ;
wire \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_10_U.facout_s1 ;
wire \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_10_U.facout_s2 ;
wire [15:0] \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_10_U.fas_s1 ;
wire [15:0] \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_10_U.fas_s2 ;
wire \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_10_U.reset ;
wire [31:0] \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_10_U.s ;
wire [15:0] \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_10_U.u1.a ;
wire [15:0] \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_10_U.u1.b ;
wire \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_10_U.u1.cin ;
wire \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_10_U.u1.cout ;
wire [15:0] \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_10_U.u1.s ;
wire [15:0] \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_10_U.u2.a ;
wire [15:0] \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_10_U.u2.b ;
wire \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_10_U.u2.cin ;
wire \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_10_U.u2.cout ;
wire [15:0] \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_10_U.u2.s ;
wire \add_34s_34s_34_2_1_U15.ce ;
wire \add_34s_34s_34_2_1_U15.clk ;
wire [33:0] \add_34s_34s_34_2_1_U15.din0 ;
wire [33:0] \add_34s_34s_34_2_1_U15.din1 ;
wire [33:0] \add_34s_34s_34_2_1_U15.dout ;
wire \add_34s_34s_34_2_1_U15.reset ;
wire [33:0] \add_34s_34s_34_2_1_U15.top_add_34s_34s_34_2_1_Adder_11_U.a ;
wire [33:0] \add_34s_34s_34_2_1_U15.top_add_34s_34s_34_2_1_Adder_11_U.ain_s0 ;
wire [33:0] \add_34s_34s_34_2_1_U15.top_add_34s_34s_34_2_1_Adder_11_U.b ;
wire [33:0] \add_34s_34s_34_2_1_U15.top_add_34s_34s_34_2_1_Adder_11_U.bin_s0 ;
wire \add_34s_34s_34_2_1_U15.top_add_34s_34s_34_2_1_Adder_11_U.ce ;
wire \add_34s_34s_34_2_1_U15.top_add_34s_34s_34_2_1_Adder_11_U.clk ;
wire \add_34s_34s_34_2_1_U15.top_add_34s_34s_34_2_1_Adder_11_U.facout_s1 ;
wire \add_34s_34s_34_2_1_U15.top_add_34s_34s_34_2_1_Adder_11_U.facout_s2 ;
wire [16:0] \add_34s_34s_34_2_1_U15.top_add_34s_34s_34_2_1_Adder_11_U.fas_s1 ;
wire [16:0] \add_34s_34s_34_2_1_U15.top_add_34s_34s_34_2_1_Adder_11_U.fas_s2 ;
wire \add_34s_34s_34_2_1_U15.top_add_34s_34s_34_2_1_Adder_11_U.reset ;
wire [33:0] \add_34s_34s_34_2_1_U15.top_add_34s_34s_34_2_1_Adder_11_U.s ;
wire [16:0] \add_34s_34s_34_2_1_U15.top_add_34s_34s_34_2_1_Adder_11_U.u1.a ;
wire [16:0] \add_34s_34s_34_2_1_U15.top_add_34s_34s_34_2_1_Adder_11_U.u1.b ;
wire \add_34s_34s_34_2_1_U15.top_add_34s_34s_34_2_1_Adder_11_U.u1.cin ;
wire \add_34s_34s_34_2_1_U15.top_add_34s_34s_34_2_1_Adder_11_U.u1.cout ;
wire [16:0] \add_34s_34s_34_2_1_U15.top_add_34s_34s_34_2_1_Adder_11_U.u1.s ;
wire [16:0] \add_34s_34s_34_2_1_U15.top_add_34s_34s_34_2_1_Adder_11_U.u2.a ;
wire [16:0] \add_34s_34s_34_2_1_U15.top_add_34s_34s_34_2_1_Adder_11_U.u2.b ;
wire \add_34s_34s_34_2_1_U15.top_add_34s_34s_34_2_1_Adder_11_U.u2.cin ;
wire \add_34s_34s_34_2_1_U15.top_add_34s_34s_34_2_1_Adder_11_U.u2.cout ;
wire [16:0] \add_34s_34s_34_2_1_U15.top_add_34s_34s_34_2_1_Adder_11_U.u2.s ;
wire \add_35s_35s_35_2_1_U10.ce ;
wire \add_35s_35s_35_2_1_U10.clk ;
wire [34:0] \add_35s_35s_35_2_1_U10.din0 ;
wire [34:0] \add_35s_35s_35_2_1_U10.din1 ;
wire [34:0] \add_35s_35s_35_2_1_U10.dout ;
wire \add_35s_35s_35_2_1_U10.reset ;
wire [34:0] \add_35s_35s_35_2_1_U10.top_add_35s_35s_35_2_1_Adder_7_U.a ;
wire [34:0] \add_35s_35s_35_2_1_U10.top_add_35s_35s_35_2_1_Adder_7_U.ain_s0 ;
wire [34:0] \add_35s_35s_35_2_1_U10.top_add_35s_35s_35_2_1_Adder_7_U.b ;
wire [34:0] \add_35s_35s_35_2_1_U10.top_add_35s_35s_35_2_1_Adder_7_U.bin_s0 ;
wire \add_35s_35s_35_2_1_U10.top_add_35s_35s_35_2_1_Adder_7_U.ce ;
wire \add_35s_35s_35_2_1_U10.top_add_35s_35s_35_2_1_Adder_7_U.clk ;
wire \add_35s_35s_35_2_1_U10.top_add_35s_35s_35_2_1_Adder_7_U.facout_s1 ;
wire \add_35s_35s_35_2_1_U10.top_add_35s_35s_35_2_1_Adder_7_U.facout_s2 ;
wire [16:0] \add_35s_35s_35_2_1_U10.top_add_35s_35s_35_2_1_Adder_7_U.fas_s1 ;
wire [17:0] \add_35s_35s_35_2_1_U10.top_add_35s_35s_35_2_1_Adder_7_U.fas_s2 ;
wire \add_35s_35s_35_2_1_U10.top_add_35s_35s_35_2_1_Adder_7_U.reset ;
wire [34:0] \add_35s_35s_35_2_1_U10.top_add_35s_35s_35_2_1_Adder_7_U.s ;
wire [16:0] \add_35s_35s_35_2_1_U10.top_add_35s_35s_35_2_1_Adder_7_U.u1.a ;
wire [16:0] \add_35s_35s_35_2_1_U10.top_add_35s_35s_35_2_1_Adder_7_U.u1.b ;
wire \add_35s_35s_35_2_1_U10.top_add_35s_35s_35_2_1_Adder_7_U.u1.cin ;
wire \add_35s_35s_35_2_1_U10.top_add_35s_35s_35_2_1_Adder_7_U.u1.cout ;
wire [16:0] \add_35s_35s_35_2_1_U10.top_add_35s_35s_35_2_1_Adder_7_U.u1.s ;
wire [17:0] \add_35s_35s_35_2_1_U10.top_add_35s_35s_35_2_1_Adder_7_U.u2.a ;
wire [17:0] \add_35s_35s_35_2_1_U10.top_add_35s_35s_35_2_1_Adder_7_U.u2.b ;
wire \add_35s_35s_35_2_1_U10.top_add_35s_35s_35_2_1_Adder_7_U.u2.cin ;
wire \add_35s_35s_35_2_1_U10.top_add_35s_35s_35_2_1_Adder_7_U.u2.cout ;
wire [17:0] \add_35s_35s_35_2_1_U10.top_add_35s_35s_35_2_1_Adder_7_U.u2.s ;
wire \add_3s_3ns_3_2_1_U13.ce ;
wire \add_3s_3ns_3_2_1_U13.clk ;
wire [2:0] \add_3s_3ns_3_2_1_U13.din0 ;
wire [2:0] \add_3s_3ns_3_2_1_U13.din1 ;
wire [2:0] \add_3s_3ns_3_2_1_U13.dout ;
wire \add_3s_3ns_3_2_1_U13.reset ;
wire [2:0] \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_9_U.a ;
wire [2:0] \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_9_U.ain_s0 ;
wire [2:0] \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_9_U.b ;
wire [2:0] \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_9_U.bin_s0 ;
wire \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_9_U.ce ;
wire \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_9_U.clk ;
wire \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_9_U.facout_s1 ;
wire \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_9_U.facout_s2 ;
wire \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_9_U.fas_s1 ;
wire [1:0] \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_9_U.fas_s2 ;
wire \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_9_U.reset ;
wire [2:0] \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_9_U.s ;
wire \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_9_U.u1.a ;
wire \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_9_U.u1.b ;
wire \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_9_U.u1.cin ;
wire \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_9_U.u1.cout ;
wire \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_9_U.u1.s ;
wire [1:0] \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_9_U.u2.a ;
wire [1:0] \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_9_U.u2.b ;
wire \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_9_U.u2.cin ;
wire \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_9_U.u2.cout ;
wire [1:0] \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_9_U.u2.s ;
wire \add_40s_40s_40_2_1_U7.ce ;
wire \add_40s_40s_40_2_1_U7.clk ;
wire [39:0] \add_40s_40s_40_2_1_U7.din0 ;
wire [39:0] \add_40s_40s_40_2_1_U7.din1 ;
wire [39:0] \add_40s_40s_40_2_1_U7.dout ;
wire \add_40s_40s_40_2_1_U7.reset ;
wire [39:0] \add_40s_40s_40_2_1_U7.top_add_40s_40s_40_2_1_Adder_5_U.a ;
wire [39:0] \add_40s_40s_40_2_1_U7.top_add_40s_40s_40_2_1_Adder_5_U.ain_s0 ;
wire [39:0] \add_40s_40s_40_2_1_U7.top_add_40s_40s_40_2_1_Adder_5_U.b ;
wire [39:0] \add_40s_40s_40_2_1_U7.top_add_40s_40s_40_2_1_Adder_5_U.bin_s0 ;
wire \add_40s_40s_40_2_1_U7.top_add_40s_40s_40_2_1_Adder_5_U.ce ;
wire \add_40s_40s_40_2_1_U7.top_add_40s_40s_40_2_1_Adder_5_U.clk ;
wire \add_40s_40s_40_2_1_U7.top_add_40s_40s_40_2_1_Adder_5_U.facout_s1 ;
wire \add_40s_40s_40_2_1_U7.top_add_40s_40s_40_2_1_Adder_5_U.facout_s2 ;
wire [19:0] \add_40s_40s_40_2_1_U7.top_add_40s_40s_40_2_1_Adder_5_U.fas_s1 ;
wire [19:0] \add_40s_40s_40_2_1_U7.top_add_40s_40s_40_2_1_Adder_5_U.fas_s2 ;
wire \add_40s_40s_40_2_1_U7.top_add_40s_40s_40_2_1_Adder_5_U.reset ;
wire [39:0] \add_40s_40s_40_2_1_U7.top_add_40s_40s_40_2_1_Adder_5_U.s ;
wire [19:0] \add_40s_40s_40_2_1_U7.top_add_40s_40s_40_2_1_Adder_5_U.u1.a ;
wire [19:0] \add_40s_40s_40_2_1_U7.top_add_40s_40s_40_2_1_Adder_5_U.u1.b ;
wire \add_40s_40s_40_2_1_U7.top_add_40s_40s_40_2_1_Adder_5_U.u1.cin ;
wire \add_40s_40s_40_2_1_U7.top_add_40s_40s_40_2_1_Adder_5_U.u1.cout ;
wire [19:0] \add_40s_40s_40_2_1_U7.top_add_40s_40s_40_2_1_Adder_5_U.u1.s ;
wire [19:0] \add_40s_40s_40_2_1_U7.top_add_40s_40s_40_2_1_Adder_5_U.u2.a ;
wire [19:0] \add_40s_40s_40_2_1_U7.top_add_40s_40s_40_2_1_Adder_5_U.u2.b ;
wire \add_40s_40s_40_2_1_U7.top_add_40s_40s_40_2_1_Adder_5_U.u2.cin ;
wire \add_40s_40s_40_2_1_U7.top_add_40s_40s_40_2_1_Adder_5_U.u2.cout ;
wire [19:0] \add_40s_40s_40_2_1_U7.top_add_40s_40s_40_2_1_Adder_5_U.u2.s ;
wire and_ln365_fu_371_p2;
wire ap_CS_fsm_state1;
wire ap_CS_fsm_state10;
wire ap_CS_fsm_state11;
wire ap_CS_fsm_state12;
wire ap_CS_fsm_state13;
wire ap_CS_fsm_state14;
wire ap_CS_fsm_state15;
wire ap_CS_fsm_state16;
wire ap_CS_fsm_state17;
wire ap_CS_fsm_state18;
wire ap_CS_fsm_state19;
wire ap_CS_fsm_state2;
wire ap_CS_fsm_state20;
wire ap_CS_fsm_state21;
wire ap_CS_fsm_state22;
wire ap_CS_fsm_state23;
wire ap_CS_fsm_state24;
wire ap_CS_fsm_state25;
wire ap_CS_fsm_state26;
wire ap_CS_fsm_state27;
wire ap_CS_fsm_state28;
wire ap_CS_fsm_state29;
wire ap_CS_fsm_state3;
wire ap_CS_fsm_state30;
wire ap_CS_fsm_state31;
wire ap_CS_fsm_state32;
wire ap_CS_fsm_state4;
wire ap_CS_fsm_state5;
wire ap_CS_fsm_state6;
wire ap_CS_fsm_state7;
wire ap_CS_fsm_state8;
wire ap_CS_fsm_state9;
wire [31:0] ap_NS_fsm;
wire ap_clk;
wire ap_done;
wire ap_idle;
wire ap_ready;
wire ap_rst;
wire ap_start;
wire empty_fu_312_p1;
wire [16:0] grp_fu_221_p0;
wire [16:0] grp_fu_221_p1;
wire [16:0] grp_fu_221_p2;
wire [9:0] grp_fu_247_p2;
wire [10:0] grp_fu_290_p0;
wire [10:0] grp_fu_290_p2;
wire [9:0] grp_fu_306_p0;
wire [9:0] grp_fu_306_p1;
wire [9:0] grp_fu_306_p2;
wire [10:0] grp_fu_339_p0;
wire [10:0] grp_fu_339_p2;
wire [10:0] grp_fu_379_p0;
wire [10:0] grp_fu_379_p2;
wire [39:0] grp_fu_438_p0;
wire [39:0] grp_fu_438_p1;
wire [39:0] grp_fu_438_p2;
wire [31:0] grp_fu_459_p2;
wire [31:0] grp_fu_491_p2;
wire [34:0] grp_fu_510_p0;
wire [34:0] grp_fu_510_p1;
wire [34:0] grp_fu_510_p2;
wire [31:0] grp_fu_536_p2;
wire [31:0] grp_fu_575_p1;
wire [31:0] grp_fu_575_p2;
wire [2:0] grp_fu_580_p0;
wire [2:0] grp_fu_580_p2;
wire [31:0] grp_fu_612_p0;
wire [31:0] grp_fu_612_p2;
wire [33:0] grp_fu_657_p0;
wire [33:0] grp_fu_657_p1;
wire [33:0] grp_fu_657_p2;
wire [31:0] grp_fu_673_p2;
wire icmp_ln785_fu_593_p2;
wire icmp_ln851_1_fu_444_p2;
wire icmp_ln851_2_fu_520_p2;
wire icmp_ln851_fu_231_p2;
wire lhs_V_fu_348_p2;
wire [14:0] lhs_fu_205_p3;
wire [7:0] op_0;
wire [15:0] op_1;
wire [3:0] op_10;
wire op_11;
wire [7:0] op_13_V_fu_413_p3;
wire op_14;
wire [7:0] op_15;
wire [3:0] op_16;
wire [1:0] op_17;
wire [1:0] op_19_V_fu_635_p3;
wire op_2;
wire [1:0] op_3;
wire [31:0] op_31;
wire op_31_ap_vld;
wire [1:0] op_4;
wire [1:0] op_8;
wire or_ln384_fu_631_p1;
wire or_ln384_fu_631_p2;
wire or_ln785_1_fu_585_p1;
wire [1:0] or_ln785_1_fu_585_p3;
wire or_ln785_fu_344_p2;
wire overflow_fu_604_p2;
wire [7:0] p_Result_3_fu_397_p4;
wire p_Result_4_fu_464_p3;
wire p_Result_5_fu_541_p3;
wire p_Result_6_fu_678_p3;
wire p_Result_7_fu_330_p2;
wire p_Result_s_fu_252_p3;
wire [7:0] p_Val2_1_fu_384_p3;
wire [6:0] p_Val2_3_fu_391_p2;
wire p_Val2_5_fu_617_p0;
wire [1:0] p_Val2_5_fu_617_p3;
wire r_fu_316_p2;
wire [9:0] ret_V_13_fu_264_p3;
wire [31:0] ret_V_17_fu_476_p3;
wire [31:0] ret_V_19_fu_553_p3;
wire [1:0] ret_fu_271_p3;
wire [33:0] rhs_4_fu_499_p3;
wire [32:0] rhs_6_fu_646_p3;
wire [10:0] select_ln1192_fu_279_p3;
wire [1:0] select_ln384_fu_624_p3;
wire [2:0] select_ln69_1_fu_560_p3;
wire [31:0] select_ln69_fu_483_p3;
wire [7:0] select_ln785_fu_406_p3;
wire [31:0] select_ln850_1_fu_471_p3;
wire [31:0] select_ln850_2_fu_548_p3;
wire [31:0] select_ln850_3_fu_688_p3;
wire [9:0] select_ln850_fu_259_p3;
wire [7:0] sext_ln69_fu_295_p1;
wire [7:0] sext_ln703_2_fu_495_p0;
wire [15:0] sext_ln703_fu_217_p0;
wire tmp_1_fu_353_p3;
wire [17:0] tmp_3_fu_427_p3;
wire tmp_fu_322_p3;
wire [6:0] trunc_ln851_1_fu_420_p1;
wire [7:0] trunc_ln851_2_fu_516_p0;
wire [1:0] trunc_ln851_2_fu_516_p1;
wire trunc_ln851_3_fu_685_p1;
wire [15:0] trunc_ln851_fu_227_p0;
wire [6:0] trunc_ln851_fu_227_p1;
wire xor_ln365_1_fu_366_p2;
wire xor_ln365_fu_360_p2;
wire xor_ln785_fu_599_p0;
wire xor_ln785_fu_599_p2;


assign _043_ = icmp_ln851_2_reg_905 & ap_CS_fsm[21];
assign _044_ = ap_CS_fsm[14] & icmp_ln851_1_reg_858;
assign _045_ = _048_ & ap_CS_fsm[3];
assign _046_ = _049_ & ap_CS_fsm[0];
assign _047_ = ap_start & ap_CS_fsm[0];
assign and_ln365_fu_371_p2 = xor_ln365_1_fu_366_p2 & or_ln785_reg_807;
assign overflow_fu_604_p2 = xor_ln785_fu_599_p2 & icmp_ln785_reg_954;
assign p_Result_7_fu_330_p2 = ~ op_8[1];
assign lhs_V_fu_348_p2 = ~ op_2;
assign xor_ln785_fu_599_p2 = ~ op_11;
assign r_fu_316_p2 = ~ op_8[0];
assign _048_ = ~ icmp_ln851_reg_712;
assign _049_ = ~ ap_start;
assign _050_ = ! op_1[6:0];
always @(posedge \add_10ns_10ns_10_2_1_U2.top_add_10ns_10ns_10_2_1_Adder_1_U.clk )
\add_10ns_10ns_10_2_1_U2.top_add_10ns_10ns_10_2_1_Adder_1_U.bin_s1  <= _052_;
always @(posedge \add_10ns_10ns_10_2_1_U2.top_add_10ns_10ns_10_2_1_Adder_1_U.clk )
\add_10ns_10ns_10_2_1_U2.top_add_10ns_10ns_10_2_1_Adder_1_U.ain_s1  <= _051_;
always @(posedge \add_10ns_10ns_10_2_1_U2.top_add_10ns_10ns_10_2_1_Adder_1_U.clk )
\add_10ns_10ns_10_2_1_U2.top_add_10ns_10ns_10_2_1_Adder_1_U.sum_s1  <= _054_;
always @(posedge \add_10ns_10ns_10_2_1_U2.top_add_10ns_10ns_10_2_1_Adder_1_U.clk )
\add_10ns_10ns_10_2_1_U2.top_add_10ns_10ns_10_2_1_Adder_1_U.carry_s1  <= _053_;
assign _052_ = \add_10ns_10ns_10_2_1_U2.top_add_10ns_10ns_10_2_1_Adder_1_U.ce  ? \add_10ns_10ns_10_2_1_U2.top_add_10ns_10ns_10_2_1_Adder_1_U.b [9:5] : \add_10ns_10ns_10_2_1_U2.top_add_10ns_10ns_10_2_1_Adder_1_U.bin_s1 ;
assign _051_ = \add_10ns_10ns_10_2_1_U2.top_add_10ns_10ns_10_2_1_Adder_1_U.ce  ? \add_10ns_10ns_10_2_1_U2.top_add_10ns_10ns_10_2_1_Adder_1_U.a [9:5] : \add_10ns_10ns_10_2_1_U2.top_add_10ns_10ns_10_2_1_Adder_1_U.ain_s1 ;
assign _053_ = \add_10ns_10ns_10_2_1_U2.top_add_10ns_10ns_10_2_1_Adder_1_U.ce  ? \add_10ns_10ns_10_2_1_U2.top_add_10ns_10ns_10_2_1_Adder_1_U.facout_s1  : \add_10ns_10ns_10_2_1_U2.top_add_10ns_10ns_10_2_1_Adder_1_U.carry_s1 ;
assign _054_ = \add_10ns_10ns_10_2_1_U2.top_add_10ns_10ns_10_2_1_Adder_1_U.ce  ? \add_10ns_10ns_10_2_1_U2.top_add_10ns_10ns_10_2_1_Adder_1_U.fas_s1  : \add_10ns_10ns_10_2_1_U2.top_add_10ns_10ns_10_2_1_Adder_1_U.sum_s1 ;
assign _055_ = \add_10ns_10ns_10_2_1_U2.top_add_10ns_10ns_10_2_1_Adder_1_U.u1.a  + \add_10ns_10ns_10_2_1_U2.top_add_10ns_10ns_10_2_1_Adder_1_U.u1.b ;
assign { \add_10ns_10ns_10_2_1_U2.top_add_10ns_10ns_10_2_1_Adder_1_U.u1.cout , \add_10ns_10ns_10_2_1_U2.top_add_10ns_10ns_10_2_1_Adder_1_U.u1.s  } = _055_ + \add_10ns_10ns_10_2_1_U2.top_add_10ns_10ns_10_2_1_Adder_1_U.u1.cin ;
assign _056_ = \add_10ns_10ns_10_2_1_U2.top_add_10ns_10ns_10_2_1_Adder_1_U.u2.a  + \add_10ns_10ns_10_2_1_U2.top_add_10ns_10ns_10_2_1_Adder_1_U.u2.b ;
assign { \add_10ns_10ns_10_2_1_U2.top_add_10ns_10ns_10_2_1_Adder_1_U.u2.cout , \add_10ns_10ns_10_2_1_U2.top_add_10ns_10ns_10_2_1_Adder_1_U.u2.s  } = _056_ + \add_10ns_10ns_10_2_1_U2.top_add_10ns_10ns_10_2_1_Adder_1_U.u2.cin ;
always @(posedge \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.clk )
\add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.bin_s1  <= _058_;
always @(posedge \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.clk )
\add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.ain_s1  <= _057_;
always @(posedge \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.clk )
\add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.sum_s1  <= _060_;
always @(posedge \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.clk )
\add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.carry_s1  <= _059_;
assign _058_ = \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.ce  ? \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.b [9:5] : \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.bin_s1 ;
assign _057_ = \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.ce  ? \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.a [9:5] : \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.ain_s1 ;
assign _059_ = \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.ce  ? \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.facout_s1  : \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.carry_s1 ;
assign _060_ = \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.ce  ? \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.fas_s1  : \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.sum_s1 ;
assign _061_ = \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.u1.a  + \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.u1.b ;
assign { \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.u1.cout , \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.u1.s  } = _061_ + \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.u1.cin ;
assign _062_ = \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.u2.a  + \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.u2.b ;
assign { \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.u2.cout , \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.u2.s  } = _062_ + \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.u2.cin ;
always @(posedge \add_11ns_11ns_11_2_1_U6.top_add_11ns_11ns_11_2_1_Adder_4_U.clk )
\add_11ns_11ns_11_2_1_U6.top_add_11ns_11ns_11_2_1_Adder_4_U.bin_s1  <= _064_;
always @(posedge \add_11ns_11ns_11_2_1_U6.top_add_11ns_11ns_11_2_1_Adder_4_U.clk )
\add_11ns_11ns_11_2_1_U6.top_add_11ns_11ns_11_2_1_Adder_4_U.ain_s1  <= _063_;
always @(posedge \add_11ns_11ns_11_2_1_U6.top_add_11ns_11ns_11_2_1_Adder_4_U.clk )
\add_11ns_11ns_11_2_1_U6.top_add_11ns_11ns_11_2_1_Adder_4_U.sum_s1  <= _066_;
always @(posedge \add_11ns_11ns_11_2_1_U6.top_add_11ns_11ns_11_2_1_Adder_4_U.clk )
\add_11ns_11ns_11_2_1_U6.top_add_11ns_11ns_11_2_1_Adder_4_U.carry_s1  <= _065_;
assign _064_ = \add_11ns_11ns_11_2_1_U6.top_add_11ns_11ns_11_2_1_Adder_4_U.ce  ? \add_11ns_11ns_11_2_1_U6.top_add_11ns_11ns_11_2_1_Adder_4_U.b [10:5] : \add_11ns_11ns_11_2_1_U6.top_add_11ns_11ns_11_2_1_Adder_4_U.bin_s1 ;
assign _063_ = \add_11ns_11ns_11_2_1_U6.top_add_11ns_11ns_11_2_1_Adder_4_U.ce  ? \add_11ns_11ns_11_2_1_U6.top_add_11ns_11ns_11_2_1_Adder_4_U.a [10:5] : \add_11ns_11ns_11_2_1_U6.top_add_11ns_11ns_11_2_1_Adder_4_U.ain_s1 ;
assign _065_ = \add_11ns_11ns_11_2_1_U6.top_add_11ns_11ns_11_2_1_Adder_4_U.ce  ? \add_11ns_11ns_11_2_1_U6.top_add_11ns_11ns_11_2_1_Adder_4_U.facout_s1  : \add_11ns_11ns_11_2_1_U6.top_add_11ns_11ns_11_2_1_Adder_4_U.carry_s1 ;
assign _066_ = \add_11ns_11ns_11_2_1_U6.top_add_11ns_11ns_11_2_1_Adder_4_U.ce  ? \add_11ns_11ns_11_2_1_U6.top_add_11ns_11ns_11_2_1_Adder_4_U.fas_s1  : \add_11ns_11ns_11_2_1_U6.top_add_11ns_11ns_11_2_1_Adder_4_U.sum_s1 ;
assign _067_ = \add_11ns_11ns_11_2_1_U6.top_add_11ns_11ns_11_2_1_Adder_4_U.u1.a  + \add_11ns_11ns_11_2_1_U6.top_add_11ns_11ns_11_2_1_Adder_4_U.u1.b ;
assign { \add_11ns_11ns_11_2_1_U6.top_add_11ns_11ns_11_2_1_Adder_4_U.u1.cout , \add_11ns_11ns_11_2_1_U6.top_add_11ns_11ns_11_2_1_Adder_4_U.u1.s  } = _067_ + \add_11ns_11ns_11_2_1_U6.top_add_11ns_11ns_11_2_1_Adder_4_U.u1.cin ;
assign _068_ = \add_11ns_11ns_11_2_1_U6.top_add_11ns_11ns_11_2_1_Adder_4_U.u2.a  + \add_11ns_11ns_11_2_1_U6.top_add_11ns_11ns_11_2_1_Adder_4_U.u2.b ;
assign { \add_11ns_11ns_11_2_1_U6.top_add_11ns_11ns_11_2_1_Adder_4_U.u2.cout , \add_11ns_11ns_11_2_1_U6.top_add_11ns_11ns_11_2_1_Adder_4_U.u2.s  } = _068_ + \add_11ns_11ns_11_2_1_U6.top_add_11ns_11ns_11_2_1_Adder_4_U.u2.cin ;
always @(posedge \add_11s_11ns_11_2_1_U3.top_add_11s_11ns_11_2_1_Adder_2_U.clk )
\add_11s_11ns_11_2_1_U3.top_add_11s_11ns_11_2_1_Adder_2_U.bin_s1  <= _070_;
always @(posedge \add_11s_11ns_11_2_1_U3.top_add_11s_11ns_11_2_1_Adder_2_U.clk )
\add_11s_11ns_11_2_1_U3.top_add_11s_11ns_11_2_1_Adder_2_U.ain_s1  <= _069_;
always @(posedge \add_11s_11ns_11_2_1_U3.top_add_11s_11ns_11_2_1_Adder_2_U.clk )
\add_11s_11ns_11_2_1_U3.top_add_11s_11ns_11_2_1_Adder_2_U.sum_s1  <= _072_;
always @(posedge \add_11s_11ns_11_2_1_U3.top_add_11s_11ns_11_2_1_Adder_2_U.clk )
\add_11s_11ns_11_2_1_U3.top_add_11s_11ns_11_2_1_Adder_2_U.carry_s1  <= _071_;
assign _070_ = \add_11s_11ns_11_2_1_U3.top_add_11s_11ns_11_2_1_Adder_2_U.ce  ? \add_11s_11ns_11_2_1_U3.top_add_11s_11ns_11_2_1_Adder_2_U.b [10:5] : \add_11s_11ns_11_2_1_U3.top_add_11s_11ns_11_2_1_Adder_2_U.bin_s1 ;
assign _069_ = \add_11s_11ns_11_2_1_U3.top_add_11s_11ns_11_2_1_Adder_2_U.ce  ? \add_11s_11ns_11_2_1_U3.top_add_11s_11ns_11_2_1_Adder_2_U.a [10:5] : \add_11s_11ns_11_2_1_U3.top_add_11s_11ns_11_2_1_Adder_2_U.ain_s1 ;
assign _071_ = \add_11s_11ns_11_2_1_U3.top_add_11s_11ns_11_2_1_Adder_2_U.ce  ? \add_11s_11ns_11_2_1_U3.top_add_11s_11ns_11_2_1_Adder_2_U.facout_s1  : \add_11s_11ns_11_2_1_U3.top_add_11s_11ns_11_2_1_Adder_2_U.carry_s1 ;
assign _072_ = \add_11s_11ns_11_2_1_U3.top_add_11s_11ns_11_2_1_Adder_2_U.ce  ? \add_11s_11ns_11_2_1_U3.top_add_11s_11ns_11_2_1_Adder_2_U.fas_s1  : \add_11s_11ns_11_2_1_U3.top_add_11s_11ns_11_2_1_Adder_2_U.sum_s1 ;
assign _073_ = \add_11s_11ns_11_2_1_U3.top_add_11s_11ns_11_2_1_Adder_2_U.u1.a  + \add_11s_11ns_11_2_1_U3.top_add_11s_11ns_11_2_1_Adder_2_U.u1.b ;
assign { \add_11s_11ns_11_2_1_U3.top_add_11s_11ns_11_2_1_Adder_2_U.u1.cout , \add_11s_11ns_11_2_1_U3.top_add_11s_11ns_11_2_1_Adder_2_U.u1.s  } = _073_ + \add_11s_11ns_11_2_1_U3.top_add_11s_11ns_11_2_1_Adder_2_U.u1.cin ;
assign _074_ = \add_11s_11ns_11_2_1_U3.top_add_11s_11ns_11_2_1_Adder_2_U.u2.a  + \add_11s_11ns_11_2_1_U3.top_add_11s_11ns_11_2_1_Adder_2_U.u2.b ;
assign { \add_11s_11ns_11_2_1_U3.top_add_11s_11ns_11_2_1_Adder_2_U.u2.cout , \add_11s_11ns_11_2_1_U3.top_add_11s_11ns_11_2_1_Adder_2_U.u2.s  } = _074_ + \add_11s_11ns_11_2_1_U3.top_add_11s_11ns_11_2_1_Adder_2_U.u2.cin ;
always @(posedge \add_11s_11ns_11_2_1_U5.top_add_11s_11ns_11_2_1_Adder_2_U.clk )
\add_11s_11ns_11_2_1_U5.top_add_11s_11ns_11_2_1_Adder_2_U.bin_s1  <= _076_;
always @(posedge \add_11s_11ns_11_2_1_U5.top_add_11s_11ns_11_2_1_Adder_2_U.clk )
\add_11s_11ns_11_2_1_U5.top_add_11s_11ns_11_2_1_Adder_2_U.ain_s1  <= _075_;
always @(posedge \add_11s_11ns_11_2_1_U5.top_add_11s_11ns_11_2_1_Adder_2_U.clk )
\add_11s_11ns_11_2_1_U5.top_add_11s_11ns_11_2_1_Adder_2_U.sum_s1  <= _078_;
always @(posedge \add_11s_11ns_11_2_1_U5.top_add_11s_11ns_11_2_1_Adder_2_U.clk )
\add_11s_11ns_11_2_1_U5.top_add_11s_11ns_11_2_1_Adder_2_U.carry_s1  <= _077_;
assign _076_ = \add_11s_11ns_11_2_1_U5.top_add_11s_11ns_11_2_1_Adder_2_U.ce  ? \add_11s_11ns_11_2_1_U5.top_add_11s_11ns_11_2_1_Adder_2_U.b [10:5] : \add_11s_11ns_11_2_1_U5.top_add_11s_11ns_11_2_1_Adder_2_U.bin_s1 ;
assign _075_ = \add_11s_11ns_11_2_1_U5.top_add_11s_11ns_11_2_1_Adder_2_U.ce  ? \add_11s_11ns_11_2_1_U5.top_add_11s_11ns_11_2_1_Adder_2_U.a [10:5] : \add_11s_11ns_11_2_1_U5.top_add_11s_11ns_11_2_1_Adder_2_U.ain_s1 ;
assign _077_ = \add_11s_11ns_11_2_1_U5.top_add_11s_11ns_11_2_1_Adder_2_U.ce  ? \add_11s_11ns_11_2_1_U5.top_add_11s_11ns_11_2_1_Adder_2_U.facout_s1  : \add_11s_11ns_11_2_1_U5.top_add_11s_11ns_11_2_1_Adder_2_U.carry_s1 ;
assign _078_ = \add_11s_11ns_11_2_1_U5.top_add_11s_11ns_11_2_1_Adder_2_U.ce  ? \add_11s_11ns_11_2_1_U5.top_add_11s_11ns_11_2_1_Adder_2_U.fas_s1  : \add_11s_11ns_11_2_1_U5.top_add_11s_11ns_11_2_1_Adder_2_U.sum_s1 ;
assign _079_ = \add_11s_11ns_11_2_1_U5.top_add_11s_11ns_11_2_1_Adder_2_U.u1.a  + \add_11s_11ns_11_2_1_U5.top_add_11s_11ns_11_2_1_Adder_2_U.u1.b ;
assign { \add_11s_11ns_11_2_1_U5.top_add_11s_11ns_11_2_1_Adder_2_U.u1.cout , \add_11s_11ns_11_2_1_U5.top_add_11s_11ns_11_2_1_Adder_2_U.u1.s  } = _079_ + \add_11s_11ns_11_2_1_U5.top_add_11s_11ns_11_2_1_Adder_2_U.u1.cin ;
assign _080_ = \add_11s_11ns_11_2_1_U5.top_add_11s_11ns_11_2_1_Adder_2_U.u2.a  + \add_11s_11ns_11_2_1_U5.top_add_11s_11ns_11_2_1_Adder_2_U.u2.b ;
assign { \add_11s_11ns_11_2_1_U5.top_add_11s_11ns_11_2_1_Adder_2_U.u2.cout , \add_11s_11ns_11_2_1_U5.top_add_11s_11ns_11_2_1_Adder_2_U.u2.s  } = _080_ + \add_11s_11ns_11_2_1_U5.top_add_11s_11ns_11_2_1_Adder_2_U.u2.cin ;
always @(posedge \add_17s_17s_17_2_1_U1.top_add_17s_17s_17_2_1_Adder_0_U.clk )
\add_17s_17s_17_2_1_U1.top_add_17s_17s_17_2_1_Adder_0_U.bin_s1  <= _082_;
always @(posedge \add_17s_17s_17_2_1_U1.top_add_17s_17s_17_2_1_Adder_0_U.clk )
\add_17s_17s_17_2_1_U1.top_add_17s_17s_17_2_1_Adder_0_U.ain_s1  <= _081_;
always @(posedge \add_17s_17s_17_2_1_U1.top_add_17s_17s_17_2_1_Adder_0_U.clk )
\add_17s_17s_17_2_1_U1.top_add_17s_17s_17_2_1_Adder_0_U.sum_s1  <= _084_;
always @(posedge \add_17s_17s_17_2_1_U1.top_add_17s_17s_17_2_1_Adder_0_U.clk )
\add_17s_17s_17_2_1_U1.top_add_17s_17s_17_2_1_Adder_0_U.carry_s1  <= _083_;
assign _082_ = \add_17s_17s_17_2_1_U1.top_add_17s_17s_17_2_1_Adder_0_U.ce  ? \add_17s_17s_17_2_1_U1.top_add_17s_17s_17_2_1_Adder_0_U.b [16:8] : \add_17s_17s_17_2_1_U1.top_add_17s_17s_17_2_1_Adder_0_U.bin_s1 ;
assign _081_ = \add_17s_17s_17_2_1_U1.top_add_17s_17s_17_2_1_Adder_0_U.ce  ? \add_17s_17s_17_2_1_U1.top_add_17s_17s_17_2_1_Adder_0_U.a [16:8] : \add_17s_17s_17_2_1_U1.top_add_17s_17s_17_2_1_Adder_0_U.ain_s1 ;
assign _083_ = \add_17s_17s_17_2_1_U1.top_add_17s_17s_17_2_1_Adder_0_U.ce  ? \add_17s_17s_17_2_1_U1.top_add_17s_17s_17_2_1_Adder_0_U.facout_s1  : \add_17s_17s_17_2_1_U1.top_add_17s_17s_17_2_1_Adder_0_U.carry_s1 ;
assign _084_ = \add_17s_17s_17_2_1_U1.top_add_17s_17s_17_2_1_Adder_0_U.ce  ? \add_17s_17s_17_2_1_U1.top_add_17s_17s_17_2_1_Adder_0_U.fas_s1  : \add_17s_17s_17_2_1_U1.top_add_17s_17s_17_2_1_Adder_0_U.sum_s1 ;
assign _085_ = \add_17s_17s_17_2_1_U1.top_add_17s_17s_17_2_1_Adder_0_U.u1.a  + \add_17s_17s_17_2_1_U1.top_add_17s_17s_17_2_1_Adder_0_U.u1.b ;
assign { \add_17s_17s_17_2_1_U1.top_add_17s_17s_17_2_1_Adder_0_U.u1.cout , \add_17s_17s_17_2_1_U1.top_add_17s_17s_17_2_1_Adder_0_U.u1.s  } = _085_ + \add_17s_17s_17_2_1_U1.top_add_17s_17s_17_2_1_Adder_0_U.u1.cin ;
assign _086_ = \add_17s_17s_17_2_1_U1.top_add_17s_17s_17_2_1_Adder_0_U.u2.a  + \add_17s_17s_17_2_1_U1.top_add_17s_17s_17_2_1_Adder_0_U.u2.b ;
assign { \add_17s_17s_17_2_1_U1.top_add_17s_17s_17_2_1_Adder_0_U.u2.cout , \add_17s_17s_17_2_1_U1.top_add_17s_17s_17_2_1_Adder_0_U.u2.s  } = _086_ + \add_17s_17s_17_2_1_U1.top_add_17s_17s_17_2_1_Adder_0_U.u2.cin ;
always @(posedge \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_6_U.clk )
\add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s1  <= _088_;
always @(posedge \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_6_U.clk )
\add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s1  <= _087_;
always @(posedge \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_6_U.clk )
\add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_6_U.sum_s1  <= _090_;
always @(posedge \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_6_U.clk )
\add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_6_U.carry_s1  <= _089_;
assign _088_ = \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  ? \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_6_U.b [31:16] : \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s1 ;
assign _087_ = \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  ? \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_6_U.a [31:16] : \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s1 ;
assign _089_ = \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  ? \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s1  : \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_6_U.carry_s1 ;
assign _090_ = \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  ? \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s1  : \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_6_U.sum_s1 ;
assign _091_ = \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.a  + \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.b ;
assign { \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cout , \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.s  } = _091_ + \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cin ;
assign _092_ = \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.a  + \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.b ;
assign { \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cout , \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.s  } = _092_ + \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cin ;
always @(posedge \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.clk )
\add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s1  <= _094_;
always @(posedge \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.clk )
\add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s1  <= _093_;
always @(posedge \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.clk )
\add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.sum_s1  <= _096_;
always @(posedge \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.clk )
\add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.carry_s1  <= _095_;
assign _094_ = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  ? \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.b [31:16] : \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s1 ;
assign _093_ = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  ? \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.a [31:16] : \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s1 ;
assign _095_ = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  ? \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s1  : \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.carry_s1 ;
assign _096_ = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  ? \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s1  : \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.sum_s1 ;
assign _097_ = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.a  + \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.b ;
assign { \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cout , \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.s  } = _097_ + \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cin ;
assign _098_ = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.a  + \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.b ;
assign { \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cout , \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.s  } = _098_ + \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cin ;
always @(posedge \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.clk )
\add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s1  <= _100_;
always @(posedge \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.clk )
\add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s1  <= _099_;
always @(posedge \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.clk )
\add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.sum_s1  <= _102_;
always @(posedge \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.clk )
\add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.carry_s1  <= _101_;
assign _100_ = \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  ? \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.b [31:16] : \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s1 ;
assign _099_ = \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  ? \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.a [31:16] : \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s1 ;
assign _101_ = \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  ? \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s1  : \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.carry_s1 ;
assign _102_ = \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  ? \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s1  : \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.sum_s1 ;
assign _103_ = \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.a  + \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.b ;
assign { \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cout , \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.s  } = _103_ + \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cin ;
assign _104_ = \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.a  + \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.b ;
assign { \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cout , \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.s  } = _104_ + \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cin ;
always @(posedge \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.clk )
\add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s1  <= _106_;
always @(posedge \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.clk )
\add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s1  <= _105_;
always @(posedge \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.clk )
\add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.sum_s1  <= _108_;
always @(posedge \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.clk )
\add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.carry_s1  <= _107_;
assign _106_ = \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  ? \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.b [31:16] : \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s1 ;
assign _105_ = \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  ? \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.a [31:16] : \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s1 ;
assign _107_ = \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  ? \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s1  : \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.carry_s1 ;
assign _108_ = \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  ? \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s1  : \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.sum_s1 ;
assign _109_ = \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.a  + \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.b ;
assign { \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cout , \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.s  } = _109_ + \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cin ;
assign _110_ = \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.a  + \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.b ;
assign { \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cout , \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.s  } = _110_ + \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cin ;
always @(posedge \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.clk )
\add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.bin_s1  <= _112_;
always @(posedge \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.clk )
\add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.ain_s1  <= _111_;
always @(posedge \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.clk )
\add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.sum_s1  <= _114_;
always @(posedge \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.clk )
\add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.carry_s1  <= _113_;
assign _112_ = \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.ce  ? \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.b [31:16] : \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.bin_s1 ;
assign _111_ = \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.ce  ? \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.a [31:16] : \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.ain_s1 ;
assign _113_ = \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.ce  ? \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.facout_s1  : \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.carry_s1 ;
assign _114_ = \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.ce  ? \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.fas_s1  : \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.sum_s1 ;
assign _115_ = \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.u1.a  + \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.u1.b ;
assign { \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.u1.cout , \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.u1.s  } = _115_ + \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.u1.cin ;
assign _116_ = \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.u2.a  + \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.u2.b ;
assign { \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.u2.cout , \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.u2.s  } = _116_ + \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.u2.cin ;
always @(posedge \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_10_U.clk )
\add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_10_U.bin_s1  <= _118_;
always @(posedge \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_10_U.clk )
\add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_10_U.ain_s1  <= _117_;
always @(posedge \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_10_U.clk )
\add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_10_U.sum_s1  <= _120_;
always @(posedge \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_10_U.clk )
\add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_10_U.carry_s1  <= _119_;
assign _118_ = \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_10_U.ce  ? \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_10_U.b [31:16] : \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_10_U.bin_s1 ;
assign _117_ = \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_10_U.ce  ? \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_10_U.a [31:16] : \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_10_U.ain_s1 ;
assign _119_ = \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_10_U.ce  ? \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_10_U.facout_s1  : \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_10_U.carry_s1 ;
assign _120_ = \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_10_U.ce  ? \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_10_U.fas_s1  : \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_10_U.sum_s1 ;
assign _121_ = \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_10_U.u1.a  + \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_10_U.u1.b ;
assign { \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_10_U.u1.cout , \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_10_U.u1.s  } = _121_ + \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_10_U.u1.cin ;
assign _122_ = \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_10_U.u2.a  + \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_10_U.u2.b ;
assign { \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_10_U.u2.cout , \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_10_U.u2.s  } = _122_ + \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_10_U.u2.cin ;
always @(posedge \add_34s_34s_34_2_1_U15.top_add_34s_34s_34_2_1_Adder_11_U.clk )
\add_34s_34s_34_2_1_U15.top_add_34s_34s_34_2_1_Adder_11_U.bin_s1  <= _124_;
always @(posedge \add_34s_34s_34_2_1_U15.top_add_34s_34s_34_2_1_Adder_11_U.clk )
\add_34s_34s_34_2_1_U15.top_add_34s_34s_34_2_1_Adder_11_U.ain_s1  <= _123_;
always @(posedge \add_34s_34s_34_2_1_U15.top_add_34s_34s_34_2_1_Adder_11_U.clk )
\add_34s_34s_34_2_1_U15.top_add_34s_34s_34_2_1_Adder_11_U.sum_s1  <= _126_;
always @(posedge \add_34s_34s_34_2_1_U15.top_add_34s_34s_34_2_1_Adder_11_U.clk )
\add_34s_34s_34_2_1_U15.top_add_34s_34s_34_2_1_Adder_11_U.carry_s1  <= _125_;
assign _124_ = \add_34s_34s_34_2_1_U15.top_add_34s_34s_34_2_1_Adder_11_U.ce  ? \add_34s_34s_34_2_1_U15.top_add_34s_34s_34_2_1_Adder_11_U.b [33:17] : \add_34s_34s_34_2_1_U15.top_add_34s_34s_34_2_1_Adder_11_U.bin_s1 ;
assign _123_ = \add_34s_34s_34_2_1_U15.top_add_34s_34s_34_2_1_Adder_11_U.ce  ? \add_34s_34s_34_2_1_U15.top_add_34s_34s_34_2_1_Adder_11_U.a [33:17] : \add_34s_34s_34_2_1_U15.top_add_34s_34s_34_2_1_Adder_11_U.ain_s1 ;
assign _125_ = \add_34s_34s_34_2_1_U15.top_add_34s_34s_34_2_1_Adder_11_U.ce  ? \add_34s_34s_34_2_1_U15.top_add_34s_34s_34_2_1_Adder_11_U.facout_s1  : \add_34s_34s_34_2_1_U15.top_add_34s_34s_34_2_1_Adder_11_U.carry_s1 ;
assign _126_ = \add_34s_34s_34_2_1_U15.top_add_34s_34s_34_2_1_Adder_11_U.ce  ? \add_34s_34s_34_2_1_U15.top_add_34s_34s_34_2_1_Adder_11_U.fas_s1  : \add_34s_34s_34_2_1_U15.top_add_34s_34s_34_2_1_Adder_11_U.sum_s1 ;
assign _127_ = \add_34s_34s_34_2_1_U15.top_add_34s_34s_34_2_1_Adder_11_U.u1.a  + \add_34s_34s_34_2_1_U15.top_add_34s_34s_34_2_1_Adder_11_U.u1.b ;
assign { \add_34s_34s_34_2_1_U15.top_add_34s_34s_34_2_1_Adder_11_U.u1.cout , \add_34s_34s_34_2_1_U15.top_add_34s_34s_34_2_1_Adder_11_U.u1.s  } = _127_ + \add_34s_34s_34_2_1_U15.top_add_34s_34s_34_2_1_Adder_11_U.u1.cin ;
assign _128_ = \add_34s_34s_34_2_1_U15.top_add_34s_34s_34_2_1_Adder_11_U.u2.a  + \add_34s_34s_34_2_1_U15.top_add_34s_34s_34_2_1_Adder_11_U.u2.b ;
assign { \add_34s_34s_34_2_1_U15.top_add_34s_34s_34_2_1_Adder_11_U.u2.cout , \add_34s_34s_34_2_1_U15.top_add_34s_34s_34_2_1_Adder_11_U.u2.s  } = _128_ + \add_34s_34s_34_2_1_U15.top_add_34s_34s_34_2_1_Adder_11_U.u2.cin ;
always @(posedge \add_35s_35s_35_2_1_U10.top_add_35s_35s_35_2_1_Adder_7_U.clk )
\add_35s_35s_35_2_1_U10.top_add_35s_35s_35_2_1_Adder_7_U.bin_s1  <= _130_;
always @(posedge \add_35s_35s_35_2_1_U10.top_add_35s_35s_35_2_1_Adder_7_U.clk )
\add_35s_35s_35_2_1_U10.top_add_35s_35s_35_2_1_Adder_7_U.ain_s1  <= _129_;
always @(posedge \add_35s_35s_35_2_1_U10.top_add_35s_35s_35_2_1_Adder_7_U.clk )
\add_35s_35s_35_2_1_U10.top_add_35s_35s_35_2_1_Adder_7_U.sum_s1  <= _132_;
always @(posedge \add_35s_35s_35_2_1_U10.top_add_35s_35s_35_2_1_Adder_7_U.clk )
\add_35s_35s_35_2_1_U10.top_add_35s_35s_35_2_1_Adder_7_U.carry_s1  <= _131_;
assign _130_ = \add_35s_35s_35_2_1_U10.top_add_35s_35s_35_2_1_Adder_7_U.ce  ? \add_35s_35s_35_2_1_U10.top_add_35s_35s_35_2_1_Adder_7_U.b [34:17] : \add_35s_35s_35_2_1_U10.top_add_35s_35s_35_2_1_Adder_7_U.bin_s1 ;
assign _129_ = \add_35s_35s_35_2_1_U10.top_add_35s_35s_35_2_1_Adder_7_U.ce  ? \add_35s_35s_35_2_1_U10.top_add_35s_35s_35_2_1_Adder_7_U.a [34:17] : \add_35s_35s_35_2_1_U10.top_add_35s_35s_35_2_1_Adder_7_U.ain_s1 ;
assign _131_ = \add_35s_35s_35_2_1_U10.top_add_35s_35s_35_2_1_Adder_7_U.ce  ? \add_35s_35s_35_2_1_U10.top_add_35s_35s_35_2_1_Adder_7_U.facout_s1  : \add_35s_35s_35_2_1_U10.top_add_35s_35s_35_2_1_Adder_7_U.carry_s1 ;
assign _132_ = \add_35s_35s_35_2_1_U10.top_add_35s_35s_35_2_1_Adder_7_U.ce  ? \add_35s_35s_35_2_1_U10.top_add_35s_35s_35_2_1_Adder_7_U.fas_s1  : \add_35s_35s_35_2_1_U10.top_add_35s_35s_35_2_1_Adder_7_U.sum_s1 ;
assign _133_ = \add_35s_35s_35_2_1_U10.top_add_35s_35s_35_2_1_Adder_7_U.u1.a  + \add_35s_35s_35_2_1_U10.top_add_35s_35s_35_2_1_Adder_7_U.u1.b ;
assign { \add_35s_35s_35_2_1_U10.top_add_35s_35s_35_2_1_Adder_7_U.u1.cout , \add_35s_35s_35_2_1_U10.top_add_35s_35s_35_2_1_Adder_7_U.u1.s  } = _133_ + \add_35s_35s_35_2_1_U10.top_add_35s_35s_35_2_1_Adder_7_U.u1.cin ;
assign _134_ = \add_35s_35s_35_2_1_U10.top_add_35s_35s_35_2_1_Adder_7_U.u2.a  + \add_35s_35s_35_2_1_U10.top_add_35s_35s_35_2_1_Adder_7_U.u2.b ;
assign { \add_35s_35s_35_2_1_U10.top_add_35s_35s_35_2_1_Adder_7_U.u2.cout , \add_35s_35s_35_2_1_U10.top_add_35s_35s_35_2_1_Adder_7_U.u2.s  } = _134_ + \add_35s_35s_35_2_1_U10.top_add_35s_35s_35_2_1_Adder_7_U.u2.cin ;
always @(posedge \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_9_U.clk )
\add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_9_U.bin_s1  <= _136_;
always @(posedge \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_9_U.clk )
\add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_9_U.ain_s1  <= _135_;
always @(posedge \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_9_U.clk )
\add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_9_U.sum_s1  <= _138_;
always @(posedge \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_9_U.clk )
\add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_9_U.carry_s1  <= _137_;
assign _136_ = \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_9_U.ce  ? \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_9_U.b [2:1] : \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_9_U.bin_s1 ;
assign _135_ = \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_9_U.ce  ? \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_9_U.a [2:1] : \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_9_U.ain_s1 ;
assign _137_ = \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_9_U.ce  ? \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_9_U.facout_s1  : \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_9_U.carry_s1 ;
assign _138_ = \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_9_U.ce  ? \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_9_U.fas_s1  : \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_9_U.sum_s1 ;
assign _139_ = \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_9_U.u1.a  + \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_9_U.u1.b ;
assign { \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_9_U.u1.cout , \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_9_U.u1.s  } = _139_ + \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_9_U.u1.cin ;
assign _140_ = \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_9_U.u2.a  + \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_9_U.u2.b ;
assign { \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_9_U.u2.cout , \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_9_U.u2.s  } = _140_ + \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_9_U.u2.cin ;
always @(posedge \add_40s_40s_40_2_1_U7.top_add_40s_40s_40_2_1_Adder_5_U.clk )
\add_40s_40s_40_2_1_U7.top_add_40s_40s_40_2_1_Adder_5_U.bin_s1  <= _142_;
always @(posedge \add_40s_40s_40_2_1_U7.top_add_40s_40s_40_2_1_Adder_5_U.clk )
\add_40s_40s_40_2_1_U7.top_add_40s_40s_40_2_1_Adder_5_U.ain_s1  <= _141_;
always @(posedge \add_40s_40s_40_2_1_U7.top_add_40s_40s_40_2_1_Adder_5_U.clk )
\add_40s_40s_40_2_1_U7.top_add_40s_40s_40_2_1_Adder_5_U.sum_s1  <= _144_;
always @(posedge \add_40s_40s_40_2_1_U7.top_add_40s_40s_40_2_1_Adder_5_U.clk )
\add_40s_40s_40_2_1_U7.top_add_40s_40s_40_2_1_Adder_5_U.carry_s1  <= _143_;
assign _142_ = \add_40s_40s_40_2_1_U7.top_add_40s_40s_40_2_1_Adder_5_U.ce  ? \add_40s_40s_40_2_1_U7.top_add_40s_40s_40_2_1_Adder_5_U.b [39:20] : \add_40s_40s_40_2_1_U7.top_add_40s_40s_40_2_1_Adder_5_U.bin_s1 ;
assign _141_ = \add_40s_40s_40_2_1_U7.top_add_40s_40s_40_2_1_Adder_5_U.ce  ? \add_40s_40s_40_2_1_U7.top_add_40s_40s_40_2_1_Adder_5_U.a [39:20] : \add_40s_40s_40_2_1_U7.top_add_40s_40s_40_2_1_Adder_5_U.ain_s1 ;
assign _143_ = \add_40s_40s_40_2_1_U7.top_add_40s_40s_40_2_1_Adder_5_U.ce  ? \add_40s_40s_40_2_1_U7.top_add_40s_40s_40_2_1_Adder_5_U.facout_s1  : \add_40s_40s_40_2_1_U7.top_add_40s_40s_40_2_1_Adder_5_U.carry_s1 ;
assign _144_ = \add_40s_40s_40_2_1_U7.top_add_40s_40s_40_2_1_Adder_5_U.ce  ? \add_40s_40s_40_2_1_U7.top_add_40s_40s_40_2_1_Adder_5_U.fas_s1  : \add_40s_40s_40_2_1_U7.top_add_40s_40s_40_2_1_Adder_5_U.sum_s1 ;
assign _145_ = \add_40s_40s_40_2_1_U7.top_add_40s_40s_40_2_1_Adder_5_U.u1.a  + \add_40s_40s_40_2_1_U7.top_add_40s_40s_40_2_1_Adder_5_U.u1.b ;
assign { \add_40s_40s_40_2_1_U7.top_add_40s_40s_40_2_1_Adder_5_U.u1.cout , \add_40s_40s_40_2_1_U7.top_add_40s_40s_40_2_1_Adder_5_U.u1.s  } = _145_ + \add_40s_40s_40_2_1_U7.top_add_40s_40s_40_2_1_Adder_5_U.u1.cin ;
assign _146_ = \add_40s_40s_40_2_1_U7.top_add_40s_40s_40_2_1_Adder_5_U.u2.a  + \add_40s_40s_40_2_1_U7.top_add_40s_40s_40_2_1_Adder_5_U.u2.b ;
assign { \add_40s_40s_40_2_1_U7.top_add_40s_40s_40_2_1_Adder_5_U.u2.cout , \add_40s_40s_40_2_1_U7.top_add_40s_40s_40_2_1_Adder_5_U.u2.s  } = _146_ + \add_40s_40s_40_2_1_U7.top_add_40s_40s_40_2_1_Adder_5_U.u2.cin ;
assign _147_ = | trunc_ln851_1_reg_843;
assign _148_ = | op_15[1:0];
assign or_ln384_fu_631_p2 = overflow_reg_969 | op_11;
assign or_ln785_fu_344_p2 = r_reg_790 | p_Result_7_reg_796;
always @(posedge ap_clk)
ret_V_2_reg_729 <= _033_;
always @(posedge ap_clk)
ret_V_19_reg_927 <= _031_;
always @(posedge ap_clk)
select_ln69_1_reg_932 <= _039_;
always @(posedge ap_clk)
ret_V_18_reg_910 <= _030_;
always @(posedge ap_clk)
ret_V_9_cast_reg_915 <= _035_;
always @(posedge ap_clk)
ret_V_17_reg_880 <= _029_;
always @(posedge ap_clk)
select_ln69_reg_885 <= _040_;
always @(posedge ap_clk)
ret_V_16_reg_863 <= _028_;
always @(posedge ap_clk)
ret_V_6_cast_reg_868 <= _034_;
always @(posedge ap_clk)
ret_V_20_reg_1001 <= _032_;
always @(posedge ap_clk)
ret_V_16_cast_reg_1006 <= _027_;
always @(posedge ap_clk)
ret_V_13_reg_740 <= _024_;
always @(posedge ap_clk)
ret_reg_745 <= _037_;
always @(posedge ap_clk)
select_ln1192_reg_750 <= _038_;
always @(posedge ap_clk)
ret_V_12_reg_717 <= _023_;
always @(posedge ap_clk)
ret_V_reg_722 <= _036_;
always @(posedge ap_clk)
overflow_reg_969 <= _020_;
always @(posedge ap_clk)
op_26_V_reg_890 <= _017_;
always @(posedge ap_clk)
op_19_V_reg_980 <= _015_;
always @(posedge ap_clk)
op_30_V_reg_986 <= _018_;
always @(posedge ap_clk)
op_13_V_reg_833 <= _014_;
always @(posedge ap_clk)
ret_V_15_reg_838 <= _026_;
always @(posedge ap_clk)
trunc_ln851_1_reg_843 <= _041_;
always @(posedge ap_clk)
or_ln785_reg_807 <= _019_;
always @(posedge ap_clk)
op_23_V_reg_813 <= _016_;
always @(posedge ap_clk)
lhs_V_reg_818 <= _013_;
always @(posedge ap_clk)
icmp_ln851_reg_712 <= _012_;
always @(posedge ap_clk)
icmp_ln851_2_reg_905 <= _011_;
always @(posedge ap_clk)
icmp_ln851_1_reg_858 <= _010_;
always @(posedge ap_clk)
empty_reg_785 <= _008_;
always @(posedge ap_clk)
r_reg_790 <= _022_;
always @(posedge ap_clk)
p_Result_7_reg_796 <= _021_;
always @(posedge ap_clk)
and_ln365_reg_823 <= _006_;
always @(posedge ap_clk)
ret_V_14_reg_770 <= _025_;
always @(posedge ap_clk)
add_ln69_reg_775 <= _005_;
always @(posedge ap_clk)
icmp_ln785_reg_954 <= _009_;
always @(posedge ap_clk)
add_ln69_3_reg_959 <= _003_;
always @(posedge ap_clk)
add_ln69_4_reg_964 <= _004_;
always @(posedge ap_clk)
add_ln691_reg_875 <= _002_;
always @(posedge ap_clk)
add_ln691_2_reg_1013 <= _001_;
always @(posedge ap_clk)
add_ln691_1_reg_922 <= _000_;
always @(posedge ap_clk)
ap_CS_fsm <= _007_;
assign _042_ = _047_ ? 2'h2 : 2'h1;
assign _149_ = ap_CS_fsm == 1'h1;
function [31:0] _435_;
input [31:0] a;
input [1023:0] b;
input [31:0] s;
case (s)
32'b00000000000000000000000000000001:
_435_ = b[31:0];
32'b00000000000000000000000000000010:
_435_ = b[63:32];
32'b00000000000000000000000000000100:
_435_ = b[95:64];
32'b00000000000000000000000000001000:
_435_ = b[127:96];
32'b00000000000000000000000000010000:
_435_ = b[159:128];
32'b00000000000000000000000000100000:
_435_ = b[191:160];
32'b00000000000000000000000001000000:
_435_ = b[223:192];
32'b00000000000000000000000010000000:
_435_ = b[255:224];
32'b00000000000000000000000100000000:
_435_ = b[287:256];
32'b00000000000000000000001000000000:
_435_ = b[319:288];
32'b00000000000000000000010000000000:
_435_ = b[351:320];
32'b00000000000000000000100000000000:
_435_ = b[383:352];
32'b00000000000000000001000000000000:
_435_ = b[415:384];
32'b00000000000000000010000000000000:
_435_ = b[447:416];
32'b00000000000000000100000000000000:
_435_ = b[479:448];
32'b00000000000000001000000000000000:
_435_ = b[511:480];
32'b00000000000000010000000000000000:
_435_ = b[543:512];
32'b00000000000000100000000000000000:
_435_ = b[575:544];
32'b00000000000001000000000000000000:
_435_ = b[607:576];
32'b00000000000010000000000000000000:
_435_ = b[639:608];
32'b00000000000100000000000000000000:
_435_ = b[671:640];
32'b00000000001000000000000000000000:
_435_ = b[703:672];
32'b00000000010000000000000000000000:
_435_ = b[735:704];
32'b00000000100000000000000000000000:
_435_ = b[767:736];
32'b00000001000000000000000000000000:
_435_ = b[799:768];
32'b00000010000000000000000000000000:
_435_ = b[831:800];
32'b00000100000000000000000000000000:
_435_ = b[863:832];
32'b00001000000000000000000000000000:
_435_ = b[895:864];
32'b00010000000000000000000000000000:
_435_ = b[927:896];
32'b00100000000000000000000000000000:
_435_ = b[959:928];
32'b01000000000000000000000000000000:
_435_ = b[991:960];
32'b10000000000000000000000000000000:
_435_ = b[1023:992];
32'b00000000000000000000000000000000:
_435_ = a;
default:
_435_ = 32'bx;
endcase
endfunction
assign ap_NS_fsm = _435_(32'hxxxxxxxx, { 30'h00000000, _042_, 992'h00000004000000080000001000000020000000400000008000000100000002000000040000000800000010000000200000004000000080000001000000020000000400000008000000100000002000000040000000800000010000000200000004000000080000001000000020000000400000008000000000000001 }, { _149_, _180_, _179_, _178_, _177_, _176_, _175_, _174_, _173_, _172_, _171_, _170_, _169_, _168_, _167_, _166_, _165_, _164_, _163_, _162_, _161_, _160_, _159_, _158_, _157_, _156_, _155_, _154_, _153_, _152_, _151_, _150_ });
assign _150_ = ap_CS_fsm == 32'd2147483648;
assign _151_ = ap_CS_fsm == 31'h40000000;
assign _152_ = ap_CS_fsm == 30'h20000000;
assign _153_ = ap_CS_fsm == 29'h10000000;
assign _154_ = ap_CS_fsm == 28'h8000000;
assign _155_ = ap_CS_fsm == 27'h4000000;
assign _156_ = ap_CS_fsm == 26'h2000000;
assign _157_ = ap_CS_fsm == 25'h1000000;
assign _158_ = ap_CS_fsm == 24'h800000;
assign _159_ = ap_CS_fsm == 23'h400000;
assign _160_ = ap_CS_fsm == 22'h200000;
assign _161_ = ap_CS_fsm == 21'h100000;
assign _162_ = ap_CS_fsm == 20'h80000;
assign _163_ = ap_CS_fsm == 19'h40000;
assign _164_ = ap_CS_fsm == 18'h20000;
assign _165_ = ap_CS_fsm == 17'h10000;
assign _166_ = ap_CS_fsm == 16'h8000;
assign _167_ = ap_CS_fsm == 15'h4000;
assign _168_ = ap_CS_fsm == 14'h2000;
assign _169_ = ap_CS_fsm == 13'h1000;
assign _170_ = ap_CS_fsm == 12'h800;
assign _171_ = ap_CS_fsm == 11'h400;
assign _172_ = ap_CS_fsm == 10'h200;
assign _173_ = ap_CS_fsm == 9'h100;
assign _174_ = ap_CS_fsm == 8'h80;
assign _175_ = ap_CS_fsm == 7'h40;
assign _176_ = ap_CS_fsm == 6'h20;
assign _177_ = ap_CS_fsm == 5'h10;
assign _178_ = ap_CS_fsm == 4'h8;
assign _179_ = ap_CS_fsm == 3'h4;
assign _180_ = ap_CS_fsm == 2'h2;
assign op_31_ap_vld = ap_CS_fsm[31] ? 1'h1 : 1'h0;
assign ap_idle = _046_ ? 1'h1 : 1'h0;
assign _033_ = _045_ ? grp_fu_247_p2 : ret_V_2_reg_729;
assign _039_ = ap_CS_fsm[22] ? select_ln69_1_fu_560_p3 : select_ln69_1_reg_932;
assign _031_ = ap_CS_fsm[22] ? ret_V_19_fu_553_p3 : ret_V_19_reg_927;
assign _035_ = ap_CS_fsm[19] ? grp_fu_510_p2[33:2] : ret_V_9_cast_reg_915;
assign _030_ = ap_CS_fsm[19] ? grp_fu_510_p2 : ret_V_18_reg_910;
assign _040_ = ap_CS_fsm[15] ? select_ln69_fu_483_p3 : select_ln69_reg_885;
assign _029_ = ap_CS_fsm[15] ? ret_V_17_fu_476_p3 : ret_V_17_reg_880;
assign _034_ = ap_CS_fsm[12] ? grp_fu_438_p2[38:7] : ret_V_6_cast_reg_868;
assign _028_ = ap_CS_fsm[12] ? grp_fu_438_p2 : ret_V_16_reg_863;
assign _027_ = ap_CS_fsm[28] ? grp_fu_657_p2[32:1] : ret_V_16_cast_reg_1006;
assign _032_ = ap_CS_fsm[28] ? grp_fu_657_p2 : ret_V_20_reg_1001;
assign _038_ = ap_CS_fsm[4] ? select_ln1192_fu_279_p3 : select_ln1192_reg_750;
assign _037_ = ap_CS_fsm[4] ? ret_fu_271_p3 : ret_reg_745;
assign _024_ = ap_CS_fsm[4] ? ret_V_13_fu_264_p3 : ret_V_13_reg_740;
assign _036_ = ap_CS_fsm[1] ? grp_fu_221_p2[16:7] : ret_V_reg_722;
assign _023_ = ap_CS_fsm[1] ? grp_fu_221_p2 : ret_V_12_reg_717;
assign _020_ = ap_CS_fsm[25] ? overflow_fu_604_p2 : overflow_reg_969;
assign _017_ = ap_CS_fsm[17] ? grp_fu_491_p2 : op_26_V_reg_890;
assign _018_ = ap_CS_fsm[26] ? grp_fu_612_p2 : op_30_V_reg_986;
assign _015_ = ap_CS_fsm[26] ? op_19_V_fu_635_p3 : op_19_V_reg_980;
assign _041_ = ap_CS_fsm[10] ? op_13_V_fu_413_p3[6:0] : trunc_ln851_1_reg_843;
assign _026_ = ap_CS_fsm[10] ? grp_fu_379_p2 : ret_V_15_reg_838;
assign _014_ = ap_CS_fsm[10] ? op_13_V_fu_413_p3 : op_13_V_reg_833;
assign _013_ = ap_CS_fsm[8] ? lhs_V_fu_348_p2 : lhs_V_reg_818;
assign _016_ = ap_CS_fsm[8] ? grp_fu_339_p2 : op_23_V_reg_813;
assign _019_ = ap_CS_fsm[8] ? or_ln785_fu_344_p2 : or_ln785_reg_807;
assign _012_ = ap_CS_fsm[0] ? icmp_ln851_fu_231_p2 : icmp_ln851_reg_712;
assign _011_ = ap_CS_fsm[18] ? icmp_ln851_2_fu_520_p2 : icmp_ln851_2_reg_905;
assign _010_ = ap_CS_fsm[11] ? icmp_ln851_1_fu_444_p2 : icmp_ln851_1_reg_858;
assign _021_ = ap_CS_fsm[7] ? p_Result_7_fu_330_p2 : p_Result_7_reg_796;
assign _022_ = ap_CS_fsm[7] ? r_fu_316_p2 : r_reg_790;
assign _008_ = ap_CS_fsm[7] ? op_8[0] : empty_reg_785;
assign _006_ = ap_CS_fsm[9] ? and_ln365_fu_371_p2 : and_ln365_reg_823;
assign _005_ = ap_CS_fsm[6] ? grp_fu_306_p2 : add_ln69_reg_775;
assign _025_ = ap_CS_fsm[6] ? grp_fu_290_p2 : ret_V_14_reg_770;
assign _004_ = ap_CS_fsm[24] ? grp_fu_580_p2 : add_ln69_4_reg_964;
assign _003_ = ap_CS_fsm[24] ? grp_fu_575_p2 : add_ln69_3_reg_959;
assign _009_ = ap_CS_fsm[24] ? icmp_ln785_fu_593_p2 : icmp_ln785_reg_954;
assign _002_ = _044_ ? grp_fu_459_p2 : add_ln691_reg_875;
assign _001_ = ap_CS_fsm[30] ? grp_fu_673_p2 : add_ln691_2_reg_1013;
assign _000_ = _043_ ? grp_fu_536_p2 : add_ln691_1_reg_922;
assign _007_ = ap_rst ? 32'd1 : ap_NS_fsm;
assign icmp_ln785_fu_593_p2 = op_11 ? 1'h1 : 1'h0;
assign icmp_ln851_1_fu_444_p2 = _147_ ? 1'h1 : 1'h0;
assign icmp_ln851_2_fu_520_p2 = _148_ ? 1'h1 : 1'h0;
assign icmp_ln851_fu_231_p2 = _050_ ? 1'h1 : 1'h0;
assign op_13_V_fu_413_p3 = and_ln365_reg_823 ? { r_reg_790, 7'h00 } : select_ln785_fu_406_p3;
assign op_19_V_fu_635_p3 = or_ln384_fu_631_p2 ? select_ln384_fu_624_p3 : p_Val2_5_fu_617_p3;
assign op_31 = ret_V_20_reg_1001[33] ? select_ln850_3_fu_688_p3 : ret_V_16_cast_reg_1006;
assign p_Val2_5_fu_617_p3 = op_11 ? 2'h2 : 2'h0;
assign ret_V_13_fu_264_p3 = ret_V_12_reg_717[16] ? select_ln850_fu_259_p3 : ret_V_reg_722;
assign ret_V_17_fu_476_p3 = ret_V_16_reg_863[39] ? select_ln850_1_fu_471_p3 : ret_V_6_cast_reg_868;
assign ret_V_19_fu_553_p3 = ret_V_18_reg_910[34] ? select_ln850_2_fu_548_p3 : ret_V_9_cast_reg_915;
assign ret_fu_271_p3 = op_2 ? 2'h3 : op_4;
assign select_ln1192_fu_279_p3 = op_2 ? 11'h7ff : 11'h000;
assign select_ln384_fu_624_p3 = overflow_reg_969 ? 2'h1 : 2'h3;
assign select_ln69_1_fu_560_p3 = op_2 ? 3'h7 : 3'h0;
assign select_ln69_fu_483_p3 = op_14 ? 32'd4294967295 : 32'd0;
assign select_ln785_fu_406_p3 = or_ln785_reg_807 ? { p_Result_7_reg_796, 7'h7f } : 8'h00;
assign select_ln850_1_fu_471_p3 = icmp_ln851_1_reg_858 ? add_ln691_reg_875 : ret_V_6_cast_reg_868;
assign select_ln850_2_fu_548_p3 = icmp_ln851_2_reg_905 ? add_ln691_1_reg_922 : ret_V_9_cast_reg_915;
assign select_ln850_3_fu_688_p3 = op_19_V_reg_980[0] ? add_ln691_2_reg_1013 : ret_V_16_cast_reg_1006;
assign select_ln850_fu_259_p3 = icmp_ln851_reg_712 ? ret_V_reg_722 : ret_V_2_reg_729;
assign xor_ln365_1_fu_366_p2 = p_Result_7_fu_330_p2 ^ empty_reg_785;
assign ap_CS_fsm_state1 = ap_CS_fsm[0];
assign ap_CS_fsm_state10 = ap_CS_fsm[9];
assign ap_CS_fsm_state11 = ap_CS_fsm[10];
assign ap_CS_fsm_state12 = ap_CS_fsm[11];
assign ap_CS_fsm_state13 = ap_CS_fsm[12];
assign ap_CS_fsm_state14 = ap_CS_fsm[13];
assign ap_CS_fsm_state15 = ap_CS_fsm[14];
assign ap_CS_fsm_state16 = ap_CS_fsm[15];
assign ap_CS_fsm_state17 = ap_CS_fsm[16];
assign ap_CS_fsm_state18 = ap_CS_fsm[17];
assign ap_CS_fsm_state19 = ap_CS_fsm[18];
assign ap_CS_fsm_state2 = ap_CS_fsm[1];
assign ap_CS_fsm_state20 = ap_CS_fsm[19];
assign ap_CS_fsm_state21 = ap_CS_fsm[20];
assign ap_CS_fsm_state22 = ap_CS_fsm[21];
assign ap_CS_fsm_state23 = ap_CS_fsm[22];
assign ap_CS_fsm_state24 = ap_CS_fsm[23];
assign ap_CS_fsm_state25 = ap_CS_fsm[24];
assign ap_CS_fsm_state26 = ap_CS_fsm[25];
assign ap_CS_fsm_state27 = ap_CS_fsm[26];
assign ap_CS_fsm_state28 = ap_CS_fsm[27];
assign ap_CS_fsm_state29 = ap_CS_fsm[28];
assign ap_CS_fsm_state3 = ap_CS_fsm[2];
assign ap_CS_fsm_state30 = ap_CS_fsm[29];
assign ap_CS_fsm_state31 = ap_CS_fsm[30];
assign ap_CS_fsm_state32 = ap_CS_fsm[31];
assign ap_CS_fsm_state4 = ap_CS_fsm[3];
assign ap_CS_fsm_state5 = ap_CS_fsm[4];
assign ap_CS_fsm_state6 = ap_CS_fsm[5];
assign ap_CS_fsm_state7 = ap_CS_fsm[6];
assign ap_CS_fsm_state8 = ap_CS_fsm[7];
assign ap_CS_fsm_state9 = ap_CS_fsm[8];
assign ap_done = op_31_ap_vld;
assign ap_ready = op_31_ap_vld;
assign empty_fu_312_p1 = op_8[0];
assign grp_fu_221_p0 = { op_0[7], op_0[7], op_0, 7'h00 };
assign grp_fu_221_p1 = { op_1[15], op_1 };
assign grp_fu_290_p0 = { ret_V_13_reg_740[9], ret_V_13_reg_740 };
assign grp_fu_306_p0 = { 2'h0, ret_reg_745[1], ret_reg_745[1], ret_reg_745[1], ret_reg_745[1], ret_reg_745[1], ret_reg_745[1], ret_reg_745 };
assign grp_fu_306_p1 = { op_10[3], op_10[3], op_10[3], op_10[3], op_10[3], op_10[3], op_10 };
assign grp_fu_339_p0 = { add_ln69_reg_775[9], add_ln69_reg_775 };
assign grp_fu_379_p0 = { 10'h000, lhs_V_reg_818 };
assign grp_fu_438_p0 = { ret_V_15_reg_838[10], ret_V_15_reg_838[10], ret_V_15_reg_838[10], ret_V_15_reg_838[10], ret_V_15_reg_838[10], ret_V_15_reg_838[10], ret_V_15_reg_838[10], ret_V_15_reg_838[10], ret_V_15_reg_838[10], ret_V_15_reg_838[10], ret_V_15_reg_838[10], ret_V_15_reg_838[10], ret_V_15_reg_838[10], ret_V_15_reg_838[10], ret_V_15_reg_838[10], ret_V_15_reg_838[10], ret_V_15_reg_838[10], ret_V_15_reg_838[10], ret_V_15_reg_838[10], ret_V_15_reg_838[10], ret_V_15_reg_838[10], ret_V_15_reg_838[10], ret_V_15_reg_838, 7'h00 };
assign grp_fu_438_p1 = { op_13_V_reg_833[7], op_13_V_reg_833[7], op_13_V_reg_833[7], op_13_V_reg_833[7], op_13_V_reg_833[7], op_13_V_reg_833[7], op_13_V_reg_833[7], op_13_V_reg_833[7], op_13_V_reg_833[7], op_13_V_reg_833[7], op_13_V_reg_833[7], op_13_V_reg_833[7], op_13_V_reg_833[7], op_13_V_reg_833[7], op_13_V_reg_833[7], op_13_V_reg_833[7], op_13_V_reg_833[7], op_13_V_reg_833[7], op_13_V_reg_833[7], op_13_V_reg_833[7], op_13_V_reg_833[7], op_13_V_reg_833[7], op_13_V_reg_833[7], op_13_V_reg_833[7], op_13_V_reg_833[7], op_13_V_reg_833[7], op_13_V_reg_833[7], op_13_V_reg_833[7], op_13_V_reg_833[7], op_13_V_reg_833[7], op_13_V_reg_833[7], op_13_V_reg_833[7], op_13_V_reg_833 };
assign grp_fu_510_p0 = { op_26_V_reg_890[31], op_26_V_reg_890, 2'h0 };
assign grp_fu_510_p1 = { op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15 };
assign grp_fu_575_p1 = { op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16 };
assign grp_fu_580_p0 = { op_17[1], op_17 };
assign grp_fu_612_p0 = { add_ln69_4_reg_964[2], add_ln69_4_reg_964[2], add_ln69_4_reg_964[2], add_ln69_4_reg_964[2], add_ln69_4_reg_964[2], add_ln69_4_reg_964[2], add_ln69_4_reg_964[2], add_ln69_4_reg_964[2], add_ln69_4_reg_964[2], add_ln69_4_reg_964[2], add_ln69_4_reg_964[2], add_ln69_4_reg_964[2], add_ln69_4_reg_964[2], add_ln69_4_reg_964[2], add_ln69_4_reg_964[2], add_ln69_4_reg_964[2], add_ln69_4_reg_964[2], add_ln69_4_reg_964[2], add_ln69_4_reg_964[2], add_ln69_4_reg_964[2], add_ln69_4_reg_964[2], add_ln69_4_reg_964[2], add_ln69_4_reg_964[2], add_ln69_4_reg_964[2], add_ln69_4_reg_964[2], add_ln69_4_reg_964[2], add_ln69_4_reg_964[2], add_ln69_4_reg_964[2], add_ln69_4_reg_964[2], add_ln69_4_reg_964 };
assign grp_fu_657_p0 = { op_30_V_reg_986[31], op_30_V_reg_986, 1'h0 };
assign grp_fu_657_p1 = { op_19_V_reg_980[1], op_19_V_reg_980[1], op_19_V_reg_980[1], op_19_V_reg_980[1], op_19_V_reg_980[1], op_19_V_reg_980[1], op_19_V_reg_980[1], op_19_V_reg_980[1], op_19_V_reg_980[1], op_19_V_reg_980[1], op_19_V_reg_980[1], op_19_V_reg_980[1], op_19_V_reg_980[1], op_19_V_reg_980[1], op_19_V_reg_980[1], op_19_V_reg_980[1], op_19_V_reg_980[1], op_19_V_reg_980[1], op_19_V_reg_980[1], op_19_V_reg_980[1], op_19_V_reg_980[1], op_19_V_reg_980[1], op_19_V_reg_980[1], op_19_V_reg_980[1], op_19_V_reg_980[1], op_19_V_reg_980[1], op_19_V_reg_980[1], op_19_V_reg_980[1], op_19_V_reg_980[1], op_19_V_reg_980[1], op_19_V_reg_980[1], op_19_V_reg_980[1], op_19_V_reg_980 };
assign lhs_fu_205_p3 = { op_0, 7'h00 };
assign or_ln384_fu_631_p1 = op_11;
assign or_ln785_1_fu_585_p1 = op_11;
assign or_ln785_1_fu_585_p3 = { op_11, 1'h0 };
assign p_Result_3_fu_397_p4 = { p_Result_7_reg_796, 7'h7f };
assign p_Result_4_fu_464_p3 = ret_V_16_reg_863[39];
assign p_Result_5_fu_541_p3 = ret_V_18_reg_910[34];
assign p_Result_6_fu_678_p3 = ret_V_20_reg_1001[33];
assign p_Result_s_fu_252_p3 = ret_V_12_reg_717[16];
assign p_Val2_1_fu_384_p3 = { r_reg_790, 7'h00 };
assign p_Val2_3_fu_391_p2 = 7'h7f;
assign p_Val2_5_fu_617_p0 = op_11;
assign rhs_4_fu_499_p3 = { op_26_V_reg_890, 2'h0 };
assign rhs_6_fu_646_p3 = { op_30_V_reg_986, 1'h0 };
assign sext_ln69_fu_295_p1 = { ret_reg_745[1], ret_reg_745[1], ret_reg_745[1], ret_reg_745[1], ret_reg_745[1], ret_reg_745[1], ret_reg_745 };
assign sext_ln703_2_fu_495_p0 = op_15;
assign sext_ln703_fu_217_p0 = op_1;
assign tmp_1_fu_353_p3 = op_8[1];
assign tmp_3_fu_427_p3 = { ret_V_15_reg_838, 7'h00 };
assign tmp_fu_322_p3 = op_8[1];
assign trunc_ln851_1_fu_420_p1 = op_13_V_fu_413_p3[6:0];
assign trunc_ln851_2_fu_516_p0 = op_15;
assign trunc_ln851_2_fu_516_p1 = op_15[1:0];
assign trunc_ln851_3_fu_685_p1 = op_19_V_reg_980[0];
assign trunc_ln851_fu_227_p0 = op_1;
assign trunc_ln851_fu_227_p1 = op_1[6:0];
assign xor_ln365_fu_360_p2 = p_Result_7_fu_330_p2;
assign xor_ln785_fu_599_p0 = op_11;
assign \add_40s_40s_40_2_1_U7.top_add_40s_40s_40_2_1_Adder_5_U.ain_s0  = \add_40s_40s_40_2_1_U7.top_add_40s_40s_40_2_1_Adder_5_U.a ;
assign \add_40s_40s_40_2_1_U7.top_add_40s_40s_40_2_1_Adder_5_U.bin_s0  = \add_40s_40s_40_2_1_U7.top_add_40s_40s_40_2_1_Adder_5_U.b ;
assign \add_40s_40s_40_2_1_U7.top_add_40s_40s_40_2_1_Adder_5_U.s  = { \add_40s_40s_40_2_1_U7.top_add_40s_40s_40_2_1_Adder_5_U.fas_s2 , \add_40s_40s_40_2_1_U7.top_add_40s_40s_40_2_1_Adder_5_U.sum_s1  };
assign \add_40s_40s_40_2_1_U7.top_add_40s_40s_40_2_1_Adder_5_U.u2.a  = \add_40s_40s_40_2_1_U7.top_add_40s_40s_40_2_1_Adder_5_U.ain_s1 ;
assign \add_40s_40s_40_2_1_U7.top_add_40s_40s_40_2_1_Adder_5_U.u2.b  = \add_40s_40s_40_2_1_U7.top_add_40s_40s_40_2_1_Adder_5_U.bin_s1 ;
assign \add_40s_40s_40_2_1_U7.top_add_40s_40s_40_2_1_Adder_5_U.u2.cin  = \add_40s_40s_40_2_1_U7.top_add_40s_40s_40_2_1_Adder_5_U.carry_s1 ;
assign \add_40s_40s_40_2_1_U7.top_add_40s_40s_40_2_1_Adder_5_U.facout_s2  = \add_40s_40s_40_2_1_U7.top_add_40s_40s_40_2_1_Adder_5_U.u2.cout ;
assign \add_40s_40s_40_2_1_U7.top_add_40s_40s_40_2_1_Adder_5_U.fas_s2  = \add_40s_40s_40_2_1_U7.top_add_40s_40s_40_2_1_Adder_5_U.u2.s ;
assign \add_40s_40s_40_2_1_U7.top_add_40s_40s_40_2_1_Adder_5_U.u1.a  = \add_40s_40s_40_2_1_U7.top_add_40s_40s_40_2_1_Adder_5_U.a [19:0];
assign \add_40s_40s_40_2_1_U7.top_add_40s_40s_40_2_1_Adder_5_U.u1.b  = \add_40s_40s_40_2_1_U7.top_add_40s_40s_40_2_1_Adder_5_U.b [19:0];
assign \add_40s_40s_40_2_1_U7.top_add_40s_40s_40_2_1_Adder_5_U.u1.cin  = 1'h0;
assign \add_40s_40s_40_2_1_U7.top_add_40s_40s_40_2_1_Adder_5_U.facout_s1  = \add_40s_40s_40_2_1_U7.top_add_40s_40s_40_2_1_Adder_5_U.u1.cout ;
assign \add_40s_40s_40_2_1_U7.top_add_40s_40s_40_2_1_Adder_5_U.fas_s1  = \add_40s_40s_40_2_1_U7.top_add_40s_40s_40_2_1_Adder_5_U.u1.s ;
assign \add_40s_40s_40_2_1_U7.top_add_40s_40s_40_2_1_Adder_5_U.a  = \add_40s_40s_40_2_1_U7.din0 ;
assign \add_40s_40s_40_2_1_U7.top_add_40s_40s_40_2_1_Adder_5_U.b  = \add_40s_40s_40_2_1_U7.din1 ;
assign \add_40s_40s_40_2_1_U7.top_add_40s_40s_40_2_1_Adder_5_U.ce  = \add_40s_40s_40_2_1_U7.ce ;
assign \add_40s_40s_40_2_1_U7.top_add_40s_40s_40_2_1_Adder_5_U.clk  = \add_40s_40s_40_2_1_U7.clk ;
assign \add_40s_40s_40_2_1_U7.top_add_40s_40s_40_2_1_Adder_5_U.reset  = \add_40s_40s_40_2_1_U7.reset ;
assign \add_40s_40s_40_2_1_U7.dout  = \add_40s_40s_40_2_1_U7.top_add_40s_40s_40_2_1_Adder_5_U.s ;
assign \add_40s_40s_40_2_1_U7.ce  = 1'h1;
assign \add_40s_40s_40_2_1_U7.clk  = ap_clk;
assign \add_40s_40s_40_2_1_U7.din0  = { ret_V_15_reg_838[10], ret_V_15_reg_838[10], ret_V_15_reg_838[10], ret_V_15_reg_838[10], ret_V_15_reg_838[10], ret_V_15_reg_838[10], ret_V_15_reg_838[10], ret_V_15_reg_838[10], ret_V_15_reg_838[10], ret_V_15_reg_838[10], ret_V_15_reg_838[10], ret_V_15_reg_838[10], ret_V_15_reg_838[10], ret_V_15_reg_838[10], ret_V_15_reg_838[10], ret_V_15_reg_838[10], ret_V_15_reg_838[10], ret_V_15_reg_838[10], ret_V_15_reg_838[10], ret_V_15_reg_838[10], ret_V_15_reg_838[10], ret_V_15_reg_838[10], ret_V_15_reg_838, 7'h00 };
assign \add_40s_40s_40_2_1_U7.din1  = { op_13_V_reg_833[7], op_13_V_reg_833[7], op_13_V_reg_833[7], op_13_V_reg_833[7], op_13_V_reg_833[7], op_13_V_reg_833[7], op_13_V_reg_833[7], op_13_V_reg_833[7], op_13_V_reg_833[7], op_13_V_reg_833[7], op_13_V_reg_833[7], op_13_V_reg_833[7], op_13_V_reg_833[7], op_13_V_reg_833[7], op_13_V_reg_833[7], op_13_V_reg_833[7], op_13_V_reg_833[7], op_13_V_reg_833[7], op_13_V_reg_833[7], op_13_V_reg_833[7], op_13_V_reg_833[7], op_13_V_reg_833[7], op_13_V_reg_833[7], op_13_V_reg_833[7], op_13_V_reg_833[7], op_13_V_reg_833[7], op_13_V_reg_833[7], op_13_V_reg_833[7], op_13_V_reg_833[7], op_13_V_reg_833[7], op_13_V_reg_833[7], op_13_V_reg_833[7], op_13_V_reg_833 };
assign grp_fu_438_p2 = \add_40s_40s_40_2_1_U7.dout ;
assign \add_40s_40s_40_2_1_U7.reset  = ap_rst;
assign \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_9_U.ain_s0  = \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_9_U.a ;
assign \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_9_U.bin_s0  = \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_9_U.b ;
assign \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_9_U.s  = { \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_9_U.fas_s2 , \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_9_U.sum_s1  };
assign \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_9_U.u2.a  = \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_9_U.ain_s1 ;
assign \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_9_U.u2.b  = \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_9_U.bin_s1 ;
assign \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_9_U.u2.cin  = \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_9_U.carry_s1 ;
assign \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_9_U.facout_s2  = \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_9_U.u2.cout ;
assign \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_9_U.fas_s2  = \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_9_U.u2.s ;
assign \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_9_U.u1.a  = \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_9_U.a [0];
assign \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_9_U.u1.b  = \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_9_U.b [0];
assign \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_9_U.u1.cin  = 1'h0;
assign \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_9_U.facout_s1  = \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_9_U.u1.cout ;
assign \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_9_U.fas_s1  = \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_9_U.u1.s ;
assign \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_9_U.a  = \add_3s_3ns_3_2_1_U13.din0 ;
assign \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_9_U.b  = \add_3s_3ns_3_2_1_U13.din1 ;
assign \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_9_U.ce  = \add_3s_3ns_3_2_1_U13.ce ;
assign \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_9_U.clk  = \add_3s_3ns_3_2_1_U13.clk ;
assign \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_9_U.reset  = \add_3s_3ns_3_2_1_U13.reset ;
assign \add_3s_3ns_3_2_1_U13.dout  = \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_9_U.s ;
assign \add_3s_3ns_3_2_1_U13.ce  = 1'h1;
assign \add_3s_3ns_3_2_1_U13.clk  = ap_clk;
assign \add_3s_3ns_3_2_1_U13.din0  = { op_17[1], op_17 };
assign \add_3s_3ns_3_2_1_U13.din1  = select_ln69_1_reg_932;
assign grp_fu_580_p2 = \add_3s_3ns_3_2_1_U13.dout ;
assign \add_3s_3ns_3_2_1_U13.reset  = ap_rst;
assign \add_35s_35s_35_2_1_U10.top_add_35s_35s_35_2_1_Adder_7_U.ain_s0  = \add_35s_35s_35_2_1_U10.top_add_35s_35s_35_2_1_Adder_7_U.a ;
assign \add_35s_35s_35_2_1_U10.top_add_35s_35s_35_2_1_Adder_7_U.bin_s0  = \add_35s_35s_35_2_1_U10.top_add_35s_35s_35_2_1_Adder_7_U.b ;
assign \add_35s_35s_35_2_1_U10.top_add_35s_35s_35_2_1_Adder_7_U.s  = { \add_35s_35s_35_2_1_U10.top_add_35s_35s_35_2_1_Adder_7_U.fas_s2 , \add_35s_35s_35_2_1_U10.top_add_35s_35s_35_2_1_Adder_7_U.sum_s1  };
assign \add_35s_35s_35_2_1_U10.top_add_35s_35s_35_2_1_Adder_7_U.u2.a  = \add_35s_35s_35_2_1_U10.top_add_35s_35s_35_2_1_Adder_7_U.ain_s1 ;
assign \add_35s_35s_35_2_1_U10.top_add_35s_35s_35_2_1_Adder_7_U.u2.b  = \add_35s_35s_35_2_1_U10.top_add_35s_35s_35_2_1_Adder_7_U.bin_s1 ;
assign \add_35s_35s_35_2_1_U10.top_add_35s_35s_35_2_1_Adder_7_U.u2.cin  = \add_35s_35s_35_2_1_U10.top_add_35s_35s_35_2_1_Adder_7_U.carry_s1 ;
assign \add_35s_35s_35_2_1_U10.top_add_35s_35s_35_2_1_Adder_7_U.facout_s2  = \add_35s_35s_35_2_1_U10.top_add_35s_35s_35_2_1_Adder_7_U.u2.cout ;
assign \add_35s_35s_35_2_1_U10.top_add_35s_35s_35_2_1_Adder_7_U.fas_s2  = \add_35s_35s_35_2_1_U10.top_add_35s_35s_35_2_1_Adder_7_U.u2.s ;
assign \add_35s_35s_35_2_1_U10.top_add_35s_35s_35_2_1_Adder_7_U.u1.a  = \add_35s_35s_35_2_1_U10.top_add_35s_35s_35_2_1_Adder_7_U.a [16:0];
assign \add_35s_35s_35_2_1_U10.top_add_35s_35s_35_2_1_Adder_7_U.u1.b  = \add_35s_35s_35_2_1_U10.top_add_35s_35s_35_2_1_Adder_7_U.b [16:0];
assign \add_35s_35s_35_2_1_U10.top_add_35s_35s_35_2_1_Adder_7_U.u1.cin  = 1'h0;
assign \add_35s_35s_35_2_1_U10.top_add_35s_35s_35_2_1_Adder_7_U.facout_s1  = \add_35s_35s_35_2_1_U10.top_add_35s_35s_35_2_1_Adder_7_U.u1.cout ;
assign \add_35s_35s_35_2_1_U10.top_add_35s_35s_35_2_1_Adder_7_U.fas_s1  = \add_35s_35s_35_2_1_U10.top_add_35s_35s_35_2_1_Adder_7_U.u1.s ;
assign \add_35s_35s_35_2_1_U10.top_add_35s_35s_35_2_1_Adder_7_U.a  = \add_35s_35s_35_2_1_U10.din0 ;
assign \add_35s_35s_35_2_1_U10.top_add_35s_35s_35_2_1_Adder_7_U.b  = \add_35s_35s_35_2_1_U10.din1 ;
assign \add_35s_35s_35_2_1_U10.top_add_35s_35s_35_2_1_Adder_7_U.ce  = \add_35s_35s_35_2_1_U10.ce ;
assign \add_35s_35s_35_2_1_U10.top_add_35s_35s_35_2_1_Adder_7_U.clk  = \add_35s_35s_35_2_1_U10.clk ;
assign \add_35s_35s_35_2_1_U10.top_add_35s_35s_35_2_1_Adder_7_U.reset  = \add_35s_35s_35_2_1_U10.reset ;
assign \add_35s_35s_35_2_1_U10.dout  = \add_35s_35s_35_2_1_U10.top_add_35s_35s_35_2_1_Adder_7_U.s ;
assign \add_35s_35s_35_2_1_U10.ce  = 1'h1;
assign \add_35s_35s_35_2_1_U10.clk  = ap_clk;
assign \add_35s_35s_35_2_1_U10.din0  = { op_26_V_reg_890[31], op_26_V_reg_890, 2'h0 };
assign \add_35s_35s_35_2_1_U10.din1  = { op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15 };
assign grp_fu_510_p2 = \add_35s_35s_35_2_1_U10.dout ;
assign \add_35s_35s_35_2_1_U10.reset  = ap_rst;
assign \add_34s_34s_34_2_1_U15.top_add_34s_34s_34_2_1_Adder_11_U.ain_s0  = \add_34s_34s_34_2_1_U15.top_add_34s_34s_34_2_1_Adder_11_U.a ;
assign \add_34s_34s_34_2_1_U15.top_add_34s_34s_34_2_1_Adder_11_U.bin_s0  = \add_34s_34s_34_2_1_U15.top_add_34s_34s_34_2_1_Adder_11_U.b ;
assign \add_34s_34s_34_2_1_U15.top_add_34s_34s_34_2_1_Adder_11_U.s  = { \add_34s_34s_34_2_1_U15.top_add_34s_34s_34_2_1_Adder_11_U.fas_s2 , \add_34s_34s_34_2_1_U15.top_add_34s_34s_34_2_1_Adder_11_U.sum_s1  };
assign \add_34s_34s_34_2_1_U15.top_add_34s_34s_34_2_1_Adder_11_U.u2.a  = \add_34s_34s_34_2_1_U15.top_add_34s_34s_34_2_1_Adder_11_U.ain_s1 ;
assign \add_34s_34s_34_2_1_U15.top_add_34s_34s_34_2_1_Adder_11_U.u2.b  = \add_34s_34s_34_2_1_U15.top_add_34s_34s_34_2_1_Adder_11_U.bin_s1 ;
assign \add_34s_34s_34_2_1_U15.top_add_34s_34s_34_2_1_Adder_11_U.u2.cin  = \add_34s_34s_34_2_1_U15.top_add_34s_34s_34_2_1_Adder_11_U.carry_s1 ;
assign \add_34s_34s_34_2_1_U15.top_add_34s_34s_34_2_1_Adder_11_U.facout_s2  = \add_34s_34s_34_2_1_U15.top_add_34s_34s_34_2_1_Adder_11_U.u2.cout ;
assign \add_34s_34s_34_2_1_U15.top_add_34s_34s_34_2_1_Adder_11_U.fas_s2  = \add_34s_34s_34_2_1_U15.top_add_34s_34s_34_2_1_Adder_11_U.u2.s ;
assign \add_34s_34s_34_2_1_U15.top_add_34s_34s_34_2_1_Adder_11_U.u1.a  = \add_34s_34s_34_2_1_U15.top_add_34s_34s_34_2_1_Adder_11_U.a [16:0];
assign \add_34s_34s_34_2_1_U15.top_add_34s_34s_34_2_1_Adder_11_U.u1.b  = \add_34s_34s_34_2_1_U15.top_add_34s_34s_34_2_1_Adder_11_U.b [16:0];
assign \add_34s_34s_34_2_1_U15.top_add_34s_34s_34_2_1_Adder_11_U.u1.cin  = 1'h0;
assign \add_34s_34s_34_2_1_U15.top_add_34s_34s_34_2_1_Adder_11_U.facout_s1  = \add_34s_34s_34_2_1_U15.top_add_34s_34s_34_2_1_Adder_11_U.u1.cout ;
assign \add_34s_34s_34_2_1_U15.top_add_34s_34s_34_2_1_Adder_11_U.fas_s1  = \add_34s_34s_34_2_1_U15.top_add_34s_34s_34_2_1_Adder_11_U.u1.s ;
assign \add_34s_34s_34_2_1_U15.top_add_34s_34s_34_2_1_Adder_11_U.a  = \add_34s_34s_34_2_1_U15.din0 ;
assign \add_34s_34s_34_2_1_U15.top_add_34s_34s_34_2_1_Adder_11_U.b  = \add_34s_34s_34_2_1_U15.din1 ;
assign \add_34s_34s_34_2_1_U15.top_add_34s_34s_34_2_1_Adder_11_U.ce  = \add_34s_34s_34_2_1_U15.ce ;
assign \add_34s_34s_34_2_1_U15.top_add_34s_34s_34_2_1_Adder_11_U.clk  = \add_34s_34s_34_2_1_U15.clk ;
assign \add_34s_34s_34_2_1_U15.top_add_34s_34s_34_2_1_Adder_11_U.reset  = \add_34s_34s_34_2_1_U15.reset ;
assign \add_34s_34s_34_2_1_U15.dout  = \add_34s_34s_34_2_1_U15.top_add_34s_34s_34_2_1_Adder_11_U.s ;
assign \add_34s_34s_34_2_1_U15.ce  = 1'h1;
assign \add_34s_34s_34_2_1_U15.clk  = ap_clk;
assign \add_34s_34s_34_2_1_U15.din0  = { op_30_V_reg_986[31], op_30_V_reg_986, 1'h0 };
assign \add_34s_34s_34_2_1_U15.din1  = { op_19_V_reg_980[1], op_19_V_reg_980[1], op_19_V_reg_980[1], op_19_V_reg_980[1], op_19_V_reg_980[1], op_19_V_reg_980[1], op_19_V_reg_980[1], op_19_V_reg_980[1], op_19_V_reg_980[1], op_19_V_reg_980[1], op_19_V_reg_980[1], op_19_V_reg_980[1], op_19_V_reg_980[1], op_19_V_reg_980[1], op_19_V_reg_980[1], op_19_V_reg_980[1], op_19_V_reg_980[1], op_19_V_reg_980[1], op_19_V_reg_980[1], op_19_V_reg_980[1], op_19_V_reg_980[1], op_19_V_reg_980[1], op_19_V_reg_980[1], op_19_V_reg_980[1], op_19_V_reg_980[1], op_19_V_reg_980[1], op_19_V_reg_980[1], op_19_V_reg_980[1], op_19_V_reg_980[1], op_19_V_reg_980[1], op_19_V_reg_980[1], op_19_V_reg_980[1], op_19_V_reg_980 };
assign grp_fu_657_p2 = \add_34s_34s_34_2_1_U15.dout ;
assign \add_34s_34s_34_2_1_U15.reset  = ap_rst;
assign \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_10_U.ain_s0  = \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_10_U.a ;
assign \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_10_U.bin_s0  = \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_10_U.b ;
assign \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_10_U.s  = { \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_10_U.fas_s2 , \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_10_U.sum_s1  };
assign \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_10_U.u2.a  = \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_10_U.ain_s1 ;
assign \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_10_U.u2.b  = \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_10_U.bin_s1 ;
assign \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_10_U.u2.cin  = \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_10_U.carry_s1 ;
assign \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_10_U.facout_s2  = \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_10_U.u2.cout ;
assign \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_10_U.fas_s2  = \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_10_U.u2.s ;
assign \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_10_U.u1.a  = \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_10_U.a [15:0];
assign \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_10_U.u1.b  = \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_10_U.b [15:0];
assign \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_10_U.u1.cin  = 1'h0;
assign \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_10_U.facout_s1  = \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_10_U.u1.cout ;
assign \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_10_U.fas_s1  = \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_10_U.u1.s ;
assign \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_10_U.a  = \add_32s_32ns_32_2_1_U14.din0 ;
assign \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_10_U.b  = \add_32s_32ns_32_2_1_U14.din1 ;
assign \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_10_U.ce  = \add_32s_32ns_32_2_1_U14.ce ;
assign \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_10_U.clk  = \add_32s_32ns_32_2_1_U14.clk ;
assign \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_10_U.reset  = \add_32s_32ns_32_2_1_U14.reset ;
assign \add_32s_32ns_32_2_1_U14.dout  = \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_10_U.s ;
assign \add_32s_32ns_32_2_1_U14.ce  = 1'h1;
assign \add_32s_32ns_32_2_1_U14.clk  = ap_clk;
assign \add_32s_32ns_32_2_1_U14.din0  = { add_ln69_4_reg_964[2], add_ln69_4_reg_964[2], add_ln69_4_reg_964[2], add_ln69_4_reg_964[2], add_ln69_4_reg_964[2], add_ln69_4_reg_964[2], add_ln69_4_reg_964[2], add_ln69_4_reg_964[2], add_ln69_4_reg_964[2], add_ln69_4_reg_964[2], add_ln69_4_reg_964[2], add_ln69_4_reg_964[2], add_ln69_4_reg_964[2], add_ln69_4_reg_964[2], add_ln69_4_reg_964[2], add_ln69_4_reg_964[2], add_ln69_4_reg_964[2], add_ln69_4_reg_964[2], add_ln69_4_reg_964[2], add_ln69_4_reg_964[2], add_ln69_4_reg_964[2], add_ln69_4_reg_964[2], add_ln69_4_reg_964[2], add_ln69_4_reg_964[2], add_ln69_4_reg_964[2], add_ln69_4_reg_964[2], add_ln69_4_reg_964[2], add_ln69_4_reg_964[2], add_ln69_4_reg_964[2], add_ln69_4_reg_964 };
assign \add_32s_32ns_32_2_1_U14.din1  = add_ln69_3_reg_959;
assign grp_fu_612_p2 = \add_32s_32ns_32_2_1_U14.dout ;
assign \add_32s_32ns_32_2_1_U14.reset  = ap_rst;
assign \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.ain_s0  = \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.a ;
assign \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.bin_s0  = \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.b ;
assign \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.s  = { \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.fas_s2 , \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.sum_s1  };
assign \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.u2.a  = \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.ain_s1 ;
assign \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.u2.b  = \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.bin_s1 ;
assign \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.u2.cin  = \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.carry_s1 ;
assign \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.facout_s2  = \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.u2.cout ;
assign \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.fas_s2  = \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.u2.s ;
assign \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.u1.a  = \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.a [15:0];
assign \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.u1.b  = \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.b [15:0];
assign \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.u1.cin  = 1'h0;
assign \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.facout_s1  = \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.u1.cout ;
assign \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.fas_s1  = \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.u1.s ;
assign \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.a  = \add_32ns_32s_32_2_1_U12.din0 ;
assign \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.b  = \add_32ns_32s_32_2_1_U12.din1 ;
assign \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.ce  = \add_32ns_32s_32_2_1_U12.ce ;
assign \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.clk  = \add_32ns_32s_32_2_1_U12.clk ;
assign \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.reset  = \add_32ns_32s_32_2_1_U12.reset ;
assign \add_32ns_32s_32_2_1_U12.dout  = \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.s ;
assign \add_32ns_32s_32_2_1_U12.ce  = 1'h1;
assign \add_32ns_32s_32_2_1_U12.clk  = ap_clk;
assign \add_32ns_32s_32_2_1_U12.din0  = ret_V_19_reg_927;
assign \add_32ns_32s_32_2_1_U12.din1  = { op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16 };
assign grp_fu_575_p2 = \add_32ns_32s_32_2_1_U12.dout ;
assign \add_32ns_32s_32_2_1_U12.reset  = ap_rst;
assign \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s0  = \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.a ;
assign \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s0  = \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.b ;
assign \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.s  = { \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s2 , \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.sum_s1  };
assign \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.a  = \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s1 ;
assign \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.b  = \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s1 ;
assign \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cin  = \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.carry_s1 ;
assign \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s2  = \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cout ;
assign \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s2  = \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.s ;
assign \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.a  = \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.a [15:0];
assign \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.b  = \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.b [15:0];
assign \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cin  = 1'h0;
assign \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s1  = \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cout ;
assign \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s1  = \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.s ;
assign \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.a  = \add_32ns_32ns_32_2_1_U9.din0 ;
assign \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.b  = \add_32ns_32ns_32_2_1_U9.din1 ;
assign \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  = \add_32ns_32ns_32_2_1_U9.ce ;
assign \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.clk  = \add_32ns_32ns_32_2_1_U9.clk ;
assign \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.reset  = \add_32ns_32ns_32_2_1_U9.reset ;
assign \add_32ns_32ns_32_2_1_U9.dout  = \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.s ;
assign \add_32ns_32ns_32_2_1_U9.ce  = 1'h1;
assign \add_32ns_32ns_32_2_1_U9.clk  = ap_clk;
assign \add_32ns_32ns_32_2_1_U9.din0  = ret_V_17_reg_880;
assign \add_32ns_32ns_32_2_1_U9.din1  = select_ln69_reg_885;
assign grp_fu_491_p2 = \add_32ns_32ns_32_2_1_U9.dout ;
assign \add_32ns_32ns_32_2_1_U9.reset  = ap_rst;
assign \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s0  = \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.a ;
assign \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s0  = \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.b ;
assign \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.s  = { \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s2 , \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.sum_s1  };
assign \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.a  = \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s1 ;
assign \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.b  = \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s1 ;
assign \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cin  = \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.carry_s1 ;
assign \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s2  = \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cout ;
assign \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s2  = \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.s ;
assign \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.a  = \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.a [15:0];
assign \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.b  = \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.b [15:0];
assign \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cin  = 1'h0;
assign \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s1  = \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cout ;
assign \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s1  = \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.s ;
assign \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.a  = \add_32ns_32ns_32_2_1_U8.din0 ;
assign \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.b  = \add_32ns_32ns_32_2_1_U8.din1 ;
assign \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  = \add_32ns_32ns_32_2_1_U8.ce ;
assign \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.clk  = \add_32ns_32ns_32_2_1_U8.clk ;
assign \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.reset  = \add_32ns_32ns_32_2_1_U8.reset ;
assign \add_32ns_32ns_32_2_1_U8.dout  = \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.s ;
assign \add_32ns_32ns_32_2_1_U8.ce  = 1'h1;
assign \add_32ns_32ns_32_2_1_U8.clk  = ap_clk;
assign \add_32ns_32ns_32_2_1_U8.din0  = ret_V_6_cast_reg_868;
assign \add_32ns_32ns_32_2_1_U8.din1  = 32'd1;
assign grp_fu_459_p2 = \add_32ns_32ns_32_2_1_U8.dout ;
assign \add_32ns_32ns_32_2_1_U8.reset  = ap_rst;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s0  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.a ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s0  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.b ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.s  = { \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s2 , \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.sum_s1  };
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.a  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s1 ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.b  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s1 ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cin  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.carry_s1 ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s2  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cout ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s2  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.s ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.a  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.a [15:0];
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.b  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.b [15:0];
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cin  = 1'h0;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s1  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cout ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s1  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.s ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.a  = \add_32ns_32ns_32_2_1_U16.din0 ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.b  = \add_32ns_32ns_32_2_1_U16.din1 ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  = \add_32ns_32ns_32_2_1_U16.ce ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.clk  = \add_32ns_32ns_32_2_1_U16.clk ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.reset  = \add_32ns_32ns_32_2_1_U16.reset ;
assign \add_32ns_32ns_32_2_1_U16.dout  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.s ;
assign \add_32ns_32ns_32_2_1_U16.ce  = 1'h1;
assign \add_32ns_32ns_32_2_1_U16.clk  = ap_clk;
assign \add_32ns_32ns_32_2_1_U16.din0  = ret_V_16_cast_reg_1006;
assign \add_32ns_32ns_32_2_1_U16.din1  = 32'd1;
assign grp_fu_673_p2 = \add_32ns_32ns_32_2_1_U16.dout ;
assign \add_32ns_32ns_32_2_1_U16.reset  = ap_rst;
assign \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s0  = \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_6_U.a ;
assign \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s0  = \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_6_U.b ;
assign \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_6_U.s  = { \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s2 , \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_6_U.sum_s1  };
assign \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.a  = \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s1 ;
assign \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.b  = \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s1 ;
assign \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cin  = \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_6_U.carry_s1 ;
assign \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s2  = \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cout ;
assign \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s2  = \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.s ;
assign \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.a  = \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_6_U.a [15:0];
assign \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.b  = \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_6_U.b [15:0];
assign \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cin  = 1'h0;
assign \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s1  = \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cout ;
assign \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s1  = \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.s ;
assign \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_6_U.a  = \add_32ns_32ns_32_2_1_U11.din0 ;
assign \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_6_U.b  = \add_32ns_32ns_32_2_1_U11.din1 ;
assign \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  = \add_32ns_32ns_32_2_1_U11.ce ;
assign \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_6_U.clk  = \add_32ns_32ns_32_2_1_U11.clk ;
assign \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_6_U.reset  = \add_32ns_32ns_32_2_1_U11.reset ;
assign \add_32ns_32ns_32_2_1_U11.dout  = \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_6_U.s ;
assign \add_32ns_32ns_32_2_1_U11.ce  = 1'h1;
assign \add_32ns_32ns_32_2_1_U11.clk  = ap_clk;
assign \add_32ns_32ns_32_2_1_U11.din0  = ret_V_9_cast_reg_915;
assign \add_32ns_32ns_32_2_1_U11.din1  = 32'd1;
assign grp_fu_536_p2 = \add_32ns_32ns_32_2_1_U11.dout ;
assign \add_32ns_32ns_32_2_1_U11.reset  = ap_rst;
assign \add_17s_17s_17_2_1_U1.top_add_17s_17s_17_2_1_Adder_0_U.ain_s0  = \add_17s_17s_17_2_1_U1.top_add_17s_17s_17_2_1_Adder_0_U.a ;
assign \add_17s_17s_17_2_1_U1.top_add_17s_17s_17_2_1_Adder_0_U.bin_s0  = \add_17s_17s_17_2_1_U1.top_add_17s_17s_17_2_1_Adder_0_U.b ;
assign \add_17s_17s_17_2_1_U1.top_add_17s_17s_17_2_1_Adder_0_U.s  = { \add_17s_17s_17_2_1_U1.top_add_17s_17s_17_2_1_Adder_0_U.fas_s2 , \add_17s_17s_17_2_1_U1.top_add_17s_17s_17_2_1_Adder_0_U.sum_s1  };
assign \add_17s_17s_17_2_1_U1.top_add_17s_17s_17_2_1_Adder_0_U.u2.a  = \add_17s_17s_17_2_1_U1.top_add_17s_17s_17_2_1_Adder_0_U.ain_s1 ;
assign \add_17s_17s_17_2_1_U1.top_add_17s_17s_17_2_1_Adder_0_U.u2.b  = \add_17s_17s_17_2_1_U1.top_add_17s_17s_17_2_1_Adder_0_U.bin_s1 ;
assign \add_17s_17s_17_2_1_U1.top_add_17s_17s_17_2_1_Adder_0_U.u2.cin  = \add_17s_17s_17_2_1_U1.top_add_17s_17s_17_2_1_Adder_0_U.carry_s1 ;
assign \add_17s_17s_17_2_1_U1.top_add_17s_17s_17_2_1_Adder_0_U.facout_s2  = \add_17s_17s_17_2_1_U1.top_add_17s_17s_17_2_1_Adder_0_U.u2.cout ;
assign \add_17s_17s_17_2_1_U1.top_add_17s_17s_17_2_1_Adder_0_U.fas_s2  = \add_17s_17s_17_2_1_U1.top_add_17s_17s_17_2_1_Adder_0_U.u2.s ;
assign \add_17s_17s_17_2_1_U1.top_add_17s_17s_17_2_1_Adder_0_U.u1.a  = \add_17s_17s_17_2_1_U1.top_add_17s_17s_17_2_1_Adder_0_U.a [7:0];
assign \add_17s_17s_17_2_1_U1.top_add_17s_17s_17_2_1_Adder_0_U.u1.b  = \add_17s_17s_17_2_1_U1.top_add_17s_17s_17_2_1_Adder_0_U.b [7:0];
assign \add_17s_17s_17_2_1_U1.top_add_17s_17s_17_2_1_Adder_0_U.u1.cin  = 1'h0;
assign \add_17s_17s_17_2_1_U1.top_add_17s_17s_17_2_1_Adder_0_U.facout_s1  = \add_17s_17s_17_2_1_U1.top_add_17s_17s_17_2_1_Adder_0_U.u1.cout ;
assign \add_17s_17s_17_2_1_U1.top_add_17s_17s_17_2_1_Adder_0_U.fas_s1  = \add_17s_17s_17_2_1_U1.top_add_17s_17s_17_2_1_Adder_0_U.u1.s ;
assign \add_17s_17s_17_2_1_U1.top_add_17s_17s_17_2_1_Adder_0_U.a  = \add_17s_17s_17_2_1_U1.din0 ;
assign \add_17s_17s_17_2_1_U1.top_add_17s_17s_17_2_1_Adder_0_U.b  = \add_17s_17s_17_2_1_U1.din1 ;
assign \add_17s_17s_17_2_1_U1.top_add_17s_17s_17_2_1_Adder_0_U.ce  = \add_17s_17s_17_2_1_U1.ce ;
assign \add_17s_17s_17_2_1_U1.top_add_17s_17s_17_2_1_Adder_0_U.clk  = \add_17s_17s_17_2_1_U1.clk ;
assign \add_17s_17s_17_2_1_U1.top_add_17s_17s_17_2_1_Adder_0_U.reset  = \add_17s_17s_17_2_1_U1.reset ;
assign \add_17s_17s_17_2_1_U1.dout  = \add_17s_17s_17_2_1_U1.top_add_17s_17s_17_2_1_Adder_0_U.s ;
assign \add_17s_17s_17_2_1_U1.ce  = 1'h1;
assign \add_17s_17s_17_2_1_U1.clk  = ap_clk;
assign \add_17s_17s_17_2_1_U1.din0  = { op_0[7], op_0[7], op_0, 7'h00 };
assign \add_17s_17s_17_2_1_U1.din1  = { op_1[15], op_1 };
assign grp_fu_221_p2 = \add_17s_17s_17_2_1_U1.dout ;
assign \add_17s_17s_17_2_1_U1.reset  = ap_rst;
assign \add_11s_11ns_11_2_1_U5.top_add_11s_11ns_11_2_1_Adder_2_U.ain_s0  = \add_11s_11ns_11_2_1_U5.top_add_11s_11ns_11_2_1_Adder_2_U.a ;
assign \add_11s_11ns_11_2_1_U5.top_add_11s_11ns_11_2_1_Adder_2_U.bin_s0  = \add_11s_11ns_11_2_1_U5.top_add_11s_11ns_11_2_1_Adder_2_U.b ;
assign \add_11s_11ns_11_2_1_U5.top_add_11s_11ns_11_2_1_Adder_2_U.s  = { \add_11s_11ns_11_2_1_U5.top_add_11s_11ns_11_2_1_Adder_2_U.fas_s2 , \add_11s_11ns_11_2_1_U5.top_add_11s_11ns_11_2_1_Adder_2_U.sum_s1  };
assign \add_11s_11ns_11_2_1_U5.top_add_11s_11ns_11_2_1_Adder_2_U.u2.a  = \add_11s_11ns_11_2_1_U5.top_add_11s_11ns_11_2_1_Adder_2_U.ain_s1 ;
assign \add_11s_11ns_11_2_1_U5.top_add_11s_11ns_11_2_1_Adder_2_U.u2.b  = \add_11s_11ns_11_2_1_U5.top_add_11s_11ns_11_2_1_Adder_2_U.bin_s1 ;
assign \add_11s_11ns_11_2_1_U5.top_add_11s_11ns_11_2_1_Adder_2_U.u2.cin  = \add_11s_11ns_11_2_1_U5.top_add_11s_11ns_11_2_1_Adder_2_U.carry_s1 ;
assign \add_11s_11ns_11_2_1_U5.top_add_11s_11ns_11_2_1_Adder_2_U.facout_s2  = \add_11s_11ns_11_2_1_U5.top_add_11s_11ns_11_2_1_Adder_2_U.u2.cout ;
assign \add_11s_11ns_11_2_1_U5.top_add_11s_11ns_11_2_1_Adder_2_U.fas_s2  = \add_11s_11ns_11_2_1_U5.top_add_11s_11ns_11_2_1_Adder_2_U.u2.s ;
assign \add_11s_11ns_11_2_1_U5.top_add_11s_11ns_11_2_1_Adder_2_U.u1.a  = \add_11s_11ns_11_2_1_U5.top_add_11s_11ns_11_2_1_Adder_2_U.a [4:0];
assign \add_11s_11ns_11_2_1_U5.top_add_11s_11ns_11_2_1_Adder_2_U.u1.b  = \add_11s_11ns_11_2_1_U5.top_add_11s_11ns_11_2_1_Adder_2_U.b [4:0];
assign \add_11s_11ns_11_2_1_U5.top_add_11s_11ns_11_2_1_Adder_2_U.u1.cin  = 1'h0;
assign \add_11s_11ns_11_2_1_U5.top_add_11s_11ns_11_2_1_Adder_2_U.facout_s1  = \add_11s_11ns_11_2_1_U5.top_add_11s_11ns_11_2_1_Adder_2_U.u1.cout ;
assign \add_11s_11ns_11_2_1_U5.top_add_11s_11ns_11_2_1_Adder_2_U.fas_s1  = \add_11s_11ns_11_2_1_U5.top_add_11s_11ns_11_2_1_Adder_2_U.u1.s ;
assign \add_11s_11ns_11_2_1_U5.top_add_11s_11ns_11_2_1_Adder_2_U.a  = \add_11s_11ns_11_2_1_U5.din0 ;
assign \add_11s_11ns_11_2_1_U5.top_add_11s_11ns_11_2_1_Adder_2_U.b  = \add_11s_11ns_11_2_1_U5.din1 ;
assign \add_11s_11ns_11_2_1_U5.top_add_11s_11ns_11_2_1_Adder_2_U.ce  = \add_11s_11ns_11_2_1_U5.ce ;
assign \add_11s_11ns_11_2_1_U5.top_add_11s_11ns_11_2_1_Adder_2_U.clk  = \add_11s_11ns_11_2_1_U5.clk ;
assign \add_11s_11ns_11_2_1_U5.top_add_11s_11ns_11_2_1_Adder_2_U.reset  = \add_11s_11ns_11_2_1_U5.reset ;
assign \add_11s_11ns_11_2_1_U5.dout  = \add_11s_11ns_11_2_1_U5.top_add_11s_11ns_11_2_1_Adder_2_U.s ;
assign \add_11s_11ns_11_2_1_U5.ce  = 1'h1;
assign \add_11s_11ns_11_2_1_U5.clk  = ap_clk;
assign \add_11s_11ns_11_2_1_U5.din0  = { add_ln69_reg_775[9], add_ln69_reg_775 };
assign \add_11s_11ns_11_2_1_U5.din1  = ret_V_14_reg_770;
assign grp_fu_339_p2 = \add_11s_11ns_11_2_1_U5.dout ;
assign \add_11s_11ns_11_2_1_U5.reset  = ap_rst;
assign \add_11s_11ns_11_2_1_U3.top_add_11s_11ns_11_2_1_Adder_2_U.ain_s0  = \add_11s_11ns_11_2_1_U3.top_add_11s_11ns_11_2_1_Adder_2_U.a ;
assign \add_11s_11ns_11_2_1_U3.top_add_11s_11ns_11_2_1_Adder_2_U.bin_s0  = \add_11s_11ns_11_2_1_U3.top_add_11s_11ns_11_2_1_Adder_2_U.b ;
assign \add_11s_11ns_11_2_1_U3.top_add_11s_11ns_11_2_1_Adder_2_U.s  = { \add_11s_11ns_11_2_1_U3.top_add_11s_11ns_11_2_1_Adder_2_U.fas_s2 , \add_11s_11ns_11_2_1_U3.top_add_11s_11ns_11_2_1_Adder_2_U.sum_s1  };
assign \add_11s_11ns_11_2_1_U3.top_add_11s_11ns_11_2_1_Adder_2_U.u2.a  = \add_11s_11ns_11_2_1_U3.top_add_11s_11ns_11_2_1_Adder_2_U.ain_s1 ;
assign \add_11s_11ns_11_2_1_U3.top_add_11s_11ns_11_2_1_Adder_2_U.u2.b  = \add_11s_11ns_11_2_1_U3.top_add_11s_11ns_11_2_1_Adder_2_U.bin_s1 ;
assign \add_11s_11ns_11_2_1_U3.top_add_11s_11ns_11_2_1_Adder_2_U.u2.cin  = \add_11s_11ns_11_2_1_U3.top_add_11s_11ns_11_2_1_Adder_2_U.carry_s1 ;
assign \add_11s_11ns_11_2_1_U3.top_add_11s_11ns_11_2_1_Adder_2_U.facout_s2  = \add_11s_11ns_11_2_1_U3.top_add_11s_11ns_11_2_1_Adder_2_U.u2.cout ;
assign \add_11s_11ns_11_2_1_U3.top_add_11s_11ns_11_2_1_Adder_2_U.fas_s2  = \add_11s_11ns_11_2_1_U3.top_add_11s_11ns_11_2_1_Adder_2_U.u2.s ;
assign \add_11s_11ns_11_2_1_U3.top_add_11s_11ns_11_2_1_Adder_2_U.u1.a  = \add_11s_11ns_11_2_1_U3.top_add_11s_11ns_11_2_1_Adder_2_U.a [4:0];
assign \add_11s_11ns_11_2_1_U3.top_add_11s_11ns_11_2_1_Adder_2_U.u1.b  = \add_11s_11ns_11_2_1_U3.top_add_11s_11ns_11_2_1_Adder_2_U.b [4:0];
assign \add_11s_11ns_11_2_1_U3.top_add_11s_11ns_11_2_1_Adder_2_U.u1.cin  = 1'h0;
assign \add_11s_11ns_11_2_1_U3.top_add_11s_11ns_11_2_1_Adder_2_U.facout_s1  = \add_11s_11ns_11_2_1_U3.top_add_11s_11ns_11_2_1_Adder_2_U.u1.cout ;
assign \add_11s_11ns_11_2_1_U3.top_add_11s_11ns_11_2_1_Adder_2_U.fas_s1  = \add_11s_11ns_11_2_1_U3.top_add_11s_11ns_11_2_1_Adder_2_U.u1.s ;
assign \add_11s_11ns_11_2_1_U3.top_add_11s_11ns_11_2_1_Adder_2_U.a  = \add_11s_11ns_11_2_1_U3.din0 ;
assign \add_11s_11ns_11_2_1_U3.top_add_11s_11ns_11_2_1_Adder_2_U.b  = \add_11s_11ns_11_2_1_U3.din1 ;
assign \add_11s_11ns_11_2_1_U3.top_add_11s_11ns_11_2_1_Adder_2_U.ce  = \add_11s_11ns_11_2_1_U3.ce ;
assign \add_11s_11ns_11_2_1_U3.top_add_11s_11ns_11_2_1_Adder_2_U.clk  = \add_11s_11ns_11_2_1_U3.clk ;
assign \add_11s_11ns_11_2_1_U3.top_add_11s_11ns_11_2_1_Adder_2_U.reset  = \add_11s_11ns_11_2_1_U3.reset ;
assign \add_11s_11ns_11_2_1_U3.dout  = \add_11s_11ns_11_2_1_U3.top_add_11s_11ns_11_2_1_Adder_2_U.s ;
assign \add_11s_11ns_11_2_1_U3.ce  = 1'h1;
assign \add_11s_11ns_11_2_1_U3.clk  = ap_clk;
assign \add_11s_11ns_11_2_1_U3.din0  = { ret_V_13_reg_740[9], ret_V_13_reg_740 };
assign \add_11s_11ns_11_2_1_U3.din1  = select_ln1192_reg_750;
assign grp_fu_290_p2 = \add_11s_11ns_11_2_1_U3.dout ;
assign \add_11s_11ns_11_2_1_U3.reset  = ap_rst;
assign \add_11ns_11ns_11_2_1_U6.top_add_11ns_11ns_11_2_1_Adder_4_U.ain_s0  = \add_11ns_11ns_11_2_1_U6.top_add_11ns_11ns_11_2_1_Adder_4_U.a ;
assign \add_11ns_11ns_11_2_1_U6.top_add_11ns_11ns_11_2_1_Adder_4_U.bin_s0  = \add_11ns_11ns_11_2_1_U6.top_add_11ns_11ns_11_2_1_Adder_4_U.b ;
assign \add_11ns_11ns_11_2_1_U6.top_add_11ns_11ns_11_2_1_Adder_4_U.s  = { \add_11ns_11ns_11_2_1_U6.top_add_11ns_11ns_11_2_1_Adder_4_U.fas_s2 , \add_11ns_11ns_11_2_1_U6.top_add_11ns_11ns_11_2_1_Adder_4_U.sum_s1  };
assign \add_11ns_11ns_11_2_1_U6.top_add_11ns_11ns_11_2_1_Adder_4_U.u2.a  = \add_11ns_11ns_11_2_1_U6.top_add_11ns_11ns_11_2_1_Adder_4_U.ain_s1 ;
assign \add_11ns_11ns_11_2_1_U6.top_add_11ns_11ns_11_2_1_Adder_4_U.u2.b  = \add_11ns_11ns_11_2_1_U6.top_add_11ns_11ns_11_2_1_Adder_4_U.bin_s1 ;
assign \add_11ns_11ns_11_2_1_U6.top_add_11ns_11ns_11_2_1_Adder_4_U.u2.cin  = \add_11ns_11ns_11_2_1_U6.top_add_11ns_11ns_11_2_1_Adder_4_U.carry_s1 ;
assign \add_11ns_11ns_11_2_1_U6.top_add_11ns_11ns_11_2_1_Adder_4_U.facout_s2  = \add_11ns_11ns_11_2_1_U6.top_add_11ns_11ns_11_2_1_Adder_4_U.u2.cout ;
assign \add_11ns_11ns_11_2_1_U6.top_add_11ns_11ns_11_2_1_Adder_4_U.fas_s2  = \add_11ns_11ns_11_2_1_U6.top_add_11ns_11ns_11_2_1_Adder_4_U.u2.s ;
assign \add_11ns_11ns_11_2_1_U6.top_add_11ns_11ns_11_2_1_Adder_4_U.u1.a  = \add_11ns_11ns_11_2_1_U6.top_add_11ns_11ns_11_2_1_Adder_4_U.a [4:0];
assign \add_11ns_11ns_11_2_1_U6.top_add_11ns_11ns_11_2_1_Adder_4_U.u1.b  = \add_11ns_11ns_11_2_1_U6.top_add_11ns_11ns_11_2_1_Adder_4_U.b [4:0];
assign \add_11ns_11ns_11_2_1_U6.top_add_11ns_11ns_11_2_1_Adder_4_U.u1.cin  = 1'h0;
assign \add_11ns_11ns_11_2_1_U6.top_add_11ns_11ns_11_2_1_Adder_4_U.facout_s1  = \add_11ns_11ns_11_2_1_U6.top_add_11ns_11ns_11_2_1_Adder_4_U.u1.cout ;
assign \add_11ns_11ns_11_2_1_U6.top_add_11ns_11ns_11_2_1_Adder_4_U.fas_s1  = \add_11ns_11ns_11_2_1_U6.top_add_11ns_11ns_11_2_1_Adder_4_U.u1.s ;
assign \add_11ns_11ns_11_2_1_U6.top_add_11ns_11ns_11_2_1_Adder_4_U.a  = \add_11ns_11ns_11_2_1_U6.din0 ;
assign \add_11ns_11ns_11_2_1_U6.top_add_11ns_11ns_11_2_1_Adder_4_U.b  = \add_11ns_11ns_11_2_1_U6.din1 ;
assign \add_11ns_11ns_11_2_1_U6.top_add_11ns_11ns_11_2_1_Adder_4_U.ce  = \add_11ns_11ns_11_2_1_U6.ce ;
assign \add_11ns_11ns_11_2_1_U6.top_add_11ns_11ns_11_2_1_Adder_4_U.clk  = \add_11ns_11ns_11_2_1_U6.clk ;
assign \add_11ns_11ns_11_2_1_U6.top_add_11ns_11ns_11_2_1_Adder_4_U.reset  = \add_11ns_11ns_11_2_1_U6.reset ;
assign \add_11ns_11ns_11_2_1_U6.dout  = \add_11ns_11ns_11_2_1_U6.top_add_11ns_11ns_11_2_1_Adder_4_U.s ;
assign \add_11ns_11ns_11_2_1_U6.ce  = 1'h1;
assign \add_11ns_11ns_11_2_1_U6.clk  = ap_clk;
assign \add_11ns_11ns_11_2_1_U6.din0  = { 10'h000, lhs_V_reg_818 };
assign \add_11ns_11ns_11_2_1_U6.din1  = op_23_V_reg_813;
assign grp_fu_379_p2 = \add_11ns_11ns_11_2_1_U6.dout ;
assign \add_11ns_11ns_11_2_1_U6.reset  = ap_rst;
assign \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.ain_s0  = \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.a ;
assign \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.bin_s0  = \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.b ;
assign \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.s  = { \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.fas_s2 , \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.sum_s1  };
assign \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.u2.a  = \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.ain_s1 ;
assign \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.u2.b  = \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.bin_s1 ;
assign \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.u2.cin  = \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.carry_s1 ;
assign \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.facout_s2  = \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.u2.cout ;
assign \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.fas_s2  = \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.u2.s ;
assign \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.u1.a  = \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.a [4:0];
assign \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.u1.b  = \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.b [4:0];
assign \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.u1.cin  = 1'h0;
assign \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.facout_s1  = \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.u1.cout ;
assign \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.fas_s1  = \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.u1.s ;
assign \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.a  = \add_10ns_10s_10_2_1_U4.din0 ;
assign \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.b  = \add_10ns_10s_10_2_1_U4.din1 ;
assign \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.ce  = \add_10ns_10s_10_2_1_U4.ce ;
assign \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.clk  = \add_10ns_10s_10_2_1_U4.clk ;
assign \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.reset  = \add_10ns_10s_10_2_1_U4.reset ;
assign \add_10ns_10s_10_2_1_U4.dout  = \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.s ;
assign \add_10ns_10s_10_2_1_U4.ce  = 1'h1;
assign \add_10ns_10s_10_2_1_U4.clk  = ap_clk;
assign \add_10ns_10s_10_2_1_U4.din0  = { 2'h0, ret_reg_745[1], ret_reg_745[1], ret_reg_745[1], ret_reg_745[1], ret_reg_745[1], ret_reg_745[1], ret_reg_745 };
assign \add_10ns_10s_10_2_1_U4.din1  = { op_10[3], op_10[3], op_10[3], op_10[3], op_10[3], op_10[3], op_10 };
assign grp_fu_306_p2 = \add_10ns_10s_10_2_1_U4.dout ;
assign \add_10ns_10s_10_2_1_U4.reset  = ap_rst;
assign \add_10ns_10ns_10_2_1_U2.top_add_10ns_10ns_10_2_1_Adder_1_U.ain_s0  = \add_10ns_10ns_10_2_1_U2.top_add_10ns_10ns_10_2_1_Adder_1_U.a ;
assign \add_10ns_10ns_10_2_1_U2.top_add_10ns_10ns_10_2_1_Adder_1_U.bin_s0  = \add_10ns_10ns_10_2_1_U2.top_add_10ns_10ns_10_2_1_Adder_1_U.b ;
assign \add_10ns_10ns_10_2_1_U2.top_add_10ns_10ns_10_2_1_Adder_1_U.s  = { \add_10ns_10ns_10_2_1_U2.top_add_10ns_10ns_10_2_1_Adder_1_U.fas_s2 , \add_10ns_10ns_10_2_1_U2.top_add_10ns_10ns_10_2_1_Adder_1_U.sum_s1  };
assign \add_10ns_10ns_10_2_1_U2.top_add_10ns_10ns_10_2_1_Adder_1_U.u2.a  = \add_10ns_10ns_10_2_1_U2.top_add_10ns_10ns_10_2_1_Adder_1_U.ain_s1 ;
assign \add_10ns_10ns_10_2_1_U2.top_add_10ns_10ns_10_2_1_Adder_1_U.u2.b  = \add_10ns_10ns_10_2_1_U2.top_add_10ns_10ns_10_2_1_Adder_1_U.bin_s1 ;
assign \add_10ns_10ns_10_2_1_U2.top_add_10ns_10ns_10_2_1_Adder_1_U.u2.cin  = \add_10ns_10ns_10_2_1_U2.top_add_10ns_10ns_10_2_1_Adder_1_U.carry_s1 ;
assign \add_10ns_10ns_10_2_1_U2.top_add_10ns_10ns_10_2_1_Adder_1_U.facout_s2  = \add_10ns_10ns_10_2_1_U2.top_add_10ns_10ns_10_2_1_Adder_1_U.u2.cout ;
assign \add_10ns_10ns_10_2_1_U2.top_add_10ns_10ns_10_2_1_Adder_1_U.fas_s2  = \add_10ns_10ns_10_2_1_U2.top_add_10ns_10ns_10_2_1_Adder_1_U.u2.s ;
assign \add_10ns_10ns_10_2_1_U2.top_add_10ns_10ns_10_2_1_Adder_1_U.u1.a  = \add_10ns_10ns_10_2_1_U2.top_add_10ns_10ns_10_2_1_Adder_1_U.a [4:0];
assign \add_10ns_10ns_10_2_1_U2.top_add_10ns_10ns_10_2_1_Adder_1_U.u1.b  = \add_10ns_10ns_10_2_1_U2.top_add_10ns_10ns_10_2_1_Adder_1_U.b [4:0];
assign \add_10ns_10ns_10_2_1_U2.top_add_10ns_10ns_10_2_1_Adder_1_U.u1.cin  = 1'h0;
assign \add_10ns_10ns_10_2_1_U2.top_add_10ns_10ns_10_2_1_Adder_1_U.facout_s1  = \add_10ns_10ns_10_2_1_U2.top_add_10ns_10ns_10_2_1_Adder_1_U.u1.cout ;
assign \add_10ns_10ns_10_2_1_U2.top_add_10ns_10ns_10_2_1_Adder_1_U.fas_s1  = \add_10ns_10ns_10_2_1_U2.top_add_10ns_10ns_10_2_1_Adder_1_U.u1.s ;
assign \add_10ns_10ns_10_2_1_U2.top_add_10ns_10ns_10_2_1_Adder_1_U.a  = \add_10ns_10ns_10_2_1_U2.din0 ;
assign \add_10ns_10ns_10_2_1_U2.top_add_10ns_10ns_10_2_1_Adder_1_U.b  = \add_10ns_10ns_10_2_1_U2.din1 ;
assign \add_10ns_10ns_10_2_1_U2.top_add_10ns_10ns_10_2_1_Adder_1_U.ce  = \add_10ns_10ns_10_2_1_U2.ce ;
assign \add_10ns_10ns_10_2_1_U2.top_add_10ns_10ns_10_2_1_Adder_1_U.clk  = \add_10ns_10ns_10_2_1_U2.clk ;
assign \add_10ns_10ns_10_2_1_U2.top_add_10ns_10ns_10_2_1_Adder_1_U.reset  = \add_10ns_10ns_10_2_1_U2.reset ;
assign \add_10ns_10ns_10_2_1_U2.dout  = \add_10ns_10ns_10_2_1_U2.top_add_10ns_10ns_10_2_1_Adder_1_U.s ;
assign \add_10ns_10ns_10_2_1_U2.ce  = 1'h1;
assign \add_10ns_10ns_10_2_1_U2.clk  = ap_clk;
assign \add_10ns_10ns_10_2_1_U2.din0  = ret_V_reg_722;
assign \add_10ns_10ns_10_2_1_U2.din1  = 10'h001;
assign grp_fu_247_p2 = \add_10ns_10ns_10_2_1_U2.dout ;
assign \add_10ns_10ns_10_2_1_U2.reset  = ap_rst;
endmodule


// Product machine:
module top_A_times_top_B (ap_start, op_0, op_1, op_10, op_11, op_14, op_15, op_16, op_17, op_2, op_3, op_4, op_8, ap_clk, unsafe_signal);
input ap_start;
input [7:0] op_0;
input [15:0] op_1;
input [3:0] op_10;
input op_11;
input op_14;
input [7:0] op_15;
input [3:0] op_16;
input [1:0] op_17;
input op_2;
input [1:0] op_3;
input [1:0] op_4;
input [1:0] op_8;
input ap_clk;
output unsafe_signal;
reg _setup;
initial _setup = 1'b0;
always @ (posedge ap_clk) _setup <= 1'b1;
reg ap_start_internal;
always @ (posedge ap_clk) if (!_setup) ap_start_internal <= ap_start;
reg [7:0] op_0_internal;
always @ (posedge ap_clk) if (!_setup) op_0_internal <= op_0;
reg [15:0] op_1_internal;
always @ (posedge ap_clk) if (!_setup) op_1_internal <= op_1;
reg [3:0] op_10_internal;
always @ (posedge ap_clk) if (!_setup) op_10_internal <= op_10;
reg op_11_internal;
always @ (posedge ap_clk) if (!_setup) op_11_internal <= op_11;
reg op_14_internal;
always @ (posedge ap_clk) if (!_setup) op_14_internal <= op_14;
reg [7:0] op_15_internal;
always @ (posedge ap_clk) if (!_setup) op_15_internal <= op_15;
reg [3:0] op_16_internal;
always @ (posedge ap_clk) if (!_setup) op_16_internal <= op_16;
reg [1:0] op_17_internal;
always @ (posedge ap_clk) if (!_setup) op_17_internal <= op_17;
reg op_2_internal;
always @ (posedge ap_clk) if (!_setup) op_2_internal <= op_2;
reg [1:0] op_3_internal;
always @ (posedge ap_clk) if (!_setup) op_3_internal <= op_3;
reg [1:0] op_4_internal;
always @ (posedge ap_clk) if (!_setup) op_4_internal <= op_4;
reg [1:0] op_8_internal;
always @ (posedge ap_clk) if (!_setup) op_8_internal <= op_8;
wire ap_done_A;
wire ap_done_B;
wire ap_done_eq;
assign ap_done_eq = ap_done_A == ap_done_B;
wire ap_idle_A;
wire ap_idle_B;
wire ap_idle_eq;
assign ap_idle_eq = ap_idle_A == ap_idle_B;
wire ap_ready_A;
wire ap_ready_B;
wire ap_ready_eq;
assign ap_ready_eq = ap_ready_A == ap_ready_B;
wire [31:0] op_31_A;
wire [31:0] op_31_B;
wire op_31_eq;
assign op_31_eq = op_31_A == op_31_B;
wire op_31_ap_vld_A;
wire op_31_ap_vld_B;
wire clk_enable_A;
wire clk_enable_B;
assign clk_enable_A = _setup & (~op_31_ap_vld_A | op_31_ap_vld_B);
assign clk_enable_B = _setup;
wire divergent;
assign divergent = ~(ap_done_eq & ap_idle_eq & ap_ready_eq & op_31_eq);
assign unsafe_signal = op_31_ap_vld_A & op_31_ap_vld_B & divergent;
top_A instance_A (
    .ap_clk(ap_clk),
    .clk_enable(clk_enable_A),
    .ap_start(ap_start_internal),
    .op_0(op_0_internal),
    .op_1(op_1_internal),
    .op_10(op_10_internal),
    .op_11(op_11_internal),
    .op_14(op_14_internal),
    .op_15(op_15_internal),
    .op_16(op_16_internal),
    .op_17(op_17_internal),
    .op_2(op_2_internal),
    .op_3(op_3_internal),
    .op_4(op_4_internal),
    .op_8(op_8_internal),
    .ap_done(ap_done_A),
    .ap_idle(ap_idle_A),
    .ap_ready(ap_ready_A),
    .op_31(op_31_A),
    .op_31_ap_vld(op_31_ap_vld_A)
);
top_B instance_B (
    .ap_clk(ap_clk),
    .clk_enable(clk_enable_B),
    .ap_start(ap_start_internal),
    .op_0(op_0_internal),
    .op_1(op_1_internal),
    .op_10(op_10_internal),
    .op_11(op_11_internal),
    .op_14(op_14_internal),
    .op_15(op_15_internal),
    .op_16(op_16_internal),
    .op_17(op_17_internal),
    .op_2(op_2_internal),
    .op_3(op_3_internal),
    .op_4(op_4_internal),
    .op_8(op_8_internal),
    .ap_done(ap_done_B),
    .ap_idle(ap_idle_B),
    .ap_ready(ap_ready_B),
    .op_31(op_31_B),
    .op_31_ap_vld(op_31_ap_vld_B)
);
endmodule
