// Processed by function `construct_kairos` in `verilog_tricks.py`.
// Machine A:
// Processed by function `add_clk_enable_signal` in `verilog_tricks.py`.
// Processed by function `remove_reset_signal` in `verilog_tricks.py`.
module top_A (
  ap_clk,
  ap_start,
  ap_done,
  ap_idle,
  ap_ready,
  op_0,
  op_1,
  op_3,
  op_4,
  op_11,
  op_12,
  op_15,
  op_17,
  op_18,
  op_19,
  op_31,
  op_31_ap_vld,
clk_enable
);
input clk_enable;


input ap_clk;
wire ap_rst;
assign ap_rst = op_31_ap_vld;
input ap_start;
input [7:0] op_0;
input [3:0] op_1;
input [3:0] op_11;
input [3:0] op_12;
input [3:0] op_15;
input [3:0] op_17;
input [1:0] op_18;
input [3:0] op_19;
input op_3;
input [1:0] op_4;
output ap_done;
output ap_idle;
output ap_ready;
output [31:0] op_31;
output op_31_ap_vld;


reg \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_6_U.ain_s1 ;
reg \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_6_U.bin_s1 ;
reg \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_6_U.carry_s1 ;
reg \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_6_U.sum_s1 ;
reg \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.ain_s1 ;
reg \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.bin_s1 ;
reg \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.carry_s1 ;
reg \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.sum_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_13_U.ain_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_13_U.bin_s1 ;
reg \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_13_U.carry_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_13_U.sum_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_13_U.ain_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_13_U.bin_s1 ;
reg \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_13_U.carry_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_13_U.sum_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_13_U.ain_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_13_U.bin_s1 ;
reg \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_13_U.carry_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_13_U.sum_s1 ;
reg [15:0] \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_15_U.ain_s1 ;
reg [15:0] \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_15_U.bin_s1 ;
reg \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_15_U.carry_s1 ;
reg [15:0] \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_15_U.sum_s1 ;
reg [15:0] \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_15_U.ain_s1 ;
reg [15:0] \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_15_U.bin_s1 ;
reg \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_15_U.carry_s1 ;
reg [15:0] \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_15_U.sum_s1 ;
reg [17:0] \add_35s_35s_35_2_1_U17.top_add_35s_35s_35_2_1_Adder_12_U.ain_s1 ;
reg [17:0] \add_35s_35s_35_2_1_U17.top_add_35s_35s_35_2_1_Adder_12_U.bin_s1 ;
reg \add_35s_35s_35_2_1_U17.top_add_35s_35s_35_2_1_Adder_12_U.carry_s1 ;
reg [16:0] \add_35s_35s_35_2_1_U17.top_add_35s_35s_35_2_1_Adder_12_U.sum_s1 ;
reg [17:0] \add_36s_36s_36_2_1_U20.top_add_36s_36s_36_2_1_Adder_14_U.ain_s1 ;
reg [17:0] \add_36s_36s_36_2_1_U20.top_add_36s_36s_36_2_1_Adder_14_U.bin_s1 ;
reg \add_36s_36s_36_2_1_U20.top_add_36s_36s_36_2_1_Adder_14_U.carry_s1 ;
reg [17:0] \add_36s_36s_36_2_1_U20.top_add_36s_36s_36_2_1_Adder_14_U.sum_s1 ;
reg [1:0] \add_3s_3s_3_2_1_U15.top_add_3s_3s_3_2_1_Adder_11_U.ain_s1 ;
reg [1:0] \add_3s_3s_3_2_1_U15.top_add_3s_3s_3_2_1_Adder_11_U.bin_s1 ;
reg \add_3s_3s_3_2_1_U15.top_add_3s_3s_3_2_1_Adder_11_U.carry_s1 ;
reg \add_3s_3s_3_2_1_U15.top_add_3s_3s_3_2_1_Adder_11_U.sum_s1 ;
reg [1:0] \add_4s_4ns_4_2_1_U8.top_add_4s_4ns_4_2_1_Adder_5_U.ain_s1 ;
reg [1:0] \add_4s_4ns_4_2_1_U8.top_add_4s_4ns_4_2_1_Adder_5_U.bin_s1 ;
reg \add_4s_4ns_4_2_1_U8.top_add_4s_4ns_4_2_1_Adder_5_U.carry_s1 ;
reg [1:0] \add_4s_4ns_4_2_1_U8.top_add_4s_4ns_4_2_1_Adder_5_U.sum_s1 ;
reg [2:0] \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_4_U.ain_s1 ;
reg [2:0] \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_4_U.bin_s1 ;
reg \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_4_U.carry_s1 ;
reg [2:0] \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_4_U.sum_s1 ;
reg [2:0] \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.ain_s1 ;
reg [2:0] \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.bin_s1 ;
reg \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.carry_s1 ;
reg [2:0] \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.sum_s1 ;
reg [3:0] \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_10_U.ain_s1 ;
reg [3:0] \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_10_U.bin_s1 ;
reg \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_10_U.carry_s1 ;
reg [2:0] \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_10_U.sum_s1 ;
reg [3:0] \add_7s_7ns_7_2_1_U16.top_add_7s_7ns_7_2_1_Adder_10_U.ain_s1 ;
reg [3:0] \add_7s_7ns_7_2_1_U16.top_add_7s_7ns_7_2_1_Adder_10_U.bin_s1 ;
reg \add_7s_7ns_7_2_1_U16.top_add_7s_7ns_7_2_1_Adder_10_U.carry_s1 ;
reg [2:0] \add_7s_7ns_7_2_1_U16.top_add_7s_7ns_7_2_1_Adder_10_U.sum_s1 ;
reg [3:0] \add_7s_7s_7_2_1_U11.top_add_7s_7s_7_2_1_Adder_8_U.ain_s1 ;
reg [3:0] \add_7s_7s_7_2_1_U11.top_add_7s_7s_7_2_1_Adder_8_U.bin_s1 ;
reg \add_7s_7s_7_2_1_U11.top_add_7s_7s_7_2_1_Adder_8_U.carry_s1 ;
reg [2:0] \add_7s_7s_7_2_1_U11.top_add_7s_7s_7_2_1_Adder_8_U.sum_s1 ;
reg [4:0] \add_9s_9ns_9_2_1_U6.top_add_9s_9ns_9_2_1_Adder_3_U.ain_s1 ;
reg [4:0] \add_9s_9ns_9_2_1_U6.top_add_9s_9ns_9_2_1_Adder_3_U.bin_s1 ;
reg \add_9s_9ns_9_2_1_U6.top_add_9s_9ns_9_2_1_Adder_3_U.carry_s1 ;
reg [3:0] \add_9s_9ns_9_2_1_U6.top_add_9s_9ns_9_2_1_Adder_3_U.sum_s1 ;
reg [31:0] add_ln691_1_reg_1377;
reg [31:0] add_ln691_reg_1330;
reg [6:0] add_ln69_1_reg_1267;
reg [1:0] add_ln69_2_reg_1247;
reg [2:0] add_ln69_3_reg_1272;
reg [5:0] add_ln69_reg_1242;
reg and_ln410_reg_1124;
reg [37:0] ap_CS_fsm = 38'h0000000001;
reg [1:0] \ashr_4s_2ns_4_7_1_U3.din1_cast_array[0] ;
reg [1:0] \ashr_4s_2ns_4_7_1_U3.din1_cast_array[1] ;
reg [1:0] \ashr_4s_2ns_4_7_1_U3.din1_cast_array[2] ;
reg [1:0] \ashr_4s_2ns_4_7_1_U3.din1_cast_array[3] ;
reg [1:0] \ashr_4s_2ns_4_7_1_U3.din1_cast_array[4] ;
reg [1:0] \ashr_4s_2ns_4_7_1_U3.din1_cast_array[5] ;
reg [3:0] \ashr_4s_2ns_4_7_1_U3.dout_array[0] ;
reg [3:0] \ashr_4s_2ns_4_7_1_U3.dout_array[1] ;
reg [3:0] \ashr_4s_2ns_4_7_1_U3.dout_array[2] ;
reg [3:0] \ashr_4s_2ns_4_7_1_U3.dout_array[3] ;
reg [3:0] \ashr_4s_2ns_4_7_1_U3.dout_array[4] ;
reg [3:0] \ashr_4s_2ns_4_7_1_U3.dout_array[5] ;
reg [3:0] ashr_ln1297_reg_1109;
reg [31:0] conv_i389_reg_954;
reg icmp_ln1494_reg_1192;
reg icmp_ln768_reg_1002;
reg icmp_ln850_1_reg_1172;
reg icmp_ln850_reg_1325;
reg icmp_ln851_1_reg_1141;
reg icmp_ln851_2_reg_1297;
reg icmp_ln851_3_reg_1360;
reg icmp_ln851_reg_1129;
reg isNeg_reg_986;
reg [6:0] op_26_V_reg_1282;
reg [31:0] op_28_V_reg_1345;
reg [1:0] op_6_V_reg_1177;
reg [1:0] op_7_V_reg_1232;
reg [3:0] op_8_V_reg_1018;
reg overflow_reg_1007;
reg p_Result_7_reg_964;
reg p_Result_8_reg_997;
reg [1:0] p_Result_s_reg_975;
reg [3:0] p_Val2_2_reg_992;
reg [1:0] r_2_reg_980;
reg [3:0] r_V_1_reg_1146;
reg [26:0] r_V_reg_1094;
reg r_reg_1072;
reg [3:0] ret_V_18_reg_1047;
reg [8:0] ret_V_19_reg_1077;
reg [5:0] ret_V_20_reg_1182;
reg [3:0] ret_V_21_reg_1187;
reg [3:0] ret_V_22_reg_1314;
reg [6:0] ret_V_23_reg_1237;
reg [34:0] ret_V_24_reg_1302;
reg [31:0] ret_V_25_reg_1335;
reg [35:0] ret_V_26_reg_1365;
reg [31:0] ret_V_27_reg_1382;
reg [31:0] ret_V_28_reg_1392;
reg [31:0] ret_V_29_cast_reg_1307;
reg [31:0] ret_V_31_cast_reg_1370;
reg [5:0] ret_V_3_reg_1162;
reg [3:0] ret_V_5_reg_1167;
reg [5:0] ret_V_reg_1082;
reg [2:0] select_ln1347_reg_929;
reg select_ln13_reg_934;
reg [31:0] select_ln1497_reg_959;
reg [31:0] select_ln69_1_reg_1340;
reg [1:0] select_ln69_reg_1197;
reg [1:0] select_ln708_reg_1119;
reg [3:0] sext_ln850_reg_1134;
reg [1:0] \shl_4s_2ns_4_7_1_U4.din1_cast_array[0] ;
reg [1:0] \shl_4s_2ns_4_7_1_U4.din1_cast_array[1] ;
reg [1:0] \shl_4s_2ns_4_7_1_U4.din1_cast_array[2] ;
reg [1:0] \shl_4s_2ns_4_7_1_U4.din1_cast_array[3] ;
reg [1:0] \shl_4s_2ns_4_7_1_U4.din1_cast_array[4] ;
reg [1:0] \shl_4s_2ns_4_7_1_U4.din1_cast_array[5] ;
reg [3:0] \shl_4s_2ns_4_7_1_U4.dout_array[0] ;
reg [3:0] \shl_4s_2ns_4_7_1_U4.dout_array[1] ;
reg [3:0] \shl_4s_2ns_4_7_1_U4.dout_array[2] ;
reg [3:0] \shl_4s_2ns_4_7_1_U4.dout_array[3] ;
reg [3:0] \shl_4s_2ns_4_7_1_U4.dout_array[4] ;
reg [3:0] \shl_4s_2ns_4_7_1_U4.dout_array[5] ;
reg [3:0] shl_ln1358_reg_1114;
reg [13:0] \sub_27ns_27s_27_2_1_U5.top_sub_27ns_27s_27_2_1_Adder_2_U.ain_s1 ;
reg [13:0] \sub_27ns_27s_27_2_1_U5.top_sub_27ns_27s_27_2_1_Adder_2_U.bin_s1 ;
reg \sub_27ns_27s_27_2_1_U5.top_sub_27ns_27s_27_2_1_Adder_2_U.carry_s1 ;
reg [12:0] \sub_27ns_27s_27_2_1_U5.top_sub_27ns_27s_27_2_1_Adder_2_U.sum_s1 ;
reg \sub_2ns_2ns_2_2_1_U2.top_sub_2ns_2ns_2_2_1_Adder_1_U.ain_s1 ;
reg \sub_2ns_2ns_2_2_1_U2.top_sub_2ns_2ns_2_2_1_Adder_1_U.bin_s1 ;
reg \sub_2ns_2ns_2_2_1_U2.top_sub_2ns_2ns_2_2_1_Adder_1_U.carry_s1 ;
reg \sub_2ns_2ns_2_2_1_U2.top_sub_2ns_2ns_2_2_1_Adder_1_U.sum_s1 ;
reg \sub_2ns_2s_2_2_1_U10.top_sub_2ns_2s_2_2_1_Adder_7_U.ain_s1 ;
reg \sub_2ns_2s_2_2_1_U10.top_sub_2ns_2s_2_2_1_Adder_7_U.bin_s1 ;
reg \sub_2ns_2s_2_2_1_U10.top_sub_2ns_2s_2_2_1_Adder_7_U.carry_s1 ;
reg \sub_2ns_2s_2_2_1_U10.top_sub_2ns_2s_2_2_1_Adder_7_U.sum_s1 ;
reg [1:0] \sub_3ns_3s_3_2_1_U1.top_sub_3ns_3s_3_2_1_Adder_0_U.ain_s1 ;
reg [1:0] \sub_3ns_3s_3_2_1_U1.top_sub_3ns_3s_3_2_1_Adder_0_U.bin_s1 ;
reg \sub_3ns_3s_3_2_1_U1.top_sub_3ns_3s_3_2_1_Adder_0_U.carry_s1 ;
reg \sub_3ns_3s_3_2_1_U1.top_sub_3ns_3s_3_2_1_Adder_0_U.sum_s1 ;
reg [26:0] sub_ln1118_reg_1067;
reg [1:0] sub_ln1357_reg_1013;
reg [1:0] sub_ln69_reg_1202;
reg [2:0] tmp_2_reg_1099;
reg tmp_reg_1052;
reg [1:0] trunc_ln718_reg_1057;
reg trunc_ln728_reg_970;
reg [23:0] trunc_ln851_1_reg_1104;
reg [2:0] trunc_ln851_2_reg_1320;
reg [2:0] trunc_ln851_3_reg_1152;
reg [2:0] trunc_ln851_reg_1089;
reg [1:0] ush_reg_1026;
wire [31:0] _000_;
wire [31:0] _001_;
wire [6:0] _002_;
wire [1:0] _003_;
wire [2:0] _004_;
wire [5:0] _005_;
wire _006_;
wire [37:0] _007_;
wire [3:0] _008_;
wire [31:0] _009_;
wire _010_;
wire _011_;
wire _012_;
wire _013_;
wire _014_;
wire _015_;
wire _016_;
wire _017_;
wire _018_;
wire [6:0] _019_;
wire [31:0] _020_;
wire [1:0] _021_;
wire [1:0] _022_;
wire [3:0] _023_;
wire _024_;
wire _025_;
wire _026_;
wire [1:0] _027_;
wire _028_;
wire [1:0] _029_;
wire [3:0] _030_;
wire [26:0] _031_;
wire _032_;
wire [3:0] _033_;
wire [8:0] _034_;
wire [5:0] _035_;
wire [3:0] _036_;
wire [3:0] _037_;
wire [6:0] _038_;
wire [34:0] _039_;
wire [31:0] _040_;
wire [35:0] _041_;
wire [31:0] _042_;
wire [31:0] _043_;
wire [31:0] _044_;
wire [31:0] _045_;
wire [5:0] _046_;
wire [3:0] _047_;
wire [5:0] _048_;
wire [2:0] _049_;
wire _050_;
wire [31:0] _051_;
wire [31:0] _052_;
wire [1:0] _053_;
wire [1:0] _054_;
wire [3:0] _055_;
wire [3:0] _056_;
wire [26:0] _057_;
wire [1:0] _058_;
wire [1:0] _059_;
wire [2:0] _060_;
wire _061_;
wire [1:0] _062_;
wire _063_;
wire [23:0] _064_;
wire [2:0] _065_;
wire [2:0] _066_;
wire [2:0] _067_;
wire [1:0] _068_;
wire [1:0] _069_;
wire _070_;
wire _071_;
wire _072_;
wire _073_;
wire _074_;
wire _075_;
wire _076_;
wire _077_;
wire _078_;
wire _079_;
wire _080_;
wire _081_;
wire _082_;
wire _083_;
wire _084_;
wire _085_;
wire _086_;
wire [1:0] _087_;
wire [1:0] _088_;
wire _089_;
wire _090_;
wire _091_;
wire _092_;
wire [1:0] _093_;
wire [1:0] _094_;
wire [15:0] _095_;
wire [15:0] _096_;
wire _097_;
wire [15:0] _098_;
wire [16:0] _099_;
wire [16:0] _100_;
wire [15:0] _101_;
wire [15:0] _102_;
wire _103_;
wire [15:0] _104_;
wire [16:0] _105_;
wire [16:0] _106_;
wire [15:0] _107_;
wire [15:0] _108_;
wire _109_;
wire [15:0] _110_;
wire [16:0] _111_;
wire [16:0] _112_;
wire [15:0] _113_;
wire [15:0] _114_;
wire _115_;
wire [15:0] _116_;
wire [16:0] _117_;
wire [16:0] _118_;
wire [15:0] _119_;
wire [15:0] _120_;
wire _121_;
wire [15:0] _122_;
wire [16:0] _123_;
wire [16:0] _124_;
wire [17:0] _125_;
wire [17:0] _126_;
wire _127_;
wire [16:0] _128_;
wire [17:0] _129_;
wire [18:0] _130_;
wire [17:0] _131_;
wire [17:0] _132_;
wire _133_;
wire [17:0] _134_;
wire [18:0] _135_;
wire [18:0] _136_;
wire [1:0] _137_;
wire [1:0] _138_;
wire _139_;
wire _140_;
wire [1:0] _141_;
wire [2:0] _142_;
wire [1:0] _143_;
wire [1:0] _144_;
wire _145_;
wire [1:0] _146_;
wire [2:0] _147_;
wire [2:0] _148_;
wire [2:0] _149_;
wire [2:0] _150_;
wire _151_;
wire [2:0] _152_;
wire [3:0] _153_;
wire [3:0] _154_;
wire [2:0] _155_;
wire [2:0] _156_;
wire _157_;
wire [2:0] _158_;
wire [3:0] _159_;
wire [3:0] _160_;
wire [3:0] _161_;
wire [3:0] _162_;
wire _163_;
wire [2:0] _164_;
wire [3:0] _165_;
wire [4:0] _166_;
wire [3:0] _167_;
wire [3:0] _168_;
wire _169_;
wire [2:0] _170_;
wire [3:0] _171_;
wire [4:0] _172_;
wire [3:0] _173_;
wire [3:0] _174_;
wire _175_;
wire [2:0] _176_;
wire [3:0] _177_;
wire [4:0] _178_;
wire [4:0] _179_;
wire [4:0] _180_;
wire _181_;
wire [3:0] _182_;
wire [4:0] _183_;
wire [5:0] _184_;
wire [1:0] _185_;
wire [1:0] _186_;
wire [1:0] _187_;
wire [1:0] _188_;
wire [1:0] _189_;
wire [1:0] _190_;
wire [3:0] _191_;
wire [3:0] _192_;
wire [3:0] _193_;
wire [3:0] _194_;
wire [3:0] _195_;
wire [3:0] _196_;
wire [1:0] _197_;
wire [3:0] _198_;
wire [1:0] _199_;
wire [3:0] _200_;
wire [1:0] _201_;
wire [3:0] _202_;
wire [1:0] _203_;
wire [3:0] _204_;
wire [1:0] _205_;
wire [3:0] _206_;
wire [1:0] _207_;
wire [3:0] _208_;
wire [3:0] _209_;
wire [1:0] _210_;
wire [1:0] _211_;
wire [1:0] _212_;
wire [1:0] _213_;
wire [1:0] _214_;
wire [1:0] _215_;
wire [3:0] _216_;
wire [3:0] _217_;
wire [3:0] _218_;
wire [3:0] _219_;
wire [3:0] _220_;
wire [3:0] _221_;
wire [1:0] _222_;
wire [3:0] _223_;
wire [1:0] _224_;
wire [3:0] _225_;
wire [1:0] _226_;
wire [3:0] _227_;
wire [1:0] _228_;
wire [3:0] _229_;
wire [1:0] _230_;
wire [3:0] _231_;
wire [1:0] _232_;
wire [3:0] _233_;
wire [3:0] _234_;
wire [13:0] _235_;
wire [13:0] _236_;
wire _237_;
wire [12:0] _238_;
wire [13:0] _239_;
wire [14:0] _240_;
wire _241_;
wire _242_;
wire _243_;
wire _244_;
wire [1:0] _245_;
wire [1:0] _246_;
wire _247_;
wire _248_;
wire _249_;
wire _250_;
wire [1:0] _251_;
wire [1:0] _252_;
wire [1:0] _253_;
wire [1:0] _254_;
wire _255_;
wire _256_;
wire [1:0] _257_;
wire [2:0] _258_;
wire _259_;
wire _260_;
wire _261_;
wire _262_;
wire _263_;
wire _264_;
wire _265_;
wire _266_;
wire _267_;
wire _268_;
wire _269_;
wire _270_;
wire _271_;
wire _272_;
wire _273_;
wire _274_;
wire _275_;
wire _276_;
wire _277_;
wire _278_;
wire _279_;
wire _280_;
wire _281_;
wire _282_;
wire _283_;
wire _284_;
wire _285_;
wire _286_;
wire _287_;
wire _288_;
wire _289_;
wire _290_;
wire _291_;
wire _292_;
wire _293_;
wire _294_;
wire _295_;
wire _296_;
wire _297_;
wire _298_;
wire _299_;
wire _300_;
wire _301_;
wire _302_;
wire _303_;
wire \add_2ns_2ns_2_2_1_U13.ce ;
wire \add_2ns_2ns_2_2_1_U13.clk ;
wire [1:0] \add_2ns_2ns_2_2_1_U13.din0 ;
wire [1:0] \add_2ns_2ns_2_2_1_U13.din1 ;
wire [1:0] \add_2ns_2ns_2_2_1_U13.dout ;
wire \add_2ns_2ns_2_2_1_U13.reset ;
wire [1:0] \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_6_U.a ;
wire [1:0] \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_6_U.ain_s0 ;
wire [1:0] \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_6_U.b ;
wire [1:0] \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_6_U.bin_s0 ;
wire \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_6_U.ce ;
wire \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_6_U.clk ;
wire \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_6_U.facout_s1 ;
wire \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_6_U.facout_s2 ;
wire \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_6_U.fas_s1 ;
wire \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_6_U.fas_s2 ;
wire \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_6_U.reset ;
wire [1:0] \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_6_U.s ;
wire \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_6_U.u1.a ;
wire \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_6_U.u1.b ;
wire \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_6_U.u1.cin ;
wire \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_6_U.u1.cout ;
wire \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_6_U.u1.s ;
wire \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_6_U.u2.a ;
wire \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_6_U.u2.b ;
wire \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_6_U.u2.cin ;
wire \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_6_U.u2.cout ;
wire \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_6_U.u2.s ;
wire \add_2ns_2ns_2_2_1_U9.ce ;
wire \add_2ns_2ns_2_2_1_U9.clk ;
wire [1:0] \add_2ns_2ns_2_2_1_U9.din0 ;
wire [1:0] \add_2ns_2ns_2_2_1_U9.din1 ;
wire [1:0] \add_2ns_2ns_2_2_1_U9.dout ;
wire \add_2ns_2ns_2_2_1_U9.reset ;
wire [1:0] \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.a ;
wire [1:0] \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.ain_s0 ;
wire [1:0] \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.b ;
wire [1:0] \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.bin_s0 ;
wire \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.ce ;
wire \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.clk ;
wire \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.facout_s1 ;
wire \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.facout_s2 ;
wire \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.fas_s1 ;
wire \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.fas_s2 ;
wire \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.reset ;
wire [1:0] \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.s ;
wire \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.u1.a ;
wire \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.u1.b ;
wire \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.u1.cin ;
wire \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.u1.cout ;
wire \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.u1.s ;
wire \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.u2.a ;
wire \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.u2.b ;
wire \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.u2.cin ;
wire \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.u2.cout ;
wire \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.u2.s ;
wire \add_32ns_32ns_32_2_1_U18.ce ;
wire \add_32ns_32ns_32_2_1_U18.clk ;
wire [31:0] \add_32ns_32ns_32_2_1_U18.din0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U18.din1 ;
wire [31:0] \add_32ns_32ns_32_2_1_U18.dout ;
wire \add_32ns_32ns_32_2_1_U18.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_13_U.a ;
wire [31:0] \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_13_U.ain_s0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_13_U.b ;
wire [31:0] \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_13_U.bin_s0 ;
wire \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_13_U.ce ;
wire \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_13_U.clk ;
wire \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_13_U.facout_s1 ;
wire \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_13_U.facout_s2 ;
wire [15:0] \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_13_U.fas_s1 ;
wire [15:0] \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_13_U.fas_s2 ;
wire \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_13_U.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_13_U.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_13_U.u1.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_13_U.u1.b ;
wire \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_13_U.u1.cin ;
wire \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_13_U.u1.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_13_U.u1.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_13_U.u2.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_13_U.u2.b ;
wire \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_13_U.u2.cin ;
wire \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_13_U.u2.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_13_U.u2.s ;
wire \add_32ns_32ns_32_2_1_U19.ce ;
wire \add_32ns_32ns_32_2_1_U19.clk ;
wire [31:0] \add_32ns_32ns_32_2_1_U19.din0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U19.din1 ;
wire [31:0] \add_32ns_32ns_32_2_1_U19.dout ;
wire \add_32ns_32ns_32_2_1_U19.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_13_U.a ;
wire [31:0] \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_13_U.ain_s0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_13_U.b ;
wire [31:0] \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_13_U.bin_s0 ;
wire \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_13_U.ce ;
wire \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_13_U.clk ;
wire \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_13_U.facout_s1 ;
wire \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_13_U.facout_s2 ;
wire [15:0] \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_13_U.fas_s1 ;
wire [15:0] \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_13_U.fas_s2 ;
wire \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_13_U.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_13_U.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_13_U.u1.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_13_U.u1.b ;
wire \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_13_U.u1.cin ;
wire \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_13_U.u1.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_13_U.u1.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_13_U.u2.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_13_U.u2.b ;
wire \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_13_U.u2.cin ;
wire \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_13_U.u2.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_13_U.u2.s ;
wire \add_32ns_32ns_32_2_1_U21.ce ;
wire \add_32ns_32ns_32_2_1_U21.clk ;
wire [31:0] \add_32ns_32ns_32_2_1_U21.din0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U21.din1 ;
wire [31:0] \add_32ns_32ns_32_2_1_U21.dout ;
wire \add_32ns_32ns_32_2_1_U21.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_13_U.a ;
wire [31:0] \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_13_U.ain_s0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_13_U.b ;
wire [31:0] \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_13_U.bin_s0 ;
wire \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_13_U.ce ;
wire \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_13_U.clk ;
wire \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_13_U.facout_s1 ;
wire \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_13_U.facout_s2 ;
wire [15:0] \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_13_U.fas_s1 ;
wire [15:0] \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_13_U.fas_s2 ;
wire \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_13_U.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_13_U.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_13_U.u1.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_13_U.u1.b ;
wire \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_13_U.u1.cin ;
wire \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_13_U.u1.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_13_U.u1.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_13_U.u2.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_13_U.u2.b ;
wire \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_13_U.u2.cin ;
wire \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_13_U.u2.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_13_U.u2.s ;
wire \add_32ns_32s_32_2_1_U22.ce ;
wire \add_32ns_32s_32_2_1_U22.clk ;
wire [31:0] \add_32ns_32s_32_2_1_U22.din0 ;
wire [31:0] \add_32ns_32s_32_2_1_U22.din1 ;
wire [31:0] \add_32ns_32s_32_2_1_U22.dout ;
wire \add_32ns_32s_32_2_1_U22.reset ;
wire [31:0] \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_15_U.a ;
wire [31:0] \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_15_U.ain_s0 ;
wire [31:0] \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_15_U.b ;
wire [31:0] \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_15_U.bin_s0 ;
wire \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_15_U.ce ;
wire \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_15_U.clk ;
wire \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_15_U.facout_s1 ;
wire \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_15_U.facout_s2 ;
wire [15:0] \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_15_U.fas_s1 ;
wire [15:0] \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_15_U.fas_s2 ;
wire \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_15_U.reset ;
wire [31:0] \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_15_U.s ;
wire [15:0] \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_15_U.u1.a ;
wire [15:0] \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_15_U.u1.b ;
wire \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_15_U.u1.cin ;
wire \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_15_U.u1.cout ;
wire [15:0] \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_15_U.u1.s ;
wire [15:0] \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_15_U.u2.a ;
wire [15:0] \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_15_U.u2.b ;
wire \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_15_U.u2.cin ;
wire \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_15_U.u2.cout ;
wire [15:0] \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_15_U.u2.s ;
wire \add_32ns_32s_32_2_1_U23.ce ;
wire \add_32ns_32s_32_2_1_U23.clk ;
wire [31:0] \add_32ns_32s_32_2_1_U23.din0 ;
wire [31:0] \add_32ns_32s_32_2_1_U23.din1 ;
wire [31:0] \add_32ns_32s_32_2_1_U23.dout ;
wire \add_32ns_32s_32_2_1_U23.reset ;
wire [31:0] \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_15_U.a ;
wire [31:0] \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_15_U.ain_s0 ;
wire [31:0] \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_15_U.b ;
wire [31:0] \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_15_U.bin_s0 ;
wire \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_15_U.ce ;
wire \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_15_U.clk ;
wire \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_15_U.facout_s1 ;
wire \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_15_U.facout_s2 ;
wire [15:0] \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_15_U.fas_s1 ;
wire [15:0] \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_15_U.fas_s2 ;
wire \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_15_U.reset ;
wire [31:0] \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_15_U.s ;
wire [15:0] \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_15_U.u1.a ;
wire [15:0] \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_15_U.u1.b ;
wire \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_15_U.u1.cin ;
wire \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_15_U.u1.cout ;
wire [15:0] \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_15_U.u1.s ;
wire [15:0] \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_15_U.u2.a ;
wire [15:0] \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_15_U.u2.b ;
wire \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_15_U.u2.cin ;
wire \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_15_U.u2.cout ;
wire [15:0] \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_15_U.u2.s ;
wire \add_35s_35s_35_2_1_U17.ce ;
wire \add_35s_35s_35_2_1_U17.clk ;
wire [34:0] \add_35s_35s_35_2_1_U17.din0 ;
wire [34:0] \add_35s_35s_35_2_1_U17.din1 ;
wire [34:0] \add_35s_35s_35_2_1_U17.dout ;
wire \add_35s_35s_35_2_1_U17.reset ;
wire [34:0] \add_35s_35s_35_2_1_U17.top_add_35s_35s_35_2_1_Adder_12_U.a ;
wire [34:0] \add_35s_35s_35_2_1_U17.top_add_35s_35s_35_2_1_Adder_12_U.ain_s0 ;
wire [34:0] \add_35s_35s_35_2_1_U17.top_add_35s_35s_35_2_1_Adder_12_U.b ;
wire [34:0] \add_35s_35s_35_2_1_U17.top_add_35s_35s_35_2_1_Adder_12_U.bin_s0 ;
wire \add_35s_35s_35_2_1_U17.top_add_35s_35s_35_2_1_Adder_12_U.ce ;
wire \add_35s_35s_35_2_1_U17.top_add_35s_35s_35_2_1_Adder_12_U.clk ;
wire \add_35s_35s_35_2_1_U17.top_add_35s_35s_35_2_1_Adder_12_U.facout_s1 ;
wire \add_35s_35s_35_2_1_U17.top_add_35s_35s_35_2_1_Adder_12_U.facout_s2 ;
wire [16:0] \add_35s_35s_35_2_1_U17.top_add_35s_35s_35_2_1_Adder_12_U.fas_s1 ;
wire [17:0] \add_35s_35s_35_2_1_U17.top_add_35s_35s_35_2_1_Adder_12_U.fas_s2 ;
wire \add_35s_35s_35_2_1_U17.top_add_35s_35s_35_2_1_Adder_12_U.reset ;
wire [34:0] \add_35s_35s_35_2_1_U17.top_add_35s_35s_35_2_1_Adder_12_U.s ;
wire [16:0] \add_35s_35s_35_2_1_U17.top_add_35s_35s_35_2_1_Adder_12_U.u1.a ;
wire [16:0] \add_35s_35s_35_2_1_U17.top_add_35s_35s_35_2_1_Adder_12_U.u1.b ;
wire \add_35s_35s_35_2_1_U17.top_add_35s_35s_35_2_1_Adder_12_U.u1.cin ;
wire \add_35s_35s_35_2_1_U17.top_add_35s_35s_35_2_1_Adder_12_U.u1.cout ;
wire [16:0] \add_35s_35s_35_2_1_U17.top_add_35s_35s_35_2_1_Adder_12_U.u1.s ;
wire [17:0] \add_35s_35s_35_2_1_U17.top_add_35s_35s_35_2_1_Adder_12_U.u2.a ;
wire [17:0] \add_35s_35s_35_2_1_U17.top_add_35s_35s_35_2_1_Adder_12_U.u2.b ;
wire \add_35s_35s_35_2_1_U17.top_add_35s_35s_35_2_1_Adder_12_U.u2.cin ;
wire \add_35s_35s_35_2_1_U17.top_add_35s_35s_35_2_1_Adder_12_U.u2.cout ;
wire [17:0] \add_35s_35s_35_2_1_U17.top_add_35s_35s_35_2_1_Adder_12_U.u2.s ;
wire \add_36s_36s_36_2_1_U20.ce ;
wire \add_36s_36s_36_2_1_U20.clk ;
wire [35:0] \add_36s_36s_36_2_1_U20.din0 ;
wire [35:0] \add_36s_36s_36_2_1_U20.din1 ;
wire [35:0] \add_36s_36s_36_2_1_U20.dout ;
wire \add_36s_36s_36_2_1_U20.reset ;
wire [35:0] \add_36s_36s_36_2_1_U20.top_add_36s_36s_36_2_1_Adder_14_U.a ;
wire [35:0] \add_36s_36s_36_2_1_U20.top_add_36s_36s_36_2_1_Adder_14_U.ain_s0 ;
wire [35:0] \add_36s_36s_36_2_1_U20.top_add_36s_36s_36_2_1_Adder_14_U.b ;
wire [35:0] \add_36s_36s_36_2_1_U20.top_add_36s_36s_36_2_1_Adder_14_U.bin_s0 ;
wire \add_36s_36s_36_2_1_U20.top_add_36s_36s_36_2_1_Adder_14_U.ce ;
wire \add_36s_36s_36_2_1_U20.top_add_36s_36s_36_2_1_Adder_14_U.clk ;
wire \add_36s_36s_36_2_1_U20.top_add_36s_36s_36_2_1_Adder_14_U.facout_s1 ;
wire \add_36s_36s_36_2_1_U20.top_add_36s_36s_36_2_1_Adder_14_U.facout_s2 ;
wire [17:0] \add_36s_36s_36_2_1_U20.top_add_36s_36s_36_2_1_Adder_14_U.fas_s1 ;
wire [17:0] \add_36s_36s_36_2_1_U20.top_add_36s_36s_36_2_1_Adder_14_U.fas_s2 ;
wire \add_36s_36s_36_2_1_U20.top_add_36s_36s_36_2_1_Adder_14_U.reset ;
wire [35:0] \add_36s_36s_36_2_1_U20.top_add_36s_36s_36_2_1_Adder_14_U.s ;
wire [17:0] \add_36s_36s_36_2_1_U20.top_add_36s_36s_36_2_1_Adder_14_U.u1.a ;
wire [17:0] \add_36s_36s_36_2_1_U20.top_add_36s_36s_36_2_1_Adder_14_U.u1.b ;
wire \add_36s_36s_36_2_1_U20.top_add_36s_36s_36_2_1_Adder_14_U.u1.cin ;
wire \add_36s_36s_36_2_1_U20.top_add_36s_36s_36_2_1_Adder_14_U.u1.cout ;
wire [17:0] \add_36s_36s_36_2_1_U20.top_add_36s_36s_36_2_1_Adder_14_U.u1.s ;
wire [17:0] \add_36s_36s_36_2_1_U20.top_add_36s_36s_36_2_1_Adder_14_U.u2.a ;
wire [17:0] \add_36s_36s_36_2_1_U20.top_add_36s_36s_36_2_1_Adder_14_U.u2.b ;
wire \add_36s_36s_36_2_1_U20.top_add_36s_36s_36_2_1_Adder_14_U.u2.cin ;
wire \add_36s_36s_36_2_1_U20.top_add_36s_36s_36_2_1_Adder_14_U.u2.cout ;
wire [17:0] \add_36s_36s_36_2_1_U20.top_add_36s_36s_36_2_1_Adder_14_U.u2.s ;
wire \add_3s_3s_3_2_1_U15.ce ;
wire \add_3s_3s_3_2_1_U15.clk ;
wire [2:0] \add_3s_3s_3_2_1_U15.din0 ;
wire [2:0] \add_3s_3s_3_2_1_U15.din1 ;
wire [2:0] \add_3s_3s_3_2_1_U15.dout ;
wire \add_3s_3s_3_2_1_U15.reset ;
wire [2:0] \add_3s_3s_3_2_1_U15.top_add_3s_3s_3_2_1_Adder_11_U.a ;
wire [2:0] \add_3s_3s_3_2_1_U15.top_add_3s_3s_3_2_1_Adder_11_U.ain_s0 ;
wire [2:0] \add_3s_3s_3_2_1_U15.top_add_3s_3s_3_2_1_Adder_11_U.b ;
wire [2:0] \add_3s_3s_3_2_1_U15.top_add_3s_3s_3_2_1_Adder_11_U.bin_s0 ;
wire \add_3s_3s_3_2_1_U15.top_add_3s_3s_3_2_1_Adder_11_U.ce ;
wire \add_3s_3s_3_2_1_U15.top_add_3s_3s_3_2_1_Adder_11_U.clk ;
wire \add_3s_3s_3_2_1_U15.top_add_3s_3s_3_2_1_Adder_11_U.facout_s1 ;
wire \add_3s_3s_3_2_1_U15.top_add_3s_3s_3_2_1_Adder_11_U.facout_s2 ;
wire \add_3s_3s_3_2_1_U15.top_add_3s_3s_3_2_1_Adder_11_U.fas_s1 ;
wire [1:0] \add_3s_3s_3_2_1_U15.top_add_3s_3s_3_2_1_Adder_11_U.fas_s2 ;
wire \add_3s_3s_3_2_1_U15.top_add_3s_3s_3_2_1_Adder_11_U.reset ;
wire [2:0] \add_3s_3s_3_2_1_U15.top_add_3s_3s_3_2_1_Adder_11_U.s ;
wire \add_3s_3s_3_2_1_U15.top_add_3s_3s_3_2_1_Adder_11_U.u1.a ;
wire \add_3s_3s_3_2_1_U15.top_add_3s_3s_3_2_1_Adder_11_U.u1.b ;
wire \add_3s_3s_3_2_1_U15.top_add_3s_3s_3_2_1_Adder_11_U.u1.cin ;
wire \add_3s_3s_3_2_1_U15.top_add_3s_3s_3_2_1_Adder_11_U.u1.cout ;
wire \add_3s_3s_3_2_1_U15.top_add_3s_3s_3_2_1_Adder_11_U.u1.s ;
wire [1:0] \add_3s_3s_3_2_1_U15.top_add_3s_3s_3_2_1_Adder_11_U.u2.a ;
wire [1:0] \add_3s_3s_3_2_1_U15.top_add_3s_3s_3_2_1_Adder_11_U.u2.b ;
wire \add_3s_3s_3_2_1_U15.top_add_3s_3s_3_2_1_Adder_11_U.u2.cin ;
wire \add_3s_3s_3_2_1_U15.top_add_3s_3s_3_2_1_Adder_11_U.u2.cout ;
wire [1:0] \add_3s_3s_3_2_1_U15.top_add_3s_3s_3_2_1_Adder_11_U.u2.s ;
wire \add_4s_4ns_4_2_1_U8.ce ;
wire \add_4s_4ns_4_2_1_U8.clk ;
wire [3:0] \add_4s_4ns_4_2_1_U8.din0 ;
wire [3:0] \add_4s_4ns_4_2_1_U8.din1 ;
wire [3:0] \add_4s_4ns_4_2_1_U8.dout ;
wire \add_4s_4ns_4_2_1_U8.reset ;
wire [3:0] \add_4s_4ns_4_2_1_U8.top_add_4s_4ns_4_2_1_Adder_5_U.a ;
wire [3:0] \add_4s_4ns_4_2_1_U8.top_add_4s_4ns_4_2_1_Adder_5_U.ain_s0 ;
wire [3:0] \add_4s_4ns_4_2_1_U8.top_add_4s_4ns_4_2_1_Adder_5_U.b ;
wire [3:0] \add_4s_4ns_4_2_1_U8.top_add_4s_4ns_4_2_1_Adder_5_U.bin_s0 ;
wire \add_4s_4ns_4_2_1_U8.top_add_4s_4ns_4_2_1_Adder_5_U.ce ;
wire \add_4s_4ns_4_2_1_U8.top_add_4s_4ns_4_2_1_Adder_5_U.clk ;
wire \add_4s_4ns_4_2_1_U8.top_add_4s_4ns_4_2_1_Adder_5_U.facout_s1 ;
wire \add_4s_4ns_4_2_1_U8.top_add_4s_4ns_4_2_1_Adder_5_U.facout_s2 ;
wire [1:0] \add_4s_4ns_4_2_1_U8.top_add_4s_4ns_4_2_1_Adder_5_U.fas_s1 ;
wire [1:0] \add_4s_4ns_4_2_1_U8.top_add_4s_4ns_4_2_1_Adder_5_U.fas_s2 ;
wire \add_4s_4ns_4_2_1_U8.top_add_4s_4ns_4_2_1_Adder_5_U.reset ;
wire [3:0] \add_4s_4ns_4_2_1_U8.top_add_4s_4ns_4_2_1_Adder_5_U.s ;
wire [1:0] \add_4s_4ns_4_2_1_U8.top_add_4s_4ns_4_2_1_Adder_5_U.u1.a ;
wire [1:0] \add_4s_4ns_4_2_1_U8.top_add_4s_4ns_4_2_1_Adder_5_U.u1.b ;
wire \add_4s_4ns_4_2_1_U8.top_add_4s_4ns_4_2_1_Adder_5_U.u1.cin ;
wire \add_4s_4ns_4_2_1_U8.top_add_4s_4ns_4_2_1_Adder_5_U.u1.cout ;
wire [1:0] \add_4s_4ns_4_2_1_U8.top_add_4s_4ns_4_2_1_Adder_5_U.u1.s ;
wire [1:0] \add_4s_4ns_4_2_1_U8.top_add_4s_4ns_4_2_1_Adder_5_U.u2.a ;
wire [1:0] \add_4s_4ns_4_2_1_U8.top_add_4s_4ns_4_2_1_Adder_5_U.u2.b ;
wire \add_4s_4ns_4_2_1_U8.top_add_4s_4ns_4_2_1_Adder_5_U.u2.cin ;
wire \add_4s_4ns_4_2_1_U8.top_add_4s_4ns_4_2_1_Adder_5_U.u2.cout ;
wire [1:0] \add_4s_4ns_4_2_1_U8.top_add_4s_4ns_4_2_1_Adder_5_U.u2.s ;
wire \add_6ns_6ns_6_2_1_U7.ce ;
wire \add_6ns_6ns_6_2_1_U7.clk ;
wire [5:0] \add_6ns_6ns_6_2_1_U7.din0 ;
wire [5:0] \add_6ns_6ns_6_2_1_U7.din1 ;
wire [5:0] \add_6ns_6ns_6_2_1_U7.dout ;
wire \add_6ns_6ns_6_2_1_U7.reset ;
wire [5:0] \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_4_U.a ;
wire [5:0] \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_4_U.ain_s0 ;
wire [5:0] \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_4_U.b ;
wire [5:0] \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_4_U.bin_s0 ;
wire \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_4_U.ce ;
wire \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_4_U.clk ;
wire \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_4_U.facout_s1 ;
wire \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_4_U.facout_s2 ;
wire [2:0] \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_4_U.fas_s1 ;
wire [2:0] \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_4_U.fas_s2 ;
wire \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_4_U.reset ;
wire [5:0] \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_4_U.s ;
wire [2:0] \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_4_U.u1.a ;
wire [2:0] \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_4_U.u1.b ;
wire \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_4_U.u1.cin ;
wire \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_4_U.u1.cout ;
wire [2:0] \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_4_U.u1.s ;
wire [2:0] \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_4_U.u2.a ;
wire [2:0] \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_4_U.u2.b ;
wire \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_4_U.u2.cin ;
wire \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_4_U.u2.cout ;
wire [2:0] \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_4_U.u2.s ;
wire \add_6s_6ns_6_2_1_U12.ce ;
wire \add_6s_6ns_6_2_1_U12.clk ;
wire [5:0] \add_6s_6ns_6_2_1_U12.din0 ;
wire [5:0] \add_6s_6ns_6_2_1_U12.din1 ;
wire [5:0] \add_6s_6ns_6_2_1_U12.dout ;
wire \add_6s_6ns_6_2_1_U12.reset ;
wire [5:0] \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.a ;
wire [5:0] \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.ain_s0 ;
wire [5:0] \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.b ;
wire [5:0] \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.bin_s0 ;
wire \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.ce ;
wire \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.clk ;
wire \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.facout_s1 ;
wire \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.facout_s2 ;
wire [2:0] \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.fas_s1 ;
wire [2:0] \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.fas_s2 ;
wire \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.reset ;
wire [5:0] \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.s ;
wire [2:0] \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.u1.a ;
wire [2:0] \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.u1.b ;
wire \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.u1.cin ;
wire \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.u1.cout ;
wire [2:0] \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.u1.s ;
wire [2:0] \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.u2.a ;
wire [2:0] \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.u2.b ;
wire \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.u2.cin ;
wire \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.u2.cout ;
wire [2:0] \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.u2.s ;
wire \add_7s_7ns_7_2_1_U14.ce ;
wire \add_7s_7ns_7_2_1_U14.clk ;
wire [6:0] \add_7s_7ns_7_2_1_U14.din0 ;
wire [6:0] \add_7s_7ns_7_2_1_U14.din1 ;
wire [6:0] \add_7s_7ns_7_2_1_U14.dout ;
wire \add_7s_7ns_7_2_1_U14.reset ;
wire [6:0] \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_10_U.a ;
wire [6:0] \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_10_U.ain_s0 ;
wire [6:0] \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_10_U.b ;
wire [6:0] \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_10_U.bin_s0 ;
wire \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_10_U.ce ;
wire \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_10_U.clk ;
wire \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_10_U.facout_s1 ;
wire \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_10_U.facout_s2 ;
wire [2:0] \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_10_U.fas_s1 ;
wire [3:0] \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_10_U.fas_s2 ;
wire \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_10_U.reset ;
wire [6:0] \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_10_U.s ;
wire [2:0] \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_10_U.u1.a ;
wire [2:0] \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_10_U.u1.b ;
wire \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_10_U.u1.cin ;
wire \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_10_U.u1.cout ;
wire [2:0] \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_10_U.u1.s ;
wire [3:0] \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_10_U.u2.a ;
wire [3:0] \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_10_U.u2.b ;
wire \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_10_U.u2.cin ;
wire \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_10_U.u2.cout ;
wire [3:0] \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_10_U.u2.s ;
wire \add_7s_7ns_7_2_1_U16.ce ;
wire \add_7s_7ns_7_2_1_U16.clk ;
wire [6:0] \add_7s_7ns_7_2_1_U16.din0 ;
wire [6:0] \add_7s_7ns_7_2_1_U16.din1 ;
wire [6:0] \add_7s_7ns_7_2_1_U16.dout ;
wire \add_7s_7ns_7_2_1_U16.reset ;
wire [6:0] \add_7s_7ns_7_2_1_U16.top_add_7s_7ns_7_2_1_Adder_10_U.a ;
wire [6:0] \add_7s_7ns_7_2_1_U16.top_add_7s_7ns_7_2_1_Adder_10_U.ain_s0 ;
wire [6:0] \add_7s_7ns_7_2_1_U16.top_add_7s_7ns_7_2_1_Adder_10_U.b ;
wire [6:0] \add_7s_7ns_7_2_1_U16.top_add_7s_7ns_7_2_1_Adder_10_U.bin_s0 ;
wire \add_7s_7ns_7_2_1_U16.top_add_7s_7ns_7_2_1_Adder_10_U.ce ;
wire \add_7s_7ns_7_2_1_U16.top_add_7s_7ns_7_2_1_Adder_10_U.clk ;
wire \add_7s_7ns_7_2_1_U16.top_add_7s_7ns_7_2_1_Adder_10_U.facout_s1 ;
wire \add_7s_7ns_7_2_1_U16.top_add_7s_7ns_7_2_1_Adder_10_U.facout_s2 ;
wire [2:0] \add_7s_7ns_7_2_1_U16.top_add_7s_7ns_7_2_1_Adder_10_U.fas_s1 ;
wire [3:0] \add_7s_7ns_7_2_1_U16.top_add_7s_7ns_7_2_1_Adder_10_U.fas_s2 ;
wire \add_7s_7ns_7_2_1_U16.top_add_7s_7ns_7_2_1_Adder_10_U.reset ;
wire [6:0] \add_7s_7ns_7_2_1_U16.top_add_7s_7ns_7_2_1_Adder_10_U.s ;
wire [2:0] \add_7s_7ns_7_2_1_U16.top_add_7s_7ns_7_2_1_Adder_10_U.u1.a ;
wire [2:0] \add_7s_7ns_7_2_1_U16.top_add_7s_7ns_7_2_1_Adder_10_U.u1.b ;
wire \add_7s_7ns_7_2_1_U16.top_add_7s_7ns_7_2_1_Adder_10_U.u1.cin ;
wire \add_7s_7ns_7_2_1_U16.top_add_7s_7ns_7_2_1_Adder_10_U.u1.cout ;
wire [2:0] \add_7s_7ns_7_2_1_U16.top_add_7s_7ns_7_2_1_Adder_10_U.u1.s ;
wire [3:0] \add_7s_7ns_7_2_1_U16.top_add_7s_7ns_7_2_1_Adder_10_U.u2.a ;
wire [3:0] \add_7s_7ns_7_2_1_U16.top_add_7s_7ns_7_2_1_Adder_10_U.u2.b ;
wire \add_7s_7ns_7_2_1_U16.top_add_7s_7ns_7_2_1_Adder_10_U.u2.cin ;
wire \add_7s_7ns_7_2_1_U16.top_add_7s_7ns_7_2_1_Adder_10_U.u2.cout ;
wire [3:0] \add_7s_7ns_7_2_1_U16.top_add_7s_7ns_7_2_1_Adder_10_U.u2.s ;
wire \add_7s_7s_7_2_1_U11.ce ;
wire \add_7s_7s_7_2_1_U11.clk ;
wire [6:0] \add_7s_7s_7_2_1_U11.din0 ;
wire [6:0] \add_7s_7s_7_2_1_U11.din1 ;
wire [6:0] \add_7s_7s_7_2_1_U11.dout ;
wire \add_7s_7s_7_2_1_U11.reset ;
wire [6:0] \add_7s_7s_7_2_1_U11.top_add_7s_7s_7_2_1_Adder_8_U.a ;
wire [6:0] \add_7s_7s_7_2_1_U11.top_add_7s_7s_7_2_1_Adder_8_U.ain_s0 ;
wire [6:0] \add_7s_7s_7_2_1_U11.top_add_7s_7s_7_2_1_Adder_8_U.b ;
wire [6:0] \add_7s_7s_7_2_1_U11.top_add_7s_7s_7_2_1_Adder_8_U.bin_s0 ;
wire \add_7s_7s_7_2_1_U11.top_add_7s_7s_7_2_1_Adder_8_U.ce ;
wire \add_7s_7s_7_2_1_U11.top_add_7s_7s_7_2_1_Adder_8_U.clk ;
wire \add_7s_7s_7_2_1_U11.top_add_7s_7s_7_2_1_Adder_8_U.facout_s1 ;
wire \add_7s_7s_7_2_1_U11.top_add_7s_7s_7_2_1_Adder_8_U.facout_s2 ;
wire [2:0] \add_7s_7s_7_2_1_U11.top_add_7s_7s_7_2_1_Adder_8_U.fas_s1 ;
wire [3:0] \add_7s_7s_7_2_1_U11.top_add_7s_7s_7_2_1_Adder_8_U.fas_s2 ;
wire \add_7s_7s_7_2_1_U11.top_add_7s_7s_7_2_1_Adder_8_U.reset ;
wire [6:0] \add_7s_7s_7_2_1_U11.top_add_7s_7s_7_2_1_Adder_8_U.s ;
wire [2:0] \add_7s_7s_7_2_1_U11.top_add_7s_7s_7_2_1_Adder_8_U.u1.a ;
wire [2:0] \add_7s_7s_7_2_1_U11.top_add_7s_7s_7_2_1_Adder_8_U.u1.b ;
wire \add_7s_7s_7_2_1_U11.top_add_7s_7s_7_2_1_Adder_8_U.u1.cin ;
wire \add_7s_7s_7_2_1_U11.top_add_7s_7s_7_2_1_Adder_8_U.u1.cout ;
wire [2:0] \add_7s_7s_7_2_1_U11.top_add_7s_7s_7_2_1_Adder_8_U.u1.s ;
wire [3:0] \add_7s_7s_7_2_1_U11.top_add_7s_7s_7_2_1_Adder_8_U.u2.a ;
wire [3:0] \add_7s_7s_7_2_1_U11.top_add_7s_7s_7_2_1_Adder_8_U.u2.b ;
wire \add_7s_7s_7_2_1_U11.top_add_7s_7s_7_2_1_Adder_8_U.u2.cin ;
wire \add_7s_7s_7_2_1_U11.top_add_7s_7s_7_2_1_Adder_8_U.u2.cout ;
wire [3:0] \add_7s_7s_7_2_1_U11.top_add_7s_7s_7_2_1_Adder_8_U.u2.s ;
wire \add_9s_9ns_9_2_1_U6.ce ;
wire \add_9s_9ns_9_2_1_U6.clk ;
wire [8:0] \add_9s_9ns_9_2_1_U6.din0 ;
wire [8:0] \add_9s_9ns_9_2_1_U6.din1 ;
wire [8:0] \add_9s_9ns_9_2_1_U6.dout ;
wire \add_9s_9ns_9_2_1_U6.reset ;
wire [8:0] \add_9s_9ns_9_2_1_U6.top_add_9s_9ns_9_2_1_Adder_3_U.a ;
wire [8:0] \add_9s_9ns_9_2_1_U6.top_add_9s_9ns_9_2_1_Adder_3_U.ain_s0 ;
wire [8:0] \add_9s_9ns_9_2_1_U6.top_add_9s_9ns_9_2_1_Adder_3_U.b ;
wire [8:0] \add_9s_9ns_9_2_1_U6.top_add_9s_9ns_9_2_1_Adder_3_U.bin_s0 ;
wire \add_9s_9ns_9_2_1_U6.top_add_9s_9ns_9_2_1_Adder_3_U.ce ;
wire \add_9s_9ns_9_2_1_U6.top_add_9s_9ns_9_2_1_Adder_3_U.clk ;
wire \add_9s_9ns_9_2_1_U6.top_add_9s_9ns_9_2_1_Adder_3_U.facout_s1 ;
wire \add_9s_9ns_9_2_1_U6.top_add_9s_9ns_9_2_1_Adder_3_U.facout_s2 ;
wire [3:0] \add_9s_9ns_9_2_1_U6.top_add_9s_9ns_9_2_1_Adder_3_U.fas_s1 ;
wire [4:0] \add_9s_9ns_9_2_1_U6.top_add_9s_9ns_9_2_1_Adder_3_U.fas_s2 ;
wire \add_9s_9ns_9_2_1_U6.top_add_9s_9ns_9_2_1_Adder_3_U.reset ;
wire [8:0] \add_9s_9ns_9_2_1_U6.top_add_9s_9ns_9_2_1_Adder_3_U.s ;
wire [3:0] \add_9s_9ns_9_2_1_U6.top_add_9s_9ns_9_2_1_Adder_3_U.u1.a ;
wire [3:0] \add_9s_9ns_9_2_1_U6.top_add_9s_9ns_9_2_1_Adder_3_U.u1.b ;
wire \add_9s_9ns_9_2_1_U6.top_add_9s_9ns_9_2_1_Adder_3_U.u1.cin ;
wire \add_9s_9ns_9_2_1_U6.top_add_9s_9ns_9_2_1_Adder_3_U.u1.cout ;
wire [3:0] \add_9s_9ns_9_2_1_U6.top_add_9s_9ns_9_2_1_Adder_3_U.u1.s ;
wire [4:0] \add_9s_9ns_9_2_1_U6.top_add_9s_9ns_9_2_1_Adder_3_U.u2.a ;
wire [4:0] \add_9s_9ns_9_2_1_U6.top_add_9s_9ns_9_2_1_Adder_3_U.u2.b ;
wire \add_9s_9ns_9_2_1_U6.top_add_9s_9ns_9_2_1_Adder_3_U.u2.cin ;
wire \add_9s_9ns_9_2_1_U6.top_add_9s_9ns_9_2_1_Adder_3_U.u2.cout ;
wire [4:0] \add_9s_9ns_9_2_1_U6.top_add_9s_9ns_9_2_1_Adder_3_U.u2.s ;
wire and_ln410_fu_511_p2;
wire and_ln850_1_fu_636_p2;
wire and_ln850_fu_796_p2;
wire ap_CS_fsm_state1;
wire ap_CS_fsm_state11;
wire ap_CS_fsm_state12;
wire ap_CS_fsm_state13;
wire ap_CS_fsm_state14;
wire ap_CS_fsm_state15;
wire ap_CS_fsm_state16;
wire ap_CS_fsm_state17;
wire ap_CS_fsm_state18;
wire ap_CS_fsm_state19;
wire ap_CS_fsm_state2;
wire ap_CS_fsm_state20;
wire ap_CS_fsm_state21;
wire ap_CS_fsm_state22;
wire ap_CS_fsm_state23;
wire ap_CS_fsm_state24;
wire ap_CS_fsm_state25;
wire ap_CS_fsm_state26;
wire ap_CS_fsm_state27;
wire ap_CS_fsm_state28;
wire ap_CS_fsm_state29;
wire ap_CS_fsm_state3;
wire ap_CS_fsm_state30;
wire ap_CS_fsm_state31;
wire ap_CS_fsm_state32;
wire ap_CS_fsm_state33;
wire ap_CS_fsm_state34;
wire ap_CS_fsm_state35;
wire ap_CS_fsm_state36;
wire ap_CS_fsm_state37;
wire ap_CS_fsm_state38;
wire ap_CS_fsm_state4;
wire ap_CS_fsm_state5;
wire ap_CS_fsm_state6;
wire ap_CS_fsm_state7;
wire [37:0] ap_NS_fsm;
wire ap_clk;
wire ap_done;
wire ap_idle;
wire ap_ready;
wire ap_rst;
wire ap_start;
wire \ashr_4s_2ns_4_7_1_U3.ce ;
wire \ashr_4s_2ns_4_7_1_U3.clk ;
wire [3:0] \ashr_4s_2ns_4_7_1_U3.din0 ;
wire [3:0] \ashr_4s_2ns_4_7_1_U3.din1 ;
wire [1:0] \ashr_4s_2ns_4_7_1_U3.din1_cast ;
wire [1:0] \ashr_4s_2ns_4_7_1_U3.din1_mask ;
wire [3:0] \ashr_4s_2ns_4_7_1_U3.dout ;
wire \ashr_4s_2ns_4_7_1_U3.reset ;
wire [31:0] ashr_ln1497_1_fu_283_p2;
wire [1:0] conv_i389_fu_222_p0;
wire [31:0] conv_i389_fu_222_p1;
wire [2:0] grp_fu_217_p1;
wire [2:0] grp_fu_217_p2;
wire [1:0] grp_fu_332_p2;
wire [3:0] grp_fu_378_p2;
wire [3:0] grp_fu_383_p2;
wire [26:0] grp_fu_399_p1;
wire [26:0] grp_fu_399_p2;
wire [8:0] grp_fu_434_p0;
wire [8:0] grp_fu_434_p2;
wire [5:0] grp_fu_522_p2;
wire [3:0] grp_fu_535_p0;
wire [3:0] grp_fu_535_p2;
wire [1:0] grp_fu_553_p0;
wire [1:0] grp_fu_553_p2;
wire [1:0] grp_fu_563_p2;
wire [6:0] grp_fu_661_p0;
wire [6:0] grp_fu_661_p1;
wire [6:0] grp_fu_661_p2;
wire [5:0] grp_fu_677_p0;
wire [5:0] grp_fu_677_p1;
wire [5:0] grp_fu_677_p2;
wire [1:0] grp_fu_683_p1;
wire [1:0] grp_fu_683_p2;
wire [6:0] grp_fu_700_p0;
wire [6:0] grp_fu_700_p2;
wire [2:0] grp_fu_708_p0;
wire [2:0] grp_fu_708_p1;
wire [2:0] grp_fu_708_p2;
wire [6:0] grp_fu_717_p0;
wire [6:0] grp_fu_717_p2;
wire [34:0] grp_fu_737_p0;
wire [34:0] grp_fu_737_p1;
wire [34:0] grp_fu_737_p2;
wire [31:0] grp_fu_772_p2;
wire [31:0] grp_fu_834_p2;
wire [35:0] grp_fu_853_p0;
wire [35:0] grp_fu_853_p1;
wire [35:0] grp_fu_853_p2;
wire [31:0] grp_fu_879_p2;
wire [31:0] grp_fu_907_p1;
wire [31:0] grp_fu_907_p2;
wire [31:0] grp_fu_916_p1;
wire [31:0] grp_fu_916_p2;
wire icmp_ln1494_fu_616_p2;
wire icmp_ln768_fu_327_p2;
wire icmp_ln850_1_fu_558_p2;
wire icmp_ln850_fu_777_p2;
wire icmp_ln851_1_fu_530_p2;
wire icmp_ln851_2_fu_747_p2;
wire icmp_ln851_3_fu_863_p2;
wire icmp_ln851_fu_517_p2;
wire [7:0] op_0;
wire [3:0] op_1;
wire [3:0] op_11;
wire [3:0] op_12;
wire [3:0] op_15;
wire [3:0] op_17;
wire [1:0] op_18;
wire [3:0] op_19;
wire op_3;
wire [31:0] op_31;
wire op_31_ap_vld;
wire op_3_read_read_fu_130_p2;
wire [1:0] op_4;
wire op_7_V_fu_688_p0;
wire [1:0] op_7_V_fu_688_p3;
wire [3:0] op_8_V_fu_363_p3;
wire or_ln384_fu_359_p2;
wire or_ln410_fu_506_p2;
wire or_ln785_fu_337_p2;
wire overflow_fu_346_p2;
wire p_Result_1_fu_587_p3;
wire p_Result_2_fu_789_p3;
wire p_Result_3_fu_629_p3;
wire p_Result_4_fu_807_p3;
wire p_Result_5_fu_884_p3;
wire p_Result_6_fu_486_p3;
wire p_Result_8_fu_321_p2;
wire p_Result_s_14_fu_568_p3;
wire [3:0] p_Val2_2_fu_314_p3;
wire [1:0] r_2_fu_302_p1;
wire [3:0] r_V_1_fu_541_p3;
wire r_V_fu_459_p0;
wire [26:0] r_V_fu_459_p3;
wire r_fu_440_p2;
wire ret_V_11_fu_622_p3;
wire ret_V_12_fu_641_p2;
wire [3:0] ret_V_18_fu_412_p2;
wire [5:0] ret_V_20_fu_580_p3;
wire [3:0] ret_V_21_fu_599_p3;
wire [3:0] ret_V_22_fu_763_p2;
wire [31:0] ret_V_25_fu_819_p3;
wire [31:0] ret_V_27_fu_896_p3;
wire ret_V_8_fu_782_p3;
wire ret_V_9_fu_801_p2;
wire [34:0] rhs_4_fu_842_p3;
wire rhs_fu_405_p1;
wire [3:0] rhs_fu_405_p3;
wire select_ln1347_fu_197_p0;
wire [2:0] select_ln1347_fu_197_p3;
wire select_ln13_fu_205_p0;
wire select_ln13_fu_205_p3;
wire [1:0] select_ln1497_1_fu_275_p3;
wire [1:0] select_ln1497_2_fu_288_p3;
wire [31:0] select_ln1497_3_fu_295_p3;
wire [31:0] select_ln1497_fu_232_p3;
wire [3:0] select_ln384_fu_352_p3;
wire [31:0] select_ln69_1_fu_826_p3;
wire [1:0] select_ln69_fu_647_p3;
wire [1:0] select_ln708_fu_479_p3;
wire select_ln835_fu_261_p3;
wire [3:0] select_ln850_2_fu_594_p3;
wire [31:0] select_ln850_3_fu_814_p3;
wire [31:0] select_ln850_4_fu_891_p3;
wire [5:0] select_ln850_fu_575_p3;
wire [1:0] sext_ln1347_fu_213_p0;
wire [4:0] sext_ln1494_fu_613_p1;
wire [3:0] sext_ln703_1_fu_722_p0;
wire [3:0] sext_ln703_2_fu_838_p0;
wire [3:0] sext_ln850_fu_527_p1;
wire \shl_4s_2ns_4_7_1_U4.ce ;
wire \shl_4s_2ns_4_7_1_U4.clk ;
wire [3:0] \shl_4s_2ns_4_7_1_U4.din0 ;
wire [3:0] \shl_4s_2ns_4_7_1_U4.din1 ;
wire [1:0] \shl_4s_2ns_4_7_1_U4.din1_cast ;
wire [1:0] \shl_4s_2ns_4_7_1_U4.din1_mask ;
wire [3:0] \shl_4s_2ns_4_7_1_U4.dout ;
wire \shl_4s_2ns_4_7_1_U4.reset ;
wire [30:0] shl_ln1497_1_fu_226_p2;
wire [1:0] shl_ln1_fu_606_p1;
wire [4:0] shl_ln1_fu_606_p3;
wire [1:0] shl_ln_fu_388_p1;
wire [25:0] shl_ln_fu_388_p3;
wire \sub_27ns_27s_27_2_1_U5.ce ;
wire \sub_27ns_27s_27_2_1_U5.clk ;
wire [26:0] \sub_27ns_27s_27_2_1_U5.din0 ;
wire [26:0] \sub_27ns_27s_27_2_1_U5.din1 ;
wire [26:0] \sub_27ns_27s_27_2_1_U5.dout ;
wire \sub_27ns_27s_27_2_1_U5.reset ;
wire [26:0] \sub_27ns_27s_27_2_1_U5.top_sub_27ns_27s_27_2_1_Adder_2_U.a ;
wire [26:0] \sub_27ns_27s_27_2_1_U5.top_sub_27ns_27s_27_2_1_Adder_2_U.ain_s0 ;
wire [26:0] \sub_27ns_27s_27_2_1_U5.top_sub_27ns_27s_27_2_1_Adder_2_U.b ;
wire [26:0] \sub_27ns_27s_27_2_1_U5.top_sub_27ns_27s_27_2_1_Adder_2_U.bin_s0 ;
wire \sub_27ns_27s_27_2_1_U5.top_sub_27ns_27s_27_2_1_Adder_2_U.ce ;
wire \sub_27ns_27s_27_2_1_U5.top_sub_27ns_27s_27_2_1_Adder_2_U.clk ;
wire \sub_27ns_27s_27_2_1_U5.top_sub_27ns_27s_27_2_1_Adder_2_U.facout_s1 ;
wire \sub_27ns_27s_27_2_1_U5.top_sub_27ns_27s_27_2_1_Adder_2_U.facout_s2 ;
wire [12:0] \sub_27ns_27s_27_2_1_U5.top_sub_27ns_27s_27_2_1_Adder_2_U.fas_s1 ;
wire [13:0] \sub_27ns_27s_27_2_1_U5.top_sub_27ns_27s_27_2_1_Adder_2_U.fas_s2 ;
wire \sub_27ns_27s_27_2_1_U5.top_sub_27ns_27s_27_2_1_Adder_2_U.reset ;
wire [26:0] \sub_27ns_27s_27_2_1_U5.top_sub_27ns_27s_27_2_1_Adder_2_U.s ;
wire [12:0] \sub_27ns_27s_27_2_1_U5.top_sub_27ns_27s_27_2_1_Adder_2_U.u1.a ;
wire [12:0] \sub_27ns_27s_27_2_1_U5.top_sub_27ns_27s_27_2_1_Adder_2_U.u1.b ;
wire \sub_27ns_27s_27_2_1_U5.top_sub_27ns_27s_27_2_1_Adder_2_U.u1.cin ;
wire \sub_27ns_27s_27_2_1_U5.top_sub_27ns_27s_27_2_1_Adder_2_U.u1.cout ;
wire [12:0] \sub_27ns_27s_27_2_1_U5.top_sub_27ns_27s_27_2_1_Adder_2_U.u1.s ;
wire [13:0] \sub_27ns_27s_27_2_1_U5.top_sub_27ns_27s_27_2_1_Adder_2_U.u2.a ;
wire [13:0] \sub_27ns_27s_27_2_1_U5.top_sub_27ns_27s_27_2_1_Adder_2_U.u2.b ;
wire \sub_27ns_27s_27_2_1_U5.top_sub_27ns_27s_27_2_1_Adder_2_U.u2.cin ;
wire \sub_27ns_27s_27_2_1_U5.top_sub_27ns_27s_27_2_1_Adder_2_U.u2.cout ;
wire [13:0] \sub_27ns_27s_27_2_1_U5.top_sub_27ns_27s_27_2_1_Adder_2_U.u2.s ;
wire \sub_2ns_2ns_2_2_1_U2.ce ;
wire \sub_2ns_2ns_2_2_1_U2.clk ;
wire [1:0] \sub_2ns_2ns_2_2_1_U2.din0 ;
wire [1:0] \sub_2ns_2ns_2_2_1_U2.din1 ;
wire [1:0] \sub_2ns_2ns_2_2_1_U2.dout ;
wire \sub_2ns_2ns_2_2_1_U2.reset ;
wire [1:0] \sub_2ns_2ns_2_2_1_U2.top_sub_2ns_2ns_2_2_1_Adder_1_U.a ;
wire [1:0] \sub_2ns_2ns_2_2_1_U2.top_sub_2ns_2ns_2_2_1_Adder_1_U.ain_s0 ;
wire [1:0] \sub_2ns_2ns_2_2_1_U2.top_sub_2ns_2ns_2_2_1_Adder_1_U.b ;
wire [1:0] \sub_2ns_2ns_2_2_1_U2.top_sub_2ns_2ns_2_2_1_Adder_1_U.bin_s0 ;
wire \sub_2ns_2ns_2_2_1_U2.top_sub_2ns_2ns_2_2_1_Adder_1_U.ce ;
wire \sub_2ns_2ns_2_2_1_U2.top_sub_2ns_2ns_2_2_1_Adder_1_U.clk ;
wire \sub_2ns_2ns_2_2_1_U2.top_sub_2ns_2ns_2_2_1_Adder_1_U.facout_s1 ;
wire \sub_2ns_2ns_2_2_1_U2.top_sub_2ns_2ns_2_2_1_Adder_1_U.facout_s2 ;
wire \sub_2ns_2ns_2_2_1_U2.top_sub_2ns_2ns_2_2_1_Adder_1_U.fas_s1 ;
wire \sub_2ns_2ns_2_2_1_U2.top_sub_2ns_2ns_2_2_1_Adder_1_U.fas_s2 ;
wire \sub_2ns_2ns_2_2_1_U2.top_sub_2ns_2ns_2_2_1_Adder_1_U.reset ;
wire [1:0] \sub_2ns_2ns_2_2_1_U2.top_sub_2ns_2ns_2_2_1_Adder_1_U.s ;
wire \sub_2ns_2ns_2_2_1_U2.top_sub_2ns_2ns_2_2_1_Adder_1_U.u1.a ;
wire \sub_2ns_2ns_2_2_1_U2.top_sub_2ns_2ns_2_2_1_Adder_1_U.u1.b ;
wire \sub_2ns_2ns_2_2_1_U2.top_sub_2ns_2ns_2_2_1_Adder_1_U.u1.cin ;
wire \sub_2ns_2ns_2_2_1_U2.top_sub_2ns_2ns_2_2_1_Adder_1_U.u1.cout ;
wire \sub_2ns_2ns_2_2_1_U2.top_sub_2ns_2ns_2_2_1_Adder_1_U.u1.s ;
wire \sub_2ns_2ns_2_2_1_U2.top_sub_2ns_2ns_2_2_1_Adder_1_U.u2.a ;
wire \sub_2ns_2ns_2_2_1_U2.top_sub_2ns_2ns_2_2_1_Adder_1_U.u2.b ;
wire \sub_2ns_2ns_2_2_1_U2.top_sub_2ns_2ns_2_2_1_Adder_1_U.u2.cin ;
wire \sub_2ns_2ns_2_2_1_U2.top_sub_2ns_2ns_2_2_1_Adder_1_U.u2.cout ;
wire \sub_2ns_2ns_2_2_1_U2.top_sub_2ns_2ns_2_2_1_Adder_1_U.u2.s ;
wire \sub_2ns_2s_2_2_1_U10.ce ;
wire \sub_2ns_2s_2_2_1_U10.clk ;
wire [1:0] \sub_2ns_2s_2_2_1_U10.din0 ;
wire [1:0] \sub_2ns_2s_2_2_1_U10.din1 ;
wire [1:0] \sub_2ns_2s_2_2_1_U10.dout ;
wire \sub_2ns_2s_2_2_1_U10.reset ;
wire [1:0] \sub_2ns_2s_2_2_1_U10.top_sub_2ns_2s_2_2_1_Adder_7_U.a ;
wire [1:0] \sub_2ns_2s_2_2_1_U10.top_sub_2ns_2s_2_2_1_Adder_7_U.ain_s0 ;
wire [1:0] \sub_2ns_2s_2_2_1_U10.top_sub_2ns_2s_2_2_1_Adder_7_U.b ;
wire [1:0] \sub_2ns_2s_2_2_1_U10.top_sub_2ns_2s_2_2_1_Adder_7_U.bin_s0 ;
wire \sub_2ns_2s_2_2_1_U10.top_sub_2ns_2s_2_2_1_Adder_7_U.ce ;
wire \sub_2ns_2s_2_2_1_U10.top_sub_2ns_2s_2_2_1_Adder_7_U.clk ;
wire \sub_2ns_2s_2_2_1_U10.top_sub_2ns_2s_2_2_1_Adder_7_U.facout_s1 ;
wire \sub_2ns_2s_2_2_1_U10.top_sub_2ns_2s_2_2_1_Adder_7_U.facout_s2 ;
wire \sub_2ns_2s_2_2_1_U10.top_sub_2ns_2s_2_2_1_Adder_7_U.fas_s1 ;
wire \sub_2ns_2s_2_2_1_U10.top_sub_2ns_2s_2_2_1_Adder_7_U.fas_s2 ;
wire \sub_2ns_2s_2_2_1_U10.top_sub_2ns_2s_2_2_1_Adder_7_U.reset ;
wire [1:0] \sub_2ns_2s_2_2_1_U10.top_sub_2ns_2s_2_2_1_Adder_7_U.s ;
wire \sub_2ns_2s_2_2_1_U10.top_sub_2ns_2s_2_2_1_Adder_7_U.u1.a ;
wire \sub_2ns_2s_2_2_1_U10.top_sub_2ns_2s_2_2_1_Adder_7_U.u1.b ;
wire \sub_2ns_2s_2_2_1_U10.top_sub_2ns_2s_2_2_1_Adder_7_U.u1.cin ;
wire \sub_2ns_2s_2_2_1_U10.top_sub_2ns_2s_2_2_1_Adder_7_U.u1.cout ;
wire \sub_2ns_2s_2_2_1_U10.top_sub_2ns_2s_2_2_1_Adder_7_U.u1.s ;
wire \sub_2ns_2s_2_2_1_U10.top_sub_2ns_2s_2_2_1_Adder_7_U.u2.a ;
wire \sub_2ns_2s_2_2_1_U10.top_sub_2ns_2s_2_2_1_Adder_7_U.u2.b ;
wire \sub_2ns_2s_2_2_1_U10.top_sub_2ns_2s_2_2_1_Adder_7_U.u2.cin ;
wire \sub_2ns_2s_2_2_1_U10.top_sub_2ns_2s_2_2_1_Adder_7_U.u2.cout ;
wire \sub_2ns_2s_2_2_1_U10.top_sub_2ns_2s_2_2_1_Adder_7_U.u2.s ;
wire \sub_3ns_3s_3_2_1_U1.ce ;
wire \sub_3ns_3s_3_2_1_U1.clk ;
wire [2:0] \sub_3ns_3s_3_2_1_U1.din0 ;
wire [2:0] \sub_3ns_3s_3_2_1_U1.din1 ;
wire [2:0] \sub_3ns_3s_3_2_1_U1.dout ;
wire \sub_3ns_3s_3_2_1_U1.reset ;
wire [2:0] \sub_3ns_3s_3_2_1_U1.top_sub_3ns_3s_3_2_1_Adder_0_U.a ;
wire [2:0] \sub_3ns_3s_3_2_1_U1.top_sub_3ns_3s_3_2_1_Adder_0_U.ain_s0 ;
wire [2:0] \sub_3ns_3s_3_2_1_U1.top_sub_3ns_3s_3_2_1_Adder_0_U.b ;
wire [2:0] \sub_3ns_3s_3_2_1_U1.top_sub_3ns_3s_3_2_1_Adder_0_U.bin_s0 ;
wire \sub_3ns_3s_3_2_1_U1.top_sub_3ns_3s_3_2_1_Adder_0_U.ce ;
wire \sub_3ns_3s_3_2_1_U1.top_sub_3ns_3s_3_2_1_Adder_0_U.clk ;
wire \sub_3ns_3s_3_2_1_U1.top_sub_3ns_3s_3_2_1_Adder_0_U.facout_s1 ;
wire \sub_3ns_3s_3_2_1_U1.top_sub_3ns_3s_3_2_1_Adder_0_U.facout_s2 ;
wire \sub_3ns_3s_3_2_1_U1.top_sub_3ns_3s_3_2_1_Adder_0_U.fas_s1 ;
wire [1:0] \sub_3ns_3s_3_2_1_U1.top_sub_3ns_3s_3_2_1_Adder_0_U.fas_s2 ;
wire \sub_3ns_3s_3_2_1_U1.top_sub_3ns_3s_3_2_1_Adder_0_U.reset ;
wire [2:0] \sub_3ns_3s_3_2_1_U1.top_sub_3ns_3s_3_2_1_Adder_0_U.s ;
wire \sub_3ns_3s_3_2_1_U1.top_sub_3ns_3s_3_2_1_Adder_0_U.u1.a ;
wire \sub_3ns_3s_3_2_1_U1.top_sub_3ns_3s_3_2_1_Adder_0_U.u1.b ;
wire \sub_3ns_3s_3_2_1_U1.top_sub_3ns_3s_3_2_1_Adder_0_U.u1.cin ;
wire \sub_3ns_3s_3_2_1_U1.top_sub_3ns_3s_3_2_1_Adder_0_U.u1.cout ;
wire \sub_3ns_3s_3_2_1_U1.top_sub_3ns_3s_3_2_1_Adder_0_U.u1.s ;
wire [1:0] \sub_3ns_3s_3_2_1_U1.top_sub_3ns_3s_3_2_1_Adder_0_U.u2.a ;
wire [1:0] \sub_3ns_3s_3_2_1_U1.top_sub_3ns_3s_3_2_1_Adder_0_U.u2.b ;
wire \sub_3ns_3s_3_2_1_U1.top_sub_3ns_3s_3_2_1_Adder_0_U.u2.cin ;
wire \sub_3ns_3s_3_2_1_U1.top_sub_3ns_3s_3_2_1_Adder_0_U.u2.cout ;
wire [1:0] \sub_3ns_3s_3_2_1_U1.top_sub_3ns_3s_3_2_1_Adder_0_U.u2.s ;
wire [8:0] tmp_14_fu_726_p3;
wire tmp_3_fu_493_p3;
wire [1:0] tmp_7_fu_268_p1;
wire tmp_7_fu_268_p3;
wire [1:0] trunc_ln718_fu_426_p1;
wire trunc_ln728_fu_247_p1;
wire [23:0] trunc_ln851_1_fu_475_p1;
wire [2:0] trunc_ln851_2_fu_768_p1;
wire [2:0] trunc_ln851_3_fu_546_p1;
wire [3:0] trunc_ln851_4_fu_743_p0;
wire [1:0] trunc_ln851_4_fu_743_p1;
wire [3:0] trunc_ln851_5_fu_859_p0;
wire [2:0] trunc_ln851_5_fu_859_p1;
wire [2:0] trunc_ln851_fu_455_p1;
wire [1:0] ush_fu_370_p3;
wire xor_ln410_fu_500_p2;
wire xor_ln785_fu_341_p2;
wire [3:0] zext_ln1357_fu_375_p1;


assign _070_ = icmp_ln851_3_reg_1360 & ap_CS_fsm[32];
assign _071_ = icmp_ln851_2_reg_1297 & ap_CS_fsm[25];
assign _072_ = ap_CS_fsm[12] & isNeg_reg_986;
assign _073_ = ap_CS_fsm[12] & _079_;
assign _074_ = op_3 & ap_CS_fsm[11];
assign _075_ = ap_CS_fsm[4] & isNeg_reg_986;
assign _076_ = op_3 & ap_CS_fsm[16];
assign _077_ = _080_ & ap_CS_fsm[0];
assign _078_ = ap_start & ap_CS_fsm[0];
assign and_ln410_fu_511_p2 = op_1[2] & or_ln410_fu_506_p2;
assign and_ln850_1_fu_636_p2 = r_V_1_reg_1146[3] & icmp_ln850_1_reg_1172;
assign and_ln850_fu_796_p2 = ret_V_22_reg_1314[3] & icmp_ln850_reg_1325;
assign overflow_fu_346_p2 = xor_ln785_fu_341_p2 & or_ln785_fu_337_p2;
assign xor_ln410_fu_500_p2 = ~ ret_V_18_reg_1047[3];
assign xor_ln785_fu_341_p2 = ~ p_Result_7_reg_964;
assign _079_ = ~ isNeg_reg_986;
assign _080_ = ~ ap_start;
assign _081_ = ! trunc_ln851_1_reg_1104;
assign _082_ = ! trunc_ln851_reg_1089;
always @(posedge \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_6_U.clk )
\add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_6_U.bin_s1  <= _084_;
always @(posedge \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_6_U.clk )
\add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_6_U.ain_s1  <= _083_;
always @(posedge \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_6_U.clk )
\add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_6_U.sum_s1  <= _086_;
always @(posedge \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_6_U.clk )
\add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_6_U.carry_s1  <= _085_;
assign _084_ = \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_6_U.ce  ? \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_6_U.b [1] : \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_6_U.bin_s1 ;
assign _083_ = \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_6_U.ce  ? \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_6_U.a [1] : \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_6_U.ain_s1 ;
assign _085_ = \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_6_U.ce  ? \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_6_U.facout_s1  : \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_6_U.carry_s1 ;
assign _086_ = \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_6_U.ce  ? \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_6_U.fas_s1  : \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_6_U.sum_s1 ;
assign _087_ = \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_6_U.u1.a  + \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_6_U.u1.b ;
assign { \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_6_U.u1.cout , \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_6_U.u1.s  } = _087_ + \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_6_U.u1.cin ;
assign _088_ = \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_6_U.u2.a  + \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_6_U.u2.b ;
assign { \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_6_U.u2.cout , \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_6_U.u2.s  } = _088_ + \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_6_U.u2.cin ;
always @(posedge \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.clk )
\add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.bin_s1  <= _090_;
always @(posedge \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.clk )
\add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.ain_s1  <= _089_;
always @(posedge \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.clk )
\add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.sum_s1  <= _092_;
always @(posedge \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.clk )
\add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.carry_s1  <= _091_;
assign _090_ = \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.ce  ? \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.b [1] : \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.bin_s1 ;
assign _089_ = \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.ce  ? \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.a [1] : \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.ain_s1 ;
assign _091_ = \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.ce  ? \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.facout_s1  : \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.carry_s1 ;
assign _092_ = \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.ce  ? \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.fas_s1  : \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.sum_s1 ;
assign _093_ = \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.u1.a  + \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.u1.b ;
assign { \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.u1.cout , \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.u1.s  } = _093_ + \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.u1.cin ;
assign _094_ = \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.u2.a  + \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.u2.b ;
assign { \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.u2.cout , \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.u2.s  } = _094_ + \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.u2.cin ;
always @(posedge \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_13_U.clk )
\add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_13_U.bin_s1  <= _096_;
always @(posedge \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_13_U.clk )
\add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_13_U.ain_s1  <= _095_;
always @(posedge \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_13_U.clk )
\add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_13_U.sum_s1  <= _098_;
always @(posedge \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_13_U.clk )
\add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_13_U.carry_s1  <= _097_;
assign _096_ = \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_13_U.ce  ? \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_13_U.b [31:16] : \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_13_U.bin_s1 ;
assign _095_ = \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_13_U.ce  ? \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_13_U.a [31:16] : \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_13_U.ain_s1 ;
assign _097_ = \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_13_U.ce  ? \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_13_U.facout_s1  : \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_13_U.carry_s1 ;
assign _098_ = \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_13_U.ce  ? \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_13_U.fas_s1  : \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_13_U.sum_s1 ;
assign _099_ = \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_13_U.u1.a  + \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_13_U.u1.b ;
assign { \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_13_U.u1.cout , \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_13_U.u1.s  } = _099_ + \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_13_U.u1.cin ;
assign _100_ = \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_13_U.u2.a  + \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_13_U.u2.b ;
assign { \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_13_U.u2.cout , \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_13_U.u2.s  } = _100_ + \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_13_U.u2.cin ;
always @(posedge \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_13_U.clk )
\add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_13_U.bin_s1  <= _102_;
always @(posedge \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_13_U.clk )
\add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_13_U.ain_s1  <= _101_;
always @(posedge \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_13_U.clk )
\add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_13_U.sum_s1  <= _104_;
always @(posedge \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_13_U.clk )
\add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_13_U.carry_s1  <= _103_;
assign _102_ = \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_13_U.ce  ? \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_13_U.b [31:16] : \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_13_U.bin_s1 ;
assign _101_ = \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_13_U.ce  ? \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_13_U.a [31:16] : \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_13_U.ain_s1 ;
assign _103_ = \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_13_U.ce  ? \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_13_U.facout_s1  : \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_13_U.carry_s1 ;
assign _104_ = \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_13_U.ce  ? \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_13_U.fas_s1  : \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_13_U.sum_s1 ;
assign _105_ = \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_13_U.u1.a  + \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_13_U.u1.b ;
assign { \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_13_U.u1.cout , \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_13_U.u1.s  } = _105_ + \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_13_U.u1.cin ;
assign _106_ = \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_13_U.u2.a  + \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_13_U.u2.b ;
assign { \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_13_U.u2.cout , \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_13_U.u2.s  } = _106_ + \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_13_U.u2.cin ;
always @(posedge \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_13_U.clk )
\add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_13_U.bin_s1  <= _108_;
always @(posedge \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_13_U.clk )
\add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_13_U.ain_s1  <= _107_;
always @(posedge \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_13_U.clk )
\add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_13_U.sum_s1  <= _110_;
always @(posedge \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_13_U.clk )
\add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_13_U.carry_s1  <= _109_;
assign _108_ = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_13_U.ce  ? \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_13_U.b [31:16] : \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_13_U.bin_s1 ;
assign _107_ = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_13_U.ce  ? \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_13_U.a [31:16] : \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_13_U.ain_s1 ;
assign _109_ = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_13_U.ce  ? \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_13_U.facout_s1  : \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_13_U.carry_s1 ;
assign _110_ = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_13_U.ce  ? \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_13_U.fas_s1  : \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_13_U.sum_s1 ;
assign _111_ = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_13_U.u1.a  + \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_13_U.u1.b ;
assign { \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_13_U.u1.cout , \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_13_U.u1.s  } = _111_ + \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_13_U.u1.cin ;
assign _112_ = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_13_U.u2.a  + \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_13_U.u2.b ;
assign { \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_13_U.u2.cout , \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_13_U.u2.s  } = _112_ + \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_13_U.u2.cin ;
always @(posedge \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_15_U.clk )
\add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_15_U.bin_s1  <= _114_;
always @(posedge \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_15_U.clk )
\add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_15_U.ain_s1  <= _113_;
always @(posedge \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_15_U.clk )
\add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_15_U.sum_s1  <= _116_;
always @(posedge \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_15_U.clk )
\add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_15_U.carry_s1  <= _115_;
assign _114_ = \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_15_U.ce  ? \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_15_U.b [31:16] : \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_15_U.bin_s1 ;
assign _113_ = \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_15_U.ce  ? \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_15_U.a [31:16] : \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_15_U.ain_s1 ;
assign _115_ = \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_15_U.ce  ? \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_15_U.facout_s1  : \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_15_U.carry_s1 ;
assign _116_ = \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_15_U.ce  ? \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_15_U.fas_s1  : \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_15_U.sum_s1 ;
assign _117_ = \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_15_U.u1.a  + \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_15_U.u1.b ;
assign { \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_15_U.u1.cout , \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_15_U.u1.s  } = _117_ + \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_15_U.u1.cin ;
assign _118_ = \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_15_U.u2.a  + \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_15_U.u2.b ;
assign { \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_15_U.u2.cout , \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_15_U.u2.s  } = _118_ + \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_15_U.u2.cin ;
always @(posedge \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_15_U.clk )
\add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_15_U.bin_s1  <= _120_;
always @(posedge \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_15_U.clk )
\add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_15_U.ain_s1  <= _119_;
always @(posedge \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_15_U.clk )
\add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_15_U.sum_s1  <= _122_;
always @(posedge \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_15_U.clk )
\add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_15_U.carry_s1  <= _121_;
assign _120_ = \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_15_U.ce  ? \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_15_U.b [31:16] : \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_15_U.bin_s1 ;
assign _119_ = \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_15_U.ce  ? \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_15_U.a [31:16] : \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_15_U.ain_s1 ;
assign _121_ = \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_15_U.ce  ? \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_15_U.facout_s1  : \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_15_U.carry_s1 ;
assign _122_ = \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_15_U.ce  ? \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_15_U.fas_s1  : \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_15_U.sum_s1 ;
assign _123_ = \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_15_U.u1.a  + \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_15_U.u1.b ;
assign { \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_15_U.u1.cout , \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_15_U.u1.s  } = _123_ + \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_15_U.u1.cin ;
assign _124_ = \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_15_U.u2.a  + \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_15_U.u2.b ;
assign { \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_15_U.u2.cout , \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_15_U.u2.s  } = _124_ + \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_15_U.u2.cin ;
always @(posedge \add_35s_35s_35_2_1_U17.top_add_35s_35s_35_2_1_Adder_12_U.clk )
\add_35s_35s_35_2_1_U17.top_add_35s_35s_35_2_1_Adder_12_U.bin_s1  <= _126_;
always @(posedge \add_35s_35s_35_2_1_U17.top_add_35s_35s_35_2_1_Adder_12_U.clk )
\add_35s_35s_35_2_1_U17.top_add_35s_35s_35_2_1_Adder_12_U.ain_s1  <= _125_;
always @(posedge \add_35s_35s_35_2_1_U17.top_add_35s_35s_35_2_1_Adder_12_U.clk )
\add_35s_35s_35_2_1_U17.top_add_35s_35s_35_2_1_Adder_12_U.sum_s1  <= _128_;
always @(posedge \add_35s_35s_35_2_1_U17.top_add_35s_35s_35_2_1_Adder_12_U.clk )
\add_35s_35s_35_2_1_U17.top_add_35s_35s_35_2_1_Adder_12_U.carry_s1  <= _127_;
assign _126_ = \add_35s_35s_35_2_1_U17.top_add_35s_35s_35_2_1_Adder_12_U.ce  ? \add_35s_35s_35_2_1_U17.top_add_35s_35s_35_2_1_Adder_12_U.b [34:17] : \add_35s_35s_35_2_1_U17.top_add_35s_35s_35_2_1_Adder_12_U.bin_s1 ;
assign _125_ = \add_35s_35s_35_2_1_U17.top_add_35s_35s_35_2_1_Adder_12_U.ce  ? \add_35s_35s_35_2_1_U17.top_add_35s_35s_35_2_1_Adder_12_U.a [34:17] : \add_35s_35s_35_2_1_U17.top_add_35s_35s_35_2_1_Adder_12_U.ain_s1 ;
assign _127_ = \add_35s_35s_35_2_1_U17.top_add_35s_35s_35_2_1_Adder_12_U.ce  ? \add_35s_35s_35_2_1_U17.top_add_35s_35s_35_2_1_Adder_12_U.facout_s1  : \add_35s_35s_35_2_1_U17.top_add_35s_35s_35_2_1_Adder_12_U.carry_s1 ;
assign _128_ = \add_35s_35s_35_2_1_U17.top_add_35s_35s_35_2_1_Adder_12_U.ce  ? \add_35s_35s_35_2_1_U17.top_add_35s_35s_35_2_1_Adder_12_U.fas_s1  : \add_35s_35s_35_2_1_U17.top_add_35s_35s_35_2_1_Adder_12_U.sum_s1 ;
assign _129_ = \add_35s_35s_35_2_1_U17.top_add_35s_35s_35_2_1_Adder_12_U.u1.a  + \add_35s_35s_35_2_1_U17.top_add_35s_35s_35_2_1_Adder_12_U.u1.b ;
assign { \add_35s_35s_35_2_1_U17.top_add_35s_35s_35_2_1_Adder_12_U.u1.cout , \add_35s_35s_35_2_1_U17.top_add_35s_35s_35_2_1_Adder_12_U.u1.s  } = _129_ + \add_35s_35s_35_2_1_U17.top_add_35s_35s_35_2_1_Adder_12_U.u1.cin ;
assign _130_ = \add_35s_35s_35_2_1_U17.top_add_35s_35s_35_2_1_Adder_12_U.u2.a  + \add_35s_35s_35_2_1_U17.top_add_35s_35s_35_2_1_Adder_12_U.u2.b ;
assign { \add_35s_35s_35_2_1_U17.top_add_35s_35s_35_2_1_Adder_12_U.u2.cout , \add_35s_35s_35_2_1_U17.top_add_35s_35s_35_2_1_Adder_12_U.u2.s  } = _130_ + \add_35s_35s_35_2_1_U17.top_add_35s_35s_35_2_1_Adder_12_U.u2.cin ;
always @(posedge \add_36s_36s_36_2_1_U20.top_add_36s_36s_36_2_1_Adder_14_U.clk )
\add_36s_36s_36_2_1_U20.top_add_36s_36s_36_2_1_Adder_14_U.bin_s1  <= _132_;
always @(posedge \add_36s_36s_36_2_1_U20.top_add_36s_36s_36_2_1_Adder_14_U.clk )
\add_36s_36s_36_2_1_U20.top_add_36s_36s_36_2_1_Adder_14_U.ain_s1  <= _131_;
always @(posedge \add_36s_36s_36_2_1_U20.top_add_36s_36s_36_2_1_Adder_14_U.clk )
\add_36s_36s_36_2_1_U20.top_add_36s_36s_36_2_1_Adder_14_U.sum_s1  <= _134_;
always @(posedge \add_36s_36s_36_2_1_U20.top_add_36s_36s_36_2_1_Adder_14_U.clk )
\add_36s_36s_36_2_1_U20.top_add_36s_36s_36_2_1_Adder_14_U.carry_s1  <= _133_;
assign _132_ = \add_36s_36s_36_2_1_U20.top_add_36s_36s_36_2_1_Adder_14_U.ce  ? \add_36s_36s_36_2_1_U20.top_add_36s_36s_36_2_1_Adder_14_U.b [35:18] : \add_36s_36s_36_2_1_U20.top_add_36s_36s_36_2_1_Adder_14_U.bin_s1 ;
assign _131_ = \add_36s_36s_36_2_1_U20.top_add_36s_36s_36_2_1_Adder_14_U.ce  ? \add_36s_36s_36_2_1_U20.top_add_36s_36s_36_2_1_Adder_14_U.a [35:18] : \add_36s_36s_36_2_1_U20.top_add_36s_36s_36_2_1_Adder_14_U.ain_s1 ;
assign _133_ = \add_36s_36s_36_2_1_U20.top_add_36s_36s_36_2_1_Adder_14_U.ce  ? \add_36s_36s_36_2_1_U20.top_add_36s_36s_36_2_1_Adder_14_U.facout_s1  : \add_36s_36s_36_2_1_U20.top_add_36s_36s_36_2_1_Adder_14_U.carry_s1 ;
assign _134_ = \add_36s_36s_36_2_1_U20.top_add_36s_36s_36_2_1_Adder_14_U.ce  ? \add_36s_36s_36_2_1_U20.top_add_36s_36s_36_2_1_Adder_14_U.fas_s1  : \add_36s_36s_36_2_1_U20.top_add_36s_36s_36_2_1_Adder_14_U.sum_s1 ;
assign _135_ = \add_36s_36s_36_2_1_U20.top_add_36s_36s_36_2_1_Adder_14_U.u1.a  + \add_36s_36s_36_2_1_U20.top_add_36s_36s_36_2_1_Adder_14_U.u1.b ;
assign { \add_36s_36s_36_2_1_U20.top_add_36s_36s_36_2_1_Adder_14_U.u1.cout , \add_36s_36s_36_2_1_U20.top_add_36s_36s_36_2_1_Adder_14_U.u1.s  } = _135_ + \add_36s_36s_36_2_1_U20.top_add_36s_36s_36_2_1_Adder_14_U.u1.cin ;
assign _136_ = \add_36s_36s_36_2_1_U20.top_add_36s_36s_36_2_1_Adder_14_U.u2.a  + \add_36s_36s_36_2_1_U20.top_add_36s_36s_36_2_1_Adder_14_U.u2.b ;
assign { \add_36s_36s_36_2_1_U20.top_add_36s_36s_36_2_1_Adder_14_U.u2.cout , \add_36s_36s_36_2_1_U20.top_add_36s_36s_36_2_1_Adder_14_U.u2.s  } = _136_ + \add_36s_36s_36_2_1_U20.top_add_36s_36s_36_2_1_Adder_14_U.u2.cin ;
always @(posedge \add_3s_3s_3_2_1_U15.top_add_3s_3s_3_2_1_Adder_11_U.clk )
\add_3s_3s_3_2_1_U15.top_add_3s_3s_3_2_1_Adder_11_U.bin_s1  <= _138_;
always @(posedge \add_3s_3s_3_2_1_U15.top_add_3s_3s_3_2_1_Adder_11_U.clk )
\add_3s_3s_3_2_1_U15.top_add_3s_3s_3_2_1_Adder_11_U.ain_s1  <= _137_;
always @(posedge \add_3s_3s_3_2_1_U15.top_add_3s_3s_3_2_1_Adder_11_U.clk )
\add_3s_3s_3_2_1_U15.top_add_3s_3s_3_2_1_Adder_11_U.sum_s1  <= _140_;
always @(posedge \add_3s_3s_3_2_1_U15.top_add_3s_3s_3_2_1_Adder_11_U.clk )
\add_3s_3s_3_2_1_U15.top_add_3s_3s_3_2_1_Adder_11_U.carry_s1  <= _139_;
assign _138_ = \add_3s_3s_3_2_1_U15.top_add_3s_3s_3_2_1_Adder_11_U.ce  ? \add_3s_3s_3_2_1_U15.top_add_3s_3s_3_2_1_Adder_11_U.b [2:1] : \add_3s_3s_3_2_1_U15.top_add_3s_3s_3_2_1_Adder_11_U.bin_s1 ;
assign _137_ = \add_3s_3s_3_2_1_U15.top_add_3s_3s_3_2_1_Adder_11_U.ce  ? \add_3s_3s_3_2_1_U15.top_add_3s_3s_3_2_1_Adder_11_U.a [2:1] : \add_3s_3s_3_2_1_U15.top_add_3s_3s_3_2_1_Adder_11_U.ain_s1 ;
assign _139_ = \add_3s_3s_3_2_1_U15.top_add_3s_3s_3_2_1_Adder_11_U.ce  ? \add_3s_3s_3_2_1_U15.top_add_3s_3s_3_2_1_Adder_11_U.facout_s1  : \add_3s_3s_3_2_1_U15.top_add_3s_3s_3_2_1_Adder_11_U.carry_s1 ;
assign _140_ = \add_3s_3s_3_2_1_U15.top_add_3s_3s_3_2_1_Adder_11_U.ce  ? \add_3s_3s_3_2_1_U15.top_add_3s_3s_3_2_1_Adder_11_U.fas_s1  : \add_3s_3s_3_2_1_U15.top_add_3s_3s_3_2_1_Adder_11_U.sum_s1 ;
assign _141_ = \add_3s_3s_3_2_1_U15.top_add_3s_3s_3_2_1_Adder_11_U.u1.a  + \add_3s_3s_3_2_1_U15.top_add_3s_3s_3_2_1_Adder_11_U.u1.b ;
assign { \add_3s_3s_3_2_1_U15.top_add_3s_3s_3_2_1_Adder_11_U.u1.cout , \add_3s_3s_3_2_1_U15.top_add_3s_3s_3_2_1_Adder_11_U.u1.s  } = _141_ + \add_3s_3s_3_2_1_U15.top_add_3s_3s_3_2_1_Adder_11_U.u1.cin ;
assign _142_ = \add_3s_3s_3_2_1_U15.top_add_3s_3s_3_2_1_Adder_11_U.u2.a  + \add_3s_3s_3_2_1_U15.top_add_3s_3s_3_2_1_Adder_11_U.u2.b ;
assign { \add_3s_3s_3_2_1_U15.top_add_3s_3s_3_2_1_Adder_11_U.u2.cout , \add_3s_3s_3_2_1_U15.top_add_3s_3s_3_2_1_Adder_11_U.u2.s  } = _142_ + \add_3s_3s_3_2_1_U15.top_add_3s_3s_3_2_1_Adder_11_U.u2.cin ;
always @(posedge \add_4s_4ns_4_2_1_U8.top_add_4s_4ns_4_2_1_Adder_5_U.clk )
\add_4s_4ns_4_2_1_U8.top_add_4s_4ns_4_2_1_Adder_5_U.bin_s1  <= _144_;
always @(posedge \add_4s_4ns_4_2_1_U8.top_add_4s_4ns_4_2_1_Adder_5_U.clk )
\add_4s_4ns_4_2_1_U8.top_add_4s_4ns_4_2_1_Adder_5_U.ain_s1  <= _143_;
always @(posedge \add_4s_4ns_4_2_1_U8.top_add_4s_4ns_4_2_1_Adder_5_U.clk )
\add_4s_4ns_4_2_1_U8.top_add_4s_4ns_4_2_1_Adder_5_U.sum_s1  <= _146_;
always @(posedge \add_4s_4ns_4_2_1_U8.top_add_4s_4ns_4_2_1_Adder_5_U.clk )
\add_4s_4ns_4_2_1_U8.top_add_4s_4ns_4_2_1_Adder_5_U.carry_s1  <= _145_;
assign _144_ = \add_4s_4ns_4_2_1_U8.top_add_4s_4ns_4_2_1_Adder_5_U.ce  ? \add_4s_4ns_4_2_1_U8.top_add_4s_4ns_4_2_1_Adder_5_U.b [3:2] : \add_4s_4ns_4_2_1_U8.top_add_4s_4ns_4_2_1_Adder_5_U.bin_s1 ;
assign _143_ = \add_4s_4ns_4_2_1_U8.top_add_4s_4ns_4_2_1_Adder_5_U.ce  ? \add_4s_4ns_4_2_1_U8.top_add_4s_4ns_4_2_1_Adder_5_U.a [3:2] : \add_4s_4ns_4_2_1_U8.top_add_4s_4ns_4_2_1_Adder_5_U.ain_s1 ;
assign _145_ = \add_4s_4ns_4_2_1_U8.top_add_4s_4ns_4_2_1_Adder_5_U.ce  ? \add_4s_4ns_4_2_1_U8.top_add_4s_4ns_4_2_1_Adder_5_U.facout_s1  : \add_4s_4ns_4_2_1_U8.top_add_4s_4ns_4_2_1_Adder_5_U.carry_s1 ;
assign _146_ = \add_4s_4ns_4_2_1_U8.top_add_4s_4ns_4_2_1_Adder_5_U.ce  ? \add_4s_4ns_4_2_1_U8.top_add_4s_4ns_4_2_1_Adder_5_U.fas_s1  : \add_4s_4ns_4_2_1_U8.top_add_4s_4ns_4_2_1_Adder_5_U.sum_s1 ;
assign _147_ = \add_4s_4ns_4_2_1_U8.top_add_4s_4ns_4_2_1_Adder_5_U.u1.a  + \add_4s_4ns_4_2_1_U8.top_add_4s_4ns_4_2_1_Adder_5_U.u1.b ;
assign { \add_4s_4ns_4_2_1_U8.top_add_4s_4ns_4_2_1_Adder_5_U.u1.cout , \add_4s_4ns_4_2_1_U8.top_add_4s_4ns_4_2_1_Adder_5_U.u1.s  } = _147_ + \add_4s_4ns_4_2_1_U8.top_add_4s_4ns_4_2_1_Adder_5_U.u1.cin ;
assign _148_ = \add_4s_4ns_4_2_1_U8.top_add_4s_4ns_4_2_1_Adder_5_U.u2.a  + \add_4s_4ns_4_2_1_U8.top_add_4s_4ns_4_2_1_Adder_5_U.u2.b ;
assign { \add_4s_4ns_4_2_1_U8.top_add_4s_4ns_4_2_1_Adder_5_U.u2.cout , \add_4s_4ns_4_2_1_U8.top_add_4s_4ns_4_2_1_Adder_5_U.u2.s  } = _148_ + \add_4s_4ns_4_2_1_U8.top_add_4s_4ns_4_2_1_Adder_5_U.u2.cin ;
always @(posedge \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_4_U.clk )
\add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_4_U.bin_s1  <= _150_;
always @(posedge \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_4_U.clk )
\add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_4_U.ain_s1  <= _149_;
always @(posedge \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_4_U.clk )
\add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_4_U.sum_s1  <= _152_;
always @(posedge \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_4_U.clk )
\add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_4_U.carry_s1  <= _151_;
assign _150_ = \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_4_U.ce  ? \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_4_U.b [5:3] : \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_4_U.bin_s1 ;
assign _149_ = \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_4_U.ce  ? \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_4_U.a [5:3] : \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_4_U.ain_s1 ;
assign _151_ = \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_4_U.ce  ? \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_4_U.facout_s1  : \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_4_U.carry_s1 ;
assign _152_ = \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_4_U.ce  ? \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_4_U.fas_s1  : \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_4_U.sum_s1 ;
assign _153_ = \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_4_U.u1.a  + \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_4_U.u1.b ;
assign { \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_4_U.u1.cout , \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_4_U.u1.s  } = _153_ + \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_4_U.u1.cin ;
assign _154_ = \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_4_U.u2.a  + \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_4_U.u2.b ;
assign { \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_4_U.u2.cout , \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_4_U.u2.s  } = _154_ + \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_4_U.u2.cin ;
always @(posedge \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.clk )
\add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.bin_s1  <= _156_;
always @(posedge \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.clk )
\add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.ain_s1  <= _155_;
always @(posedge \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.clk )
\add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.sum_s1  <= _158_;
always @(posedge \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.clk )
\add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.carry_s1  <= _157_;
assign _156_ = \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.ce  ? \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.b [5:3] : \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.bin_s1 ;
assign _155_ = \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.ce  ? \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.a [5:3] : \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.ain_s1 ;
assign _157_ = \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.ce  ? \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.facout_s1  : \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.carry_s1 ;
assign _158_ = \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.ce  ? \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.fas_s1  : \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.sum_s1 ;
assign _159_ = \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.u1.a  + \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.u1.b ;
assign { \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.u1.cout , \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.u1.s  } = _159_ + \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.u1.cin ;
assign _160_ = \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.u2.a  + \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.u2.b ;
assign { \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.u2.cout , \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.u2.s  } = _160_ + \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.u2.cin ;
always @(posedge \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_10_U.clk )
\add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_10_U.bin_s1  <= _162_;
always @(posedge \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_10_U.clk )
\add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_10_U.ain_s1  <= _161_;
always @(posedge \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_10_U.clk )
\add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_10_U.sum_s1  <= _164_;
always @(posedge \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_10_U.clk )
\add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_10_U.carry_s1  <= _163_;
assign _162_ = \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_10_U.ce  ? \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_10_U.b [6:3] : \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_10_U.bin_s1 ;
assign _161_ = \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_10_U.ce  ? \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_10_U.a [6:3] : \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_10_U.ain_s1 ;
assign _163_ = \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_10_U.ce  ? \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_10_U.facout_s1  : \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_10_U.carry_s1 ;
assign _164_ = \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_10_U.ce  ? \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_10_U.fas_s1  : \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_10_U.sum_s1 ;
assign _165_ = \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_10_U.u1.a  + \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_10_U.u1.b ;
assign { \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_10_U.u1.cout , \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_10_U.u1.s  } = _165_ + \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_10_U.u1.cin ;
assign _166_ = \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_10_U.u2.a  + \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_10_U.u2.b ;
assign { \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_10_U.u2.cout , \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_10_U.u2.s  } = _166_ + \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_10_U.u2.cin ;
always @(posedge \add_7s_7ns_7_2_1_U16.top_add_7s_7ns_7_2_1_Adder_10_U.clk )
\add_7s_7ns_7_2_1_U16.top_add_7s_7ns_7_2_1_Adder_10_U.bin_s1  <= _168_;
always @(posedge \add_7s_7ns_7_2_1_U16.top_add_7s_7ns_7_2_1_Adder_10_U.clk )
\add_7s_7ns_7_2_1_U16.top_add_7s_7ns_7_2_1_Adder_10_U.ain_s1  <= _167_;
always @(posedge \add_7s_7ns_7_2_1_U16.top_add_7s_7ns_7_2_1_Adder_10_U.clk )
\add_7s_7ns_7_2_1_U16.top_add_7s_7ns_7_2_1_Adder_10_U.sum_s1  <= _170_;
always @(posedge \add_7s_7ns_7_2_1_U16.top_add_7s_7ns_7_2_1_Adder_10_U.clk )
\add_7s_7ns_7_2_1_U16.top_add_7s_7ns_7_2_1_Adder_10_U.carry_s1  <= _169_;
assign _168_ = \add_7s_7ns_7_2_1_U16.top_add_7s_7ns_7_2_1_Adder_10_U.ce  ? \add_7s_7ns_7_2_1_U16.top_add_7s_7ns_7_2_1_Adder_10_U.b [6:3] : \add_7s_7ns_7_2_1_U16.top_add_7s_7ns_7_2_1_Adder_10_U.bin_s1 ;
assign _167_ = \add_7s_7ns_7_2_1_U16.top_add_7s_7ns_7_2_1_Adder_10_U.ce  ? \add_7s_7ns_7_2_1_U16.top_add_7s_7ns_7_2_1_Adder_10_U.a [6:3] : \add_7s_7ns_7_2_1_U16.top_add_7s_7ns_7_2_1_Adder_10_U.ain_s1 ;
assign _169_ = \add_7s_7ns_7_2_1_U16.top_add_7s_7ns_7_2_1_Adder_10_U.ce  ? \add_7s_7ns_7_2_1_U16.top_add_7s_7ns_7_2_1_Adder_10_U.facout_s1  : \add_7s_7ns_7_2_1_U16.top_add_7s_7ns_7_2_1_Adder_10_U.carry_s1 ;
assign _170_ = \add_7s_7ns_7_2_1_U16.top_add_7s_7ns_7_2_1_Adder_10_U.ce  ? \add_7s_7ns_7_2_1_U16.top_add_7s_7ns_7_2_1_Adder_10_U.fas_s1  : \add_7s_7ns_7_2_1_U16.top_add_7s_7ns_7_2_1_Adder_10_U.sum_s1 ;
assign _171_ = \add_7s_7ns_7_2_1_U16.top_add_7s_7ns_7_2_1_Adder_10_U.u1.a  + \add_7s_7ns_7_2_1_U16.top_add_7s_7ns_7_2_1_Adder_10_U.u1.b ;
assign { \add_7s_7ns_7_2_1_U16.top_add_7s_7ns_7_2_1_Adder_10_U.u1.cout , \add_7s_7ns_7_2_1_U16.top_add_7s_7ns_7_2_1_Adder_10_U.u1.s  } = _171_ + \add_7s_7ns_7_2_1_U16.top_add_7s_7ns_7_2_1_Adder_10_U.u1.cin ;
assign _172_ = \add_7s_7ns_7_2_1_U16.top_add_7s_7ns_7_2_1_Adder_10_U.u2.a  + \add_7s_7ns_7_2_1_U16.top_add_7s_7ns_7_2_1_Adder_10_U.u2.b ;
assign { \add_7s_7ns_7_2_1_U16.top_add_7s_7ns_7_2_1_Adder_10_U.u2.cout , \add_7s_7ns_7_2_1_U16.top_add_7s_7ns_7_2_1_Adder_10_U.u2.s  } = _172_ + \add_7s_7ns_7_2_1_U16.top_add_7s_7ns_7_2_1_Adder_10_U.u2.cin ;
always @(posedge \add_7s_7s_7_2_1_U11.top_add_7s_7s_7_2_1_Adder_8_U.clk )
\add_7s_7s_7_2_1_U11.top_add_7s_7s_7_2_1_Adder_8_U.bin_s1  <= _174_;
always @(posedge \add_7s_7s_7_2_1_U11.top_add_7s_7s_7_2_1_Adder_8_U.clk )
\add_7s_7s_7_2_1_U11.top_add_7s_7s_7_2_1_Adder_8_U.ain_s1  <= _173_;
always @(posedge \add_7s_7s_7_2_1_U11.top_add_7s_7s_7_2_1_Adder_8_U.clk )
\add_7s_7s_7_2_1_U11.top_add_7s_7s_7_2_1_Adder_8_U.sum_s1  <= _176_;
always @(posedge \add_7s_7s_7_2_1_U11.top_add_7s_7s_7_2_1_Adder_8_U.clk )
\add_7s_7s_7_2_1_U11.top_add_7s_7s_7_2_1_Adder_8_U.carry_s1  <= _175_;
assign _174_ = \add_7s_7s_7_2_1_U11.top_add_7s_7s_7_2_1_Adder_8_U.ce  ? \add_7s_7s_7_2_1_U11.top_add_7s_7s_7_2_1_Adder_8_U.b [6:3] : \add_7s_7s_7_2_1_U11.top_add_7s_7s_7_2_1_Adder_8_U.bin_s1 ;
assign _173_ = \add_7s_7s_7_2_1_U11.top_add_7s_7s_7_2_1_Adder_8_U.ce  ? \add_7s_7s_7_2_1_U11.top_add_7s_7s_7_2_1_Adder_8_U.a [6:3] : \add_7s_7s_7_2_1_U11.top_add_7s_7s_7_2_1_Adder_8_U.ain_s1 ;
assign _175_ = \add_7s_7s_7_2_1_U11.top_add_7s_7s_7_2_1_Adder_8_U.ce  ? \add_7s_7s_7_2_1_U11.top_add_7s_7s_7_2_1_Adder_8_U.facout_s1  : \add_7s_7s_7_2_1_U11.top_add_7s_7s_7_2_1_Adder_8_U.carry_s1 ;
assign _176_ = \add_7s_7s_7_2_1_U11.top_add_7s_7s_7_2_1_Adder_8_U.ce  ? \add_7s_7s_7_2_1_U11.top_add_7s_7s_7_2_1_Adder_8_U.fas_s1  : \add_7s_7s_7_2_1_U11.top_add_7s_7s_7_2_1_Adder_8_U.sum_s1 ;
assign _177_ = \add_7s_7s_7_2_1_U11.top_add_7s_7s_7_2_1_Adder_8_U.u1.a  + \add_7s_7s_7_2_1_U11.top_add_7s_7s_7_2_1_Adder_8_U.u1.b ;
assign { \add_7s_7s_7_2_1_U11.top_add_7s_7s_7_2_1_Adder_8_U.u1.cout , \add_7s_7s_7_2_1_U11.top_add_7s_7s_7_2_1_Adder_8_U.u1.s  } = _177_ + \add_7s_7s_7_2_1_U11.top_add_7s_7s_7_2_1_Adder_8_U.u1.cin ;
assign _178_ = \add_7s_7s_7_2_1_U11.top_add_7s_7s_7_2_1_Adder_8_U.u2.a  + \add_7s_7s_7_2_1_U11.top_add_7s_7s_7_2_1_Adder_8_U.u2.b ;
assign { \add_7s_7s_7_2_1_U11.top_add_7s_7s_7_2_1_Adder_8_U.u2.cout , \add_7s_7s_7_2_1_U11.top_add_7s_7s_7_2_1_Adder_8_U.u2.s  } = _178_ + \add_7s_7s_7_2_1_U11.top_add_7s_7s_7_2_1_Adder_8_U.u2.cin ;
always @(posedge \add_9s_9ns_9_2_1_U6.top_add_9s_9ns_9_2_1_Adder_3_U.clk )
\add_9s_9ns_9_2_1_U6.top_add_9s_9ns_9_2_1_Adder_3_U.bin_s1  <= _180_;
always @(posedge \add_9s_9ns_9_2_1_U6.top_add_9s_9ns_9_2_1_Adder_3_U.clk )
\add_9s_9ns_9_2_1_U6.top_add_9s_9ns_9_2_1_Adder_3_U.ain_s1  <= _179_;
always @(posedge \add_9s_9ns_9_2_1_U6.top_add_9s_9ns_9_2_1_Adder_3_U.clk )
\add_9s_9ns_9_2_1_U6.top_add_9s_9ns_9_2_1_Adder_3_U.sum_s1  <= _182_;
always @(posedge \add_9s_9ns_9_2_1_U6.top_add_9s_9ns_9_2_1_Adder_3_U.clk )
\add_9s_9ns_9_2_1_U6.top_add_9s_9ns_9_2_1_Adder_3_U.carry_s1  <= _181_;
assign _180_ = \add_9s_9ns_9_2_1_U6.top_add_9s_9ns_9_2_1_Adder_3_U.ce  ? \add_9s_9ns_9_2_1_U6.top_add_9s_9ns_9_2_1_Adder_3_U.b [8:4] : \add_9s_9ns_9_2_1_U6.top_add_9s_9ns_9_2_1_Adder_3_U.bin_s1 ;
assign _179_ = \add_9s_9ns_9_2_1_U6.top_add_9s_9ns_9_2_1_Adder_3_U.ce  ? \add_9s_9ns_9_2_1_U6.top_add_9s_9ns_9_2_1_Adder_3_U.a [8:4] : \add_9s_9ns_9_2_1_U6.top_add_9s_9ns_9_2_1_Adder_3_U.ain_s1 ;
assign _181_ = \add_9s_9ns_9_2_1_U6.top_add_9s_9ns_9_2_1_Adder_3_U.ce  ? \add_9s_9ns_9_2_1_U6.top_add_9s_9ns_9_2_1_Adder_3_U.facout_s1  : \add_9s_9ns_9_2_1_U6.top_add_9s_9ns_9_2_1_Adder_3_U.carry_s1 ;
assign _182_ = \add_9s_9ns_9_2_1_U6.top_add_9s_9ns_9_2_1_Adder_3_U.ce  ? \add_9s_9ns_9_2_1_U6.top_add_9s_9ns_9_2_1_Adder_3_U.fas_s1  : \add_9s_9ns_9_2_1_U6.top_add_9s_9ns_9_2_1_Adder_3_U.sum_s1 ;
assign _183_ = \add_9s_9ns_9_2_1_U6.top_add_9s_9ns_9_2_1_Adder_3_U.u1.a  + \add_9s_9ns_9_2_1_U6.top_add_9s_9ns_9_2_1_Adder_3_U.u1.b ;
assign { \add_9s_9ns_9_2_1_U6.top_add_9s_9ns_9_2_1_Adder_3_U.u1.cout , \add_9s_9ns_9_2_1_U6.top_add_9s_9ns_9_2_1_Adder_3_U.u1.s  } = _183_ + \add_9s_9ns_9_2_1_U6.top_add_9s_9ns_9_2_1_Adder_3_U.u1.cin ;
assign _184_ = \add_9s_9ns_9_2_1_U6.top_add_9s_9ns_9_2_1_Adder_3_U.u2.a  + \add_9s_9ns_9_2_1_U6.top_add_9s_9ns_9_2_1_Adder_3_U.u2.b ;
assign { \add_9s_9ns_9_2_1_U6.top_add_9s_9ns_9_2_1_Adder_3_U.u2.cout , \add_9s_9ns_9_2_1_U6.top_add_9s_9ns_9_2_1_Adder_3_U.u2.s  } = _184_ + \add_9s_9ns_9_2_1_U6.top_add_9s_9ns_9_2_1_Adder_3_U.u2.cin ;
always @(posedge \ashr_4s_2ns_4_7_1_U3.clk )
\ashr_4s_2ns_4_7_1_U3.dout_array[5]  <= _196_;
always @(posedge \ashr_4s_2ns_4_7_1_U3.clk )
\ashr_4s_2ns_4_7_1_U3.din1_cast_array[5]  <= _190_;
always @(posedge \ashr_4s_2ns_4_7_1_U3.clk )
\ashr_4s_2ns_4_7_1_U3.dout_array[4]  <= _195_;
always @(posedge \ashr_4s_2ns_4_7_1_U3.clk )
\ashr_4s_2ns_4_7_1_U3.din1_cast_array[4]  <= _189_;
always @(posedge \ashr_4s_2ns_4_7_1_U3.clk )
\ashr_4s_2ns_4_7_1_U3.dout_array[3]  <= _194_;
always @(posedge \ashr_4s_2ns_4_7_1_U3.clk )
\ashr_4s_2ns_4_7_1_U3.din1_cast_array[3]  <= _188_;
always @(posedge \ashr_4s_2ns_4_7_1_U3.clk )
\ashr_4s_2ns_4_7_1_U3.dout_array[2]  <= _193_;
always @(posedge \ashr_4s_2ns_4_7_1_U3.clk )
\ashr_4s_2ns_4_7_1_U3.din1_cast_array[2]  <= _187_;
always @(posedge \ashr_4s_2ns_4_7_1_U3.clk )
\ashr_4s_2ns_4_7_1_U3.dout_array[1]  <= _192_;
always @(posedge \ashr_4s_2ns_4_7_1_U3.clk )
\ashr_4s_2ns_4_7_1_U3.din1_cast_array[1]  <= _186_;
always @(posedge \ashr_4s_2ns_4_7_1_U3.clk )
\ashr_4s_2ns_4_7_1_U3.dout_array[0]  <= _191_;
always @(posedge \ashr_4s_2ns_4_7_1_U3.clk )
\ashr_4s_2ns_4_7_1_U3.din1_cast_array[0]  <= _185_;
assign _197_ = \ashr_4s_2ns_4_7_1_U3.ce  ? \ashr_4s_2ns_4_7_1_U3.din1_cast_array[4]  : \ashr_4s_2ns_4_7_1_U3.din1_cast_array[5] ;
assign _190_ = \ashr_4s_2ns_4_7_1_U3.reset  ? 2'h0 : _197_;
assign _198_ = \ashr_4s_2ns_4_7_1_U3.ce  ? _209_ : \ashr_4s_2ns_4_7_1_U3.dout_array[5] ;
assign _196_ = \ashr_4s_2ns_4_7_1_U3.reset  ? 4'h0 : _198_;
assign _199_ = \ashr_4s_2ns_4_7_1_U3.ce  ? \ashr_4s_2ns_4_7_1_U3.din1_cast_array[3]  : \ashr_4s_2ns_4_7_1_U3.din1_cast_array[4] ;
assign _189_ = \ashr_4s_2ns_4_7_1_U3.reset  ? 2'h0 : _199_;
assign _200_ = \ashr_4s_2ns_4_7_1_U3.ce  ? \ashr_4s_2ns_4_7_1_U3.dout_array[3]  : \ashr_4s_2ns_4_7_1_U3.dout_array[4] ;
assign _195_ = \ashr_4s_2ns_4_7_1_U3.reset  ? 4'h0 : _200_;
assign _201_ = \ashr_4s_2ns_4_7_1_U3.ce  ? \ashr_4s_2ns_4_7_1_U3.din1_cast_array[2]  : \ashr_4s_2ns_4_7_1_U3.din1_cast_array[3] ;
assign _188_ = \ashr_4s_2ns_4_7_1_U3.reset  ? 2'h0 : _201_;
assign _202_ = \ashr_4s_2ns_4_7_1_U3.ce  ? \ashr_4s_2ns_4_7_1_U3.dout_array[2]  : \ashr_4s_2ns_4_7_1_U3.dout_array[3] ;
assign _194_ = \ashr_4s_2ns_4_7_1_U3.reset  ? 4'h0 : _202_;
assign _203_ = \ashr_4s_2ns_4_7_1_U3.ce  ? \ashr_4s_2ns_4_7_1_U3.din1_cast_array[1]  : \ashr_4s_2ns_4_7_1_U3.din1_cast_array[2] ;
assign _187_ = \ashr_4s_2ns_4_7_1_U3.reset  ? 2'h0 : _203_;
assign _204_ = \ashr_4s_2ns_4_7_1_U3.ce  ? \ashr_4s_2ns_4_7_1_U3.dout_array[1]  : \ashr_4s_2ns_4_7_1_U3.dout_array[2] ;
assign _193_ = \ashr_4s_2ns_4_7_1_U3.reset  ? 4'h0 : _204_;
assign _205_ = \ashr_4s_2ns_4_7_1_U3.ce  ? \ashr_4s_2ns_4_7_1_U3.din1_cast_array[0]  : \ashr_4s_2ns_4_7_1_U3.din1_cast_array[1] ;
assign _186_ = \ashr_4s_2ns_4_7_1_U3.reset  ? 2'h0 : _205_;
assign _206_ = \ashr_4s_2ns_4_7_1_U3.ce  ? \ashr_4s_2ns_4_7_1_U3.dout_array[0]  : \ashr_4s_2ns_4_7_1_U3.dout_array[1] ;
assign _192_ = \ashr_4s_2ns_4_7_1_U3.reset  ? 4'h0 : _206_;
assign _207_ = \ashr_4s_2ns_4_7_1_U3.ce  ? \ashr_4s_2ns_4_7_1_U3.din1 [1:0] : \ashr_4s_2ns_4_7_1_U3.din1_cast_array[0] ;
assign _185_ = \ashr_4s_2ns_4_7_1_U3.reset  ? 2'h0 : _207_;
assign _208_ = \ashr_4s_2ns_4_7_1_U3.ce  ? \ashr_4s_2ns_4_7_1_U3.din0  : \ashr_4s_2ns_4_7_1_U3.dout_array[0] ;
assign _191_ = \ashr_4s_2ns_4_7_1_U3.reset  ? 4'h0 : _208_;
assign _209_ = $signed(\ashr_4s_2ns_4_7_1_U3.dout_array[4] ) >>> { \ashr_4s_2ns_4_7_1_U3.din1_cast_array[4] [1], 1'h0 };
assign \ashr_4s_2ns_4_7_1_U3.dout  = $signed(\ashr_4s_2ns_4_7_1_U3.dout_array[5] ) >>> \ashr_4s_2ns_4_7_1_U3.din1_cast_array[5] [0];
always @(posedge \shl_4s_2ns_4_7_1_U4.clk )
\shl_4s_2ns_4_7_1_U4.dout_array[5]  <= _221_;
always @(posedge \shl_4s_2ns_4_7_1_U4.clk )
\shl_4s_2ns_4_7_1_U4.din1_cast_array[5]  <= _215_;
always @(posedge \shl_4s_2ns_4_7_1_U4.clk )
\shl_4s_2ns_4_7_1_U4.dout_array[4]  <= _220_;
always @(posedge \shl_4s_2ns_4_7_1_U4.clk )
\shl_4s_2ns_4_7_1_U4.din1_cast_array[4]  <= _214_;
always @(posedge \shl_4s_2ns_4_7_1_U4.clk )
\shl_4s_2ns_4_7_1_U4.dout_array[3]  <= _219_;
always @(posedge \shl_4s_2ns_4_7_1_U4.clk )
\shl_4s_2ns_4_7_1_U4.din1_cast_array[3]  <= _213_;
always @(posedge \shl_4s_2ns_4_7_1_U4.clk )
\shl_4s_2ns_4_7_1_U4.dout_array[2]  <= _218_;
always @(posedge \shl_4s_2ns_4_7_1_U4.clk )
\shl_4s_2ns_4_7_1_U4.din1_cast_array[2]  <= _212_;
always @(posedge \shl_4s_2ns_4_7_1_U4.clk )
\shl_4s_2ns_4_7_1_U4.dout_array[1]  <= _217_;
always @(posedge \shl_4s_2ns_4_7_1_U4.clk )
\shl_4s_2ns_4_7_1_U4.din1_cast_array[1]  <= _211_;
always @(posedge \shl_4s_2ns_4_7_1_U4.clk )
\shl_4s_2ns_4_7_1_U4.dout_array[0]  <= _216_;
always @(posedge \shl_4s_2ns_4_7_1_U4.clk )
\shl_4s_2ns_4_7_1_U4.din1_cast_array[0]  <= _210_;
assign _222_ = \shl_4s_2ns_4_7_1_U4.ce  ? \shl_4s_2ns_4_7_1_U4.din1_cast_array[4]  : \shl_4s_2ns_4_7_1_U4.din1_cast_array[5] ;
assign _215_ = \shl_4s_2ns_4_7_1_U4.reset  ? 2'h0 : _222_;
assign _223_ = \shl_4s_2ns_4_7_1_U4.ce  ? _234_ : \shl_4s_2ns_4_7_1_U4.dout_array[5] ;
assign _221_ = \shl_4s_2ns_4_7_1_U4.reset  ? 4'h0 : _223_;
assign _224_ = \shl_4s_2ns_4_7_1_U4.ce  ? \shl_4s_2ns_4_7_1_U4.din1_cast_array[3]  : \shl_4s_2ns_4_7_1_U4.din1_cast_array[4] ;
assign _214_ = \shl_4s_2ns_4_7_1_U4.reset  ? 2'h0 : _224_;
assign _225_ = \shl_4s_2ns_4_7_1_U4.ce  ? \shl_4s_2ns_4_7_1_U4.dout_array[3]  : \shl_4s_2ns_4_7_1_U4.dout_array[4] ;
assign _220_ = \shl_4s_2ns_4_7_1_U4.reset  ? 4'h0 : _225_;
assign _226_ = \shl_4s_2ns_4_7_1_U4.ce  ? \shl_4s_2ns_4_7_1_U4.din1_cast_array[2]  : \shl_4s_2ns_4_7_1_U4.din1_cast_array[3] ;
assign _213_ = \shl_4s_2ns_4_7_1_U4.reset  ? 2'h0 : _226_;
assign _227_ = \shl_4s_2ns_4_7_1_U4.ce  ? \shl_4s_2ns_4_7_1_U4.dout_array[2]  : \shl_4s_2ns_4_7_1_U4.dout_array[3] ;
assign _219_ = \shl_4s_2ns_4_7_1_U4.reset  ? 4'h0 : _227_;
assign _228_ = \shl_4s_2ns_4_7_1_U4.ce  ? \shl_4s_2ns_4_7_1_U4.din1_cast_array[1]  : \shl_4s_2ns_4_7_1_U4.din1_cast_array[2] ;
assign _212_ = \shl_4s_2ns_4_7_1_U4.reset  ? 2'h0 : _228_;
assign _229_ = \shl_4s_2ns_4_7_1_U4.ce  ? \shl_4s_2ns_4_7_1_U4.dout_array[1]  : \shl_4s_2ns_4_7_1_U4.dout_array[2] ;
assign _218_ = \shl_4s_2ns_4_7_1_U4.reset  ? 4'h0 : _229_;
assign _230_ = \shl_4s_2ns_4_7_1_U4.ce  ? \shl_4s_2ns_4_7_1_U4.din1_cast_array[0]  : \shl_4s_2ns_4_7_1_U4.din1_cast_array[1] ;
assign _211_ = \shl_4s_2ns_4_7_1_U4.reset  ? 2'h0 : _230_;
assign _231_ = \shl_4s_2ns_4_7_1_U4.ce  ? \shl_4s_2ns_4_7_1_U4.dout_array[0]  : \shl_4s_2ns_4_7_1_U4.dout_array[1] ;
assign _217_ = \shl_4s_2ns_4_7_1_U4.reset  ? 4'h0 : _231_;
assign _232_ = \shl_4s_2ns_4_7_1_U4.ce  ? \shl_4s_2ns_4_7_1_U4.din1 [1:0] : \shl_4s_2ns_4_7_1_U4.din1_cast_array[0] ;
assign _210_ = \shl_4s_2ns_4_7_1_U4.reset  ? 2'h0 : _232_;
assign _233_ = \shl_4s_2ns_4_7_1_U4.ce  ? \shl_4s_2ns_4_7_1_U4.din0  : \shl_4s_2ns_4_7_1_U4.dout_array[0] ;
assign _216_ = \shl_4s_2ns_4_7_1_U4.reset  ? 4'h0 : _233_;
assign _234_ = \shl_4s_2ns_4_7_1_U4.dout_array[4]  << { \shl_4s_2ns_4_7_1_U4.din1_cast_array[4] [1], 1'h0 };
assign \shl_4s_2ns_4_7_1_U4.dout  = \shl_4s_2ns_4_7_1_U4.dout_array[5]  << \shl_4s_2ns_4_7_1_U4.din1_cast_array[5] [0];
assign \sub_27ns_27s_27_2_1_U5.top_sub_27ns_27s_27_2_1_Adder_2_U.bin_s0  = ~ \sub_27ns_27s_27_2_1_U5.top_sub_27ns_27s_27_2_1_Adder_2_U.b ;
always @(posedge \sub_27ns_27s_27_2_1_U5.top_sub_27ns_27s_27_2_1_Adder_2_U.clk )
\sub_27ns_27s_27_2_1_U5.top_sub_27ns_27s_27_2_1_Adder_2_U.bin_s1  <= _236_;
always @(posedge \sub_27ns_27s_27_2_1_U5.top_sub_27ns_27s_27_2_1_Adder_2_U.clk )
\sub_27ns_27s_27_2_1_U5.top_sub_27ns_27s_27_2_1_Adder_2_U.ain_s1  <= _235_;
always @(posedge \sub_27ns_27s_27_2_1_U5.top_sub_27ns_27s_27_2_1_Adder_2_U.clk )
\sub_27ns_27s_27_2_1_U5.top_sub_27ns_27s_27_2_1_Adder_2_U.sum_s1  <= _238_;
always @(posedge \sub_27ns_27s_27_2_1_U5.top_sub_27ns_27s_27_2_1_Adder_2_U.clk )
\sub_27ns_27s_27_2_1_U5.top_sub_27ns_27s_27_2_1_Adder_2_U.carry_s1  <= _237_;
assign _236_ = \sub_27ns_27s_27_2_1_U5.top_sub_27ns_27s_27_2_1_Adder_2_U.ce  ? \sub_27ns_27s_27_2_1_U5.top_sub_27ns_27s_27_2_1_Adder_2_U.bin_s0 [26:13] : \sub_27ns_27s_27_2_1_U5.top_sub_27ns_27s_27_2_1_Adder_2_U.bin_s1 ;
assign _235_ = \sub_27ns_27s_27_2_1_U5.top_sub_27ns_27s_27_2_1_Adder_2_U.ce  ? \sub_27ns_27s_27_2_1_U5.top_sub_27ns_27s_27_2_1_Adder_2_U.a [26:13] : \sub_27ns_27s_27_2_1_U5.top_sub_27ns_27s_27_2_1_Adder_2_U.ain_s1 ;
assign _237_ = \sub_27ns_27s_27_2_1_U5.top_sub_27ns_27s_27_2_1_Adder_2_U.ce  ? \sub_27ns_27s_27_2_1_U5.top_sub_27ns_27s_27_2_1_Adder_2_U.facout_s1  : \sub_27ns_27s_27_2_1_U5.top_sub_27ns_27s_27_2_1_Adder_2_U.carry_s1 ;
assign _238_ = \sub_27ns_27s_27_2_1_U5.top_sub_27ns_27s_27_2_1_Adder_2_U.ce  ? \sub_27ns_27s_27_2_1_U5.top_sub_27ns_27s_27_2_1_Adder_2_U.fas_s1  : \sub_27ns_27s_27_2_1_U5.top_sub_27ns_27s_27_2_1_Adder_2_U.sum_s1 ;
assign _239_ = \sub_27ns_27s_27_2_1_U5.top_sub_27ns_27s_27_2_1_Adder_2_U.u1.a  + \sub_27ns_27s_27_2_1_U5.top_sub_27ns_27s_27_2_1_Adder_2_U.u1.b ;
assign { \sub_27ns_27s_27_2_1_U5.top_sub_27ns_27s_27_2_1_Adder_2_U.u1.cout , \sub_27ns_27s_27_2_1_U5.top_sub_27ns_27s_27_2_1_Adder_2_U.u1.s  } = _239_ + \sub_27ns_27s_27_2_1_U5.top_sub_27ns_27s_27_2_1_Adder_2_U.u1.cin ;
assign _240_ = \sub_27ns_27s_27_2_1_U5.top_sub_27ns_27s_27_2_1_Adder_2_U.u2.a  + \sub_27ns_27s_27_2_1_U5.top_sub_27ns_27s_27_2_1_Adder_2_U.u2.b ;
assign { \sub_27ns_27s_27_2_1_U5.top_sub_27ns_27s_27_2_1_Adder_2_U.u2.cout , \sub_27ns_27s_27_2_1_U5.top_sub_27ns_27s_27_2_1_Adder_2_U.u2.s  } = _240_ + \sub_27ns_27s_27_2_1_U5.top_sub_27ns_27s_27_2_1_Adder_2_U.u2.cin ;
assign \sub_2ns_2ns_2_2_1_U2.top_sub_2ns_2ns_2_2_1_Adder_1_U.bin_s0  = ~ \sub_2ns_2ns_2_2_1_U2.top_sub_2ns_2ns_2_2_1_Adder_1_U.b ;
always @(posedge \sub_2ns_2ns_2_2_1_U2.top_sub_2ns_2ns_2_2_1_Adder_1_U.clk )
\sub_2ns_2ns_2_2_1_U2.top_sub_2ns_2ns_2_2_1_Adder_1_U.bin_s1  <= _242_;
always @(posedge \sub_2ns_2ns_2_2_1_U2.top_sub_2ns_2ns_2_2_1_Adder_1_U.clk )
\sub_2ns_2ns_2_2_1_U2.top_sub_2ns_2ns_2_2_1_Adder_1_U.ain_s1  <= _241_;
always @(posedge \sub_2ns_2ns_2_2_1_U2.top_sub_2ns_2ns_2_2_1_Adder_1_U.clk )
\sub_2ns_2ns_2_2_1_U2.top_sub_2ns_2ns_2_2_1_Adder_1_U.sum_s1  <= _244_;
always @(posedge \sub_2ns_2ns_2_2_1_U2.top_sub_2ns_2ns_2_2_1_Adder_1_U.clk )
\sub_2ns_2ns_2_2_1_U2.top_sub_2ns_2ns_2_2_1_Adder_1_U.carry_s1  <= _243_;
assign _242_ = \sub_2ns_2ns_2_2_1_U2.top_sub_2ns_2ns_2_2_1_Adder_1_U.ce  ? \sub_2ns_2ns_2_2_1_U2.top_sub_2ns_2ns_2_2_1_Adder_1_U.bin_s0 [1] : \sub_2ns_2ns_2_2_1_U2.top_sub_2ns_2ns_2_2_1_Adder_1_U.bin_s1 ;
assign _241_ = \sub_2ns_2ns_2_2_1_U2.top_sub_2ns_2ns_2_2_1_Adder_1_U.ce  ? \sub_2ns_2ns_2_2_1_U2.top_sub_2ns_2ns_2_2_1_Adder_1_U.a [1] : \sub_2ns_2ns_2_2_1_U2.top_sub_2ns_2ns_2_2_1_Adder_1_U.ain_s1 ;
assign _243_ = \sub_2ns_2ns_2_2_1_U2.top_sub_2ns_2ns_2_2_1_Adder_1_U.ce  ? \sub_2ns_2ns_2_2_1_U2.top_sub_2ns_2ns_2_2_1_Adder_1_U.facout_s1  : \sub_2ns_2ns_2_2_1_U2.top_sub_2ns_2ns_2_2_1_Adder_1_U.carry_s1 ;
assign _244_ = \sub_2ns_2ns_2_2_1_U2.top_sub_2ns_2ns_2_2_1_Adder_1_U.ce  ? \sub_2ns_2ns_2_2_1_U2.top_sub_2ns_2ns_2_2_1_Adder_1_U.fas_s1  : \sub_2ns_2ns_2_2_1_U2.top_sub_2ns_2ns_2_2_1_Adder_1_U.sum_s1 ;
assign _245_ = \sub_2ns_2ns_2_2_1_U2.top_sub_2ns_2ns_2_2_1_Adder_1_U.u1.a  + \sub_2ns_2ns_2_2_1_U2.top_sub_2ns_2ns_2_2_1_Adder_1_U.u1.b ;
assign { \sub_2ns_2ns_2_2_1_U2.top_sub_2ns_2ns_2_2_1_Adder_1_U.u1.cout , \sub_2ns_2ns_2_2_1_U2.top_sub_2ns_2ns_2_2_1_Adder_1_U.u1.s  } = _245_ + \sub_2ns_2ns_2_2_1_U2.top_sub_2ns_2ns_2_2_1_Adder_1_U.u1.cin ;
assign _246_ = \sub_2ns_2ns_2_2_1_U2.top_sub_2ns_2ns_2_2_1_Adder_1_U.u2.a  + \sub_2ns_2ns_2_2_1_U2.top_sub_2ns_2ns_2_2_1_Adder_1_U.u2.b ;
assign { \sub_2ns_2ns_2_2_1_U2.top_sub_2ns_2ns_2_2_1_Adder_1_U.u2.cout , \sub_2ns_2ns_2_2_1_U2.top_sub_2ns_2ns_2_2_1_Adder_1_U.u2.s  } = _246_ + \sub_2ns_2ns_2_2_1_U2.top_sub_2ns_2ns_2_2_1_Adder_1_U.u2.cin ;
assign \sub_2ns_2s_2_2_1_U10.top_sub_2ns_2s_2_2_1_Adder_7_U.bin_s0  = ~ \sub_2ns_2s_2_2_1_U10.top_sub_2ns_2s_2_2_1_Adder_7_U.b ;
always @(posedge \sub_2ns_2s_2_2_1_U10.top_sub_2ns_2s_2_2_1_Adder_7_U.clk )
\sub_2ns_2s_2_2_1_U10.top_sub_2ns_2s_2_2_1_Adder_7_U.bin_s1  <= _248_;
always @(posedge \sub_2ns_2s_2_2_1_U10.top_sub_2ns_2s_2_2_1_Adder_7_U.clk )
\sub_2ns_2s_2_2_1_U10.top_sub_2ns_2s_2_2_1_Adder_7_U.ain_s1  <= _247_;
always @(posedge \sub_2ns_2s_2_2_1_U10.top_sub_2ns_2s_2_2_1_Adder_7_U.clk )
\sub_2ns_2s_2_2_1_U10.top_sub_2ns_2s_2_2_1_Adder_7_U.sum_s1  <= _250_;
always @(posedge \sub_2ns_2s_2_2_1_U10.top_sub_2ns_2s_2_2_1_Adder_7_U.clk )
\sub_2ns_2s_2_2_1_U10.top_sub_2ns_2s_2_2_1_Adder_7_U.carry_s1  <= _249_;
assign _248_ = \sub_2ns_2s_2_2_1_U10.top_sub_2ns_2s_2_2_1_Adder_7_U.ce  ? \sub_2ns_2s_2_2_1_U10.top_sub_2ns_2s_2_2_1_Adder_7_U.bin_s0 [1] : \sub_2ns_2s_2_2_1_U10.top_sub_2ns_2s_2_2_1_Adder_7_U.bin_s1 ;
assign _247_ = \sub_2ns_2s_2_2_1_U10.top_sub_2ns_2s_2_2_1_Adder_7_U.ce  ? \sub_2ns_2s_2_2_1_U10.top_sub_2ns_2s_2_2_1_Adder_7_U.a [1] : \sub_2ns_2s_2_2_1_U10.top_sub_2ns_2s_2_2_1_Adder_7_U.ain_s1 ;
assign _249_ = \sub_2ns_2s_2_2_1_U10.top_sub_2ns_2s_2_2_1_Adder_7_U.ce  ? \sub_2ns_2s_2_2_1_U10.top_sub_2ns_2s_2_2_1_Adder_7_U.facout_s1  : \sub_2ns_2s_2_2_1_U10.top_sub_2ns_2s_2_2_1_Adder_7_U.carry_s1 ;
assign _250_ = \sub_2ns_2s_2_2_1_U10.top_sub_2ns_2s_2_2_1_Adder_7_U.ce  ? \sub_2ns_2s_2_2_1_U10.top_sub_2ns_2s_2_2_1_Adder_7_U.fas_s1  : \sub_2ns_2s_2_2_1_U10.top_sub_2ns_2s_2_2_1_Adder_7_U.sum_s1 ;
assign _251_ = \sub_2ns_2s_2_2_1_U10.top_sub_2ns_2s_2_2_1_Adder_7_U.u1.a  + \sub_2ns_2s_2_2_1_U10.top_sub_2ns_2s_2_2_1_Adder_7_U.u1.b ;
assign { \sub_2ns_2s_2_2_1_U10.top_sub_2ns_2s_2_2_1_Adder_7_U.u1.cout , \sub_2ns_2s_2_2_1_U10.top_sub_2ns_2s_2_2_1_Adder_7_U.u1.s  } = _251_ + \sub_2ns_2s_2_2_1_U10.top_sub_2ns_2s_2_2_1_Adder_7_U.u1.cin ;
assign _252_ = \sub_2ns_2s_2_2_1_U10.top_sub_2ns_2s_2_2_1_Adder_7_U.u2.a  + \sub_2ns_2s_2_2_1_U10.top_sub_2ns_2s_2_2_1_Adder_7_U.u2.b ;
assign { \sub_2ns_2s_2_2_1_U10.top_sub_2ns_2s_2_2_1_Adder_7_U.u2.cout , \sub_2ns_2s_2_2_1_U10.top_sub_2ns_2s_2_2_1_Adder_7_U.u2.s  } = _252_ + \sub_2ns_2s_2_2_1_U10.top_sub_2ns_2s_2_2_1_Adder_7_U.u2.cin ;
assign \sub_3ns_3s_3_2_1_U1.top_sub_3ns_3s_3_2_1_Adder_0_U.bin_s0  = ~ \sub_3ns_3s_3_2_1_U1.top_sub_3ns_3s_3_2_1_Adder_0_U.b ;
always @(posedge \sub_3ns_3s_3_2_1_U1.top_sub_3ns_3s_3_2_1_Adder_0_U.clk )
\sub_3ns_3s_3_2_1_U1.top_sub_3ns_3s_3_2_1_Adder_0_U.bin_s1  <= _254_;
always @(posedge \sub_3ns_3s_3_2_1_U1.top_sub_3ns_3s_3_2_1_Adder_0_U.clk )
\sub_3ns_3s_3_2_1_U1.top_sub_3ns_3s_3_2_1_Adder_0_U.ain_s1  <= _253_;
always @(posedge \sub_3ns_3s_3_2_1_U1.top_sub_3ns_3s_3_2_1_Adder_0_U.clk )
\sub_3ns_3s_3_2_1_U1.top_sub_3ns_3s_3_2_1_Adder_0_U.sum_s1  <= _256_;
always @(posedge \sub_3ns_3s_3_2_1_U1.top_sub_3ns_3s_3_2_1_Adder_0_U.clk )
\sub_3ns_3s_3_2_1_U1.top_sub_3ns_3s_3_2_1_Adder_0_U.carry_s1  <= _255_;
assign _254_ = \sub_3ns_3s_3_2_1_U1.top_sub_3ns_3s_3_2_1_Adder_0_U.ce  ? \sub_3ns_3s_3_2_1_U1.top_sub_3ns_3s_3_2_1_Adder_0_U.bin_s0 [2:1] : \sub_3ns_3s_3_2_1_U1.top_sub_3ns_3s_3_2_1_Adder_0_U.bin_s1 ;
assign _253_ = \sub_3ns_3s_3_2_1_U1.top_sub_3ns_3s_3_2_1_Adder_0_U.ce  ? \sub_3ns_3s_3_2_1_U1.top_sub_3ns_3s_3_2_1_Adder_0_U.a [2:1] : \sub_3ns_3s_3_2_1_U1.top_sub_3ns_3s_3_2_1_Adder_0_U.ain_s1 ;
assign _255_ = \sub_3ns_3s_3_2_1_U1.top_sub_3ns_3s_3_2_1_Adder_0_U.ce  ? \sub_3ns_3s_3_2_1_U1.top_sub_3ns_3s_3_2_1_Adder_0_U.facout_s1  : \sub_3ns_3s_3_2_1_U1.top_sub_3ns_3s_3_2_1_Adder_0_U.carry_s1 ;
assign _256_ = \sub_3ns_3s_3_2_1_U1.top_sub_3ns_3s_3_2_1_Adder_0_U.ce  ? \sub_3ns_3s_3_2_1_U1.top_sub_3ns_3s_3_2_1_Adder_0_U.fas_s1  : \sub_3ns_3s_3_2_1_U1.top_sub_3ns_3s_3_2_1_Adder_0_U.sum_s1 ;
assign _257_ = \sub_3ns_3s_3_2_1_U1.top_sub_3ns_3s_3_2_1_Adder_0_U.u1.a  + \sub_3ns_3s_3_2_1_U1.top_sub_3ns_3s_3_2_1_Adder_0_U.u1.b ;
assign { \sub_3ns_3s_3_2_1_U1.top_sub_3ns_3s_3_2_1_Adder_0_U.u1.cout , \sub_3ns_3s_3_2_1_U1.top_sub_3ns_3s_3_2_1_Adder_0_U.u1.s  } = _257_ + \sub_3ns_3s_3_2_1_U1.top_sub_3ns_3s_3_2_1_Adder_0_U.u1.cin ;
assign _258_ = \sub_3ns_3s_3_2_1_U1.top_sub_3ns_3s_3_2_1_Adder_0_U.u2.a  + \sub_3ns_3s_3_2_1_U1.top_sub_3ns_3s_3_2_1_Adder_0_U.u2.b ;
assign { \sub_3ns_3s_3_2_1_U1.top_sub_3ns_3s_3_2_1_Adder_0_U.u2.cout , \sub_3ns_3s_3_2_1_U1.top_sub_3ns_3s_3_2_1_Adder_0_U.u2.s  } = _258_ + \sub_3ns_3s_3_2_1_U1.top_sub_3ns_3s_3_2_1_Adder_0_U.u2.cin ;
assign _259_ = $signed({ op_4, 3'h0 }) > $signed(op_8_V_reg_1018);
assign _260_ = | p_Result_s_reg_975;
assign _261_ = | trunc_ln851_3_reg_1152;
assign _262_ = | trunc_ln851_2_reg_1320;
assign _263_ = | op_15[1:0];
assign _264_ = | op_17[2:0];
assign _265_ = | trunc_ln718_reg_1057;
assign or_ln384_fu_359_p2 = p_Result_7_reg_964 | overflow_reg_1007;
assign or_ln410_fu_506_p2 = xor_ln410_fu_500_p2 | r_reg_1072;
assign or_ln785_fu_337_p2 = p_Result_8_reg_997 | icmp_ln768_reg_1002;
assign ret_V_18_fu_412_p2 = { op_3, 3'h0 } | op_1;
assign ret_V_22_fu_763_p2 = op_8_V_reg_1018 | op_11;
always @(posedge ap_clk)
p_Val2_2_reg_992[2:0] <= 3'h0;
always @(posedge ap_clk)
sub_ln69_reg_1202 <= _059_;
always @(posedge ap_clk)
sub_ln1357_reg_1013 <= _058_;
always @(posedge ap_clk)
sub_ln1118_reg_1067 <= _057_;
always @(posedge ap_clk)
shl_ln1358_reg_1114 <= _056_;
always @(posedge ap_clk)
select_ln1347_reg_929 <= _049_;
always @(posedge ap_clk)
select_ln13_reg_934 <= _050_;
always @(posedge ap_clk)
ret_V_28_reg_1392 <= _043_;
always @(posedge ap_clk)
ret_V_27_reg_1382 <= _042_;
always @(posedge ap_clk)
ret_V_26_reg_1365 <= _041_;
always @(posedge ap_clk)
ret_V_31_cast_reg_1370 <= _045_;
always @(posedge ap_clk)
ret_V_25_reg_1335 <= _040_;
always @(posedge ap_clk)
select_ln69_1_reg_1340 <= _052_;
always @(posedge ap_clk)
ret_V_24_reg_1302 <= _039_;
always @(posedge ap_clk)
ret_V_29_cast_reg_1307 <= _044_;
always @(posedge ap_clk)
ret_V_22_reg_1314 <= _037_;
always @(posedge ap_clk)
trunc_ln851_2_reg_1320 <= _065_;
always @(posedge ap_clk)
ret_V_18_reg_1047 <= _033_;
always @(posedge ap_clk)
tmp_reg_1052 <= _061_;
always @(posedge ap_clk)
trunc_ln718_reg_1057 <= _062_;
always @(posedge ap_clk)
r_reg_1072 <= _032_;
always @(posedge ap_clk)
ret_V_19_reg_1077 <= _034_;
always @(posedge ap_clk)
ret_V_reg_1082 <= _048_;
always @(posedge ap_clk)
trunc_ln851_reg_1089 <= _067_;
always @(posedge ap_clk)
r_V_reg_1094 <= _031_;
always @(posedge ap_clk)
tmp_2_reg_1099 <= _060_;
always @(posedge ap_clk)
trunc_ln851_1_reg_1104 <= _064_;
always @(posedge ap_clk)
overflow_reg_1007 <= _024_;
always @(posedge ap_clk)
op_8_V_reg_1018 <= _023_;
always @(posedge ap_clk)
ush_reg_1026 <= _068_;
always @(posedge ap_clk)
op_28_V_reg_1345 <= _020_;
always @(posedge ap_clk)
op_26_V_reg_1282 <= _019_;
always @(posedge ap_clk)
p_Result_7_reg_964 <= _025_;
always @(posedge ap_clk)
trunc_ln728_reg_970 <= _063_;
always @(posedge ap_clk)
p_Result_s_reg_975 <= _027_;
always @(posedge ap_clk)
r_2_reg_980 <= _029_;
always @(posedge ap_clk)
isNeg_reg_986 <= _018_;
always @(posedge ap_clk)
icmp_ln851_3_reg_1360 <= _016_;
always @(posedge ap_clk)
icmp_ln851_2_reg_1297 <= _015_;
always @(posedge ap_clk)
icmp_ln850_reg_1325 <= _013_;
always @(posedge ap_clk)
ret_V_3_reg_1162 <= _046_;
always @(posedge ap_clk)
ret_V_5_reg_1167 <= _047_;
always @(posedge ap_clk)
icmp_ln850_1_reg_1172 <= _012_;
always @(posedge ap_clk)
p_Val2_2_reg_992[3] <= _028_;
always @(posedge ap_clk)
p_Result_8_reg_997 <= _026_;
always @(posedge ap_clk)
icmp_ln768_reg_1002 <= _011_;
always @(posedge ap_clk)
op_6_V_reg_1177 <= _021_;
always @(posedge ap_clk)
ret_V_20_reg_1182 <= _035_;
always @(posedge ap_clk)
ret_V_21_reg_1187 <= _036_;
always @(posedge ap_clk)
icmp_ln1494_reg_1192 <= _010_;
always @(posedge ap_clk)
select_ln69_reg_1197 <= _053_;
always @(posedge ap_clk)
conv_i389_reg_954 <= _009_;
always @(posedge ap_clk)
select_ln1497_reg_959 <= _051_;
always @(posedge ap_clk)
ashr_ln1297_reg_1109 <= _008_;
always @(posedge ap_clk)
select_ln708_reg_1119 <= _054_;
always @(posedge ap_clk)
and_ln410_reg_1124 <= _006_;
always @(posedge ap_clk)
icmp_ln851_reg_1129 <= _017_;
always @(posedge ap_clk)
sext_ln850_reg_1134 <= _055_;
always @(posedge ap_clk)
icmp_ln851_1_reg_1141 <= _014_;
always @(posedge ap_clk)
r_V_1_reg_1146 <= _030_;
always @(posedge ap_clk)
trunc_ln851_3_reg_1152 <= _066_;
always @(posedge ap_clk)
op_7_V_reg_1232 <= _022_;
always @(posedge ap_clk)
ret_V_23_reg_1237 <= _038_;
always @(posedge ap_clk)
add_ln69_reg_1242 <= _005_;
always @(posedge ap_clk)
add_ln69_2_reg_1247 <= _003_;
always @(posedge ap_clk)
add_ln69_1_reg_1267 <= _002_;
always @(posedge ap_clk)
add_ln69_3_reg_1272 <= _004_;
always @(posedge ap_clk)
add_ln691_reg_1330 <= _001_;
always @(posedge ap_clk)
add_ln691_1_reg_1377 <= _000_;
always @(posedge ap_clk)
ap_CS_fsm <= _007_;
assign _069_ = _078_ ? 2'h2 : 2'h1;
assign _266_ = ap_CS_fsm == 1'h1;
function [37:0] _739_;
input [37:0] a;
input [1443:0] b;
input [37:0] s;
case (s)
38'b00000000000000000000000000000000000001:
_739_ = b[37:0];
38'b00000000000000000000000000000000000010:
_739_ = b[75:38];
38'b00000000000000000000000000000000000100:
_739_ = b[113:76];
38'b00000000000000000000000000000000001000:
_739_ = b[151:114];
38'b00000000000000000000000000000000010000:
_739_ = b[189:152];
38'b00000000000000000000000000000000100000:
_739_ = b[227:190];
38'b00000000000000000000000000000001000000:
_739_ = b[265:228];
38'b00000000000000000000000000000010000000:
_739_ = b[303:266];
38'b00000000000000000000000000000100000000:
_739_ = b[341:304];
38'b00000000000000000000000000001000000000:
_739_ = b[379:342];
38'b00000000000000000000000000010000000000:
_739_ = b[417:380];
38'b00000000000000000000000000100000000000:
_739_ = b[455:418];
38'b00000000000000000000000001000000000000:
_739_ = b[493:456];
38'b00000000000000000000000010000000000000:
_739_ = b[531:494];
38'b00000000000000000000000100000000000000:
_739_ = b[569:532];
38'b00000000000000000000001000000000000000:
_739_ = b[607:570];
38'b00000000000000000000010000000000000000:
_739_ = b[645:608];
38'b00000000000000000000100000000000000000:
_739_ = b[683:646];
38'b00000000000000000001000000000000000000:
_739_ = b[721:684];
38'b00000000000000000010000000000000000000:
_739_ = b[759:722];
38'b00000000000000000100000000000000000000:
_739_ = b[797:760];
38'b00000000000000001000000000000000000000:
_739_ = b[835:798];
38'b00000000000000010000000000000000000000:
_739_ = b[873:836];
38'b00000000000000100000000000000000000000:
_739_ = b[911:874];
38'b00000000000001000000000000000000000000:
_739_ = b[949:912];
38'b00000000000010000000000000000000000000:
_739_ = b[987:950];
38'b00000000000100000000000000000000000000:
_739_ = b[1025:988];
38'b00000000001000000000000000000000000000:
_739_ = b[1063:1026];
38'b00000000010000000000000000000000000000:
_739_ = b[1101:1064];
38'b00000000100000000000000000000000000000:
_739_ = b[1139:1102];
38'b00000001000000000000000000000000000000:
_739_ = b[1177:1140];
38'b00000010000000000000000000000000000000:
_739_ = b[1215:1178];
38'b00000100000000000000000000000000000000:
_739_ = b[1253:1216];
38'b00001000000000000000000000000000000000:
_739_ = b[1291:1254];
38'b00010000000000000000000000000000000000:
_739_ = b[1329:1292];
38'b00100000000000000000000000000000000000:
_739_ = b[1367:1330];
38'b01000000000000000000000000000000000000:
_739_ = b[1405:1368];
38'b10000000000000000000000000000000000000:
_739_ = b[1443:1406];
38'b00000000000000000000000000000000000000:
_739_ = a;
default:
_739_ = 38'bx;
endcase
endfunction
assign ap_NS_fsm = _739_(38'hxxxxxxxxxx, { 36'h000000000, _069_, 1406'h0000000004000000002000000001000000000800000000400000000200000000100000000080000000040000000020000000010000000008000000004000000002000000001000000000800000000400000000200000000100000000080000000040000000020000000010000000008000000004000000002000000001000000000800000000400000000200000000100000000080000000040000000020000000010000000008000000000000000001 }, { _266_, _303_, _302_, _301_, _300_, _299_, _298_, _297_, _296_, _295_, _294_, _293_, _292_, _291_, _290_, _289_, _288_, _287_, _286_, _285_, _284_, _283_, _282_, _281_, _280_, _279_, _278_, _277_, _276_, _275_, _274_, _273_, _272_, _271_, _270_, _269_, _268_, _267_ });
assign _267_ = ap_CS_fsm == 38'h2000000000;
assign _268_ = ap_CS_fsm == 37'h1000000000;
assign _269_ = ap_CS_fsm == 36'h800000000;
assign _270_ = ap_CS_fsm == 35'h400000000;
assign _271_ = ap_CS_fsm == 34'h200000000;
assign _272_ = ap_CS_fsm == 33'h100000000;
assign _273_ = ap_CS_fsm == 32'd2147483648;
assign _274_ = ap_CS_fsm == 31'h40000000;
assign _275_ = ap_CS_fsm == 30'h20000000;
assign _276_ = ap_CS_fsm == 29'h10000000;
assign _277_ = ap_CS_fsm == 28'h8000000;
assign _278_ = ap_CS_fsm == 27'h4000000;
assign _279_ = ap_CS_fsm == 26'h2000000;
assign _280_ = ap_CS_fsm == 25'h1000000;
assign _281_ = ap_CS_fsm == 24'h800000;
assign _282_ = ap_CS_fsm == 23'h400000;
assign _283_ = ap_CS_fsm == 22'h200000;
assign _284_ = ap_CS_fsm == 21'h100000;
assign _285_ = ap_CS_fsm == 20'h80000;
assign _286_ = ap_CS_fsm == 19'h40000;
assign _287_ = ap_CS_fsm == 18'h20000;
assign _288_ = ap_CS_fsm == 17'h10000;
assign _289_ = ap_CS_fsm == 16'h8000;
assign _290_ = ap_CS_fsm == 15'h4000;
assign _291_ = ap_CS_fsm == 14'h2000;
assign _292_ = ap_CS_fsm == 13'h1000;
assign _293_ = ap_CS_fsm == 12'h800;
assign _294_ = ap_CS_fsm == 11'h400;
assign _295_ = ap_CS_fsm == 10'h200;
assign _296_ = ap_CS_fsm == 9'h100;
assign _297_ = ap_CS_fsm == 8'h80;
assign _298_ = ap_CS_fsm == 7'h40;
assign _299_ = ap_CS_fsm == 6'h20;
assign _300_ = ap_CS_fsm == 5'h10;
assign _301_ = ap_CS_fsm == 4'h8;
assign _302_ = ap_CS_fsm == 3'h4;
assign _303_ = ap_CS_fsm == 2'h2;
assign op_31_ap_vld = ap_CS_fsm[37] ? 1'h1 : 1'h0;
assign ap_idle = _077_ ? 1'h1 : 1'h0;
assign _059_ = _076_ ? grp_fu_563_p2 : sub_ln69_reg_1202;
assign _058_ = _075_ ? grp_fu_332_p2 : sub_ln1357_reg_1013;
assign _057_ = _074_ ? grp_fu_399_p2 : sub_ln1118_reg_1067;
assign _056_ = _073_ ? grp_fu_383_p2 : shl_ln1358_reg_1114;
assign _050_ = ap_CS_fsm[0] ? select_ln13_fu_205_p3 : select_ln13_reg_934;
assign _049_ = ap_CS_fsm[0] ? select_ln1347_fu_197_p3 : select_ln1347_reg_929;
assign _043_ = ap_CS_fsm[35] ? grp_fu_907_p2 : ret_V_28_reg_1392;
assign _042_ = ap_CS_fsm[33] ? ret_V_27_fu_896_p3 : ret_V_27_reg_1382;
assign _045_ = ap_CS_fsm[30] ? grp_fu_853_p2[34:3] : ret_V_31_cast_reg_1370;
assign _041_ = ap_CS_fsm[30] ? grp_fu_853_p2 : ret_V_26_reg_1365;
assign _052_ = ap_CS_fsm[26] ? select_ln69_1_fu_826_p3 : select_ln69_1_reg_1340;
assign _040_ = ap_CS_fsm[26] ? ret_V_25_fu_819_p3 : ret_V_25_reg_1335;
assign _044_ = ap_CS_fsm[23] ? grp_fu_737_p2[33:2] : ret_V_29_cast_reg_1307;
assign _039_ = ap_CS_fsm[23] ? grp_fu_737_p2 : ret_V_24_reg_1302;
assign _065_ = ap_CS_fsm[24] ? ret_V_22_fu_763_p2[2:0] : trunc_ln851_2_reg_1320;
assign _037_ = ap_CS_fsm[24] ? ret_V_22_fu_763_p2 : ret_V_22_reg_1314;
assign _062_ = ap_CS_fsm[11] ? ret_V_18_fu_412_p2[1:0] : trunc_ln718_reg_1057;
assign _061_ = ap_CS_fsm[11] ? ret_V_18_fu_412_p2[3] : tmp_reg_1052;
assign _033_ = ap_CS_fsm[11] ? ret_V_18_fu_412_p2 : ret_V_18_reg_1047;
assign _064_ = ap_CS_fsm[12] ? r_V_fu_459_p3[23:0] : trunc_ln851_1_reg_1104;
assign _060_ = ap_CS_fsm[12] ? r_V_fu_459_p3[26:24] : tmp_2_reg_1099;
assign _031_ = ap_CS_fsm[12] ? r_V_fu_459_p3 : r_V_reg_1094;
assign _067_ = ap_CS_fsm[12] ? grp_fu_434_p2[2:0] : trunc_ln851_reg_1089;
assign _048_ = ap_CS_fsm[12] ? grp_fu_434_p2[8:3] : ret_V_reg_1082;
assign _034_ = ap_CS_fsm[12] ? grp_fu_434_p2 : ret_V_19_reg_1077;
assign _032_ = ap_CS_fsm[12] ? r_fu_440_p2 : r_reg_1072;
assign _024_ = ap_CS_fsm[4] ? overflow_fu_346_p2 : overflow_reg_1007;
assign _068_ = ap_CS_fsm[5] ? ush_fu_370_p3 : ush_reg_1026;
assign _023_ = ap_CS_fsm[5] ? op_8_V_fu_363_p3 : op_8_V_reg_1018;
assign _020_ = ap_CS_fsm[28] ? grp_fu_834_p2 : op_28_V_reg_1345;
assign _019_ = ap_CS_fsm[21] ? grp_fu_717_p2 : op_26_V_reg_1282;
assign _018_ = ap_CS_fsm[2] ? r_2_fu_302_p1[1] : isNeg_reg_986;
assign _029_ = ap_CS_fsm[2] ? r_2_fu_302_p1 : r_2_reg_980;
assign _027_ = ap_CS_fsm[2] ? grp_fu_217_p2[2:1] : p_Result_s_reg_975;
assign _063_ = ap_CS_fsm[2] ? grp_fu_217_p2[0] : trunc_ln728_reg_970;
assign _025_ = ap_CS_fsm[2] ? grp_fu_217_p2[2] : p_Result_7_reg_964;
assign _016_ = ap_CS_fsm[29] ? icmp_ln851_3_fu_863_p2 : icmp_ln851_3_reg_1360;
assign _015_ = ap_CS_fsm[22] ? icmp_ln851_2_fu_747_p2 : icmp_ln851_2_reg_1297;
assign _013_ = ap_CS_fsm[25] ? icmp_ln850_fu_777_p2 : icmp_ln850_reg_1325;
assign _012_ = ap_CS_fsm[14] ? icmp_ln850_1_fu_558_p2 : icmp_ln850_1_reg_1172;
assign _047_ = ap_CS_fsm[14] ? grp_fu_535_p2 : ret_V_5_reg_1167;
assign _046_ = ap_CS_fsm[14] ? grp_fu_522_p2 : ret_V_3_reg_1162;
assign _011_ = ap_CS_fsm[3] ? icmp_ln768_fu_327_p2 : icmp_ln768_reg_1002;
assign _026_ = ap_CS_fsm[3] ? p_Result_8_fu_321_p2 : p_Result_8_reg_997;
assign _028_ = ap_CS_fsm[3] ? trunc_ln728_reg_970 : p_Val2_2_reg_992[3];
assign _053_ = ap_CS_fsm[15] ? select_ln69_fu_647_p3 : select_ln69_reg_1197;
assign _010_ = ap_CS_fsm[15] ? icmp_ln1494_fu_616_p2 : icmp_ln1494_reg_1192;
assign _036_ = ap_CS_fsm[15] ? ret_V_21_fu_599_p3 : ret_V_21_reg_1187;
assign _035_ = ap_CS_fsm[15] ? ret_V_20_fu_580_p3 : ret_V_20_reg_1182;
assign _021_ = ap_CS_fsm[15] ? grp_fu_553_p2 : op_6_V_reg_1177;
assign _051_ = ap_CS_fsm[1] ? select_ln1497_fu_232_p3 : select_ln1497_reg_959;
assign _009_ = ap_CS_fsm[1] ? { op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4 } : conv_i389_reg_954;
assign _008_ = _072_ ? grp_fu_378_p2 : ashr_ln1297_reg_1109;
assign _066_ = ap_CS_fsm[13] ? r_V_1_fu_541_p3[2:0] : trunc_ln851_3_reg_1152;
assign _030_ = ap_CS_fsm[13] ? r_V_1_fu_541_p3 : r_V_1_reg_1146;
assign _014_ = ap_CS_fsm[13] ? icmp_ln851_1_fu_530_p2 : icmp_ln851_1_reg_1141;
assign _055_ = ap_CS_fsm[13] ? { tmp_2_reg_1099[2], tmp_2_reg_1099 } : sext_ln850_reg_1134;
assign _017_ = ap_CS_fsm[13] ? icmp_ln851_fu_517_p2 : icmp_ln851_reg_1129;
assign _006_ = ap_CS_fsm[13] ? and_ln410_fu_511_p2 : and_ln410_reg_1124;
assign _054_ = ap_CS_fsm[13] ? select_ln708_fu_479_p3 : select_ln708_reg_1119;
assign _003_ = ap_CS_fsm[17] ? grp_fu_683_p2 : add_ln69_2_reg_1247;
assign _005_ = ap_CS_fsm[17] ? grp_fu_677_p2 : add_ln69_reg_1242;
assign _038_ = ap_CS_fsm[17] ? grp_fu_661_p2 : ret_V_23_reg_1237;
assign _022_ = ap_CS_fsm[17] ? op_7_V_fu_688_p3 : op_7_V_reg_1232;
assign _004_ = ap_CS_fsm[19] ? grp_fu_708_p2 : add_ln69_3_reg_1272;
assign _002_ = ap_CS_fsm[19] ? grp_fu_700_p2 : add_ln69_1_reg_1267;
assign _001_ = _071_ ? grp_fu_772_p2 : add_ln691_reg_1330;
assign _000_ = _070_ ? grp_fu_879_p2 : add_ln691_1_reg_1377;
assign _007_ = ap_rst ? 38'h0000000001 : ap_NS_fsm;
assign icmp_ln1494_fu_616_p2 = _259_ ? 1'h1 : 1'h0;
assign icmp_ln768_fu_327_p2 = _260_ ? 1'h1 : 1'h0;
assign icmp_ln850_1_fu_558_p2 = _261_ ? 1'h1 : 1'h0;
assign icmp_ln850_fu_777_p2 = _262_ ? 1'h1 : 1'h0;
assign icmp_ln851_1_fu_530_p2 = _081_ ? 1'h1 : 1'h0;
assign icmp_ln851_2_fu_747_p2 = _263_ ? 1'h1 : 1'h0;
assign icmp_ln851_3_fu_863_p2 = _264_ ? 1'h1 : 1'h0;
assign icmp_ln851_fu_517_p2 = _082_ ? 1'h1 : 1'h0;
assign op_7_V_fu_688_p3 = op_3 ? sub_ln69_reg_1202 : 2'h0;
assign op_8_V_fu_363_p3 = or_ln384_fu_359_p2 ? select_ln384_fu_352_p3 : p_Val2_2_reg_992;
assign p_Result_8_fu_321_p2 = trunc_ln728_reg_970 ? 1'h1 : 1'h0;
assign r_V_1_fu_541_p3 = isNeg_reg_986 ? ashr_ln1297_reg_1109 : shl_ln1358_reg_1114;
assign r_V_fu_459_p3 = op_3 ? sub_ln1118_reg_1067 : 27'h0000000;
assign r_fu_440_p2 = _265_ ? 1'h1 : 1'h0;
assign ret_V_20_fu_580_p3 = ret_V_19_reg_1077[8] ? select_ln850_fu_575_p3 : ret_V_reg_1082;
assign ret_V_21_fu_599_p3 = r_V_reg_1094[26] ? select_ln850_2_fu_594_p3 : sext_ln850_reg_1134;
assign ret_V_25_fu_819_p3 = ret_V_24_reg_1302[34] ? select_ln850_3_fu_814_p3 : ret_V_29_cast_reg_1307;
assign ret_V_27_fu_896_p3 = ret_V_26_reg_1365[35] ? select_ln850_4_fu_891_p3 : ret_V_31_cast_reg_1370;
assign select_ln1347_fu_197_p3 = op_3 ? 3'h7 : 3'h0;
assign select_ln13_fu_205_p3 = op_3 ? 1'h1 : 1'h0;
assign select_ln1497_1_fu_275_p3 = op_4[1] ? 2'h3 : 2'h0;
assign select_ln1497_2_fu_288_p3 = select_ln13_reg_934 ? select_ln1497_1_fu_275_p3 : conv_i389_reg_954[1:0];
assign r_2_fu_302_p1 = select_ln835_fu_261_p3 ? select_ln1497_2_fu_288_p3 : select_ln1497_reg_959[1:0];
assign select_ln1497_fu_232_p3 = select_ln13_reg_934 ? { 1'h0, op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1] } : { op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4 };
assign select_ln384_fu_352_p3 = overflow_reg_1007 ? 4'h7 : 4'h9;
assign select_ln69_1_fu_826_p3 = ret_V_9_fu_801_p2 ? 32'd4294967295 : 32'd0;
assign select_ln69_fu_647_p3 = ret_V_12_fu_641_p2 ? 2'h3 : 2'h0;
assign select_ln708_fu_479_p3 = tmp_reg_1052 ? 2'h3 : 2'h0;
assign select_ln835_fu_261_p3 = select_ln13_reg_934 ? 1'h1 : 1'h0;
assign select_ln850_2_fu_594_p3 = icmp_ln851_1_reg_1141 ? sext_ln850_reg_1134 : ret_V_5_reg_1167;
assign select_ln850_3_fu_814_p3 = icmp_ln851_2_reg_1297 ? add_ln691_reg_1330 : ret_V_29_cast_reg_1307;
assign select_ln850_4_fu_891_p3 = icmp_ln851_3_reg_1360 ? add_ln691_1_reg_1377 : ret_V_31_cast_reg_1370;
assign select_ln850_fu_575_p3 = icmp_ln851_reg_1129 ? ret_V_reg_1082 : ret_V_3_reg_1162;
assign ush_fu_370_p3 = isNeg_reg_986 ? sub_ln1357_reg_1013 : r_2_reg_980;
assign ret_V_12_fu_641_p2 = r_V_1_reg_1146[3] ^ and_ln850_1_fu_636_p2;
assign ret_V_9_fu_801_p2 = ret_V_22_reg_1314[3] ^ and_ln850_fu_796_p2;
assign ap_CS_fsm_state1 = ap_CS_fsm[0];
assign ap_CS_fsm_state11 = ap_CS_fsm[10];
assign ap_CS_fsm_state12 = ap_CS_fsm[11];
assign ap_CS_fsm_state13 = ap_CS_fsm[12];
assign ap_CS_fsm_state14 = ap_CS_fsm[13];
assign ap_CS_fsm_state15 = ap_CS_fsm[14];
assign ap_CS_fsm_state16 = ap_CS_fsm[15];
assign ap_CS_fsm_state17 = ap_CS_fsm[16];
assign ap_CS_fsm_state18 = ap_CS_fsm[17];
assign ap_CS_fsm_state19 = ap_CS_fsm[18];
assign ap_CS_fsm_state2 = ap_CS_fsm[1];
assign ap_CS_fsm_state20 = ap_CS_fsm[19];
assign ap_CS_fsm_state21 = ap_CS_fsm[20];
assign ap_CS_fsm_state22 = ap_CS_fsm[21];
assign ap_CS_fsm_state23 = ap_CS_fsm[22];
assign ap_CS_fsm_state24 = ap_CS_fsm[23];
assign ap_CS_fsm_state25 = ap_CS_fsm[24];
assign ap_CS_fsm_state26 = ap_CS_fsm[25];
assign ap_CS_fsm_state27 = ap_CS_fsm[26];
assign ap_CS_fsm_state28 = ap_CS_fsm[27];
assign ap_CS_fsm_state29 = ap_CS_fsm[28];
assign ap_CS_fsm_state3 = ap_CS_fsm[2];
assign ap_CS_fsm_state30 = ap_CS_fsm[29];
assign ap_CS_fsm_state31 = ap_CS_fsm[30];
assign ap_CS_fsm_state32 = ap_CS_fsm[31];
assign ap_CS_fsm_state33 = ap_CS_fsm[32];
assign ap_CS_fsm_state34 = ap_CS_fsm[33];
assign ap_CS_fsm_state35 = ap_CS_fsm[34];
assign ap_CS_fsm_state36 = ap_CS_fsm[35];
assign ap_CS_fsm_state37 = ap_CS_fsm[36];
assign ap_CS_fsm_state38 = ap_CS_fsm[37];
assign ap_CS_fsm_state4 = ap_CS_fsm[3];
assign ap_CS_fsm_state5 = ap_CS_fsm[4];
assign ap_CS_fsm_state6 = ap_CS_fsm[5];
assign ap_CS_fsm_state7 = ap_CS_fsm[6];
assign ap_done = op_31_ap_vld;
assign ap_ready = op_31_ap_vld;
assign ashr_ln1497_1_fu_283_p2 = conv_i389_reg_954;
assign conv_i389_fu_222_p0 = op_4;
assign conv_i389_fu_222_p1 = { op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4 };
assign grp_fu_217_p1 = { op_4[1], op_4 };
assign grp_fu_399_p1 = { op_4[1], op_4, 24'h000000 };
assign grp_fu_434_p0 = { op_0[7], op_0 };
assign grp_fu_535_p0 = { tmp_2_reg_1099[2], tmp_2_reg_1099 };
assign grp_fu_553_p0 = { 1'h0, and_ln410_reg_1124 };
assign grp_fu_661_p0 = { ret_V_20_reg_1182[5], ret_V_20_reg_1182 };
assign grp_fu_661_p1 = { op_6_V_reg_1177[1], op_6_V_reg_1177[1], op_6_V_reg_1177[1], op_6_V_reg_1177[1], op_6_V_reg_1177[1], op_6_V_reg_1177 };
assign grp_fu_677_p0 = { ret_V_21_reg_1187[3], ret_V_21_reg_1187[3], ret_V_21_reg_1187 };
assign grp_fu_677_p1 = { 2'h0, op_12 };
assign grp_fu_683_p1 = { 1'h0, icmp_ln1494_reg_1192 };
assign grp_fu_700_p0 = { add_ln69_reg_1242[5], add_ln69_reg_1242 };
assign grp_fu_708_p0 = { add_ln69_2_reg_1247[1], add_ln69_2_reg_1247 };
assign grp_fu_708_p1 = { op_7_V_reg_1232[1], op_7_V_reg_1232 };
assign grp_fu_717_p0 = { add_ln69_3_reg_1272[2], add_ln69_3_reg_1272[2], add_ln69_3_reg_1272[2], add_ln69_3_reg_1272[2], add_ln69_3_reg_1272 };
assign grp_fu_737_p0 = { op_26_V_reg_1282[6], op_26_V_reg_1282[6], op_26_V_reg_1282[6], op_26_V_reg_1282[6], op_26_V_reg_1282[6], op_26_V_reg_1282[6], op_26_V_reg_1282[6], op_26_V_reg_1282[6], op_26_V_reg_1282[6], op_26_V_reg_1282[6], op_26_V_reg_1282[6], op_26_V_reg_1282[6], op_26_V_reg_1282[6], op_26_V_reg_1282[6], op_26_V_reg_1282[6], op_26_V_reg_1282[6], op_26_V_reg_1282[6], op_26_V_reg_1282[6], op_26_V_reg_1282[6], op_26_V_reg_1282[6], op_26_V_reg_1282[6], op_26_V_reg_1282[6], op_26_V_reg_1282[6], op_26_V_reg_1282[6], op_26_V_reg_1282[6], op_26_V_reg_1282[6], op_26_V_reg_1282, 2'h0 };
assign grp_fu_737_p1 = { op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15 };
assign grp_fu_853_p0 = { op_28_V_reg_1345[31], op_28_V_reg_1345, 3'h0 };
assign grp_fu_853_p1 = { op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17 };
assign grp_fu_907_p1 = { op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18 };
assign grp_fu_916_p1 = { op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19 };
assign op_31 = grp_fu_916_p2;
assign op_3_read_read_fu_130_p2 = op_3;
assign op_7_V_fu_688_p0 = op_3;
assign p_Result_1_fu_587_p3 = r_V_reg_1094[26];
assign p_Result_2_fu_789_p3 = ret_V_22_reg_1314[3];
assign p_Result_3_fu_629_p3 = r_V_1_reg_1146[3];
assign p_Result_4_fu_807_p3 = ret_V_24_reg_1302[34];
assign p_Result_5_fu_884_p3 = ret_V_26_reg_1365[35];
assign p_Result_6_fu_486_p3 = op_1[2];
assign p_Result_s_14_fu_568_p3 = ret_V_19_reg_1077[8];
assign p_Val2_2_fu_314_p3 = { trunc_ln728_reg_970, 3'h0 };
assign r_V_fu_459_p0 = op_3;
assign ret_V_11_fu_622_p3 = r_V_1_reg_1146[3];
assign ret_V_8_fu_782_p3 = ret_V_22_reg_1314[3];
assign rhs_4_fu_842_p3 = { op_28_V_reg_1345, 3'h0 };
assign rhs_fu_405_p1 = op_3;
assign rhs_fu_405_p3 = { op_3, 3'h0 };
assign select_ln1347_fu_197_p0 = op_3;
assign select_ln13_fu_205_p0 = op_3;
assign select_ln1497_3_fu_295_p3 = { 30'hxxxxxxxx, r_2_fu_302_p1 };
assign sext_ln1347_fu_213_p0 = op_4;
assign sext_ln1494_fu_613_p1 = { op_8_V_reg_1018[3], op_8_V_reg_1018 };
assign sext_ln703_1_fu_722_p0 = op_15;
assign sext_ln703_2_fu_838_p0 = op_17;
assign sext_ln850_fu_527_p1 = { tmp_2_reg_1099[2], tmp_2_reg_1099 };
assign shl_ln1497_1_fu_226_p2 = { op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1] };
assign shl_ln1_fu_606_p1 = op_4;
assign shl_ln1_fu_606_p3 = { op_4, 3'h0 };
assign shl_ln_fu_388_p1 = op_4;
assign shl_ln_fu_388_p3 = { op_4, 24'h000000 };
assign tmp_14_fu_726_p3 = { op_26_V_reg_1282, 2'h0 };
assign tmp_3_fu_493_p3 = ret_V_18_reg_1047[3];
assign tmp_7_fu_268_p1 = op_4;
assign tmp_7_fu_268_p3 = op_4[1];
assign trunc_ln718_fu_426_p1 = ret_V_18_fu_412_p2[1:0];
assign trunc_ln728_fu_247_p1 = grp_fu_217_p2[0];
assign trunc_ln851_1_fu_475_p1 = r_V_fu_459_p3[23:0];
assign trunc_ln851_2_fu_768_p1 = ret_V_22_fu_763_p2[2:0];
assign trunc_ln851_3_fu_546_p1 = r_V_1_fu_541_p3[2:0];
assign trunc_ln851_4_fu_743_p0 = op_15;
assign trunc_ln851_4_fu_743_p1 = op_15[1:0];
assign trunc_ln851_5_fu_859_p0 = op_17;
assign trunc_ln851_5_fu_859_p1 = op_17[2:0];
assign trunc_ln851_fu_455_p1 = grp_fu_434_p2[2:0];
assign zext_ln1357_fu_375_p1 = { 2'h0, ush_reg_1026 };
assign \sub_3ns_3s_3_2_1_U1.top_sub_3ns_3s_3_2_1_Adder_0_U.ain_s0  = \sub_3ns_3s_3_2_1_U1.top_sub_3ns_3s_3_2_1_Adder_0_U.a ;
assign \sub_3ns_3s_3_2_1_U1.top_sub_3ns_3s_3_2_1_Adder_0_U.s  = { \sub_3ns_3s_3_2_1_U1.top_sub_3ns_3s_3_2_1_Adder_0_U.fas_s2 , \sub_3ns_3s_3_2_1_U1.top_sub_3ns_3s_3_2_1_Adder_0_U.sum_s1  };
assign \sub_3ns_3s_3_2_1_U1.top_sub_3ns_3s_3_2_1_Adder_0_U.u2.a  = \sub_3ns_3s_3_2_1_U1.top_sub_3ns_3s_3_2_1_Adder_0_U.ain_s1 ;
assign \sub_3ns_3s_3_2_1_U1.top_sub_3ns_3s_3_2_1_Adder_0_U.u2.b  = \sub_3ns_3s_3_2_1_U1.top_sub_3ns_3s_3_2_1_Adder_0_U.bin_s1 ;
assign \sub_3ns_3s_3_2_1_U1.top_sub_3ns_3s_3_2_1_Adder_0_U.u2.cin  = \sub_3ns_3s_3_2_1_U1.top_sub_3ns_3s_3_2_1_Adder_0_U.carry_s1 ;
assign \sub_3ns_3s_3_2_1_U1.top_sub_3ns_3s_3_2_1_Adder_0_U.facout_s2  = \sub_3ns_3s_3_2_1_U1.top_sub_3ns_3s_3_2_1_Adder_0_U.u2.cout ;
assign \sub_3ns_3s_3_2_1_U1.top_sub_3ns_3s_3_2_1_Adder_0_U.fas_s2  = \sub_3ns_3s_3_2_1_U1.top_sub_3ns_3s_3_2_1_Adder_0_U.u2.s ;
assign \sub_3ns_3s_3_2_1_U1.top_sub_3ns_3s_3_2_1_Adder_0_U.u1.a  = \sub_3ns_3s_3_2_1_U1.top_sub_3ns_3s_3_2_1_Adder_0_U.a [0];
assign \sub_3ns_3s_3_2_1_U1.top_sub_3ns_3s_3_2_1_Adder_0_U.u1.b  = \sub_3ns_3s_3_2_1_U1.top_sub_3ns_3s_3_2_1_Adder_0_U.bin_s0 [0];
assign \sub_3ns_3s_3_2_1_U1.top_sub_3ns_3s_3_2_1_Adder_0_U.u1.cin  = 1'h1;
assign \sub_3ns_3s_3_2_1_U1.top_sub_3ns_3s_3_2_1_Adder_0_U.facout_s1  = \sub_3ns_3s_3_2_1_U1.top_sub_3ns_3s_3_2_1_Adder_0_U.u1.cout ;
assign \sub_3ns_3s_3_2_1_U1.top_sub_3ns_3s_3_2_1_Adder_0_U.fas_s1  = \sub_3ns_3s_3_2_1_U1.top_sub_3ns_3s_3_2_1_Adder_0_U.u1.s ;
assign \sub_3ns_3s_3_2_1_U1.top_sub_3ns_3s_3_2_1_Adder_0_U.a  = \sub_3ns_3s_3_2_1_U1.din0 ;
assign \sub_3ns_3s_3_2_1_U1.top_sub_3ns_3s_3_2_1_Adder_0_U.b  = \sub_3ns_3s_3_2_1_U1.din1 ;
assign \sub_3ns_3s_3_2_1_U1.top_sub_3ns_3s_3_2_1_Adder_0_U.ce  = \sub_3ns_3s_3_2_1_U1.ce ;
assign \sub_3ns_3s_3_2_1_U1.top_sub_3ns_3s_3_2_1_Adder_0_U.clk  = \sub_3ns_3s_3_2_1_U1.clk ;
assign \sub_3ns_3s_3_2_1_U1.top_sub_3ns_3s_3_2_1_Adder_0_U.reset  = \sub_3ns_3s_3_2_1_U1.reset ;
assign \sub_3ns_3s_3_2_1_U1.dout  = \sub_3ns_3s_3_2_1_U1.top_sub_3ns_3s_3_2_1_Adder_0_U.s ;
assign \sub_3ns_3s_3_2_1_U1.ce  = 1'h1;
assign \sub_3ns_3s_3_2_1_U1.clk  = ap_clk;
assign \sub_3ns_3s_3_2_1_U1.din0  = select_ln1347_reg_929;
assign \sub_3ns_3s_3_2_1_U1.din1  = { op_4[1], op_4 };
assign grp_fu_217_p2 = \sub_3ns_3s_3_2_1_U1.dout ;
assign \sub_3ns_3s_3_2_1_U1.reset  = ap_rst;
assign \sub_2ns_2s_2_2_1_U10.top_sub_2ns_2s_2_2_1_Adder_7_U.ain_s0  = \sub_2ns_2s_2_2_1_U10.top_sub_2ns_2s_2_2_1_Adder_7_U.a ;
assign \sub_2ns_2s_2_2_1_U10.top_sub_2ns_2s_2_2_1_Adder_7_U.s  = { \sub_2ns_2s_2_2_1_U10.top_sub_2ns_2s_2_2_1_Adder_7_U.fas_s2 , \sub_2ns_2s_2_2_1_U10.top_sub_2ns_2s_2_2_1_Adder_7_U.sum_s1  };
assign \sub_2ns_2s_2_2_1_U10.top_sub_2ns_2s_2_2_1_Adder_7_U.u2.a  = \sub_2ns_2s_2_2_1_U10.top_sub_2ns_2s_2_2_1_Adder_7_U.ain_s1 ;
assign \sub_2ns_2s_2_2_1_U10.top_sub_2ns_2s_2_2_1_Adder_7_U.u2.b  = \sub_2ns_2s_2_2_1_U10.top_sub_2ns_2s_2_2_1_Adder_7_U.bin_s1 ;
assign \sub_2ns_2s_2_2_1_U10.top_sub_2ns_2s_2_2_1_Adder_7_U.u2.cin  = \sub_2ns_2s_2_2_1_U10.top_sub_2ns_2s_2_2_1_Adder_7_U.carry_s1 ;
assign \sub_2ns_2s_2_2_1_U10.top_sub_2ns_2s_2_2_1_Adder_7_U.facout_s2  = \sub_2ns_2s_2_2_1_U10.top_sub_2ns_2s_2_2_1_Adder_7_U.u2.cout ;
assign \sub_2ns_2s_2_2_1_U10.top_sub_2ns_2s_2_2_1_Adder_7_U.fas_s2  = \sub_2ns_2s_2_2_1_U10.top_sub_2ns_2s_2_2_1_Adder_7_U.u2.s ;
assign \sub_2ns_2s_2_2_1_U10.top_sub_2ns_2s_2_2_1_Adder_7_U.u1.a  = \sub_2ns_2s_2_2_1_U10.top_sub_2ns_2s_2_2_1_Adder_7_U.a [0];
assign \sub_2ns_2s_2_2_1_U10.top_sub_2ns_2s_2_2_1_Adder_7_U.u1.b  = \sub_2ns_2s_2_2_1_U10.top_sub_2ns_2s_2_2_1_Adder_7_U.bin_s0 [0];
assign \sub_2ns_2s_2_2_1_U10.top_sub_2ns_2s_2_2_1_Adder_7_U.u1.cin  = 1'h1;
assign \sub_2ns_2s_2_2_1_U10.top_sub_2ns_2s_2_2_1_Adder_7_U.facout_s1  = \sub_2ns_2s_2_2_1_U10.top_sub_2ns_2s_2_2_1_Adder_7_U.u1.cout ;
assign \sub_2ns_2s_2_2_1_U10.top_sub_2ns_2s_2_2_1_Adder_7_U.fas_s1  = \sub_2ns_2s_2_2_1_U10.top_sub_2ns_2s_2_2_1_Adder_7_U.u1.s ;
assign \sub_2ns_2s_2_2_1_U10.top_sub_2ns_2s_2_2_1_Adder_7_U.a  = \sub_2ns_2s_2_2_1_U10.din0 ;
assign \sub_2ns_2s_2_2_1_U10.top_sub_2ns_2s_2_2_1_Adder_7_U.b  = \sub_2ns_2s_2_2_1_U10.din1 ;
assign \sub_2ns_2s_2_2_1_U10.top_sub_2ns_2s_2_2_1_Adder_7_U.ce  = \sub_2ns_2s_2_2_1_U10.ce ;
assign \sub_2ns_2s_2_2_1_U10.top_sub_2ns_2s_2_2_1_Adder_7_U.clk  = \sub_2ns_2s_2_2_1_U10.clk ;
assign \sub_2ns_2s_2_2_1_U10.top_sub_2ns_2s_2_2_1_Adder_7_U.reset  = \sub_2ns_2s_2_2_1_U10.reset ;
assign \sub_2ns_2s_2_2_1_U10.dout  = \sub_2ns_2s_2_2_1_U10.top_sub_2ns_2s_2_2_1_Adder_7_U.s ;
assign \sub_2ns_2s_2_2_1_U10.ce  = 1'h1;
assign \sub_2ns_2s_2_2_1_U10.clk  = ap_clk;
assign \sub_2ns_2s_2_2_1_U10.din0  = 2'h0;
assign \sub_2ns_2s_2_2_1_U10.din1  = op_4;
assign grp_fu_563_p2 = \sub_2ns_2s_2_2_1_U10.dout ;
assign \sub_2ns_2s_2_2_1_U10.reset  = ap_rst;
assign \sub_2ns_2ns_2_2_1_U2.top_sub_2ns_2ns_2_2_1_Adder_1_U.ain_s0  = \sub_2ns_2ns_2_2_1_U2.top_sub_2ns_2ns_2_2_1_Adder_1_U.a ;
assign \sub_2ns_2ns_2_2_1_U2.top_sub_2ns_2ns_2_2_1_Adder_1_U.s  = { \sub_2ns_2ns_2_2_1_U2.top_sub_2ns_2ns_2_2_1_Adder_1_U.fas_s2 , \sub_2ns_2ns_2_2_1_U2.top_sub_2ns_2ns_2_2_1_Adder_1_U.sum_s1  };
assign \sub_2ns_2ns_2_2_1_U2.top_sub_2ns_2ns_2_2_1_Adder_1_U.u2.a  = \sub_2ns_2ns_2_2_1_U2.top_sub_2ns_2ns_2_2_1_Adder_1_U.ain_s1 ;
assign \sub_2ns_2ns_2_2_1_U2.top_sub_2ns_2ns_2_2_1_Adder_1_U.u2.b  = \sub_2ns_2ns_2_2_1_U2.top_sub_2ns_2ns_2_2_1_Adder_1_U.bin_s1 ;
assign \sub_2ns_2ns_2_2_1_U2.top_sub_2ns_2ns_2_2_1_Adder_1_U.u2.cin  = \sub_2ns_2ns_2_2_1_U2.top_sub_2ns_2ns_2_2_1_Adder_1_U.carry_s1 ;
assign \sub_2ns_2ns_2_2_1_U2.top_sub_2ns_2ns_2_2_1_Adder_1_U.facout_s2  = \sub_2ns_2ns_2_2_1_U2.top_sub_2ns_2ns_2_2_1_Adder_1_U.u2.cout ;
assign \sub_2ns_2ns_2_2_1_U2.top_sub_2ns_2ns_2_2_1_Adder_1_U.fas_s2  = \sub_2ns_2ns_2_2_1_U2.top_sub_2ns_2ns_2_2_1_Adder_1_U.u2.s ;
assign \sub_2ns_2ns_2_2_1_U2.top_sub_2ns_2ns_2_2_1_Adder_1_U.u1.a  = \sub_2ns_2ns_2_2_1_U2.top_sub_2ns_2ns_2_2_1_Adder_1_U.a [0];
assign \sub_2ns_2ns_2_2_1_U2.top_sub_2ns_2ns_2_2_1_Adder_1_U.u1.b  = \sub_2ns_2ns_2_2_1_U2.top_sub_2ns_2ns_2_2_1_Adder_1_U.bin_s0 [0];
assign \sub_2ns_2ns_2_2_1_U2.top_sub_2ns_2ns_2_2_1_Adder_1_U.u1.cin  = 1'h1;
assign \sub_2ns_2ns_2_2_1_U2.top_sub_2ns_2ns_2_2_1_Adder_1_U.facout_s1  = \sub_2ns_2ns_2_2_1_U2.top_sub_2ns_2ns_2_2_1_Adder_1_U.u1.cout ;
assign \sub_2ns_2ns_2_2_1_U2.top_sub_2ns_2ns_2_2_1_Adder_1_U.fas_s1  = \sub_2ns_2ns_2_2_1_U2.top_sub_2ns_2ns_2_2_1_Adder_1_U.u1.s ;
assign \sub_2ns_2ns_2_2_1_U2.top_sub_2ns_2ns_2_2_1_Adder_1_U.a  = \sub_2ns_2ns_2_2_1_U2.din0 ;
assign \sub_2ns_2ns_2_2_1_U2.top_sub_2ns_2ns_2_2_1_Adder_1_U.b  = \sub_2ns_2ns_2_2_1_U2.din1 ;
assign \sub_2ns_2ns_2_2_1_U2.top_sub_2ns_2ns_2_2_1_Adder_1_U.ce  = \sub_2ns_2ns_2_2_1_U2.ce ;
assign \sub_2ns_2ns_2_2_1_U2.top_sub_2ns_2ns_2_2_1_Adder_1_U.clk  = \sub_2ns_2ns_2_2_1_U2.clk ;
assign \sub_2ns_2ns_2_2_1_U2.top_sub_2ns_2ns_2_2_1_Adder_1_U.reset  = \sub_2ns_2ns_2_2_1_U2.reset ;
assign \sub_2ns_2ns_2_2_1_U2.dout  = \sub_2ns_2ns_2_2_1_U2.top_sub_2ns_2ns_2_2_1_Adder_1_U.s ;
assign \sub_2ns_2ns_2_2_1_U2.ce  = 1'h1;
assign \sub_2ns_2ns_2_2_1_U2.clk  = ap_clk;
assign \sub_2ns_2ns_2_2_1_U2.din0  = 2'h0;
assign \sub_2ns_2ns_2_2_1_U2.din1  = r_2_reg_980;
assign grp_fu_332_p2 = \sub_2ns_2ns_2_2_1_U2.dout ;
assign \sub_2ns_2ns_2_2_1_U2.reset  = ap_rst;
assign \sub_27ns_27s_27_2_1_U5.top_sub_27ns_27s_27_2_1_Adder_2_U.ain_s0  = \sub_27ns_27s_27_2_1_U5.top_sub_27ns_27s_27_2_1_Adder_2_U.a ;
assign \sub_27ns_27s_27_2_1_U5.top_sub_27ns_27s_27_2_1_Adder_2_U.s  = { \sub_27ns_27s_27_2_1_U5.top_sub_27ns_27s_27_2_1_Adder_2_U.fas_s2 , \sub_27ns_27s_27_2_1_U5.top_sub_27ns_27s_27_2_1_Adder_2_U.sum_s1  };
assign \sub_27ns_27s_27_2_1_U5.top_sub_27ns_27s_27_2_1_Adder_2_U.u2.a  = \sub_27ns_27s_27_2_1_U5.top_sub_27ns_27s_27_2_1_Adder_2_U.ain_s1 ;
assign \sub_27ns_27s_27_2_1_U5.top_sub_27ns_27s_27_2_1_Adder_2_U.u2.b  = \sub_27ns_27s_27_2_1_U5.top_sub_27ns_27s_27_2_1_Adder_2_U.bin_s1 ;
assign \sub_27ns_27s_27_2_1_U5.top_sub_27ns_27s_27_2_1_Adder_2_U.u2.cin  = \sub_27ns_27s_27_2_1_U5.top_sub_27ns_27s_27_2_1_Adder_2_U.carry_s1 ;
assign \sub_27ns_27s_27_2_1_U5.top_sub_27ns_27s_27_2_1_Adder_2_U.facout_s2  = \sub_27ns_27s_27_2_1_U5.top_sub_27ns_27s_27_2_1_Adder_2_U.u2.cout ;
assign \sub_27ns_27s_27_2_1_U5.top_sub_27ns_27s_27_2_1_Adder_2_U.fas_s2  = \sub_27ns_27s_27_2_1_U5.top_sub_27ns_27s_27_2_1_Adder_2_U.u2.s ;
assign \sub_27ns_27s_27_2_1_U5.top_sub_27ns_27s_27_2_1_Adder_2_U.u1.a  = \sub_27ns_27s_27_2_1_U5.top_sub_27ns_27s_27_2_1_Adder_2_U.a [12:0];
assign \sub_27ns_27s_27_2_1_U5.top_sub_27ns_27s_27_2_1_Adder_2_U.u1.b  = \sub_27ns_27s_27_2_1_U5.top_sub_27ns_27s_27_2_1_Adder_2_U.bin_s0 [12:0];
assign \sub_27ns_27s_27_2_1_U5.top_sub_27ns_27s_27_2_1_Adder_2_U.u1.cin  = 1'h1;
assign \sub_27ns_27s_27_2_1_U5.top_sub_27ns_27s_27_2_1_Adder_2_U.facout_s1  = \sub_27ns_27s_27_2_1_U5.top_sub_27ns_27s_27_2_1_Adder_2_U.u1.cout ;
assign \sub_27ns_27s_27_2_1_U5.top_sub_27ns_27s_27_2_1_Adder_2_U.fas_s1  = \sub_27ns_27s_27_2_1_U5.top_sub_27ns_27s_27_2_1_Adder_2_U.u1.s ;
assign \sub_27ns_27s_27_2_1_U5.top_sub_27ns_27s_27_2_1_Adder_2_U.a  = \sub_27ns_27s_27_2_1_U5.din0 ;
assign \sub_27ns_27s_27_2_1_U5.top_sub_27ns_27s_27_2_1_Adder_2_U.b  = \sub_27ns_27s_27_2_1_U5.din1 ;
assign \sub_27ns_27s_27_2_1_U5.top_sub_27ns_27s_27_2_1_Adder_2_U.ce  = \sub_27ns_27s_27_2_1_U5.ce ;
assign \sub_27ns_27s_27_2_1_U5.top_sub_27ns_27s_27_2_1_Adder_2_U.clk  = \sub_27ns_27s_27_2_1_U5.clk ;
assign \sub_27ns_27s_27_2_1_U5.top_sub_27ns_27s_27_2_1_Adder_2_U.reset  = \sub_27ns_27s_27_2_1_U5.reset ;
assign \sub_27ns_27s_27_2_1_U5.dout  = \sub_27ns_27s_27_2_1_U5.top_sub_27ns_27s_27_2_1_Adder_2_U.s ;
assign \sub_27ns_27s_27_2_1_U5.ce  = 1'h1;
assign \sub_27ns_27s_27_2_1_U5.clk  = ap_clk;
assign \sub_27ns_27s_27_2_1_U5.din0  = 27'h0000000;
assign \sub_27ns_27s_27_2_1_U5.din1  = { op_4[1], op_4, 24'h000000 };
assign grp_fu_399_p2 = \sub_27ns_27s_27_2_1_U5.dout ;
assign \sub_27ns_27s_27_2_1_U5.reset  = ap_rst;
assign \shl_4s_2ns_4_7_1_U4.din1_cast  = \shl_4s_2ns_4_7_1_U4.din1 [1:0];
assign \shl_4s_2ns_4_7_1_U4.din1_mask  = 2'h1;
assign \shl_4s_2ns_4_7_1_U4.ce  = 1'h1;
assign \shl_4s_2ns_4_7_1_U4.clk  = ap_clk;
assign \shl_4s_2ns_4_7_1_U4.din0  = op_8_V_reg_1018;
assign \shl_4s_2ns_4_7_1_U4.din1  = { 2'h0, ush_reg_1026 };
assign grp_fu_383_p2 = \shl_4s_2ns_4_7_1_U4.dout ;
assign \shl_4s_2ns_4_7_1_U4.reset  = ap_rst;
assign \ashr_4s_2ns_4_7_1_U3.din1_cast  = \ashr_4s_2ns_4_7_1_U3.din1 [1:0];
assign \ashr_4s_2ns_4_7_1_U3.din1_mask  = 2'h1;
assign \ashr_4s_2ns_4_7_1_U3.ce  = 1'h1;
assign \ashr_4s_2ns_4_7_1_U3.clk  = ap_clk;
assign \ashr_4s_2ns_4_7_1_U3.din0  = op_8_V_reg_1018;
assign \ashr_4s_2ns_4_7_1_U3.din1  = { 2'h0, ush_reg_1026 };
assign grp_fu_378_p2 = \ashr_4s_2ns_4_7_1_U3.dout ;
assign \ashr_4s_2ns_4_7_1_U3.reset  = ap_rst;
assign \add_9s_9ns_9_2_1_U6.top_add_9s_9ns_9_2_1_Adder_3_U.ain_s0  = \add_9s_9ns_9_2_1_U6.top_add_9s_9ns_9_2_1_Adder_3_U.a ;
assign \add_9s_9ns_9_2_1_U6.top_add_9s_9ns_9_2_1_Adder_3_U.bin_s0  = \add_9s_9ns_9_2_1_U6.top_add_9s_9ns_9_2_1_Adder_3_U.b ;
assign \add_9s_9ns_9_2_1_U6.top_add_9s_9ns_9_2_1_Adder_3_U.s  = { \add_9s_9ns_9_2_1_U6.top_add_9s_9ns_9_2_1_Adder_3_U.fas_s2 , \add_9s_9ns_9_2_1_U6.top_add_9s_9ns_9_2_1_Adder_3_U.sum_s1  };
assign \add_9s_9ns_9_2_1_U6.top_add_9s_9ns_9_2_1_Adder_3_U.u2.a  = \add_9s_9ns_9_2_1_U6.top_add_9s_9ns_9_2_1_Adder_3_U.ain_s1 ;
assign \add_9s_9ns_9_2_1_U6.top_add_9s_9ns_9_2_1_Adder_3_U.u2.b  = \add_9s_9ns_9_2_1_U6.top_add_9s_9ns_9_2_1_Adder_3_U.bin_s1 ;
assign \add_9s_9ns_9_2_1_U6.top_add_9s_9ns_9_2_1_Adder_3_U.u2.cin  = \add_9s_9ns_9_2_1_U6.top_add_9s_9ns_9_2_1_Adder_3_U.carry_s1 ;
assign \add_9s_9ns_9_2_1_U6.top_add_9s_9ns_9_2_1_Adder_3_U.facout_s2  = \add_9s_9ns_9_2_1_U6.top_add_9s_9ns_9_2_1_Adder_3_U.u2.cout ;
assign \add_9s_9ns_9_2_1_U6.top_add_9s_9ns_9_2_1_Adder_3_U.fas_s2  = \add_9s_9ns_9_2_1_U6.top_add_9s_9ns_9_2_1_Adder_3_U.u2.s ;
assign \add_9s_9ns_9_2_1_U6.top_add_9s_9ns_9_2_1_Adder_3_U.u1.a  = \add_9s_9ns_9_2_1_U6.top_add_9s_9ns_9_2_1_Adder_3_U.a [3:0];
assign \add_9s_9ns_9_2_1_U6.top_add_9s_9ns_9_2_1_Adder_3_U.u1.b  = \add_9s_9ns_9_2_1_U6.top_add_9s_9ns_9_2_1_Adder_3_U.b [3:0];
assign \add_9s_9ns_9_2_1_U6.top_add_9s_9ns_9_2_1_Adder_3_U.u1.cin  = 1'h0;
assign \add_9s_9ns_9_2_1_U6.top_add_9s_9ns_9_2_1_Adder_3_U.facout_s1  = \add_9s_9ns_9_2_1_U6.top_add_9s_9ns_9_2_1_Adder_3_U.u1.cout ;
assign \add_9s_9ns_9_2_1_U6.top_add_9s_9ns_9_2_1_Adder_3_U.fas_s1  = \add_9s_9ns_9_2_1_U6.top_add_9s_9ns_9_2_1_Adder_3_U.u1.s ;
assign \add_9s_9ns_9_2_1_U6.top_add_9s_9ns_9_2_1_Adder_3_U.a  = \add_9s_9ns_9_2_1_U6.din0 ;
assign \add_9s_9ns_9_2_1_U6.top_add_9s_9ns_9_2_1_Adder_3_U.b  = \add_9s_9ns_9_2_1_U6.din1 ;
assign \add_9s_9ns_9_2_1_U6.top_add_9s_9ns_9_2_1_Adder_3_U.ce  = \add_9s_9ns_9_2_1_U6.ce ;
assign \add_9s_9ns_9_2_1_U6.top_add_9s_9ns_9_2_1_Adder_3_U.clk  = \add_9s_9ns_9_2_1_U6.clk ;
assign \add_9s_9ns_9_2_1_U6.top_add_9s_9ns_9_2_1_Adder_3_U.reset  = \add_9s_9ns_9_2_1_U6.reset ;
assign \add_9s_9ns_9_2_1_U6.dout  = \add_9s_9ns_9_2_1_U6.top_add_9s_9ns_9_2_1_Adder_3_U.s ;
assign \add_9s_9ns_9_2_1_U6.ce  = 1'h1;
assign \add_9s_9ns_9_2_1_U6.clk  = ap_clk;
assign \add_9s_9ns_9_2_1_U6.din0  = { op_0[7], op_0 };
assign \add_9s_9ns_9_2_1_U6.din1  = 9'h008;
assign grp_fu_434_p2 = \add_9s_9ns_9_2_1_U6.dout ;
assign \add_9s_9ns_9_2_1_U6.reset  = ap_rst;
assign \add_7s_7s_7_2_1_U11.top_add_7s_7s_7_2_1_Adder_8_U.ain_s0  = \add_7s_7s_7_2_1_U11.top_add_7s_7s_7_2_1_Adder_8_U.a ;
assign \add_7s_7s_7_2_1_U11.top_add_7s_7s_7_2_1_Adder_8_U.bin_s0  = \add_7s_7s_7_2_1_U11.top_add_7s_7s_7_2_1_Adder_8_U.b ;
assign \add_7s_7s_7_2_1_U11.top_add_7s_7s_7_2_1_Adder_8_U.s  = { \add_7s_7s_7_2_1_U11.top_add_7s_7s_7_2_1_Adder_8_U.fas_s2 , \add_7s_7s_7_2_1_U11.top_add_7s_7s_7_2_1_Adder_8_U.sum_s1  };
assign \add_7s_7s_7_2_1_U11.top_add_7s_7s_7_2_1_Adder_8_U.u2.a  = \add_7s_7s_7_2_1_U11.top_add_7s_7s_7_2_1_Adder_8_U.ain_s1 ;
assign \add_7s_7s_7_2_1_U11.top_add_7s_7s_7_2_1_Adder_8_U.u2.b  = \add_7s_7s_7_2_1_U11.top_add_7s_7s_7_2_1_Adder_8_U.bin_s1 ;
assign \add_7s_7s_7_2_1_U11.top_add_7s_7s_7_2_1_Adder_8_U.u2.cin  = \add_7s_7s_7_2_1_U11.top_add_7s_7s_7_2_1_Adder_8_U.carry_s1 ;
assign \add_7s_7s_7_2_1_U11.top_add_7s_7s_7_2_1_Adder_8_U.facout_s2  = \add_7s_7s_7_2_1_U11.top_add_7s_7s_7_2_1_Adder_8_U.u2.cout ;
assign \add_7s_7s_7_2_1_U11.top_add_7s_7s_7_2_1_Adder_8_U.fas_s2  = \add_7s_7s_7_2_1_U11.top_add_7s_7s_7_2_1_Adder_8_U.u2.s ;
assign \add_7s_7s_7_2_1_U11.top_add_7s_7s_7_2_1_Adder_8_U.u1.a  = \add_7s_7s_7_2_1_U11.top_add_7s_7s_7_2_1_Adder_8_U.a [2:0];
assign \add_7s_7s_7_2_1_U11.top_add_7s_7s_7_2_1_Adder_8_U.u1.b  = \add_7s_7s_7_2_1_U11.top_add_7s_7s_7_2_1_Adder_8_U.b [2:0];
assign \add_7s_7s_7_2_1_U11.top_add_7s_7s_7_2_1_Adder_8_U.u1.cin  = 1'h0;
assign \add_7s_7s_7_2_1_U11.top_add_7s_7s_7_2_1_Adder_8_U.facout_s1  = \add_7s_7s_7_2_1_U11.top_add_7s_7s_7_2_1_Adder_8_U.u1.cout ;
assign \add_7s_7s_7_2_1_U11.top_add_7s_7s_7_2_1_Adder_8_U.fas_s1  = \add_7s_7s_7_2_1_U11.top_add_7s_7s_7_2_1_Adder_8_U.u1.s ;
assign \add_7s_7s_7_2_1_U11.top_add_7s_7s_7_2_1_Adder_8_U.a  = \add_7s_7s_7_2_1_U11.din0 ;
assign \add_7s_7s_7_2_1_U11.top_add_7s_7s_7_2_1_Adder_8_U.b  = \add_7s_7s_7_2_1_U11.din1 ;
assign \add_7s_7s_7_2_1_U11.top_add_7s_7s_7_2_1_Adder_8_U.ce  = \add_7s_7s_7_2_1_U11.ce ;
assign \add_7s_7s_7_2_1_U11.top_add_7s_7s_7_2_1_Adder_8_U.clk  = \add_7s_7s_7_2_1_U11.clk ;
assign \add_7s_7s_7_2_1_U11.top_add_7s_7s_7_2_1_Adder_8_U.reset  = \add_7s_7s_7_2_1_U11.reset ;
assign \add_7s_7s_7_2_1_U11.dout  = \add_7s_7s_7_2_1_U11.top_add_7s_7s_7_2_1_Adder_8_U.s ;
assign \add_7s_7s_7_2_1_U11.ce  = 1'h1;
assign \add_7s_7s_7_2_1_U11.clk  = ap_clk;
assign \add_7s_7s_7_2_1_U11.din0  = { ret_V_20_reg_1182[5], ret_V_20_reg_1182 };
assign \add_7s_7s_7_2_1_U11.din1  = { op_6_V_reg_1177[1], op_6_V_reg_1177[1], op_6_V_reg_1177[1], op_6_V_reg_1177[1], op_6_V_reg_1177[1], op_6_V_reg_1177 };
assign grp_fu_661_p2 = \add_7s_7s_7_2_1_U11.dout ;
assign \add_7s_7s_7_2_1_U11.reset  = ap_rst;
assign \add_7s_7ns_7_2_1_U16.top_add_7s_7ns_7_2_1_Adder_10_U.ain_s0  = \add_7s_7ns_7_2_1_U16.top_add_7s_7ns_7_2_1_Adder_10_U.a ;
assign \add_7s_7ns_7_2_1_U16.top_add_7s_7ns_7_2_1_Adder_10_U.bin_s0  = \add_7s_7ns_7_2_1_U16.top_add_7s_7ns_7_2_1_Adder_10_U.b ;
assign \add_7s_7ns_7_2_1_U16.top_add_7s_7ns_7_2_1_Adder_10_U.s  = { \add_7s_7ns_7_2_1_U16.top_add_7s_7ns_7_2_1_Adder_10_U.fas_s2 , \add_7s_7ns_7_2_1_U16.top_add_7s_7ns_7_2_1_Adder_10_U.sum_s1  };
assign \add_7s_7ns_7_2_1_U16.top_add_7s_7ns_7_2_1_Adder_10_U.u2.a  = \add_7s_7ns_7_2_1_U16.top_add_7s_7ns_7_2_1_Adder_10_U.ain_s1 ;
assign \add_7s_7ns_7_2_1_U16.top_add_7s_7ns_7_2_1_Adder_10_U.u2.b  = \add_7s_7ns_7_2_1_U16.top_add_7s_7ns_7_2_1_Adder_10_U.bin_s1 ;
assign \add_7s_7ns_7_2_1_U16.top_add_7s_7ns_7_2_1_Adder_10_U.u2.cin  = \add_7s_7ns_7_2_1_U16.top_add_7s_7ns_7_2_1_Adder_10_U.carry_s1 ;
assign \add_7s_7ns_7_2_1_U16.top_add_7s_7ns_7_2_1_Adder_10_U.facout_s2  = \add_7s_7ns_7_2_1_U16.top_add_7s_7ns_7_2_1_Adder_10_U.u2.cout ;
assign \add_7s_7ns_7_2_1_U16.top_add_7s_7ns_7_2_1_Adder_10_U.fas_s2  = \add_7s_7ns_7_2_1_U16.top_add_7s_7ns_7_2_1_Adder_10_U.u2.s ;
assign \add_7s_7ns_7_2_1_U16.top_add_7s_7ns_7_2_1_Adder_10_U.u1.a  = \add_7s_7ns_7_2_1_U16.top_add_7s_7ns_7_2_1_Adder_10_U.a [2:0];
assign \add_7s_7ns_7_2_1_U16.top_add_7s_7ns_7_2_1_Adder_10_U.u1.b  = \add_7s_7ns_7_2_1_U16.top_add_7s_7ns_7_2_1_Adder_10_U.b [2:0];
assign \add_7s_7ns_7_2_1_U16.top_add_7s_7ns_7_2_1_Adder_10_U.u1.cin  = 1'h0;
assign \add_7s_7ns_7_2_1_U16.top_add_7s_7ns_7_2_1_Adder_10_U.facout_s1  = \add_7s_7ns_7_2_1_U16.top_add_7s_7ns_7_2_1_Adder_10_U.u1.cout ;
assign \add_7s_7ns_7_2_1_U16.top_add_7s_7ns_7_2_1_Adder_10_U.fas_s1  = \add_7s_7ns_7_2_1_U16.top_add_7s_7ns_7_2_1_Adder_10_U.u1.s ;
assign \add_7s_7ns_7_2_1_U16.top_add_7s_7ns_7_2_1_Adder_10_U.a  = \add_7s_7ns_7_2_1_U16.din0 ;
assign \add_7s_7ns_7_2_1_U16.top_add_7s_7ns_7_2_1_Adder_10_U.b  = \add_7s_7ns_7_2_1_U16.din1 ;
assign \add_7s_7ns_7_2_1_U16.top_add_7s_7ns_7_2_1_Adder_10_U.ce  = \add_7s_7ns_7_2_1_U16.ce ;
assign \add_7s_7ns_7_2_1_U16.top_add_7s_7ns_7_2_1_Adder_10_U.clk  = \add_7s_7ns_7_2_1_U16.clk ;
assign \add_7s_7ns_7_2_1_U16.top_add_7s_7ns_7_2_1_Adder_10_U.reset  = \add_7s_7ns_7_2_1_U16.reset ;
assign \add_7s_7ns_7_2_1_U16.dout  = \add_7s_7ns_7_2_1_U16.top_add_7s_7ns_7_2_1_Adder_10_U.s ;
assign \add_7s_7ns_7_2_1_U16.ce  = 1'h1;
assign \add_7s_7ns_7_2_1_U16.clk  = ap_clk;
assign \add_7s_7ns_7_2_1_U16.din0  = { add_ln69_3_reg_1272[2], add_ln69_3_reg_1272[2], add_ln69_3_reg_1272[2], add_ln69_3_reg_1272[2], add_ln69_3_reg_1272 };
assign \add_7s_7ns_7_2_1_U16.din1  = add_ln69_1_reg_1267;
assign grp_fu_717_p2 = \add_7s_7ns_7_2_1_U16.dout ;
assign \add_7s_7ns_7_2_1_U16.reset  = ap_rst;
assign \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_10_U.ain_s0  = \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_10_U.a ;
assign \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_10_U.bin_s0  = \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_10_U.b ;
assign \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_10_U.s  = { \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_10_U.fas_s2 , \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_10_U.sum_s1  };
assign \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_10_U.u2.a  = \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_10_U.ain_s1 ;
assign \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_10_U.u2.b  = \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_10_U.bin_s1 ;
assign \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_10_U.u2.cin  = \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_10_U.carry_s1 ;
assign \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_10_U.facout_s2  = \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_10_U.u2.cout ;
assign \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_10_U.fas_s2  = \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_10_U.u2.s ;
assign \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_10_U.u1.a  = \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_10_U.a [2:0];
assign \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_10_U.u1.b  = \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_10_U.b [2:0];
assign \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_10_U.u1.cin  = 1'h0;
assign \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_10_U.facout_s1  = \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_10_U.u1.cout ;
assign \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_10_U.fas_s1  = \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_10_U.u1.s ;
assign \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_10_U.a  = \add_7s_7ns_7_2_1_U14.din0 ;
assign \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_10_U.b  = \add_7s_7ns_7_2_1_U14.din1 ;
assign \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_10_U.ce  = \add_7s_7ns_7_2_1_U14.ce ;
assign \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_10_U.clk  = \add_7s_7ns_7_2_1_U14.clk ;
assign \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_10_U.reset  = \add_7s_7ns_7_2_1_U14.reset ;
assign \add_7s_7ns_7_2_1_U14.dout  = \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_10_U.s ;
assign \add_7s_7ns_7_2_1_U14.ce  = 1'h1;
assign \add_7s_7ns_7_2_1_U14.clk  = ap_clk;
assign \add_7s_7ns_7_2_1_U14.din0  = { add_ln69_reg_1242[5], add_ln69_reg_1242 };
assign \add_7s_7ns_7_2_1_U14.din1  = ret_V_23_reg_1237;
assign grp_fu_700_p2 = \add_7s_7ns_7_2_1_U14.dout ;
assign \add_7s_7ns_7_2_1_U14.reset  = ap_rst;
assign \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.ain_s0  = \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.a ;
assign \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.bin_s0  = \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.b ;
assign \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.s  = { \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.fas_s2 , \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.sum_s1  };
assign \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.u2.a  = \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.ain_s1 ;
assign \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.u2.b  = \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.bin_s1 ;
assign \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.u2.cin  = \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.carry_s1 ;
assign \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.facout_s2  = \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.u2.cout ;
assign \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.fas_s2  = \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.u2.s ;
assign \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.u1.a  = \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.a [2:0];
assign \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.u1.b  = \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.b [2:0];
assign \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.u1.cin  = 1'h0;
assign \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.facout_s1  = \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.u1.cout ;
assign \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.fas_s1  = \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.u1.s ;
assign \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.a  = \add_6s_6ns_6_2_1_U12.din0 ;
assign \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.b  = \add_6s_6ns_6_2_1_U12.din1 ;
assign \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.ce  = \add_6s_6ns_6_2_1_U12.ce ;
assign \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.clk  = \add_6s_6ns_6_2_1_U12.clk ;
assign \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.reset  = \add_6s_6ns_6_2_1_U12.reset ;
assign \add_6s_6ns_6_2_1_U12.dout  = \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.s ;
assign \add_6s_6ns_6_2_1_U12.ce  = 1'h1;
assign \add_6s_6ns_6_2_1_U12.clk  = ap_clk;
assign \add_6s_6ns_6_2_1_U12.din0  = { ret_V_21_reg_1187[3], ret_V_21_reg_1187[3], ret_V_21_reg_1187 };
assign \add_6s_6ns_6_2_1_U12.din1  = { 2'h0, op_12 };
assign grp_fu_677_p2 = \add_6s_6ns_6_2_1_U12.dout ;
assign \add_6s_6ns_6_2_1_U12.reset  = ap_rst;
assign \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_4_U.ain_s0  = \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_4_U.a ;
assign \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_4_U.bin_s0  = \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_4_U.b ;
assign \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_4_U.s  = { \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_4_U.fas_s2 , \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_4_U.sum_s1  };
assign \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_4_U.u2.a  = \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_4_U.ain_s1 ;
assign \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_4_U.u2.b  = \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_4_U.bin_s1 ;
assign \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_4_U.u2.cin  = \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_4_U.carry_s1 ;
assign \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_4_U.facout_s2  = \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_4_U.u2.cout ;
assign \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_4_U.fas_s2  = \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_4_U.u2.s ;
assign \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_4_U.u1.a  = \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_4_U.a [2:0];
assign \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_4_U.u1.b  = \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_4_U.b [2:0];
assign \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_4_U.u1.cin  = 1'h0;
assign \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_4_U.facout_s1  = \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_4_U.u1.cout ;
assign \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_4_U.fas_s1  = \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_4_U.u1.s ;
assign \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_4_U.a  = \add_6ns_6ns_6_2_1_U7.din0 ;
assign \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_4_U.b  = \add_6ns_6ns_6_2_1_U7.din1 ;
assign \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_4_U.ce  = \add_6ns_6ns_6_2_1_U7.ce ;
assign \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_4_U.clk  = \add_6ns_6ns_6_2_1_U7.clk ;
assign \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_4_U.reset  = \add_6ns_6ns_6_2_1_U7.reset ;
assign \add_6ns_6ns_6_2_1_U7.dout  = \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_4_U.s ;
assign \add_6ns_6ns_6_2_1_U7.ce  = 1'h1;
assign \add_6ns_6ns_6_2_1_U7.clk  = ap_clk;
assign \add_6ns_6ns_6_2_1_U7.din0  = ret_V_reg_1082;
assign \add_6ns_6ns_6_2_1_U7.din1  = 6'h01;
assign grp_fu_522_p2 = \add_6ns_6ns_6_2_1_U7.dout ;
assign \add_6ns_6ns_6_2_1_U7.reset  = ap_rst;
assign \add_4s_4ns_4_2_1_U8.top_add_4s_4ns_4_2_1_Adder_5_U.ain_s0  = \add_4s_4ns_4_2_1_U8.top_add_4s_4ns_4_2_1_Adder_5_U.a ;
assign \add_4s_4ns_4_2_1_U8.top_add_4s_4ns_4_2_1_Adder_5_U.bin_s0  = \add_4s_4ns_4_2_1_U8.top_add_4s_4ns_4_2_1_Adder_5_U.b ;
assign \add_4s_4ns_4_2_1_U8.top_add_4s_4ns_4_2_1_Adder_5_U.s  = { \add_4s_4ns_4_2_1_U8.top_add_4s_4ns_4_2_1_Adder_5_U.fas_s2 , \add_4s_4ns_4_2_1_U8.top_add_4s_4ns_4_2_1_Adder_5_U.sum_s1  };
assign \add_4s_4ns_4_2_1_U8.top_add_4s_4ns_4_2_1_Adder_5_U.u2.a  = \add_4s_4ns_4_2_1_U8.top_add_4s_4ns_4_2_1_Adder_5_U.ain_s1 ;
assign \add_4s_4ns_4_2_1_U8.top_add_4s_4ns_4_2_1_Adder_5_U.u2.b  = \add_4s_4ns_4_2_1_U8.top_add_4s_4ns_4_2_1_Adder_5_U.bin_s1 ;
assign \add_4s_4ns_4_2_1_U8.top_add_4s_4ns_4_2_1_Adder_5_U.u2.cin  = \add_4s_4ns_4_2_1_U8.top_add_4s_4ns_4_2_1_Adder_5_U.carry_s1 ;
assign \add_4s_4ns_4_2_1_U8.top_add_4s_4ns_4_2_1_Adder_5_U.facout_s2  = \add_4s_4ns_4_2_1_U8.top_add_4s_4ns_4_2_1_Adder_5_U.u2.cout ;
assign \add_4s_4ns_4_2_1_U8.top_add_4s_4ns_4_2_1_Adder_5_U.fas_s2  = \add_4s_4ns_4_2_1_U8.top_add_4s_4ns_4_2_1_Adder_5_U.u2.s ;
assign \add_4s_4ns_4_2_1_U8.top_add_4s_4ns_4_2_1_Adder_5_U.u1.a  = \add_4s_4ns_4_2_1_U8.top_add_4s_4ns_4_2_1_Adder_5_U.a [1:0];
assign \add_4s_4ns_4_2_1_U8.top_add_4s_4ns_4_2_1_Adder_5_U.u1.b  = \add_4s_4ns_4_2_1_U8.top_add_4s_4ns_4_2_1_Adder_5_U.b [1:0];
assign \add_4s_4ns_4_2_1_U8.top_add_4s_4ns_4_2_1_Adder_5_U.u1.cin  = 1'h0;
assign \add_4s_4ns_4_2_1_U8.top_add_4s_4ns_4_2_1_Adder_5_U.facout_s1  = \add_4s_4ns_4_2_1_U8.top_add_4s_4ns_4_2_1_Adder_5_U.u1.cout ;
assign \add_4s_4ns_4_2_1_U8.top_add_4s_4ns_4_2_1_Adder_5_U.fas_s1  = \add_4s_4ns_4_2_1_U8.top_add_4s_4ns_4_2_1_Adder_5_U.u1.s ;
assign \add_4s_4ns_4_2_1_U8.top_add_4s_4ns_4_2_1_Adder_5_U.a  = \add_4s_4ns_4_2_1_U8.din0 ;
assign \add_4s_4ns_4_2_1_U8.top_add_4s_4ns_4_2_1_Adder_5_U.b  = \add_4s_4ns_4_2_1_U8.din1 ;
assign \add_4s_4ns_4_2_1_U8.top_add_4s_4ns_4_2_1_Adder_5_U.ce  = \add_4s_4ns_4_2_1_U8.ce ;
assign \add_4s_4ns_4_2_1_U8.top_add_4s_4ns_4_2_1_Adder_5_U.clk  = \add_4s_4ns_4_2_1_U8.clk ;
assign \add_4s_4ns_4_2_1_U8.top_add_4s_4ns_4_2_1_Adder_5_U.reset  = \add_4s_4ns_4_2_1_U8.reset ;
assign \add_4s_4ns_4_2_1_U8.dout  = \add_4s_4ns_4_2_1_U8.top_add_4s_4ns_4_2_1_Adder_5_U.s ;
assign \add_4s_4ns_4_2_1_U8.ce  = 1'h1;
assign \add_4s_4ns_4_2_1_U8.clk  = ap_clk;
assign \add_4s_4ns_4_2_1_U8.din0  = { tmp_2_reg_1099[2], tmp_2_reg_1099 };
assign \add_4s_4ns_4_2_1_U8.din1  = 4'h1;
assign grp_fu_535_p2 = \add_4s_4ns_4_2_1_U8.dout ;
assign \add_4s_4ns_4_2_1_U8.reset  = ap_rst;
assign \add_3s_3s_3_2_1_U15.top_add_3s_3s_3_2_1_Adder_11_U.ain_s0  = \add_3s_3s_3_2_1_U15.top_add_3s_3s_3_2_1_Adder_11_U.a ;
assign \add_3s_3s_3_2_1_U15.top_add_3s_3s_3_2_1_Adder_11_U.bin_s0  = \add_3s_3s_3_2_1_U15.top_add_3s_3s_3_2_1_Adder_11_U.b ;
assign \add_3s_3s_3_2_1_U15.top_add_3s_3s_3_2_1_Adder_11_U.s  = { \add_3s_3s_3_2_1_U15.top_add_3s_3s_3_2_1_Adder_11_U.fas_s2 , \add_3s_3s_3_2_1_U15.top_add_3s_3s_3_2_1_Adder_11_U.sum_s1  };
assign \add_3s_3s_3_2_1_U15.top_add_3s_3s_3_2_1_Adder_11_U.u2.a  = \add_3s_3s_3_2_1_U15.top_add_3s_3s_3_2_1_Adder_11_U.ain_s1 ;
assign \add_3s_3s_3_2_1_U15.top_add_3s_3s_3_2_1_Adder_11_U.u2.b  = \add_3s_3s_3_2_1_U15.top_add_3s_3s_3_2_1_Adder_11_U.bin_s1 ;
assign \add_3s_3s_3_2_1_U15.top_add_3s_3s_3_2_1_Adder_11_U.u2.cin  = \add_3s_3s_3_2_1_U15.top_add_3s_3s_3_2_1_Adder_11_U.carry_s1 ;
assign \add_3s_3s_3_2_1_U15.top_add_3s_3s_3_2_1_Adder_11_U.facout_s2  = \add_3s_3s_3_2_1_U15.top_add_3s_3s_3_2_1_Adder_11_U.u2.cout ;
assign \add_3s_3s_3_2_1_U15.top_add_3s_3s_3_2_1_Adder_11_U.fas_s2  = \add_3s_3s_3_2_1_U15.top_add_3s_3s_3_2_1_Adder_11_U.u2.s ;
assign \add_3s_3s_3_2_1_U15.top_add_3s_3s_3_2_1_Adder_11_U.u1.a  = \add_3s_3s_3_2_1_U15.top_add_3s_3s_3_2_1_Adder_11_U.a [0];
assign \add_3s_3s_3_2_1_U15.top_add_3s_3s_3_2_1_Adder_11_U.u1.b  = \add_3s_3s_3_2_1_U15.top_add_3s_3s_3_2_1_Adder_11_U.b [0];
assign \add_3s_3s_3_2_1_U15.top_add_3s_3s_3_2_1_Adder_11_U.u1.cin  = 1'h0;
assign \add_3s_3s_3_2_1_U15.top_add_3s_3s_3_2_1_Adder_11_U.facout_s1  = \add_3s_3s_3_2_1_U15.top_add_3s_3s_3_2_1_Adder_11_U.u1.cout ;
assign \add_3s_3s_3_2_1_U15.top_add_3s_3s_3_2_1_Adder_11_U.fas_s1  = \add_3s_3s_3_2_1_U15.top_add_3s_3s_3_2_1_Adder_11_U.u1.s ;
assign \add_3s_3s_3_2_1_U15.top_add_3s_3s_3_2_1_Adder_11_U.a  = \add_3s_3s_3_2_1_U15.din0 ;
assign \add_3s_3s_3_2_1_U15.top_add_3s_3s_3_2_1_Adder_11_U.b  = \add_3s_3s_3_2_1_U15.din1 ;
assign \add_3s_3s_3_2_1_U15.top_add_3s_3s_3_2_1_Adder_11_U.ce  = \add_3s_3s_3_2_1_U15.ce ;
assign \add_3s_3s_3_2_1_U15.top_add_3s_3s_3_2_1_Adder_11_U.clk  = \add_3s_3s_3_2_1_U15.clk ;
assign \add_3s_3s_3_2_1_U15.top_add_3s_3s_3_2_1_Adder_11_U.reset  = \add_3s_3s_3_2_1_U15.reset ;
assign \add_3s_3s_3_2_1_U15.dout  = \add_3s_3s_3_2_1_U15.top_add_3s_3s_3_2_1_Adder_11_U.s ;
assign \add_3s_3s_3_2_1_U15.ce  = 1'h1;
assign \add_3s_3s_3_2_1_U15.clk  = ap_clk;
assign \add_3s_3s_3_2_1_U15.din0  = { add_ln69_2_reg_1247[1], add_ln69_2_reg_1247 };
assign \add_3s_3s_3_2_1_U15.din1  = { op_7_V_reg_1232[1], op_7_V_reg_1232 };
assign grp_fu_708_p2 = \add_3s_3s_3_2_1_U15.dout ;
assign \add_3s_3s_3_2_1_U15.reset  = ap_rst;
assign \add_36s_36s_36_2_1_U20.top_add_36s_36s_36_2_1_Adder_14_U.ain_s0  = \add_36s_36s_36_2_1_U20.top_add_36s_36s_36_2_1_Adder_14_U.a ;
assign \add_36s_36s_36_2_1_U20.top_add_36s_36s_36_2_1_Adder_14_U.bin_s0  = \add_36s_36s_36_2_1_U20.top_add_36s_36s_36_2_1_Adder_14_U.b ;
assign \add_36s_36s_36_2_1_U20.top_add_36s_36s_36_2_1_Adder_14_U.s  = { \add_36s_36s_36_2_1_U20.top_add_36s_36s_36_2_1_Adder_14_U.fas_s2 , \add_36s_36s_36_2_1_U20.top_add_36s_36s_36_2_1_Adder_14_U.sum_s1  };
assign \add_36s_36s_36_2_1_U20.top_add_36s_36s_36_2_1_Adder_14_U.u2.a  = \add_36s_36s_36_2_1_U20.top_add_36s_36s_36_2_1_Adder_14_U.ain_s1 ;
assign \add_36s_36s_36_2_1_U20.top_add_36s_36s_36_2_1_Adder_14_U.u2.b  = \add_36s_36s_36_2_1_U20.top_add_36s_36s_36_2_1_Adder_14_U.bin_s1 ;
assign \add_36s_36s_36_2_1_U20.top_add_36s_36s_36_2_1_Adder_14_U.u2.cin  = \add_36s_36s_36_2_1_U20.top_add_36s_36s_36_2_1_Adder_14_U.carry_s1 ;
assign \add_36s_36s_36_2_1_U20.top_add_36s_36s_36_2_1_Adder_14_U.facout_s2  = \add_36s_36s_36_2_1_U20.top_add_36s_36s_36_2_1_Adder_14_U.u2.cout ;
assign \add_36s_36s_36_2_1_U20.top_add_36s_36s_36_2_1_Adder_14_U.fas_s2  = \add_36s_36s_36_2_1_U20.top_add_36s_36s_36_2_1_Adder_14_U.u2.s ;
assign \add_36s_36s_36_2_1_U20.top_add_36s_36s_36_2_1_Adder_14_U.u1.a  = \add_36s_36s_36_2_1_U20.top_add_36s_36s_36_2_1_Adder_14_U.a [17:0];
assign \add_36s_36s_36_2_1_U20.top_add_36s_36s_36_2_1_Adder_14_U.u1.b  = \add_36s_36s_36_2_1_U20.top_add_36s_36s_36_2_1_Adder_14_U.b [17:0];
assign \add_36s_36s_36_2_1_U20.top_add_36s_36s_36_2_1_Adder_14_U.u1.cin  = 1'h0;
assign \add_36s_36s_36_2_1_U20.top_add_36s_36s_36_2_1_Adder_14_U.facout_s1  = \add_36s_36s_36_2_1_U20.top_add_36s_36s_36_2_1_Adder_14_U.u1.cout ;
assign \add_36s_36s_36_2_1_U20.top_add_36s_36s_36_2_1_Adder_14_U.fas_s1  = \add_36s_36s_36_2_1_U20.top_add_36s_36s_36_2_1_Adder_14_U.u1.s ;
assign \add_36s_36s_36_2_1_U20.top_add_36s_36s_36_2_1_Adder_14_U.a  = \add_36s_36s_36_2_1_U20.din0 ;
assign \add_36s_36s_36_2_1_U20.top_add_36s_36s_36_2_1_Adder_14_U.b  = \add_36s_36s_36_2_1_U20.din1 ;
assign \add_36s_36s_36_2_1_U20.top_add_36s_36s_36_2_1_Adder_14_U.ce  = \add_36s_36s_36_2_1_U20.ce ;
assign \add_36s_36s_36_2_1_U20.top_add_36s_36s_36_2_1_Adder_14_U.clk  = \add_36s_36s_36_2_1_U20.clk ;
assign \add_36s_36s_36_2_1_U20.top_add_36s_36s_36_2_1_Adder_14_U.reset  = \add_36s_36s_36_2_1_U20.reset ;
assign \add_36s_36s_36_2_1_U20.dout  = \add_36s_36s_36_2_1_U20.top_add_36s_36s_36_2_1_Adder_14_U.s ;
assign \add_36s_36s_36_2_1_U20.ce  = 1'h1;
assign \add_36s_36s_36_2_1_U20.clk  = ap_clk;
assign \add_36s_36s_36_2_1_U20.din0  = { op_28_V_reg_1345[31], op_28_V_reg_1345, 3'h0 };
assign \add_36s_36s_36_2_1_U20.din1  = { op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17 };
assign grp_fu_853_p2 = \add_36s_36s_36_2_1_U20.dout ;
assign \add_36s_36s_36_2_1_U20.reset  = ap_rst;
assign \add_35s_35s_35_2_1_U17.top_add_35s_35s_35_2_1_Adder_12_U.ain_s0  = \add_35s_35s_35_2_1_U17.top_add_35s_35s_35_2_1_Adder_12_U.a ;
assign \add_35s_35s_35_2_1_U17.top_add_35s_35s_35_2_1_Adder_12_U.bin_s0  = \add_35s_35s_35_2_1_U17.top_add_35s_35s_35_2_1_Adder_12_U.b ;
assign \add_35s_35s_35_2_1_U17.top_add_35s_35s_35_2_1_Adder_12_U.s  = { \add_35s_35s_35_2_1_U17.top_add_35s_35s_35_2_1_Adder_12_U.fas_s2 , \add_35s_35s_35_2_1_U17.top_add_35s_35s_35_2_1_Adder_12_U.sum_s1  };
assign \add_35s_35s_35_2_1_U17.top_add_35s_35s_35_2_1_Adder_12_U.u2.a  = \add_35s_35s_35_2_1_U17.top_add_35s_35s_35_2_1_Adder_12_U.ain_s1 ;
assign \add_35s_35s_35_2_1_U17.top_add_35s_35s_35_2_1_Adder_12_U.u2.b  = \add_35s_35s_35_2_1_U17.top_add_35s_35s_35_2_1_Adder_12_U.bin_s1 ;
assign \add_35s_35s_35_2_1_U17.top_add_35s_35s_35_2_1_Adder_12_U.u2.cin  = \add_35s_35s_35_2_1_U17.top_add_35s_35s_35_2_1_Adder_12_U.carry_s1 ;
assign \add_35s_35s_35_2_1_U17.top_add_35s_35s_35_2_1_Adder_12_U.facout_s2  = \add_35s_35s_35_2_1_U17.top_add_35s_35s_35_2_1_Adder_12_U.u2.cout ;
assign \add_35s_35s_35_2_1_U17.top_add_35s_35s_35_2_1_Adder_12_U.fas_s2  = \add_35s_35s_35_2_1_U17.top_add_35s_35s_35_2_1_Adder_12_U.u2.s ;
assign \add_35s_35s_35_2_1_U17.top_add_35s_35s_35_2_1_Adder_12_U.u1.a  = \add_35s_35s_35_2_1_U17.top_add_35s_35s_35_2_1_Adder_12_U.a [16:0];
assign \add_35s_35s_35_2_1_U17.top_add_35s_35s_35_2_1_Adder_12_U.u1.b  = \add_35s_35s_35_2_1_U17.top_add_35s_35s_35_2_1_Adder_12_U.b [16:0];
assign \add_35s_35s_35_2_1_U17.top_add_35s_35s_35_2_1_Adder_12_U.u1.cin  = 1'h0;
assign \add_35s_35s_35_2_1_U17.top_add_35s_35s_35_2_1_Adder_12_U.facout_s1  = \add_35s_35s_35_2_1_U17.top_add_35s_35s_35_2_1_Adder_12_U.u1.cout ;
assign \add_35s_35s_35_2_1_U17.top_add_35s_35s_35_2_1_Adder_12_U.fas_s1  = \add_35s_35s_35_2_1_U17.top_add_35s_35s_35_2_1_Adder_12_U.u1.s ;
assign \add_35s_35s_35_2_1_U17.top_add_35s_35s_35_2_1_Adder_12_U.a  = \add_35s_35s_35_2_1_U17.din0 ;
assign \add_35s_35s_35_2_1_U17.top_add_35s_35s_35_2_1_Adder_12_U.b  = \add_35s_35s_35_2_1_U17.din1 ;
assign \add_35s_35s_35_2_1_U17.top_add_35s_35s_35_2_1_Adder_12_U.ce  = \add_35s_35s_35_2_1_U17.ce ;
assign \add_35s_35s_35_2_1_U17.top_add_35s_35s_35_2_1_Adder_12_U.clk  = \add_35s_35s_35_2_1_U17.clk ;
assign \add_35s_35s_35_2_1_U17.top_add_35s_35s_35_2_1_Adder_12_U.reset  = \add_35s_35s_35_2_1_U17.reset ;
assign \add_35s_35s_35_2_1_U17.dout  = \add_35s_35s_35_2_1_U17.top_add_35s_35s_35_2_1_Adder_12_U.s ;
assign \add_35s_35s_35_2_1_U17.ce  = 1'h1;
assign \add_35s_35s_35_2_1_U17.clk  = ap_clk;
assign \add_35s_35s_35_2_1_U17.din0  = { op_26_V_reg_1282[6], op_26_V_reg_1282[6], op_26_V_reg_1282[6], op_26_V_reg_1282[6], op_26_V_reg_1282[6], op_26_V_reg_1282[6], op_26_V_reg_1282[6], op_26_V_reg_1282[6], op_26_V_reg_1282[6], op_26_V_reg_1282[6], op_26_V_reg_1282[6], op_26_V_reg_1282[6], op_26_V_reg_1282[6], op_26_V_reg_1282[6], op_26_V_reg_1282[6], op_26_V_reg_1282[6], op_26_V_reg_1282[6], op_26_V_reg_1282[6], op_26_V_reg_1282[6], op_26_V_reg_1282[6], op_26_V_reg_1282[6], op_26_V_reg_1282[6], op_26_V_reg_1282[6], op_26_V_reg_1282[6], op_26_V_reg_1282[6], op_26_V_reg_1282[6], op_26_V_reg_1282, 2'h0 };
assign \add_35s_35s_35_2_1_U17.din1  = { op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15 };
assign grp_fu_737_p2 = \add_35s_35s_35_2_1_U17.dout ;
assign \add_35s_35s_35_2_1_U17.reset  = ap_rst;
assign \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_15_U.ain_s0  = \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_15_U.a ;
assign \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_15_U.bin_s0  = \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_15_U.b ;
assign \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_15_U.s  = { \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_15_U.fas_s2 , \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_15_U.sum_s1  };
assign \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_15_U.u2.a  = \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_15_U.ain_s1 ;
assign \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_15_U.u2.b  = \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_15_U.bin_s1 ;
assign \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_15_U.u2.cin  = \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_15_U.carry_s1 ;
assign \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_15_U.facout_s2  = \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_15_U.u2.cout ;
assign \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_15_U.fas_s2  = \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_15_U.u2.s ;
assign \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_15_U.u1.a  = \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_15_U.a [15:0];
assign \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_15_U.u1.b  = \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_15_U.b [15:0];
assign \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_15_U.u1.cin  = 1'h0;
assign \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_15_U.facout_s1  = \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_15_U.u1.cout ;
assign \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_15_U.fas_s1  = \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_15_U.u1.s ;
assign \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_15_U.a  = \add_32ns_32s_32_2_1_U23.din0 ;
assign \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_15_U.b  = \add_32ns_32s_32_2_1_U23.din1 ;
assign \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_15_U.ce  = \add_32ns_32s_32_2_1_U23.ce ;
assign \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_15_U.clk  = \add_32ns_32s_32_2_1_U23.clk ;
assign \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_15_U.reset  = \add_32ns_32s_32_2_1_U23.reset ;
assign \add_32ns_32s_32_2_1_U23.dout  = \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_15_U.s ;
assign \add_32ns_32s_32_2_1_U23.ce  = 1'h1;
assign \add_32ns_32s_32_2_1_U23.clk  = ap_clk;
assign \add_32ns_32s_32_2_1_U23.din0  = ret_V_28_reg_1392;
assign \add_32ns_32s_32_2_1_U23.din1  = { op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19 };
assign grp_fu_916_p2 = \add_32ns_32s_32_2_1_U23.dout ;
assign \add_32ns_32s_32_2_1_U23.reset  = ap_rst;
assign \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_15_U.ain_s0  = \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_15_U.a ;
assign \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_15_U.bin_s0  = \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_15_U.b ;
assign \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_15_U.s  = { \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_15_U.fas_s2 , \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_15_U.sum_s1  };
assign \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_15_U.u2.a  = \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_15_U.ain_s1 ;
assign \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_15_U.u2.b  = \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_15_U.bin_s1 ;
assign \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_15_U.u2.cin  = \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_15_U.carry_s1 ;
assign \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_15_U.facout_s2  = \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_15_U.u2.cout ;
assign \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_15_U.fas_s2  = \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_15_U.u2.s ;
assign \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_15_U.u1.a  = \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_15_U.a [15:0];
assign \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_15_U.u1.b  = \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_15_U.b [15:0];
assign \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_15_U.u1.cin  = 1'h0;
assign \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_15_U.facout_s1  = \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_15_U.u1.cout ;
assign \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_15_U.fas_s1  = \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_15_U.u1.s ;
assign \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_15_U.a  = \add_32ns_32s_32_2_1_U22.din0 ;
assign \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_15_U.b  = \add_32ns_32s_32_2_1_U22.din1 ;
assign \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_15_U.ce  = \add_32ns_32s_32_2_1_U22.ce ;
assign \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_15_U.clk  = \add_32ns_32s_32_2_1_U22.clk ;
assign \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_15_U.reset  = \add_32ns_32s_32_2_1_U22.reset ;
assign \add_32ns_32s_32_2_1_U22.dout  = \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_15_U.s ;
assign \add_32ns_32s_32_2_1_U22.ce  = 1'h1;
assign \add_32ns_32s_32_2_1_U22.clk  = ap_clk;
assign \add_32ns_32s_32_2_1_U22.din0  = ret_V_27_reg_1382;
assign \add_32ns_32s_32_2_1_U22.din1  = { op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18 };
assign grp_fu_907_p2 = \add_32ns_32s_32_2_1_U22.dout ;
assign \add_32ns_32s_32_2_1_U22.reset  = ap_rst;
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_13_U.ain_s0  = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_13_U.a ;
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_13_U.bin_s0  = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_13_U.b ;
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_13_U.s  = { \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_13_U.fas_s2 , \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_13_U.sum_s1  };
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_13_U.u2.a  = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_13_U.ain_s1 ;
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_13_U.u2.b  = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_13_U.bin_s1 ;
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_13_U.u2.cin  = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_13_U.carry_s1 ;
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_13_U.facout_s2  = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_13_U.u2.cout ;
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_13_U.fas_s2  = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_13_U.u2.s ;
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_13_U.u1.a  = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_13_U.a [15:0];
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_13_U.u1.b  = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_13_U.b [15:0];
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_13_U.u1.cin  = 1'h0;
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_13_U.facout_s1  = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_13_U.u1.cout ;
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_13_U.fas_s1  = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_13_U.u1.s ;
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_13_U.a  = \add_32ns_32ns_32_2_1_U21.din0 ;
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_13_U.b  = \add_32ns_32ns_32_2_1_U21.din1 ;
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_13_U.ce  = \add_32ns_32ns_32_2_1_U21.ce ;
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_13_U.clk  = \add_32ns_32ns_32_2_1_U21.clk ;
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_13_U.reset  = \add_32ns_32ns_32_2_1_U21.reset ;
assign \add_32ns_32ns_32_2_1_U21.dout  = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_13_U.s ;
assign \add_32ns_32ns_32_2_1_U21.ce  = 1'h1;
assign \add_32ns_32ns_32_2_1_U21.clk  = ap_clk;
assign \add_32ns_32ns_32_2_1_U21.din0  = ret_V_31_cast_reg_1370;
assign \add_32ns_32ns_32_2_1_U21.din1  = 32'd1;
assign grp_fu_879_p2 = \add_32ns_32ns_32_2_1_U21.dout ;
assign \add_32ns_32ns_32_2_1_U21.reset  = ap_rst;
assign \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_13_U.ain_s0  = \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_13_U.a ;
assign \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_13_U.bin_s0  = \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_13_U.b ;
assign \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_13_U.s  = { \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_13_U.fas_s2 , \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_13_U.sum_s1  };
assign \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_13_U.u2.a  = \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_13_U.ain_s1 ;
assign \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_13_U.u2.b  = \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_13_U.bin_s1 ;
assign \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_13_U.u2.cin  = \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_13_U.carry_s1 ;
assign \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_13_U.facout_s2  = \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_13_U.u2.cout ;
assign \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_13_U.fas_s2  = \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_13_U.u2.s ;
assign \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_13_U.u1.a  = \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_13_U.a [15:0];
assign \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_13_U.u1.b  = \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_13_U.b [15:0];
assign \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_13_U.u1.cin  = 1'h0;
assign \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_13_U.facout_s1  = \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_13_U.u1.cout ;
assign \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_13_U.fas_s1  = \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_13_U.u1.s ;
assign \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_13_U.a  = \add_32ns_32ns_32_2_1_U19.din0 ;
assign \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_13_U.b  = \add_32ns_32ns_32_2_1_U19.din1 ;
assign \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_13_U.ce  = \add_32ns_32ns_32_2_1_U19.ce ;
assign \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_13_U.clk  = \add_32ns_32ns_32_2_1_U19.clk ;
assign \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_13_U.reset  = \add_32ns_32ns_32_2_1_U19.reset ;
assign \add_32ns_32ns_32_2_1_U19.dout  = \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_13_U.s ;
assign \add_32ns_32ns_32_2_1_U19.ce  = 1'h1;
assign \add_32ns_32ns_32_2_1_U19.clk  = ap_clk;
assign \add_32ns_32ns_32_2_1_U19.din0  = ret_V_25_reg_1335;
assign \add_32ns_32ns_32_2_1_U19.din1  = select_ln69_1_reg_1340;
assign grp_fu_834_p2 = \add_32ns_32ns_32_2_1_U19.dout ;
assign \add_32ns_32ns_32_2_1_U19.reset  = ap_rst;
assign \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_13_U.ain_s0  = \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_13_U.a ;
assign \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_13_U.bin_s0  = \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_13_U.b ;
assign \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_13_U.s  = { \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_13_U.fas_s2 , \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_13_U.sum_s1  };
assign \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_13_U.u2.a  = \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_13_U.ain_s1 ;
assign \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_13_U.u2.b  = \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_13_U.bin_s1 ;
assign \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_13_U.u2.cin  = \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_13_U.carry_s1 ;
assign \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_13_U.facout_s2  = \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_13_U.u2.cout ;
assign \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_13_U.fas_s2  = \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_13_U.u2.s ;
assign \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_13_U.u1.a  = \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_13_U.a [15:0];
assign \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_13_U.u1.b  = \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_13_U.b [15:0];
assign \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_13_U.u1.cin  = 1'h0;
assign \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_13_U.facout_s1  = \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_13_U.u1.cout ;
assign \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_13_U.fas_s1  = \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_13_U.u1.s ;
assign \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_13_U.a  = \add_32ns_32ns_32_2_1_U18.din0 ;
assign \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_13_U.b  = \add_32ns_32ns_32_2_1_U18.din1 ;
assign \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_13_U.ce  = \add_32ns_32ns_32_2_1_U18.ce ;
assign \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_13_U.clk  = \add_32ns_32ns_32_2_1_U18.clk ;
assign \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_13_U.reset  = \add_32ns_32ns_32_2_1_U18.reset ;
assign \add_32ns_32ns_32_2_1_U18.dout  = \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_13_U.s ;
assign \add_32ns_32ns_32_2_1_U18.ce  = 1'h1;
assign \add_32ns_32ns_32_2_1_U18.clk  = ap_clk;
assign \add_32ns_32ns_32_2_1_U18.din0  = ret_V_29_cast_reg_1307;
assign \add_32ns_32ns_32_2_1_U18.din1  = 32'd1;
assign grp_fu_772_p2 = \add_32ns_32ns_32_2_1_U18.dout ;
assign \add_32ns_32ns_32_2_1_U18.reset  = ap_rst;
assign \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.ain_s0  = \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.a ;
assign \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.bin_s0  = \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.b ;
assign \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.s  = { \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.fas_s2 , \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.sum_s1  };
assign \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.u2.a  = \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.ain_s1 ;
assign \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.u2.b  = \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.bin_s1 ;
assign \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.u2.cin  = \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.carry_s1 ;
assign \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.facout_s2  = \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.u2.cout ;
assign \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.fas_s2  = \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.u2.s ;
assign \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.u1.a  = \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.a [0];
assign \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.u1.b  = \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.b [0];
assign \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.u1.cin  = 1'h0;
assign \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.facout_s1  = \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.u1.cout ;
assign \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.fas_s1  = \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.u1.s ;
assign \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.a  = \add_2ns_2ns_2_2_1_U9.din0 ;
assign \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.b  = \add_2ns_2ns_2_2_1_U9.din1 ;
assign \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.ce  = \add_2ns_2ns_2_2_1_U9.ce ;
assign \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.clk  = \add_2ns_2ns_2_2_1_U9.clk ;
assign \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.reset  = \add_2ns_2ns_2_2_1_U9.reset ;
assign \add_2ns_2ns_2_2_1_U9.dout  = \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.s ;
assign \add_2ns_2ns_2_2_1_U9.ce  = 1'h1;
assign \add_2ns_2ns_2_2_1_U9.clk  = ap_clk;
assign \add_2ns_2ns_2_2_1_U9.din0  = { 1'h0, and_ln410_reg_1124 };
assign \add_2ns_2ns_2_2_1_U9.din1  = select_ln708_reg_1119;
assign grp_fu_553_p2 = \add_2ns_2ns_2_2_1_U9.dout ;
assign \add_2ns_2ns_2_2_1_U9.reset  = ap_rst;
assign \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_6_U.ain_s0  = \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_6_U.a ;
assign \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_6_U.bin_s0  = \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_6_U.b ;
assign \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_6_U.s  = { \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_6_U.fas_s2 , \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_6_U.sum_s1  };
assign \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_6_U.u2.a  = \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_6_U.ain_s1 ;
assign \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_6_U.u2.b  = \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_6_U.bin_s1 ;
assign \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_6_U.u2.cin  = \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_6_U.carry_s1 ;
assign \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_6_U.facout_s2  = \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_6_U.u2.cout ;
assign \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_6_U.fas_s2  = \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_6_U.u2.s ;
assign \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_6_U.u1.a  = \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_6_U.a [0];
assign \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_6_U.u1.b  = \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_6_U.b [0];
assign \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_6_U.u1.cin  = 1'h0;
assign \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_6_U.facout_s1  = \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_6_U.u1.cout ;
assign \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_6_U.fas_s1  = \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_6_U.u1.s ;
assign \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_6_U.a  = \add_2ns_2ns_2_2_1_U13.din0 ;
assign \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_6_U.b  = \add_2ns_2ns_2_2_1_U13.din1 ;
assign \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_6_U.ce  = \add_2ns_2ns_2_2_1_U13.ce ;
assign \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_6_U.clk  = \add_2ns_2ns_2_2_1_U13.clk ;
assign \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_6_U.reset  = \add_2ns_2ns_2_2_1_U13.reset ;
assign \add_2ns_2ns_2_2_1_U13.dout  = \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_6_U.s ;
assign \add_2ns_2ns_2_2_1_U13.ce  = 1'h1;
assign \add_2ns_2ns_2_2_1_U13.clk  = ap_clk;
assign \add_2ns_2ns_2_2_1_U13.din0  = select_ln69_reg_1197;
assign \add_2ns_2ns_2_2_1_U13.din1  = { 1'h0, icmp_ln1494_reg_1192 };
assign grp_fu_683_p2 = \add_2ns_2ns_2_2_1_U13.dout ;
assign \add_2ns_2ns_2_2_1_U13.reset  = ap_rst;
endmodule


// Machine B:
// Processed by function `add_clk_enable_signal` in `verilog_tricks.py`.
// Processed by function `remove_reset_signal` in `verilog_tricks.py`.
module top_B (
  ap_clk,
  ap_start,
  ap_done,
  ap_idle,
  ap_ready,
  op_0,
  op_1,
  op_3,
  op_4,
  op_11,
  op_12,
  op_15,
  op_17,
  op_18,
  op_19,
  op_31,
  op_31_ap_vld,
clk_enable
);
input clk_enable;


input ap_clk;
wire ap_rst;
assign ap_rst = op_31_ap_vld;
input ap_start;
input [7:0] op_0;
input [3:0] op_1;
input [3:0] op_11;
input [3:0] op_12;
input [3:0] op_15;
input [3:0] op_17;
input [1:0] op_18;
input [3:0] op_19;
input op_3;
input [1:0] op_4;
output ap_done;
output ap_idle;
output ap_ready;
output [31:0] op_31;
output op_31_ap_vld;


reg [1:0] add_ln69_2_reg_1046;
reg [2:0] add_ln69_3_reg_1061;
reg [5:0] add_ln69_reg_1056;
reg [9:0] ap_CS_fsm = 10'h001;
reg icmp_ln851_2_reg_1083;
reg icmp_ln851_3_reg_1110;
reg icmp_ln851_reg_1036;
reg isNeg_reg_1004;
reg [6:0] op_26_V_reg_1066;
reg [31:0] op_28_V_reg_1093;
reg [1:0] op_6_V_reg_1014;
reg [3:0] op_8_V_reg_996;
reg [8:0] ret_V_19_reg_1024;
reg [6:0] ret_V_23_reg_1051;
reg [34:0] ret_V_24_reg_1071;
reg [35:0] ret_V_26_reg_1098;
reg [31:0] ret_V_27_reg_1115;
reg [31:0] ret_V_29_cast_reg_1076;
reg [31:0] ret_V_31_cast_reg_1103;
reg [5:0] ret_V_reg_1029;
reg select_ln13_reg_982;
reg [31:0] select_ln69_1_reg_1088;
reg [26:0] sub_ln1118_reg_1041;
reg [1:0] sub_ln69_reg_1019;
reg [1:0] ush_reg_1009;
wire [1:0] _000_;
wire [2:0] _001_;
wire [5:0] _002_;
wire [9:0] _003_;
wire _004_;
wire _005_;
wire _006_;
wire _007_;
wire [6:0] _008_;
wire [31:0] _009_;
wire [1:0] _010_;
wire [3:0] _011_;
wire [8:0] _012_;
wire [6:0] _013_;
wire [34:0] _014_;
wire [35:0] _015_;
wire [31:0] _016_;
wire [31:0] _017_;
wire [31:0] _018_;
wire [5:0] _019_;
wire _020_;
wire [31:0] _021_;
wire [2:0] _022_;
wire [1:0] _023_;
wire [1:0] _024_;
wire [1:0] _025_;
wire _026_;
wire _027_;
wire _028_;
wire _029_;
wire _030_;
wire _031_;
wire _032_;
wire _033_;
wire _034_;
wire _035_;
wire _036_;
wire _037_;
wire _038_;
wire _039_;
wire _040_;
wire _041_;
wire _042_;
wire _043_;
wire _044_;
wire _045_;
wire _046_;
wire _047_;
wire _048_;
wire [31:0] add_ln691_1_fu_936_p2;
wire [31:0] add_ln691_fu_865_p2;
wire [6:0] add_ln69_1_fu_752_p2;
wire [1:0] add_ln69_2_fu_612_p2;
wire [2:0] add_ln69_3_fu_743_p2;
wire [5:0] add_ln69_fu_734_p2;
wire and_ln410_fu_458_p2;
wire and_ln850_1_fu_588_p2;
wire and_ln850_fu_797_p2;
wire ap_CS_fsm_state1;
wire ap_CS_fsm_state10;
wire ap_CS_fsm_state2;
wire ap_CS_fsm_state3;
wire ap_CS_fsm_state4;
wire ap_CS_fsm_state5;
wire ap_CS_fsm_state6;
wire ap_CS_fsm_state7;
wire ap_CS_fsm_state8;
wire ap_CS_fsm_state9;
wire [9:0] ap_NS_fsm;
wire ap_clk;
wire ap_done;
wire ap_idle;
wire ap_ready;
wire ap_rst;
wire ap_start;
wire [3:0] ashr_ln1297_fu_545_p2;
wire [31:0] ashr_ln1497_1_fu_344_p2;
wire [1:0] conv_i389_fu_311_p0;
wire [31:0] conv_i389_fu_311_p1;
wire icmp_ln1494_fu_536_p2;
wire icmp_ln768_fu_258_p2;
wire icmp_ln850_1_fu_582_p2;
wire icmp_ln850_fu_791_p2;
wire icmp_ln851_1_fu_681_p2;
wire icmp_ln851_2_fu_844_p2;
wire icmp_ln851_3_fu_923_p2;
wire icmp_ln851_fu_503_p2;
wire isNeg_fu_369_p3;
wire [7:0] op_0;
wire [3:0] op_1;
wire [3:0] op_11;
wire [3:0] op_12;
wire [3:0] op_15;
wire [3:0] op_17;
wire [1:0] op_18;
wire [3:0] op_19;
wire [6:0] op_26_V_fu_760_p2;
wire [31:0] op_28_V_fu_883_p2;
wire op_3;
wire [31:0] op_31;
wire op_31_ap_vld;
wire op_3_read_read_fu_130_p2;
wire [1:0] op_4;
wire [1:0] op_6_V_fu_468_p2;
wire op_7_V_fu_618_p0;
wire [1:0] op_7_V_fu_618_p3;
wire [3:0] op_8_V_fu_296_p3;
wire or_ln384_fu_290_p2;
wire or_ln410_fu_452_p2;
wire or_ln785_fu_264_p2;
wire overflow_fu_276_p2;
wire p_Result_1_fu_669_p3;
wire p_Result_2_fu_779_p3;
wire p_Result_3_fu_570_p3;
wire p_Result_4_fu_858_p3;
wire p_Result_5_fu_929_p3;
wire p_Result_6_fu_420_p3;
wire p_Result_7_fu_222_p3;
wire p_Result_8_fu_242_p2;
wire p_Result_s_14_fu_624_p3;
wire [1:0] p_Result_s_fu_248_p4;
wire [3:0] p_Val2_2_fu_234_p3;
wire [1:0] r_2_fu_365_p1;
wire [3:0] r_V_1_fu_555_p3;
wire r_V_fu_649_p0;
wire [26:0] r_V_fu_649_p3;
wire r_fu_432_p2;
wire ret_V_11_fu_562_p3;
wire ret_V_12_fu_594_p2;
wire [3:0] ret_V_18_fu_398_p2;
wire [8:0] ret_V_19_fu_483_p2;
wire [5:0] ret_V_20_fu_642_p3;
wire [3:0] ret_V_21_fu_701_p3;
wire [3:0] ret_V_22_fu_766_p2;
wire [6:0] ret_V_23_fu_716_p2;
wire [34:0] ret_V_24_fu_824_p2;
wire [31:0] ret_V_25_fu_876_p3;
wire [35:0] ret_V_26_fu_903_p2;
wire [31:0] ret_V_27_fu_947_p3;
wire [31:0] ret_V_28_fu_958_p2;
wire [5:0] ret_V_3_fu_631_p2;
wire [3:0] ret_V_5_fu_687_p2;
wire ret_V_8_fu_771_p3;
wire ret_V_9_fu_803_p2;
wire [2:0] ret_fu_216_p2;
wire [34:0] rhs_4_fu_892_p3;
wire rhs_fu_391_p1;
wire [3:0] rhs_fu_391_p3;
wire select_ln1347_fu_205_p0;
wire [2:0] select_ln1347_fu_205_p3;
wire select_ln13_fu_197_p0;
wire select_ln13_fu_197_p3;
wire [1:0] select_ln1497_1_fu_336_p3;
wire [1:0] select_ln1497_2_fu_350_p3;
wire [31:0] select_ln1497_3_fu_357_p3;
wire [1:0] select_ln1497_fu_321_p3;
wire [3:0] select_ln384_fu_282_p3;
wire [31:0] select_ln69_1_fu_850_p3;
wire [1:0] select_ln69_fu_604_p3;
wire [1:0] select_ln708_fu_412_p3;
wire select_ln835_fu_304_p3;
wire [3:0] select_ln850_2_fu_693_p3;
wire [31:0] select_ln850_3_fu_870_p3;
wire [31:0] select_ln850_4_fu_941_p3;
wire [5:0] select_ln850_fu_636_p3;
wire [26:0] sext_ln1118_fu_516_p1;
wire [6:0] sext_ln1192_1_fu_712_p1;
wire [34:0] sext_ln1192_2_fu_820_p1;
wire [35:0] sext_ln1192_3_fu_899_p1;
wire [31:0] sext_ln1192_4_fu_954_p1;
wire [6:0] sext_ln1192_fu_709_p1;
wire [1:0] sext_ln1347_fu_212_p0;
wire [2:0] sext_ln1347_fu_212_p1;
wire [4:0] sext_ln1494_fu_533_p1;
wire [5:0] sext_ln69_1_fu_726_p1;
wire [6:0] sext_ln69_2_fu_749_p1;
wire [31:0] sext_ln69_4_fu_963_p1;
wire [2:0] sext_ln69_5_fu_740_p1;
wire [6:0] sext_ln69_6_fu_757_p1;
wire [2:0] sext_ln69_fu_722_p1;
wire [3:0] sext_ln703_1_fu_809_p0;
wire [34:0] sext_ln703_1_fu_809_p1;
wire [3:0] sext_ln703_2_fu_888_p0;
wire [35:0] sext_ln703_2_fu_888_p1;
wire [8:0] sext_ln703_fu_479_p1;
wire [3:0] sext_ln850_fu_665_p1;
wire [3:0] shl_ln1358_fu_550_p2;
wire [30:0] shl_ln1497_1_fu_315_p2;
wire [1:0] shl_ln1_fu_526_p1;
wire [4:0] shl_ln1_fu_526_p3;
wire [1:0] shl_ln_fu_509_p1;
wire [25:0] shl_ln_fu_509_p3;
wire [26:0] sub_ln1118_fu_520_p2;
wire [1:0] sub_ln1357_fu_377_p2;
wire [1:0] sub_ln69_fu_474_p1;
wire [1:0] sub_ln69_fu_474_p2;
wire [8:0] tmp_14_fu_813_p3;
wire [2:0] tmp_2_fu_655_p4;
wire tmp_3_fu_438_p3;
wire [1:0] tmp_7_fu_328_p1;
wire tmp_7_fu_328_p3;
wire tmp_fu_404_p3;
wire [1:0] trunc_ln718_fu_428_p1;
wire trunc_ln728_fu_230_p1;
wire [23:0] trunc_ln851_1_fu_677_p1;
wire [2:0] trunc_ln851_2_fu_787_p1;
wire [2:0] trunc_ln851_3_fu_578_p1;
wire [3:0] trunc_ln851_4_fu_840_p0;
wire [1:0] trunc_ln851_4_fu_840_p1;
wire [3:0] trunc_ln851_5_fu_919_p0;
wire [2:0] trunc_ln851_5_fu_919_p1;
wire [2:0] trunc_ln851_fu_499_p1;
wire [1:0] ush_fu_383_p3;
wire xor_ln410_fu_446_p2;
wire xor_ln785_fu_270_p2;
wire [3:0] zext_ln1357_fu_542_p1;
wire [1:0] zext_ln415_fu_464_p1;
wire [1:0] zext_ln69_1_fu_600_p1;
wire [5:0] zext_ln69_fu_730_p1;


assign add_ln691_1_fu_936_p2 = ret_V_31_cast_reg_1103 + 1'h1;
assign add_ln691_fu_865_p2 = ret_V_29_cast_reg_1076 + 1'h1;
assign add_ln69_1_fu_752_p2 = $signed(add_ln69_reg_1056) + $signed(ret_V_23_reg_1051);
assign add_ln69_2_fu_612_p2 = select_ln69_fu_604_p3 + icmp_ln1494_fu_536_p2;
assign add_ln69_3_fu_743_p2 = $signed(add_ln69_2_reg_1046) + $signed(op_7_V_fu_618_p3);
assign add_ln69_fu_734_p2 = $signed(ret_V_21_fu_701_p3) + $signed({ 1'h0, op_12 });
assign op_26_V_fu_760_p2 = $signed(add_ln69_3_reg_1061) + $signed(add_ln69_1_fu_752_p2);
assign op_28_V_fu_883_p2 = ret_V_25_fu_876_p3 + select_ln69_1_reg_1088;
assign op_31 = $signed(ret_V_28_fu_958_p2) + $signed(op_19);
assign op_6_V_fu_468_p2 = and_ln410_fu_458_p2 + select_ln708_fu_412_p3;
assign ret_V_19_fu_483_p2 = $signed(op_0) + $signed(5'h08);
assign ret_V_23_fu_716_p2 = $signed(ret_V_20_fu_642_p3) + $signed(op_6_V_reg_1014);
assign { ret_V_24_fu_824_p2[34], ret_V_24_fu_824_p2[8:0] } = $signed({ op_26_V_reg_1066, 2'h0 }) + $signed(op_15);
assign ret_V_26_fu_903_p2 = $signed({ op_28_V_reg_1093, 3'h0 }) + $signed(op_17);
assign ret_V_28_fu_958_p2 = $signed(ret_V_27_reg_1115) + $signed(op_18);
assign ret_V_3_fu_631_p2 = ret_V_reg_1029 + 1'h1;
assign ret_V_5_fu_687_p2 = $signed(r_V_fu_649_p3[26:24]) + $signed(2'h1);
assign _026_ = op_3 & ap_CS_fsm[2];
assign _027_ = ap_CS_fsm[0] & _029_;
assign _028_ = ap_CS_fsm[0] & ap_start;
assign and_ln410_fu_458_p2 = op_1[2] & or_ln410_fu_452_p2;
assign and_ln850_1_fu_588_p2 = r_V_1_fu_555_p3[3] & icmp_ln850_1_fu_582_p2;
assign and_ln850_fu_797_p2 = ret_V_22_fu_766_p2[3] & icmp_ln850_fu_791_p2;
assign overflow_fu_276_p2 = xor_ln785_fu_270_p2 & or_ln785_fu_264_p2;
assign xor_ln410_fu_446_p2 = ~ ret_V_18_fu_398_p2[3];
assign xor_ln785_fu_270_p2 = ~ ret_fu_216_p2[2];
assign _029_ = ~ ap_start;
assign _030_ = ! r_V_fu_649_p3[23:0];
assign _031_ = ! ret_V_19_fu_483_p2[2:0];
assign _032_ = $signed({ op_4, 3'h0 }) > $signed(op_8_V_reg_996);
assign _033_ = | ret_fu_216_p2[2:1];
assign _034_ = | r_V_1_fu_555_p3[2:0];
assign _035_ = | ret_V_22_fu_766_p2[2:0];
assign _036_ = | op_15[1:0];
assign _037_ = | op_17[2:0];
assign _038_ = | ret_V_18_fu_398_p2[1:0];
assign or_ln384_fu_290_p2 = ret_fu_216_p2[2] | overflow_fu_276_p2;
assign or_ln410_fu_452_p2 = xor_ln410_fu_446_p2 | r_fu_432_p2;
assign or_ln785_fu_264_p2 = p_Result_8_fu_242_p2 | icmp_ln768_fu_258_p2;
assign ret_V_18_fu_398_p2 = { op_3, 3'h0 } | op_1;
assign ret_V_22_fu_766_p2 = op_8_V_reg_996 | op_11;
always @(posedge ap_clk)
sub_ln1118_reg_1041[23:0] <= 24'h000000;
always @(posedge ap_clk)
sub_ln69_reg_1019 <= _023_;
always @(posedge ap_clk)
sub_ln1118_reg_1041[26:24] <= _022_;
always @(posedge ap_clk)
select_ln13_reg_982 <= _020_;
always @(posedge ap_clk)
ret_V_27_reg_1115 <= _016_;
always @(posedge ap_clk)
op_28_V_reg_1093 <= _009_;
always @(posedge ap_clk)
op_26_V_reg_1066 <= _008_;
always @(posedge ap_clk)
op_8_V_reg_996 <= _011_;
always @(posedge ap_clk)
isNeg_reg_1004 <= _007_;
always @(posedge ap_clk)
ush_reg_1009 <= _024_;
always @(posedge ap_clk)
ret_V_26_reg_1098 <= _015_;
always @(posedge ap_clk)
ret_V_31_cast_reg_1103 <= _018_;
always @(posedge ap_clk)
icmp_ln851_3_reg_1110 <= _005_;
always @(posedge ap_clk)
ret_V_24_reg_1071 <= _014_;
always @(posedge ap_clk)
ret_V_29_cast_reg_1076 <= _017_;
always @(posedge ap_clk)
icmp_ln851_2_reg_1083 <= _004_;
always @(posedge ap_clk)
select_ln69_1_reg_1088 <= _021_;
always @(posedge ap_clk)
ret_V_23_reg_1051 <= _013_;
always @(posedge ap_clk)
add_ln69_reg_1056 <= _002_;
always @(posedge ap_clk)
add_ln69_3_reg_1061 <= _001_;
always @(posedge ap_clk)
op_6_V_reg_1014 <= _010_;
always @(posedge ap_clk)
ret_V_19_reg_1024 <= _012_;
always @(posedge ap_clk)
ret_V_reg_1029 <= _019_;
always @(posedge ap_clk)
icmp_ln851_reg_1036 <= _006_;
always @(posedge ap_clk)
add_ln69_2_reg_1046 <= _000_;
always @(posedge ap_clk)
ap_CS_fsm <= _003_;
assign _025_ = _028_ ? 2'h2 : 2'h1;
assign _039_ = ap_CS_fsm == 1'h1;
function [9:0] _118_;
input [9:0] a;
input [99:0] b;
input [9:0] s;
case (s)
10'b0000000001:
_118_ = b[9:0];
10'b0000000010:
_118_ = b[19:10];
10'b0000000100:
_118_ = b[29:20];
10'b0000001000:
_118_ = b[39:30];
10'b0000010000:
_118_ = b[49:40];
10'b0000100000:
_118_ = b[59:50];
10'b0001000000:
_118_ = b[69:60];
10'b0010000000:
_118_ = b[79:70];
10'b0100000000:
_118_ = b[89:80];
10'b1000000000:
_118_ = b[99:90];
10'b0000000000:
_118_ = a;
default:
_118_ = 10'bx;
endcase
endfunction
assign ap_NS_fsm = _118_(10'hxxx, { 8'h00, _025_, 90'h00402010080402010080001 }, { _039_, _048_, _047_, _046_, _045_, _044_, _043_, _042_, _041_, _040_ });
assign _040_ = ap_CS_fsm == 10'h200;
assign _041_ = ap_CS_fsm == 9'h100;
assign _042_ = ap_CS_fsm == 8'h80;
assign _043_ = ap_CS_fsm == 7'h40;
assign _044_ = ap_CS_fsm == 6'h20;
assign _045_ = ap_CS_fsm == 5'h10;
assign _046_ = ap_CS_fsm == 4'h8;
assign _047_ = ap_CS_fsm == 3'h4;
assign _048_ = ap_CS_fsm == 2'h2;
assign op_31_ap_vld = ap_CS_fsm[9] ? 1'h1 : 1'h0;
assign ap_idle = _027_ ? 1'h1 : 1'h0;
assign _022_ = _026_ ? sub_ln1118_fu_520_p2[26:24] : sub_ln1118_reg_1041[26:24];
assign _023_ = _026_ ? sub_ln69_fu_474_p2 : sub_ln69_reg_1019;
assign _020_ = ap_CS_fsm[0] ? select_ln13_fu_197_p3 : select_ln13_reg_982;
assign _016_ = ap_CS_fsm[8] ? ret_V_27_fu_947_p3 : ret_V_27_reg_1115;
assign _009_ = ap_CS_fsm[6] ? op_28_V_fu_883_p2 : op_28_V_reg_1093;
assign _008_ = ap_CS_fsm[4] ? op_26_V_fu_760_p2 : op_26_V_reg_1066;
assign _024_ = ap_CS_fsm[1] ? ush_fu_383_p3 : ush_reg_1009;
assign _007_ = ap_CS_fsm[1] ? r_2_fu_365_p1[1] : isNeg_reg_1004;
assign _011_ = ap_CS_fsm[1] ? op_8_V_fu_296_p3 : op_8_V_reg_996;
assign _005_ = ap_CS_fsm[7] ? icmp_ln851_3_fu_923_p2 : icmp_ln851_3_reg_1110;
assign _018_ = ap_CS_fsm[7] ? ret_V_26_fu_903_p2[34:3] : ret_V_31_cast_reg_1103;
assign _015_ = ap_CS_fsm[7] ? ret_V_26_fu_903_p2 : ret_V_26_reg_1098;
assign _021_ = ap_CS_fsm[5] ? select_ln69_1_fu_850_p3 : select_ln69_1_reg_1088;
assign _004_ = ap_CS_fsm[5] ? icmp_ln851_2_fu_844_p2 : icmp_ln851_2_reg_1083;
assign _017_ = ap_CS_fsm[5] ? { ret_V_24_fu_824_p2[34], ret_V_24_fu_824_p2[34], ret_V_24_fu_824_p2[34], ret_V_24_fu_824_p2[34], ret_V_24_fu_824_p2[34], ret_V_24_fu_824_p2[34], ret_V_24_fu_824_p2[34], ret_V_24_fu_824_p2[34], ret_V_24_fu_824_p2[34], ret_V_24_fu_824_p2[34], ret_V_24_fu_824_p2[34], ret_V_24_fu_824_p2[34], ret_V_24_fu_824_p2[34], ret_V_24_fu_824_p2[34], ret_V_24_fu_824_p2[34], ret_V_24_fu_824_p2[34], ret_V_24_fu_824_p2[34], ret_V_24_fu_824_p2[34], ret_V_24_fu_824_p2[34], ret_V_24_fu_824_p2[34], ret_V_24_fu_824_p2[34], ret_V_24_fu_824_p2[34], ret_V_24_fu_824_p2[34], ret_V_24_fu_824_p2[34], ret_V_24_fu_824_p2[34], ret_V_24_fu_824_p2[8:2] } : ret_V_29_cast_reg_1076;
assign _014_ = ap_CS_fsm[5] ? { ret_V_24_fu_824_p2[34], ret_V_24_fu_824_p2[34], ret_V_24_fu_824_p2[34], ret_V_24_fu_824_p2[34], ret_V_24_fu_824_p2[34], ret_V_24_fu_824_p2[34], ret_V_24_fu_824_p2[34], ret_V_24_fu_824_p2[34], ret_V_24_fu_824_p2[34], ret_V_24_fu_824_p2[34], ret_V_24_fu_824_p2[34], ret_V_24_fu_824_p2[34], ret_V_24_fu_824_p2[34], ret_V_24_fu_824_p2[34], ret_V_24_fu_824_p2[34], ret_V_24_fu_824_p2[34], ret_V_24_fu_824_p2[34], ret_V_24_fu_824_p2[34], ret_V_24_fu_824_p2[34], ret_V_24_fu_824_p2[34], ret_V_24_fu_824_p2[34], ret_V_24_fu_824_p2[34], ret_V_24_fu_824_p2[34], ret_V_24_fu_824_p2[34], ret_V_24_fu_824_p2[34], ret_V_24_fu_824_p2[34], ret_V_24_fu_824_p2[8:0] } : ret_V_24_reg_1071;
assign _001_ = ap_CS_fsm[3] ? add_ln69_3_fu_743_p2 : add_ln69_3_reg_1061;
assign _002_ = ap_CS_fsm[3] ? add_ln69_fu_734_p2 : add_ln69_reg_1056;
assign _013_ = ap_CS_fsm[3] ? ret_V_23_fu_716_p2 : ret_V_23_reg_1051;
assign _000_ = ap_CS_fsm[2] ? add_ln69_2_fu_612_p2 : add_ln69_2_reg_1046;
assign _006_ = ap_CS_fsm[2] ? icmp_ln851_fu_503_p2 : icmp_ln851_reg_1036;
assign _019_ = ap_CS_fsm[2] ? ret_V_19_fu_483_p2[8:3] : ret_V_reg_1029;
assign _012_ = ap_CS_fsm[2] ? ret_V_19_fu_483_p2 : ret_V_19_reg_1024;
assign _010_ = ap_CS_fsm[2] ? op_6_V_fu_468_p2 : op_6_V_reg_1014;
assign _003_ = ap_rst ? 10'h001 : ap_NS_fsm;
assign shl_ln1358_fu_550_p2 = $signed(op_8_V_reg_996) << ush_reg_1009;
assign ashr_ln1297_fu_545_p2 = $signed(op_8_V_reg_996) >>> ush_reg_1009;
assign ret_fu_216_p2 = $signed(select_ln1347_fu_205_p3) - $signed(op_4);
assign sub_ln1118_fu_520_p2 = $signed(1'h0) - $signed({ op_4, 24'h000000 });
assign sub_ln1357_fu_377_p2 = 1'h0 - r_2_fu_365_p1;
assign sub_ln69_fu_474_p2 = $signed(1'h0) - $signed(op_4);
assign icmp_ln1494_fu_536_p2 = _032_ ? 1'h1 : 1'h0;
assign icmp_ln768_fu_258_p2 = _033_ ? 1'h1 : 1'h0;
assign icmp_ln850_1_fu_582_p2 = _034_ ? 1'h1 : 1'h0;
assign icmp_ln850_fu_791_p2 = _035_ ? 1'h1 : 1'h0;
assign icmp_ln851_1_fu_681_p2 = _030_ ? 1'h1 : 1'h0;
assign icmp_ln851_2_fu_844_p2 = _036_ ? 1'h1 : 1'h0;
assign icmp_ln851_3_fu_923_p2 = _037_ ? 1'h1 : 1'h0;
assign icmp_ln851_fu_503_p2 = _031_ ? 1'h1 : 1'h0;
assign op_7_V_fu_618_p3 = op_3 ? sub_ln69_reg_1019 : 2'h0;
assign op_8_V_fu_296_p3 = or_ln384_fu_290_p2 ? select_ln384_fu_282_p3 : { ret_fu_216_p2[0], 3'h0 };
assign p_Result_8_fu_242_p2 = ret_fu_216_p2[0] ? 1'h1 : 1'h0;
assign r_V_1_fu_555_p3 = isNeg_reg_1004 ? ashr_ln1297_fu_545_p2 : shl_ln1358_fu_550_p2;
assign r_V_fu_649_p3 = op_3 ? sub_ln1118_reg_1041 : 27'h0000000;
assign r_fu_432_p2 = _038_ ? 1'h1 : 1'h0;
assign ret_V_20_fu_642_p3 = ret_V_19_reg_1024[8] ? select_ln850_fu_636_p3 : ret_V_reg_1029;
assign ret_V_21_fu_701_p3 = r_V_fu_649_p3[26] ? select_ln850_2_fu_693_p3 : { 2'h0, r_V_fu_649_p3[25:24] };
assign ret_V_25_fu_876_p3 = ret_V_24_reg_1071[34] ? select_ln850_3_fu_870_p3 : ret_V_29_cast_reg_1076;
assign ret_V_27_fu_947_p3 = ret_V_26_reg_1098[35] ? select_ln850_4_fu_941_p3 : ret_V_31_cast_reg_1103;
assign select_ln1347_fu_205_p3 = op_3 ? 3'h7 : 3'h0;
assign select_ln13_fu_197_p3 = op_3 ? 1'h1 : 1'h0;
assign select_ln1497_1_fu_336_p3 = op_4[1] ? 2'h3 : 2'h0;
assign select_ln1497_2_fu_350_p3 = select_ln13_reg_982 ? select_ln1497_1_fu_336_p3 : op_4;
assign r_2_fu_365_p1 = select_ln835_fu_304_p3 ? select_ln1497_2_fu_350_p3 : { op_4[1], select_ln1497_fu_321_p3[0] };
assign select_ln1497_fu_321_p3[0] = select_ln13_reg_982 ? op_4[1] : op_4[0];
assign select_ln384_fu_282_p3 = overflow_fu_276_p2 ? 4'h7 : 4'h9;
assign select_ln69_1_fu_850_p3 = ret_V_9_fu_803_p2 ? 32'd4294967295 : 32'd0;
assign select_ln69_fu_604_p3 = ret_V_12_fu_594_p2 ? 2'h3 : 2'h0;
assign select_ln708_fu_412_p3 = ret_V_18_fu_398_p2[3] ? 2'h3 : 2'h0;
assign select_ln835_fu_304_p3 = select_ln13_reg_982 ? 1'h1 : 1'h0;
assign select_ln850_2_fu_693_p3 = icmp_ln851_1_fu_681_p2 ? { 2'h3, r_V_fu_649_p3[25:24] } : ret_V_5_fu_687_p2;
assign select_ln850_3_fu_870_p3 = icmp_ln851_2_reg_1083 ? add_ln691_fu_865_p2 : ret_V_29_cast_reg_1076;
assign select_ln850_4_fu_941_p3 = icmp_ln851_3_reg_1110 ? add_ln691_1_fu_936_p2 : ret_V_31_cast_reg_1103;
assign select_ln850_fu_636_p3 = icmp_ln851_reg_1036 ? ret_V_reg_1029 : ret_V_3_fu_631_p2;
assign ush_fu_383_p3 = r_2_fu_365_p1[1] ? sub_ln1357_fu_377_p2 : { 1'h0, r_2_fu_365_p1[0] };
assign ret_V_12_fu_594_p2 = r_V_1_fu_555_p3[3] ^ and_ln850_1_fu_588_p2;
assign ret_V_9_fu_803_p2 = ret_V_22_fu_766_p2[3] ^ and_ln850_fu_797_p2;
assign ap_CS_fsm_state1 = ap_CS_fsm[0];
assign ap_CS_fsm_state10 = ap_CS_fsm[9];
assign ap_CS_fsm_state2 = ap_CS_fsm[1];
assign ap_CS_fsm_state3 = ap_CS_fsm[2];
assign ap_CS_fsm_state4 = ap_CS_fsm[3];
assign ap_CS_fsm_state5 = ap_CS_fsm[4];
assign ap_CS_fsm_state6 = ap_CS_fsm[5];
assign ap_CS_fsm_state7 = ap_CS_fsm[6];
assign ap_CS_fsm_state8 = ap_CS_fsm[7];
assign ap_CS_fsm_state9 = ap_CS_fsm[8];
assign ap_done = op_31_ap_vld;
assign ap_ready = op_31_ap_vld;
assign ashr_ln1497_1_fu_344_p2 = { op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4 };
assign conv_i389_fu_311_p0 = op_4;
assign conv_i389_fu_311_p1 = { op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4 };
assign isNeg_fu_369_p3 = r_2_fu_365_p1[1];
assign op_3_read_read_fu_130_p2 = op_3;
assign op_7_V_fu_618_p0 = op_3;
assign p_Result_1_fu_669_p3 = r_V_fu_649_p3[26];
assign p_Result_2_fu_779_p3 = ret_V_22_fu_766_p2[3];
assign p_Result_3_fu_570_p3 = r_V_1_fu_555_p3[3];
assign p_Result_4_fu_858_p3 = ret_V_24_reg_1071[34];
assign p_Result_5_fu_929_p3 = ret_V_26_reg_1098[35];
assign p_Result_6_fu_420_p3 = op_1[2];
assign p_Result_7_fu_222_p3 = ret_fu_216_p2[2];
assign p_Result_s_14_fu_624_p3 = ret_V_19_reg_1024[8];
assign p_Result_s_fu_248_p4 = ret_fu_216_p2[2:1];
assign p_Val2_2_fu_234_p3 = { ret_fu_216_p2[0], 3'h0 };
assign r_V_fu_649_p0 = op_3;
assign ret_V_11_fu_562_p3 = r_V_1_fu_555_p3[3];
assign ret_V_24_fu_824_p2[33:9] = { ret_V_24_fu_824_p2[34], ret_V_24_fu_824_p2[34], ret_V_24_fu_824_p2[34], ret_V_24_fu_824_p2[34], ret_V_24_fu_824_p2[34], ret_V_24_fu_824_p2[34], ret_V_24_fu_824_p2[34], ret_V_24_fu_824_p2[34], ret_V_24_fu_824_p2[34], ret_V_24_fu_824_p2[34], ret_V_24_fu_824_p2[34], ret_V_24_fu_824_p2[34], ret_V_24_fu_824_p2[34], ret_V_24_fu_824_p2[34], ret_V_24_fu_824_p2[34], ret_V_24_fu_824_p2[34], ret_V_24_fu_824_p2[34], ret_V_24_fu_824_p2[34], ret_V_24_fu_824_p2[34], ret_V_24_fu_824_p2[34], ret_V_24_fu_824_p2[34], ret_V_24_fu_824_p2[34], ret_V_24_fu_824_p2[34], ret_V_24_fu_824_p2[34], ret_V_24_fu_824_p2[34] };
assign ret_V_8_fu_771_p3 = ret_V_22_fu_766_p2[3];
assign rhs_4_fu_892_p3 = { op_28_V_reg_1093, 3'h0 };
assign rhs_fu_391_p1 = op_3;
assign rhs_fu_391_p3 = { op_3, 3'h0 };
assign select_ln1347_fu_205_p0 = op_3;
assign select_ln13_fu_197_p0 = op_3;
assign select_ln1497_3_fu_357_p3 = { 30'hxxxxxxxx, r_2_fu_365_p1 };
assign select_ln1497_fu_321_p3[1] = op_4[1];
assign sext_ln1118_fu_516_p1 = { op_4[1], op_4, 24'h000000 };
assign sext_ln1192_1_fu_712_p1 = { ret_V_20_fu_642_p3[5], ret_V_20_fu_642_p3 };
assign sext_ln1192_2_fu_820_p1 = { op_26_V_reg_1066[6], op_26_V_reg_1066[6], op_26_V_reg_1066[6], op_26_V_reg_1066[6], op_26_V_reg_1066[6], op_26_V_reg_1066[6], op_26_V_reg_1066[6], op_26_V_reg_1066[6], op_26_V_reg_1066[6], op_26_V_reg_1066[6], op_26_V_reg_1066[6], op_26_V_reg_1066[6], op_26_V_reg_1066[6], op_26_V_reg_1066[6], op_26_V_reg_1066[6], op_26_V_reg_1066[6], op_26_V_reg_1066[6], op_26_V_reg_1066[6], op_26_V_reg_1066[6], op_26_V_reg_1066[6], op_26_V_reg_1066[6], op_26_V_reg_1066[6], op_26_V_reg_1066[6], op_26_V_reg_1066[6], op_26_V_reg_1066[6], op_26_V_reg_1066[6], op_26_V_reg_1066, 2'h0 };
assign sext_ln1192_3_fu_899_p1 = { op_28_V_reg_1093[31], op_28_V_reg_1093, 3'h0 };
assign sext_ln1192_4_fu_954_p1 = { op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18 };
assign sext_ln1192_fu_709_p1 = { op_6_V_reg_1014[1], op_6_V_reg_1014[1], op_6_V_reg_1014[1], op_6_V_reg_1014[1], op_6_V_reg_1014[1], op_6_V_reg_1014 };
assign sext_ln1347_fu_212_p0 = op_4;
assign sext_ln1347_fu_212_p1 = { op_4[1], op_4 };
assign sext_ln1494_fu_533_p1 = { op_8_V_reg_996[3], op_8_V_reg_996 };
assign sext_ln69_1_fu_726_p1 = { ret_V_21_fu_701_p3[3], ret_V_21_fu_701_p3[3], ret_V_21_fu_701_p3 };
assign sext_ln69_2_fu_749_p1 = { add_ln69_reg_1056[5], add_ln69_reg_1056 };
assign sext_ln69_4_fu_963_p1 = { op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19 };
assign sext_ln69_5_fu_740_p1 = { add_ln69_2_reg_1046[1], add_ln69_2_reg_1046 };
assign sext_ln69_6_fu_757_p1 = { add_ln69_3_reg_1061[2], add_ln69_3_reg_1061[2], add_ln69_3_reg_1061[2], add_ln69_3_reg_1061[2], add_ln69_3_reg_1061 };
assign sext_ln69_fu_722_p1 = { op_7_V_fu_618_p3[1], op_7_V_fu_618_p3 };
assign sext_ln703_1_fu_809_p0 = op_15;
assign sext_ln703_1_fu_809_p1 = { op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15 };
assign sext_ln703_2_fu_888_p0 = op_17;
assign sext_ln703_2_fu_888_p1 = { op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17 };
assign sext_ln703_fu_479_p1 = { op_0[7], op_0 };
assign sext_ln850_fu_665_p1 = { r_V_fu_649_p3[26], r_V_fu_649_p3[26:24] };
assign shl_ln1497_1_fu_315_p2 = { op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1], op_4[1] };
assign shl_ln1_fu_526_p1 = op_4;
assign shl_ln1_fu_526_p3 = { op_4, 3'h0 };
assign shl_ln_fu_509_p1 = op_4;
assign shl_ln_fu_509_p3 = { op_4, 24'h000000 };
assign sub_ln69_fu_474_p1 = op_4;
assign tmp_14_fu_813_p3 = { op_26_V_reg_1066, 2'h0 };
assign tmp_2_fu_655_p4 = r_V_fu_649_p3[26:24];
assign tmp_3_fu_438_p3 = ret_V_18_fu_398_p2[3];
assign tmp_7_fu_328_p1 = op_4;
assign tmp_7_fu_328_p3 = op_4[1];
assign tmp_fu_404_p3 = ret_V_18_fu_398_p2[3];
assign trunc_ln718_fu_428_p1 = ret_V_18_fu_398_p2[1:0];
assign trunc_ln728_fu_230_p1 = ret_fu_216_p2[0];
assign trunc_ln851_1_fu_677_p1 = r_V_fu_649_p3[23:0];
assign trunc_ln851_2_fu_787_p1 = ret_V_22_fu_766_p2[2:0];
assign trunc_ln851_3_fu_578_p1 = r_V_1_fu_555_p3[2:0];
assign trunc_ln851_4_fu_840_p0 = op_15;
assign trunc_ln851_4_fu_840_p1 = op_15[1:0];
assign trunc_ln851_5_fu_919_p0 = op_17;
assign trunc_ln851_5_fu_919_p1 = op_17[2:0];
assign trunc_ln851_fu_499_p1 = ret_V_19_fu_483_p2[2:0];
assign zext_ln1357_fu_542_p1 = { 2'h0, ush_reg_1009 };
assign zext_ln415_fu_464_p1 = { 1'h0, and_ln410_fu_458_p2 };
assign zext_ln69_1_fu_600_p1 = { 1'h0, icmp_ln1494_fu_536_p2 };
assign zext_ln69_fu_730_p1 = { 2'h0, op_12 };
endmodule


// Product machine:
module top_A_times_top_B (ap_start, op_0, op_1, op_11, op_12, op_15, op_17, op_18, op_19, op_3, op_4, ap_clk, unsafe_signal);
input ap_start;
input [7:0] op_0;
input [3:0] op_1;
input [3:0] op_11;
input [3:0] op_12;
input [3:0] op_15;
input [3:0] op_17;
input [1:0] op_18;
input [3:0] op_19;
input op_3;
input [1:0] op_4;
input ap_clk;
output unsafe_signal;
reg _setup;
initial _setup = 1'b0;
always @ (posedge ap_clk) _setup <= 1'b1;
reg ap_start_internal;
always @ (posedge ap_clk) if (!_setup) ap_start_internal <= ap_start;
reg [7:0] op_0_internal;
always @ (posedge ap_clk) if (!_setup) op_0_internal <= op_0;
reg [3:0] op_1_internal;
always @ (posedge ap_clk) if (!_setup) op_1_internal <= op_1;
reg [3:0] op_11_internal;
always @ (posedge ap_clk) if (!_setup) op_11_internal <= op_11;
reg [3:0] op_12_internal;
always @ (posedge ap_clk) if (!_setup) op_12_internal <= op_12;
reg [3:0] op_15_internal;
always @ (posedge ap_clk) if (!_setup) op_15_internal <= op_15;
reg [3:0] op_17_internal;
always @ (posedge ap_clk) if (!_setup) op_17_internal <= op_17;
reg [1:0] op_18_internal;
always @ (posedge ap_clk) if (!_setup) op_18_internal <= op_18;
reg [3:0] op_19_internal;
always @ (posedge ap_clk) if (!_setup) op_19_internal <= op_19;
reg op_3_internal;
always @ (posedge ap_clk) if (!_setup) op_3_internal <= op_3;
reg [1:0] op_4_internal;
always @ (posedge ap_clk) if (!_setup) op_4_internal <= op_4;
wire ap_done_A;
wire ap_done_B;
wire ap_done_eq;
assign ap_done_eq = ap_done_A == ap_done_B;
wire ap_idle_A;
wire ap_idle_B;
wire ap_idle_eq;
assign ap_idle_eq = ap_idle_A == ap_idle_B;
wire ap_ready_A;
wire ap_ready_B;
wire ap_ready_eq;
assign ap_ready_eq = ap_ready_A == ap_ready_B;
wire [31:0] op_31_A;
wire [31:0] op_31_B;
wire op_31_eq;
assign op_31_eq = op_31_A == op_31_B;
wire op_31_ap_vld_A;
wire op_31_ap_vld_B;
wire clk_enable_A;
wire clk_enable_B;
assign clk_enable_A = _setup & (~op_31_ap_vld_A | op_31_ap_vld_B);
assign clk_enable_B = _setup;
wire divergent;
assign divergent = ~(ap_done_eq & ap_idle_eq & ap_ready_eq & op_31_eq);
assign unsafe_signal = op_31_ap_vld_A & op_31_ap_vld_B & divergent;
top_A instance_A (
    .ap_clk(ap_clk),
    .clk_enable(clk_enable_A),
    .ap_start(ap_start_internal),
    .op_0(op_0_internal),
    .op_1(op_1_internal),
    .op_11(op_11_internal),
    .op_12(op_12_internal),
    .op_15(op_15_internal),
    .op_17(op_17_internal),
    .op_18(op_18_internal),
    .op_19(op_19_internal),
    .op_3(op_3_internal),
    .op_4(op_4_internal),
    .ap_done(ap_done_A),
    .ap_idle(ap_idle_A),
    .ap_ready(ap_ready_A),
    .op_31(op_31_A),
    .op_31_ap_vld(op_31_ap_vld_A)
);
top_B instance_B (
    .ap_clk(ap_clk),
    .clk_enable(clk_enable_B),
    .ap_start(ap_start_internal),
    .op_0(op_0_internal),
    .op_1(op_1_internal),
    .op_11(op_11_internal),
    .op_12(op_12_internal),
    .op_15(op_15_internal),
    .op_17(op_17_internal),
    .op_18(op_18_internal),
    .op_19(op_19_internal),
    .op_3(op_3_internal),
    .op_4(op_4_internal),
    .ap_done(ap_done_B),
    .ap_idle(ap_idle_B),
    .ap_ready(ap_ready_B),
    .op_31(op_31_B),
    .op_31_ap_vld(op_31_ap_vld_B)
);
endmodule
