// Processed by function `construct_kairos` in `verilog_tricks.py`.
// Machine A:
// Processed by function `add_clk_enable_signal` in `verilog_tricks.py`.
// Processed by function `remove_reset_signal` in `verilog_tricks.py`.
module top_A (
  ap_clk,
  ap_start,
  ap_done,
  ap_idle,
  ap_ready,
  op_0,
  op_1,
  op_4,
  op_5,
  op_6,
  op_7,
  op_10,
  op_11,
  op_18,
  op_19,
  op_29,
  op_29_ap_vld,
clk_enable
);
input clk_enable;


input ap_clk;
wire ap_rst;
assign ap_rst = op_29_ap_vld;
input ap_start;
input [3:0] op_0;
input [3:0] op_1;
input [3:0] op_10;
input [3:0] op_11;
input [1:0] op_18;
input [3:0] op_19;
input [1:0] op_4;
input [3:0] op_5;
input [3:0] op_6;
input [15:0] op_7;
output ap_done;
output ap_idle;
output ap_ready;
output [31:0] op_29;
output op_29_ap_vld;


reg [8:0] \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.ain_s1 ;
reg [8:0] \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.bin_s1 ;
reg \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.carry_s1 ;
reg [7:0] \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.sum_s1 ;
reg [8:0] \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.ain_s1 ;
reg [8:0] \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.bin_s1 ;
reg \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.carry_s1 ;
reg [7:0] \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.sum_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s1 ;
reg \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.carry_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.sum_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s1 ;
reg \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.carry_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.sum_s1 ;
reg [15:0] \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.ain_s1 ;
reg [15:0] \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.bin_s1 ;
reg \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.carry_s1 ;
reg [15:0] \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.sum_s1 ;
reg [15:0] \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.ain_s1 ;
reg [15:0] \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.bin_s1 ;
reg \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.carry_s1 ;
reg [15:0] \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.sum_s1 ;
reg [16:0] \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.ain_s1 ;
reg [16:0] \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.bin_s1 ;
reg \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.carry_s1 ;
reg [16:0] \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.sum_s1 ;
reg [17:0] \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.ain_s1 ;
reg [17:0] \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.bin_s1 ;
reg \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.carry_s1 ;
reg [17:0] \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.sum_s1 ;
reg [17:0] \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.ain_s1 ;
reg [17:0] \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.bin_s1 ;
reg \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.carry_s1 ;
reg [17:0] \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.sum_s1 ;
reg [1:0] \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.ain_s1 ;
reg [1:0] \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.bin_s1 ;
reg \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.carry_s1 ;
reg [1:0] \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.sum_s1 ;
reg [1:0] \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.ain_s1 ;
reg [1:0] \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.bin_s1 ;
reg \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.carry_s1 ;
reg [1:0] \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.sum_s1 ;
reg [1:0] \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.ain_s1 ;
reg [1:0] \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.bin_s1 ;
reg \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.carry_s1 ;
reg [1:0] \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.sum_s1 ;
reg [2:0] \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.ain_s1 ;
reg [2:0] \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.bin_s1 ;
reg \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.carry_s1 ;
reg [1:0] \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.sum_s1 ;
reg [2:0] \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.ain_s1 ;
reg [2:0] \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.bin_s1 ;
reg \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.carry_s1 ;
reg [2:0] \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.sum_s1 ;
reg [3:0] \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.ain_s1 ;
reg [3:0] \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.bin_s1 ;
reg \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.carry_s1 ;
reg [3:0] \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.sum_s1 ;
reg [31:0] add_ln691_1_reg_995;
reg [5:0] add_ln691_reg_957;
reg [31:0] add_ln69_2_reg_1100;
reg [3:0] add_ln69_3_reg_1105;
reg [16:0] add_ln69_reg_1040;
reg [36:0] ap_CS_fsm = 37'h0000000001;
reg [31:0] \ashr_32s_32s_32_7_1_U5.din1_cast_array[0] ;
reg [31:0] \ashr_32s_32s_32_7_1_U5.din1_cast_array[1] ;
reg [31:0] \ashr_32s_32s_32_7_1_U5.din1_cast_array[2] ;
reg [31:0] \ashr_32s_32s_32_7_1_U5.din1_cast_array[3] ;
reg [31:0] \ashr_32s_32s_32_7_1_U5.din1_cast_array[4] ;
reg [31:0] \ashr_32s_32s_32_7_1_U5.din1_cast_array[5] ;
reg [31:0] \ashr_32s_32s_32_7_1_U5.dout_array[0] ;
reg [31:0] \ashr_32s_32s_32_7_1_U5.dout_array[1] ;
reg [31:0] \ashr_32s_32s_32_7_1_U5.dout_array[2] ;
reg [31:0] \ashr_32s_32s_32_7_1_U5.dout_array[3] ;
reg [31:0] \ashr_32s_32s_32_7_1_U5.dout_array[4] ;
reg [31:0] \ashr_32s_32s_32_7_1_U5.dout_array[5] ;
reg icmp_ln768_reg_939;
reg icmp_ln851_1_reg_907;
reg icmp_ln851_reg_872;
reg icmp_ln890_reg_820;
reg [3:0] \mul_4s_4s_4_7_1_U2.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.a_reg0 ;
reg [3:0] \mul_4s_4s_4_7_1_U2.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.b_reg0 ;
reg [3:0] \mul_4s_4s_4_7_1_U2.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.buff0 ;
reg [3:0] \mul_4s_4s_4_7_1_U2.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.buff1 ;
reg [3:0] \mul_4s_4s_4_7_1_U2.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.buff2 ;
reg [3:0] \mul_4s_4s_4_7_1_U2.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.buff3 ;
reg [3:0] \mul_4s_4s_4_7_1_U2.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.buff4 ;
reg [1:0] op_12_V_reg_962;
reg [1:0] op_17_V_reg_1075;
reg [31:0] op_23_V_reg_1035;
reg [31:0] op_25_V_reg_1055;
reg [31:0] op_26_V_reg_1080;
reg [3:0] op_3_V_reg_793;
reg overflow_reg_951;
reg p_Result_8_reg_918;
reg p_Result_9_reg_912;
reg [4:0] ret_V_14_reg_750;
reg [3:0] ret_V_15_reg_1000;
reg [4:0] ret_V_16_reg_840;
reg [16:0] ret_V_17_reg_855;
reg [7:0] ret_V_18_reg_929;
reg [33:0] ret_V_19_reg_983;
reg [31:0] ret_V_21_cast_reg_988;
reg [3:0] ret_V_2_reg_763;
reg [3:0] ret_V_3_reg_768;
reg [3:0] ret_V_6_reg_1005;
reg [3:0] ret_V_7_reg_860;
reg [3:0] ret_V_9_reg_877;
reg [3:0] ret_V_reg_756;
reg [31:0] select_ln353_1_reg_1010;
reg [5:0] select_ln353_reg_968;
reg [3:0] select_ln850_3_reg_882;
reg [4:0] sext_ln703_3_reg_782;
reg [5:0] sext_ln850_reg_944;
reg [31:0] \shl_32s_32s_32_7_1_U6.din1_cast_array[0] ;
reg [31:0] \shl_32s_32s_32_7_1_U6.din1_cast_array[1] ;
reg [31:0] \shl_32s_32s_32_7_1_U6.din1_cast_array[2] ;
reg [31:0] \shl_32s_32s_32_7_1_U6.din1_cast_array[3] ;
reg [31:0] \shl_32s_32s_32_7_1_U6.din1_cast_array[4] ;
reg [31:0] \shl_32s_32s_32_7_1_U6.din1_cast_array[5] ;
reg [31:0] \shl_32s_32s_32_7_1_U6.dout_array[0] ;
reg [31:0] \shl_32s_32s_32_7_1_U6.dout_array[1] ;
reg [31:0] \shl_32s_32s_32_7_1_U6.dout_array[2] ;
reg [31:0] \shl_32s_32s_32_7_1_U6.dout_array[3] ;
reg [31:0] \shl_32s_32s_32_7_1_U6.dout_array[4] ;
reg [31:0] \shl_32s_32s_32_7_1_U6.dout_array[5] ;
reg signbit_reg_835;
reg \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.ain_s1 ;
reg \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.bin_s1 ;
reg \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.carry_s1 ;
reg \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.sum_s1 ;
reg [2:0] \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.ain_s1 ;
reg [2:0] \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.bin_s1 ;
reg \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.carry_s1 ;
reg [1:0] \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.sum_s1 ;
reg [4:0] sub_ln1497_reg_799;
reg [10:0] tmp_1_reg_924;
reg [4:0] tmp_2_reg_934;
reg tmp_V_reg_1050;
reg tmp_reg_788;
reg [1:0] trunc_ln1347_reg_804;
reg [11:0] trunc_ln1497_1_reg_892;
reg [3:0] trunc_ln1497_reg_887;
reg [12:0] trunc_ln851_1_reg_867;
wire [31:0] _000_;
wire [5:0] _001_;
wire [31:0] _002_;
wire [3:0] _003_;
wire [16:0] _004_;
wire [36:0] _005_;
wire _006_;
wire _007_;
wire _008_;
wire _009_;
wire [1:0] _010_;
wire [1:0] _011_;
wire [31:0] _012_;
wire [31:0] _013_;
wire [31:0] _014_;
wire [3:0] _015_;
wire _016_;
wire _017_;
wire _018_;
wire [4:0] _019_;
wire [3:0] _020_;
wire [4:0] _021_;
wire [16:0] _022_;
wire [7:0] _023_;
wire [33:0] _024_;
wire [31:0] _025_;
wire [3:0] _026_;
wire [3:0] _027_;
wire [3:0] _028_;
wire [3:0] _029_;
wire [3:0] _030_;
wire [3:0] _031_;
wire [31:0] _032_;
wire [5:0] _033_;
wire [3:0] _034_;
wire [4:0] _035_;
wire [5:0] _036_;
wire _037_;
wire [4:0] _038_;
wire [10:0] _039_;
wire [4:0] _040_;
wire _041_;
wire _042_;
wire [1:0] _043_;
wire [11:0] _044_;
wire [3:0] _045_;
wire [12:0] _046_;
wire [1:0] _047_;
wire _048_;
wire _049_;
wire _050_;
wire _051_;
wire _052_;
wire _053_;
wire _054_;
wire _055_;
wire [8:0] _056_;
wire [8:0] _057_;
wire _058_;
wire [7:0] _059_;
wire [8:0] _060_;
wire [9:0] _061_;
wire [8:0] _062_;
wire [8:0] _063_;
wire _064_;
wire [7:0] _065_;
wire [8:0] _066_;
wire [9:0] _067_;
wire [15:0] _068_;
wire [15:0] _069_;
wire _070_;
wire [15:0] _071_;
wire [16:0] _072_;
wire [16:0] _073_;
wire [15:0] _074_;
wire [15:0] _075_;
wire _076_;
wire [15:0] _077_;
wire [16:0] _078_;
wire [16:0] _079_;
wire [15:0] _080_;
wire [15:0] _081_;
wire _082_;
wire [15:0] _083_;
wire [16:0] _084_;
wire [16:0] _085_;
wire [15:0] _086_;
wire [15:0] _087_;
wire _088_;
wire [15:0] _089_;
wire [16:0] _090_;
wire [16:0] _091_;
wire [16:0] _092_;
wire [16:0] _093_;
wire _094_;
wire [16:0] _095_;
wire [17:0] _096_;
wire [17:0] _097_;
wire [17:0] _098_;
wire [17:0] _099_;
wire _100_;
wire [17:0] _101_;
wire [18:0] _102_;
wire [18:0] _103_;
wire [17:0] _104_;
wire [17:0] _105_;
wire _106_;
wire [17:0] _107_;
wire [18:0] _108_;
wire [18:0] _109_;
wire [1:0] _110_;
wire [1:0] _111_;
wire _112_;
wire [1:0] _113_;
wire [2:0] _114_;
wire [2:0] _115_;
wire [1:0] _116_;
wire [1:0] _117_;
wire _118_;
wire [1:0] _119_;
wire [2:0] _120_;
wire [2:0] _121_;
wire [1:0] _122_;
wire [1:0] _123_;
wire _124_;
wire [1:0] _125_;
wire [2:0] _126_;
wire [2:0] _127_;
wire [2:0] _128_;
wire [2:0] _129_;
wire _130_;
wire [1:0] _131_;
wire [2:0] _132_;
wire [3:0] _133_;
wire [2:0] _134_;
wire [2:0] _135_;
wire _136_;
wire [2:0] _137_;
wire [3:0] _138_;
wire [3:0] _139_;
wire [3:0] _140_;
wire [3:0] _141_;
wire _142_;
wire [3:0] _143_;
wire [4:0] _144_;
wire [4:0] _145_;
wire [31:0] _146_;
wire [31:0] _147_;
wire [31:0] _148_;
wire [31:0] _149_;
wire [31:0] _150_;
wire [31:0] _151_;
wire [31:0] _152_;
wire [31:0] _153_;
wire [31:0] _154_;
wire [31:0] _155_;
wire [31:0] _156_;
wire [31:0] _157_;
wire [31:0] _158_;
wire [31:0] _159_;
wire [31:0] _160_;
wire [31:0] _161_;
wire [31:0] _162_;
wire [31:0] _163_;
wire [31:0] _164_;
wire [31:0] _165_;
wire [31:0] _166_;
wire [31:0] _167_;
wire [31:0] _168_;
wire [31:0] _169_;
wire [31:0] _170_;
wire [31:0] _171_;
wire [31:0] _172_;
wire [31:0] _173_;
wire [31:0] _174_;
wire [31:0] _175_;
wire [3:0] _176_;
wire [3:0] _177_;
wire [3:0] _178_;
wire [3:0] _179_;
wire [3:0] _180_;
wire [3:0] _181_;
wire [3:0] _182_;
wire [31:0] _183_;
wire [31:0] _184_;
wire [31:0] _185_;
wire [31:0] _186_;
wire [31:0] _187_;
wire [31:0] _188_;
wire [31:0] _189_;
wire [31:0] _190_;
wire [31:0] _191_;
wire [31:0] _192_;
wire [31:0] _193_;
wire [31:0] _194_;
wire [31:0] _195_;
wire [31:0] _196_;
wire [31:0] _197_;
wire [31:0] _198_;
wire [31:0] _199_;
wire [31:0] _200_;
wire [31:0] _201_;
wire [31:0] _202_;
wire [31:0] _203_;
wire [31:0] _204_;
wire [31:0] _205_;
wire [31:0] _206_;
wire [31:0] _207_;
wire [31:0] _208_;
wire [31:0] _209_;
wire [31:0] _210_;
wire [31:0] _211_;
wire [31:0] _212_;
wire _213_;
wire _214_;
wire _215_;
wire _216_;
wire [1:0] _217_;
wire [1:0] _218_;
wire [2:0] _219_;
wire [2:0] _220_;
wire _221_;
wire [1:0] _222_;
wire [2:0] _223_;
wire [3:0] _224_;
wire _225_;
wire _226_;
wire _227_;
wire _228_;
wire _229_;
wire _230_;
wire _231_;
wire _232_;
wire _233_;
wire _234_;
wire _235_;
wire _236_;
wire _237_;
wire _238_;
wire _239_;
wire _240_;
wire _241_;
wire _242_;
wire _243_;
wire _244_;
wire _245_;
wire _246_;
wire _247_;
wire _248_;
wire _249_;
wire _250_;
wire _251_;
wire _252_;
wire _253_;
wire _254_;
wire _255_;
wire _256_;
wire _257_;
wire _258_;
wire _259_;
wire _260_;
wire _261_;
wire _262_;
wire _263_;
wire _264_;
wire _265_;
wire \add_17ns_17ns_17_2_1_U14.ce ;
wire \add_17ns_17ns_17_2_1_U14.clk ;
wire [16:0] \add_17ns_17ns_17_2_1_U14.din0 ;
wire [16:0] \add_17ns_17ns_17_2_1_U14.din1 ;
wire [16:0] \add_17ns_17ns_17_2_1_U14.dout ;
wire \add_17ns_17ns_17_2_1_U14.reset ;
wire [16:0] \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.a ;
wire [16:0] \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.ain_s0 ;
wire [16:0] \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.b ;
wire [16:0] \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.bin_s0 ;
wire \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.ce ;
wire \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.clk ;
wire \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.facout_s1 ;
wire \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.facout_s2 ;
wire [7:0] \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.fas_s1 ;
wire [8:0] \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.fas_s2 ;
wire \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.reset ;
wire [16:0] \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.s ;
wire [7:0] \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.u1.a ;
wire [7:0] \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.u1.b ;
wire \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.u1.cin ;
wire \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.u1.cout ;
wire [7:0] \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.u1.s ;
wire [8:0] \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.u2.a ;
wire [8:0] \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.u2.b ;
wire \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.u2.cin ;
wire \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.u2.cout ;
wire [8:0] \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.u2.s ;
wire \add_17ns_17s_17_2_1_U7.ce ;
wire \add_17ns_17s_17_2_1_U7.clk ;
wire [16:0] \add_17ns_17s_17_2_1_U7.din0 ;
wire [16:0] \add_17ns_17s_17_2_1_U7.din1 ;
wire [16:0] \add_17ns_17s_17_2_1_U7.dout ;
wire \add_17ns_17s_17_2_1_U7.reset ;
wire [16:0] \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.a ;
wire [16:0] \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.ain_s0 ;
wire [16:0] \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.b ;
wire [16:0] \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.bin_s0 ;
wire \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.ce ;
wire \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.clk ;
wire \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.facout_s1 ;
wire \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.facout_s2 ;
wire [7:0] \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.fas_s1 ;
wire [8:0] \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.fas_s2 ;
wire \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.reset ;
wire [16:0] \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.s ;
wire [7:0] \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.u1.a ;
wire [7:0] \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.u1.b ;
wire \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.u1.cin ;
wire \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.u1.cout ;
wire [7:0] \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.u1.s ;
wire [8:0] \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.u2.a ;
wire [8:0] \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.u2.b ;
wire \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.u2.cin ;
wire \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.u2.cout ;
wire [8:0] \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.u2.s ;
wire \add_32ns_32ns_32_2_1_U12.ce ;
wire \add_32ns_32ns_32_2_1_U12.clk ;
wire [31:0] \add_32ns_32ns_32_2_1_U12.din0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U12.din1 ;
wire [31:0] \add_32ns_32ns_32_2_1_U12.dout ;
wire \add_32ns_32ns_32_2_1_U12.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.a ;
wire [31:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.b ;
wire [31:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s0 ;
wire \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.ce ;
wire \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.clk ;
wire \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.facout_s1 ;
wire \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.facout_s2 ;
wire [15:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s1 ;
wire [15:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s2 ;
wire \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.b ;
wire \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cin ;
wire \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.b ;
wire \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cin ;
wire \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.s ;
wire \add_32ns_32ns_32_2_1_U15.ce ;
wire \add_32ns_32ns_32_2_1_U15.clk ;
wire [31:0] \add_32ns_32ns_32_2_1_U15.din0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U15.din1 ;
wire [31:0] \add_32ns_32ns_32_2_1_U15.dout ;
wire \add_32ns_32ns_32_2_1_U15.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.a ;
wire [31:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.b ;
wire [31:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s0 ;
wire \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.ce ;
wire \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.clk ;
wire \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.facout_s1 ;
wire \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.facout_s2 ;
wire [15:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s1 ;
wire [15:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s2 ;
wire \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.b ;
wire \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cin ;
wire \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.b ;
wire \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cin ;
wire \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.s ;
wire \add_32ns_32s_32_2_1_U18.ce ;
wire \add_32ns_32s_32_2_1_U18.clk ;
wire [31:0] \add_32ns_32s_32_2_1_U18.din0 ;
wire [31:0] \add_32ns_32s_32_2_1_U18.din1 ;
wire [31:0] \add_32ns_32s_32_2_1_U18.dout ;
wire \add_32ns_32s_32_2_1_U18.reset ;
wire [31:0] \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.a ;
wire [31:0] \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.ain_s0 ;
wire [31:0] \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.b ;
wire [31:0] \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.bin_s0 ;
wire \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.ce ;
wire \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.clk ;
wire \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.facout_s1 ;
wire \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.facout_s2 ;
wire [15:0] \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.fas_s1 ;
wire [15:0] \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.fas_s2 ;
wire \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.reset ;
wire [31:0] \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.s ;
wire [15:0] \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.u1.a ;
wire [15:0] \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.u1.b ;
wire \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.u1.cin ;
wire \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.u1.cout ;
wire [15:0] \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.u1.s ;
wire [15:0] \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.u2.a ;
wire [15:0] \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.u2.b ;
wire \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.u2.cin ;
wire \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.u2.cout ;
wire [15:0] \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.u2.s ;
wire \add_32s_32ns_32_2_1_U20.ce ;
wire \add_32s_32ns_32_2_1_U20.clk ;
wire [31:0] \add_32s_32ns_32_2_1_U20.din0 ;
wire [31:0] \add_32s_32ns_32_2_1_U20.din1 ;
wire [31:0] \add_32s_32ns_32_2_1_U20.dout ;
wire \add_32s_32ns_32_2_1_U20.reset ;
wire [31:0] \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.a ;
wire [31:0] \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.ain_s0 ;
wire [31:0] \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.b ;
wire [31:0] \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.bin_s0 ;
wire \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.ce ;
wire \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.clk ;
wire \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.facout_s1 ;
wire \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.facout_s2 ;
wire [15:0] \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.fas_s1 ;
wire [15:0] \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.fas_s2 ;
wire \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.reset ;
wire [31:0] \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.s ;
wire [15:0] \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.u1.a ;
wire [15:0] \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.u1.b ;
wire \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.u1.cin ;
wire \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.u1.cout ;
wire [15:0] \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.u1.s ;
wire [15:0] \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.u2.a ;
wire [15:0] \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.u2.b ;
wire \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.u2.cin ;
wire \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.u2.cout ;
wire [15:0] \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.u2.s ;
wire \add_34s_34s_34_2_1_U11.ce ;
wire \add_34s_34s_34_2_1_U11.clk ;
wire [33:0] \add_34s_34s_34_2_1_U11.din0 ;
wire [33:0] \add_34s_34s_34_2_1_U11.din1 ;
wire [33:0] \add_34s_34s_34_2_1_U11.dout ;
wire \add_34s_34s_34_2_1_U11.reset ;
wire [33:0] \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.a ;
wire [33:0] \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.ain_s0 ;
wire [33:0] \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.b ;
wire [33:0] \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.bin_s0 ;
wire \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.ce ;
wire \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.clk ;
wire \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.facout_s1 ;
wire \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.facout_s2 ;
wire [16:0] \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.fas_s1 ;
wire [16:0] \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.fas_s2 ;
wire \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.reset ;
wire [33:0] \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.s ;
wire [16:0] \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.u1.a ;
wire [16:0] \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.u1.b ;
wire \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.u1.cin ;
wire \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.u1.cout ;
wire [16:0] \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.u1.s ;
wire [16:0] \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.u2.a ;
wire [16:0] \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.u2.b ;
wire \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.u2.cin ;
wire \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.u2.cout ;
wire [16:0] \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.u2.s ;
wire \add_36ns_36ns_36_2_1_U17.ce ;
wire \add_36ns_36ns_36_2_1_U17.clk ;
wire [35:0] \add_36ns_36ns_36_2_1_U17.din0 ;
wire [35:0] \add_36ns_36ns_36_2_1_U17.din1 ;
wire [35:0] \add_36ns_36ns_36_2_1_U17.dout ;
wire \add_36ns_36ns_36_2_1_U17.reset ;
wire [35:0] \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.a ;
wire [35:0] \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.ain_s0 ;
wire [35:0] \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.b ;
wire [35:0] \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.bin_s0 ;
wire \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.ce ;
wire \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.clk ;
wire \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.facout_s1 ;
wire \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.facout_s2 ;
wire [17:0] \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.fas_s1 ;
wire [17:0] \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.fas_s2 ;
wire \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.reset ;
wire [35:0] \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.s ;
wire [17:0] \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.u1.a ;
wire [17:0] \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.u1.b ;
wire \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.u1.cin ;
wire \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.u1.cout ;
wire [17:0] \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.u1.s ;
wire [17:0] \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.u2.a ;
wire [17:0] \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.u2.b ;
wire \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.u2.cin ;
wire \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.u2.cout ;
wire [17:0] \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.u2.s ;
wire \add_36ns_36s_36_2_1_U13.ce ;
wire \add_36ns_36s_36_2_1_U13.clk ;
wire [35:0] \add_36ns_36s_36_2_1_U13.din0 ;
wire [35:0] \add_36ns_36s_36_2_1_U13.din1 ;
wire [35:0] \add_36ns_36s_36_2_1_U13.dout ;
wire \add_36ns_36s_36_2_1_U13.reset ;
wire [35:0] \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.a ;
wire [35:0] \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.ain_s0 ;
wire [35:0] \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.b ;
wire [35:0] \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.bin_s0 ;
wire \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.ce ;
wire \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.clk ;
wire \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.facout_s1 ;
wire \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.facout_s2 ;
wire [17:0] \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.fas_s1 ;
wire [17:0] \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.fas_s2 ;
wire \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.reset ;
wire [35:0] \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.s ;
wire [17:0] \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.u1.a ;
wire [17:0] \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.u1.b ;
wire \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.u1.cin ;
wire \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.u1.cout ;
wire [17:0] \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.u1.s ;
wire [17:0] \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.u2.a ;
wire [17:0] \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.u2.b ;
wire \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.u2.cin ;
wire \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.u2.cout ;
wire [17:0] \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.u2.s ;
wire \add_4ns_4ns_4_2_1_U1.ce ;
wire \add_4ns_4ns_4_2_1_U1.clk ;
wire [3:0] \add_4ns_4ns_4_2_1_U1.din0 ;
wire [3:0] \add_4ns_4ns_4_2_1_U1.din1 ;
wire [3:0] \add_4ns_4ns_4_2_1_U1.dout ;
wire \add_4ns_4ns_4_2_1_U1.reset ;
wire [3:0] \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.a ;
wire [3:0] \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.ain_s0 ;
wire [3:0] \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.b ;
wire [3:0] \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.bin_s0 ;
wire \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.ce ;
wire \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.clk ;
wire \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.facout_s1 ;
wire \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.facout_s2 ;
wire [1:0] \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.fas_s1 ;
wire [1:0] \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.fas_s2 ;
wire \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.reset ;
wire [3:0] \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.s ;
wire [1:0] \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.u1.a ;
wire [1:0] \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.u1.b ;
wire \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.u1.cin ;
wire \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.u1.cout ;
wire [1:0] \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.u1.s ;
wire [1:0] \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.u2.a ;
wire [1:0] \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.u2.b ;
wire \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.u2.cin ;
wire \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.u2.cout ;
wire [1:0] \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.u2.s ;
wire \add_4ns_4ns_4_2_1_U8.ce ;
wire \add_4ns_4ns_4_2_1_U8.clk ;
wire [3:0] \add_4ns_4ns_4_2_1_U8.din0 ;
wire [3:0] \add_4ns_4ns_4_2_1_U8.din1 ;
wire [3:0] \add_4ns_4ns_4_2_1_U8.dout ;
wire \add_4ns_4ns_4_2_1_U8.reset ;
wire [3:0] \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.a ;
wire [3:0] \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.ain_s0 ;
wire [3:0] \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.b ;
wire [3:0] \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.bin_s0 ;
wire \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.ce ;
wire \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.clk ;
wire \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.facout_s1 ;
wire \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.facout_s2 ;
wire [1:0] \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.fas_s1 ;
wire [1:0] \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.fas_s2 ;
wire \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.reset ;
wire [3:0] \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.s ;
wire [1:0] \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.u1.a ;
wire [1:0] \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.u1.b ;
wire \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.u1.cin ;
wire \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.u1.cout ;
wire [1:0] \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.u1.s ;
wire [1:0] \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.u2.a ;
wire [1:0] \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.u2.b ;
wire \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.u2.cin ;
wire \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.u2.cout ;
wire [1:0] \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.u2.s ;
wire \add_4ns_4s_4_2_1_U19.ce ;
wire \add_4ns_4s_4_2_1_U19.clk ;
wire [3:0] \add_4ns_4s_4_2_1_U19.din0 ;
wire [3:0] \add_4ns_4s_4_2_1_U19.din1 ;
wire [3:0] \add_4ns_4s_4_2_1_U19.dout ;
wire \add_4ns_4s_4_2_1_U19.reset ;
wire [3:0] \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.a ;
wire [3:0] \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.ain_s0 ;
wire [3:0] \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.b ;
wire [3:0] \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.bin_s0 ;
wire \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.ce ;
wire \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.clk ;
wire \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.facout_s1 ;
wire \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.facout_s2 ;
wire [1:0] \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.fas_s1 ;
wire [1:0] \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.fas_s2 ;
wire \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.reset ;
wire [3:0] \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.s ;
wire [1:0] \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.u1.a ;
wire [1:0] \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.u1.b ;
wire \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.u1.cin ;
wire \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.u1.cout ;
wire [1:0] \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.u1.s ;
wire [1:0] \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.u2.a ;
wire [1:0] \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.u2.b ;
wire \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.u2.cin ;
wire \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.u2.cout ;
wire [1:0] \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.u2.s ;
wire \add_5s_5s_5_2_1_U4.ce ;
wire \add_5s_5s_5_2_1_U4.clk ;
wire [4:0] \add_5s_5s_5_2_1_U4.din0 ;
wire [4:0] \add_5s_5s_5_2_1_U4.din1 ;
wire [4:0] \add_5s_5s_5_2_1_U4.dout ;
wire \add_5s_5s_5_2_1_U4.reset ;
wire [4:0] \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.a ;
wire [4:0] \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.ain_s0 ;
wire [4:0] \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.b ;
wire [4:0] \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.bin_s0 ;
wire \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.ce ;
wire \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.clk ;
wire \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.facout_s1 ;
wire \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.facout_s2 ;
wire [1:0] \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.fas_s1 ;
wire [2:0] \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.fas_s2 ;
wire \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.reset ;
wire [4:0] \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.s ;
wire [1:0] \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.u1.a ;
wire [1:0] \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.u1.b ;
wire \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.u1.cin ;
wire \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.u1.cout ;
wire [1:0] \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.u1.s ;
wire [2:0] \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.u2.a ;
wire [2:0] \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.u2.b ;
wire \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.u2.cin ;
wire \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.u2.cout ;
wire [2:0] \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.u2.s ;
wire \add_6s_6ns_6_2_1_U10.ce ;
wire \add_6s_6ns_6_2_1_U10.clk ;
wire [5:0] \add_6s_6ns_6_2_1_U10.din0 ;
wire [5:0] \add_6s_6ns_6_2_1_U10.din1 ;
wire [5:0] \add_6s_6ns_6_2_1_U10.dout ;
wire \add_6s_6ns_6_2_1_U10.reset ;
wire [5:0] \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.a ;
wire [5:0] \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.ain_s0 ;
wire [5:0] \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.b ;
wire [5:0] \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.bin_s0 ;
wire \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.ce ;
wire \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.clk ;
wire \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.facout_s1 ;
wire \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.facout_s2 ;
wire [2:0] \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.fas_s1 ;
wire [2:0] \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.fas_s2 ;
wire \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.reset ;
wire [5:0] \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.s ;
wire [2:0] \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.u1.a ;
wire [2:0] \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.u1.b ;
wire \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.u1.cin ;
wire \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.u1.cout ;
wire [2:0] \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.u1.s ;
wire [2:0] \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.u2.a ;
wire [2:0] \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.u2.b ;
wire \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.u2.cin ;
wire \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.u2.cout ;
wire [2:0] \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.u2.s ;
wire \add_8s_8s_8_2_1_U9.ce ;
wire \add_8s_8s_8_2_1_U9.clk ;
wire [7:0] \add_8s_8s_8_2_1_U9.din0 ;
wire [7:0] \add_8s_8s_8_2_1_U9.din1 ;
wire [7:0] \add_8s_8s_8_2_1_U9.dout ;
wire \add_8s_8s_8_2_1_U9.reset ;
wire [7:0] \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.a ;
wire [7:0] \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.ain_s0 ;
wire [7:0] \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.b ;
wire [7:0] \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.bin_s0 ;
wire \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.ce ;
wire \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.clk ;
wire \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.facout_s1 ;
wire \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.facout_s2 ;
wire [3:0] \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.fas_s1 ;
wire [3:0] \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.fas_s2 ;
wire \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.reset ;
wire [7:0] \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.s ;
wire [3:0] \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.u1.a ;
wire [3:0] \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.u1.b ;
wire \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.u1.cin ;
wire \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.u1.cout ;
wire [3:0] \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.u1.s ;
wire [3:0] \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.u2.a ;
wire [3:0] \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.u2.b ;
wire \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.u2.cin ;
wire \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.u2.cout ;
wire [3:0] \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.u2.s ;
wire ap_CS_fsm_state1;
wire ap_CS_fsm_state10;
wire ap_CS_fsm_state11;
wire ap_CS_fsm_state12;
wire ap_CS_fsm_state13;
wire ap_CS_fsm_state14;
wire ap_CS_fsm_state15;
wire ap_CS_fsm_state16;
wire ap_CS_fsm_state17;
wire ap_CS_fsm_state18;
wire ap_CS_fsm_state19;
wire ap_CS_fsm_state2;
wire ap_CS_fsm_state20;
wire ap_CS_fsm_state21;
wire ap_CS_fsm_state22;
wire ap_CS_fsm_state23;
wire ap_CS_fsm_state24;
wire ap_CS_fsm_state25;
wire ap_CS_fsm_state26;
wire ap_CS_fsm_state27;
wire ap_CS_fsm_state28;
wire ap_CS_fsm_state29;
wire ap_CS_fsm_state3;
wire ap_CS_fsm_state30;
wire ap_CS_fsm_state31;
wire ap_CS_fsm_state32;
wire ap_CS_fsm_state33;
wire ap_CS_fsm_state34;
wire ap_CS_fsm_state35;
wire ap_CS_fsm_state36;
wire ap_CS_fsm_state37;
wire ap_CS_fsm_state4;
wire ap_CS_fsm_state5;
wire [36:0] ap_NS_fsm;
wire ap_clk;
wire ap_done;
wire ap_idle;
wire ap_ready;
wire ap_rst;
wire ap_start;
wire \ashr_32s_32s_32_7_1_U5.ce ;
wire \ashr_32s_32s_32_7_1_U5.clk ;
wire [31:0] \ashr_32s_32s_32_7_1_U5.din0 ;
wire [31:0] \ashr_32s_32s_32_7_1_U5.din1 ;
wire [31:0] \ashr_32s_32s_32_7_1_U5.din1_cast ;
wire [31:0] \ashr_32s_32s_32_7_1_U5.din1_mask ;
wire [31:0] \ashr_32s_32s_32_7_1_U5.dout ;
wire \ashr_32s_32s_32_7_1_U5.reset ;
wire [3:0] grp_fu_221_p2;
wire [3:0] grp_fu_249_p2;
wire [4:0] grp_fu_265_p1;
wire [4:0] grp_fu_265_p2;
wire [4:0] grp_fu_279_p1;
wire [4:0] grp_fu_279_p2;
wire [31:0] grp_fu_295_p1;
wire [31:0] grp_fu_295_p2;
wire [31:0] grp_fu_304_p1;
wire [31:0] grp_fu_304_p2;
wire [16:0] grp_fu_330_p0;
wire [16:0] grp_fu_330_p1;
wire [16:0] grp_fu_330_p2;
wire [3:0] grp_fu_355_p2;
wire [7:0] grp_fu_402_p0;
wire [7:0] grp_fu_402_p1;
wire [7:0] grp_fu_402_p2;
wire [5:0] grp_fu_467_p0;
wire [5:0] grp_fu_467_p2;
wire [33:0] grp_fu_547_p0;
wire [33:0] grp_fu_547_p1;
wire [33:0] grp_fu_547_p2;
wire [31:0] grp_fu_563_p2;
wire [35:0] grp_fu_622_p0;
wire [35:0] grp_fu_622_p1;
wire [35:0] grp_fu_622_p2;
wire [16:0] grp_fu_642_p0;
wire [16:0] grp_fu_642_p1;
wire [16:0] grp_fu_642_p2;
wire [31:0] grp_fu_661_p0;
wire [31:0] grp_fu_661_p2;
wire [1:0] grp_fu_675_p1;
wire [1:0] grp_fu_675_p2;
wire [35:0] grp_fu_698_p0;
wire [35:0] grp_fu_698_p1;
wire [35:0] grp_fu_698_p2;
wire [31:0] grp_fu_725_p1;
wire [31:0] grp_fu_725_p2;
wire [3:0] grp_fu_730_p0;
wire [3:0] grp_fu_730_p1;
wire [3:0] grp_fu_730_p2;
wire [31:0] grp_fu_739_p0;
wire [31:0] grp_fu_739_p2;
wire icmp_ln768_fu_459_p2;
wire icmp_ln851_1_fu_412_p2;
wire icmp_ln851_fu_350_p2;
wire [3:0] icmp_ln890_fu_287_p0;
wire icmp_ln890_fu_287_p2;
wire \mul_4s_4s_4_7_1_U2.ce ;
wire \mul_4s_4s_4_7_1_U2.clk ;
wire [3:0] \mul_4s_4s_4_7_1_U2.din0 ;
wire [3:0] \mul_4s_4s_4_7_1_U2.din1 ;
wire [3:0] \mul_4s_4s_4_7_1_U2.dout ;
wire \mul_4s_4s_4_7_1_U2.reset ;
wire [3:0] \mul_4s_4s_4_7_1_U2.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.a ;
wire [3:0] \mul_4s_4s_4_7_1_U2.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.b ;
wire \mul_4s_4s_4_7_1_U2.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.ce ;
wire \mul_4s_4s_4_7_1_U2.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.clk ;
wire [3:0] \mul_4s_4s_4_7_1_U2.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.p ;
wire [3:0] \mul_4s_4s_4_7_1_U2.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.tmp_product ;
wire [3:0] op_0;
wire [3:0] op_1;
wire [3:0] op_10;
wire [3:0] op_11;
wire [1:0] op_12_V_fu_506_p3;
wire [7:0] op_13_V_fu_604_p3;
wire [1:0] op_18;
wire [3:0] op_19;
wire [31:0] op_29;
wire op_29_ap_vld;
wire [1:0] op_4;
wire [3:0] op_5;
wire [3:0] op_6;
wire [15:0] op_7;
wire or_ln384_fu_502_p2;
wire or_ln785_fu_473_p2;
wire overflow_fu_482_p2;
wire p_Result_5_fu_360_p3;
wire p_Result_6_fu_514_p3;
wire p_Result_7_fu_581_p3;
wire p_Result_9_fu_427_p1;
wire p_Result_s_fu_226_p3;
wire [1:0] p_Val2_4_fu_488_p3;
wire [4:0] p_Val2_s_fu_680_p3;
wire [11:0] r_fu_421_p3;
wire [4:0] ret_V_14_fu_205_p2;
wire [3:0] ret_V_15_fu_572_p1;
wire [3:0] ret_V_15_fu_572_p2;
wire [3:0] ret_V_3_fu_242_p3;
wire [3:0] ret_V_6_fu_577_p1;
wire [3:0] ret_V_6_fu_577_p2;
wire [13:0] rhs_1_fu_319_p3;
wire [6:0] rhs_2_fu_391_p3;
wire [3:0] rhs_fu_197_p1;
wire [4:0] rhs_fu_197_p3;
wire [31:0] select_ln353_1_fu_597_p3;
wire [5:0] select_ln353_fu_526_p3;
wire [1:0] select_ln384_fu_495_p3;
wire [3:0] select_ln850_2_fu_367_p3;
wire [3:0] select_ln850_3_fu_372_p3;
wire [5:0] select_ln850_4_fu_521_p3;
wire [31:0] select_ln850_5_fu_591_p3;
wire [3:0] select_ln850_fu_236_p3;
wire [3:0] sext_ln1192_fu_387_p0;
wire [11:0] sext_ln1497_fu_418_p1;
wire [3:0] sext_ln545_fu_292_p0;
wire [7:0] sext_ln69_2_fu_635_p1;
wire [15:0] sext_ln69_fu_628_p1;
wire [3:0] sext_ln703_1_fu_568_p1;
wire [3:0] sext_ln703_2_fu_275_p0;
wire [3:0] sext_ln703_3_fu_253_p0;
wire [4:0] sext_ln703_3_fu_253_p1;
wire [4:0] sext_ln703_fu_193_p1;
wire [5:0] sext_ln850_fu_464_p1;
wire [31:0] sext_ln890_fu_284_p1;
wire \shl_32s_32s_32_7_1_U6.ce ;
wire \shl_32s_32s_32_7_1_U6.clk ;
wire [31:0] \shl_32s_32s_32_7_1_U6.din0 ;
wire [31:0] \shl_32s_32s_32_7_1_U6.din1 ;
wire [31:0] \shl_32s_32s_32_7_1_U6.din1_cast ;
wire [31:0] \shl_32s_32s_32_7_1_U6.din1_mask ;
wire [31:0] \shl_32s_32s_32_7_1_U6.dout ;
wire \shl_32s_32s_32_7_1_U6.reset ;
wire [3:0] signbit_fu_310_p1;
wire signbit_fu_310_p2;
wire \sub_2ns_2ns_2_2_1_U16.ce ;
wire \sub_2ns_2ns_2_2_1_U16.clk ;
wire [1:0] \sub_2ns_2ns_2_2_1_U16.din0 ;
wire [1:0] \sub_2ns_2ns_2_2_1_U16.din1 ;
wire [1:0] \sub_2ns_2ns_2_2_1_U16.dout ;
wire \sub_2ns_2ns_2_2_1_U16.reset ;
wire [1:0] \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.a ;
wire [1:0] \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.ain_s0 ;
wire [1:0] \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.b ;
wire [1:0] \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.bin_s0 ;
wire \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.ce ;
wire \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.clk ;
wire \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.facout_s1 ;
wire \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.facout_s2 ;
wire \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.fas_s1 ;
wire \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.fas_s2 ;
wire \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.reset ;
wire [1:0] \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.s ;
wire \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.u1.a ;
wire \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.u1.b ;
wire \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.u1.cin ;
wire \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.u1.cout ;
wire \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.u1.s ;
wire \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.u2.a ;
wire \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.u2.b ;
wire \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.u2.cin ;
wire \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.u2.cout ;
wire \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.u2.s ;
wire \sub_5ns_5s_5_2_1_U3.ce ;
wire \sub_5ns_5s_5_2_1_U3.clk ;
wire [4:0] \sub_5ns_5s_5_2_1_U3.din0 ;
wire [4:0] \sub_5ns_5s_5_2_1_U3.din1 ;
wire [4:0] \sub_5ns_5s_5_2_1_U3.dout ;
wire \sub_5ns_5s_5_2_1_U3.reset ;
wire [4:0] \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.a ;
wire [4:0] \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.ain_s0 ;
wire [4:0] \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.b ;
wire [4:0] \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.bin_s0 ;
wire \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.ce ;
wire \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.clk ;
wire \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.facout_s1 ;
wire \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.facout_s2 ;
wire [1:0] \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.fas_s1 ;
wire [2:0] \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.fas_s2 ;
wire \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.reset ;
wire [4:0] \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.s ;
wire [1:0] \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.u1.a ;
wire [1:0] \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.u1.b ;
wire \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.u1.cin ;
wire \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.u1.cout ;
wire [1:0] \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.u1.s ;
wire [2:0] \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.u2.a ;
wire [2:0] \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.u2.b ;
wire \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.u2.cin ;
wire \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.u2.cout ;
wire [2:0] \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.u2.s ;
wire [6:0] tmp_6_fu_536_p3;
wire tmp_V_fu_666_p2;
wire [3:0] tmp_fu_257_p1;
wire [1:0] trunc_ln1347_fu_271_p1;
wire [11:0] trunc_ln1497_1_fu_383_p1;
wire [3:0] trunc_ln1497_fu_379_p1;
wire [12:0] trunc_ln851_1_fu_346_p1;
wire [3:0] trunc_ln851_2_fu_408_p0;
wire [2:0] trunc_ln851_2_fu_408_p1;
wire trunc_ln851_3_fu_588_p1;
wire trunc_ln851_fu_233_p1;
wire xor_ln785_fu_477_p2;


assign _048_ = ap_CS_fsm[20] & icmp_ln851_1_reg_907;
assign _049_ = tmp_reg_788 & ap_CS_fsm[17];
assign _050_ = _053_ & ap_CS_fsm[17];
assign _051_ = _054_ & ap_CS_fsm[0];
assign _052_ = ap_start & ap_CS_fsm[0];
assign overflow_fu_482_p2 = xor_ln785_fu_477_p2 & or_ln785_fu_473_p2;
assign ret_V_15_fu_572_p2 = $signed(op_4) & $signed(op_6);
assign xor_ln785_fu_477_p2 = ~ p_Result_8_reg_918;
assign tmp_V_fu_666_p2 = ~ icmp_ln890_reg_820;
assign _053_ = ~ tmp_reg_788;
assign _054_ = ~ ap_start;
assign _055_ = ! trunc_ln851_1_reg_867;
always @(posedge \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.clk )
\add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.bin_s1  <= _057_;
always @(posedge \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.clk )
\add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.ain_s1  <= _056_;
always @(posedge \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.clk )
\add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.sum_s1  <= _059_;
always @(posedge \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.clk )
\add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.carry_s1  <= _058_;
assign _057_ = \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.ce  ? \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.b [16:8] : \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.bin_s1 ;
assign _056_ = \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.ce  ? \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.a [16:8] : \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.ain_s1 ;
assign _058_ = \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.ce  ? \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.facout_s1  : \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.carry_s1 ;
assign _059_ = \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.ce  ? \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.fas_s1  : \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.sum_s1 ;
assign _060_ = \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.u1.a  + \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.u1.b ;
assign { \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.u1.cout , \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.u1.s  } = _060_ + \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.u1.cin ;
assign _061_ = \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.u2.a  + \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.u2.b ;
assign { \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.u2.cout , \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.u2.s  } = _061_ + \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.u2.cin ;
always @(posedge \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.clk )
\add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.bin_s1  <= _063_;
always @(posedge \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.clk )
\add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.ain_s1  <= _062_;
always @(posedge \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.clk )
\add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.sum_s1  <= _065_;
always @(posedge \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.clk )
\add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.carry_s1  <= _064_;
assign _063_ = \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.ce  ? \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.b [16:8] : \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.bin_s1 ;
assign _062_ = \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.ce  ? \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.a [16:8] : \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.ain_s1 ;
assign _064_ = \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.ce  ? \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.facout_s1  : \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.carry_s1 ;
assign _065_ = \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.ce  ? \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.fas_s1  : \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.sum_s1 ;
assign _066_ = \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.u1.a  + \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.u1.b ;
assign { \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.u1.cout , \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.u1.s  } = _066_ + \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.u1.cin ;
assign _067_ = \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.u2.a  + \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.u2.b ;
assign { \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.u2.cout , \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.u2.s  } = _067_ + \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.u2.cin ;
always @(posedge \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.clk )
\add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s1  <= _069_;
always @(posedge \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.clk )
\add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s1  <= _068_;
always @(posedge \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.clk )
\add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.sum_s1  <= _071_;
always @(posedge \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.clk )
\add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.carry_s1  <= _070_;
assign _069_ = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.ce  ? \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.b [31:16] : \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s1 ;
assign _068_ = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.ce  ? \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.a [31:16] : \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s1 ;
assign _070_ = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.ce  ? \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.facout_s1  : \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.carry_s1 ;
assign _071_ = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.ce  ? \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s1  : \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.sum_s1 ;
assign _072_ = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.a  + \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.b ;
assign { \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cout , \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.s  } = _072_ + \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cin ;
assign _073_ = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.a  + \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.b ;
assign { \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cout , \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.s  } = _073_ + \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cin ;
always @(posedge \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.clk )
\add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s1  <= _075_;
always @(posedge \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.clk )
\add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s1  <= _074_;
always @(posedge \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.clk )
\add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.sum_s1  <= _077_;
always @(posedge \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.clk )
\add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.carry_s1  <= _076_;
assign _075_ = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.ce  ? \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.b [31:16] : \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s1 ;
assign _074_ = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.ce  ? \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.a [31:16] : \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s1 ;
assign _076_ = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.ce  ? \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.facout_s1  : \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.carry_s1 ;
assign _077_ = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.ce  ? \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s1  : \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.sum_s1 ;
assign _078_ = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.a  + \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.b ;
assign { \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cout , \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.s  } = _078_ + \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cin ;
assign _079_ = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.a  + \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.b ;
assign { \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cout , \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.s  } = _079_ + \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cin ;
always @(posedge \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.clk )
\add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.bin_s1  <= _081_;
always @(posedge \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.clk )
\add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.ain_s1  <= _080_;
always @(posedge \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.clk )
\add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.sum_s1  <= _083_;
always @(posedge \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.clk )
\add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.carry_s1  <= _082_;
assign _081_ = \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.ce  ? \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.b [31:16] : \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.bin_s1 ;
assign _080_ = \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.ce  ? \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.a [31:16] : \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.ain_s1 ;
assign _082_ = \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.ce  ? \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.facout_s1  : \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.carry_s1 ;
assign _083_ = \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.ce  ? \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.fas_s1  : \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.sum_s1 ;
assign _084_ = \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.u1.a  + \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.u1.b ;
assign { \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.u1.cout , \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.u1.s  } = _084_ + \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.u1.cin ;
assign _085_ = \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.u2.a  + \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.u2.b ;
assign { \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.u2.cout , \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.u2.s  } = _085_ + \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.u2.cin ;
always @(posedge \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.clk )
\add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.bin_s1  <= _087_;
always @(posedge \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.clk )
\add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.ain_s1  <= _086_;
always @(posedge \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.clk )
\add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.sum_s1  <= _089_;
always @(posedge \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.clk )
\add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.carry_s1  <= _088_;
assign _087_ = \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.ce  ? \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.b [31:16] : \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.bin_s1 ;
assign _086_ = \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.ce  ? \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.a [31:16] : \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.ain_s1 ;
assign _088_ = \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.ce  ? \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.facout_s1  : \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.carry_s1 ;
assign _089_ = \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.ce  ? \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.fas_s1  : \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.sum_s1 ;
assign _090_ = \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.u1.a  + \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.u1.b ;
assign { \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.u1.cout , \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.u1.s  } = _090_ + \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.u1.cin ;
assign _091_ = \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.u2.a  + \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.u2.b ;
assign { \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.u2.cout , \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.u2.s  } = _091_ + \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.u2.cin ;
always @(posedge \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.clk )
\add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.bin_s1  <= _093_;
always @(posedge \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.clk )
\add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.ain_s1  <= _092_;
always @(posedge \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.clk )
\add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.sum_s1  <= _095_;
always @(posedge \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.clk )
\add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.carry_s1  <= _094_;
assign _093_ = \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.ce  ? \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.b [33:17] : \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.bin_s1 ;
assign _092_ = \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.ce  ? \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.a [33:17] : \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.ain_s1 ;
assign _094_ = \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.ce  ? \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.facout_s1  : \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.carry_s1 ;
assign _095_ = \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.ce  ? \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.fas_s1  : \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.sum_s1 ;
assign _096_ = \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.u1.a  + \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.u1.b ;
assign { \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.u1.cout , \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.u1.s  } = _096_ + \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.u1.cin ;
assign _097_ = \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.u2.a  + \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.u2.b ;
assign { \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.u2.cout , \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.u2.s  } = _097_ + \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.u2.cin ;
always @(posedge \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.clk )
\add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.bin_s1  <= _099_;
always @(posedge \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.clk )
\add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.ain_s1  <= _098_;
always @(posedge \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.clk )
\add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.sum_s1  <= _101_;
always @(posedge \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.clk )
\add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.carry_s1  <= _100_;
assign _099_ = \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.ce  ? \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.b [35:18] : \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.bin_s1 ;
assign _098_ = \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.ce  ? \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.a [35:18] : \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.ain_s1 ;
assign _100_ = \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.ce  ? \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.facout_s1  : \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.carry_s1 ;
assign _101_ = \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.ce  ? \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.fas_s1  : \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.sum_s1 ;
assign _102_ = \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.u1.a  + \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.u1.b ;
assign { \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.u1.cout , \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.u1.s  } = _102_ + \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.u1.cin ;
assign _103_ = \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.u2.a  + \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.u2.b ;
assign { \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.u2.cout , \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.u2.s  } = _103_ + \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.u2.cin ;
always @(posedge \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.clk )
\add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.bin_s1  <= _105_;
always @(posedge \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.clk )
\add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.ain_s1  <= _104_;
always @(posedge \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.clk )
\add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.sum_s1  <= _107_;
always @(posedge \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.clk )
\add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.carry_s1  <= _106_;
assign _105_ = \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.ce  ? \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.b [35:18] : \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.bin_s1 ;
assign _104_ = \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.ce  ? \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.a [35:18] : \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.ain_s1 ;
assign _106_ = \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.ce  ? \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.facout_s1  : \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.carry_s1 ;
assign _107_ = \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.ce  ? \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.fas_s1  : \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.sum_s1 ;
assign _108_ = \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.u1.a  + \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.u1.b ;
assign { \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.u1.cout , \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.u1.s  } = _108_ + \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.u1.cin ;
assign _109_ = \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.u2.a  + \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.u2.b ;
assign { \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.u2.cout , \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.u2.s  } = _109_ + \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.u2.cin ;
always @(posedge \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.clk )
\add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.bin_s1  <= _111_;
always @(posedge \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.clk )
\add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.ain_s1  <= _110_;
always @(posedge \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.clk )
\add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.sum_s1  <= _113_;
always @(posedge \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.clk )
\add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.carry_s1  <= _112_;
assign _111_ = \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.ce  ? \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.b [3:2] : \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.bin_s1 ;
assign _110_ = \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.ce  ? \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.a [3:2] : \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.ain_s1 ;
assign _112_ = \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.ce  ? \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.facout_s1  : \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.carry_s1 ;
assign _113_ = \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.ce  ? \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.fas_s1  : \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.sum_s1 ;
assign _114_ = \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.u1.a  + \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.u1.b ;
assign { \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.u1.cout , \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.u1.s  } = _114_ + \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.u1.cin ;
assign _115_ = \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.u2.a  + \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.u2.b ;
assign { \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.u2.cout , \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.u2.s  } = _115_ + \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.u2.cin ;
always @(posedge \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.clk )
\add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.bin_s1  <= _117_;
always @(posedge \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.clk )
\add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.ain_s1  <= _116_;
always @(posedge \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.clk )
\add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.sum_s1  <= _119_;
always @(posedge \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.clk )
\add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.carry_s1  <= _118_;
assign _117_ = \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.ce  ? \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.b [3:2] : \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.bin_s1 ;
assign _116_ = \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.ce  ? \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.a [3:2] : \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.ain_s1 ;
assign _118_ = \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.ce  ? \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.facout_s1  : \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.carry_s1 ;
assign _119_ = \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.ce  ? \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.fas_s1  : \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.sum_s1 ;
assign _120_ = \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.u1.a  + \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.u1.b ;
assign { \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.u1.cout , \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.u1.s  } = _120_ + \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.u1.cin ;
assign _121_ = \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.u2.a  + \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.u2.b ;
assign { \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.u2.cout , \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.u2.s  } = _121_ + \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.u2.cin ;
always @(posedge \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.clk )
\add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.bin_s1  <= _123_;
always @(posedge \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.clk )
\add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.ain_s1  <= _122_;
always @(posedge \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.clk )
\add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.sum_s1  <= _125_;
always @(posedge \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.clk )
\add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.carry_s1  <= _124_;
assign _123_ = \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.ce  ? \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.b [3:2] : \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.bin_s1 ;
assign _122_ = \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.ce  ? \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.a [3:2] : \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.ain_s1 ;
assign _124_ = \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.ce  ? \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.facout_s1  : \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.carry_s1 ;
assign _125_ = \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.ce  ? \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.fas_s1  : \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.sum_s1 ;
assign _126_ = \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.u1.a  + \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.u1.b ;
assign { \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.u1.cout , \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.u1.s  } = _126_ + \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.u1.cin ;
assign _127_ = \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.u2.a  + \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.u2.b ;
assign { \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.u2.cout , \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.u2.s  } = _127_ + \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.u2.cin ;
always @(posedge \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.clk )
\add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.bin_s1  <= _129_;
always @(posedge \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.clk )
\add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.ain_s1  <= _128_;
always @(posedge \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.clk )
\add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.sum_s1  <= _131_;
always @(posedge \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.clk )
\add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.carry_s1  <= _130_;
assign _129_ = \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.ce  ? \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.b [4:2] : \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.bin_s1 ;
assign _128_ = \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.ce  ? \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.a [4:2] : \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.ain_s1 ;
assign _130_ = \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.ce  ? \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.facout_s1  : \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.carry_s1 ;
assign _131_ = \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.ce  ? \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.fas_s1  : \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.sum_s1 ;
assign _132_ = \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.u1.a  + \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.u1.b ;
assign { \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.u1.cout , \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.u1.s  } = _132_ + \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.u1.cin ;
assign _133_ = \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.u2.a  + \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.u2.b ;
assign { \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.u2.cout , \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.u2.s  } = _133_ + \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.u2.cin ;
always @(posedge \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.clk )
\add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.bin_s1  <= _135_;
always @(posedge \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.clk )
\add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.ain_s1  <= _134_;
always @(posedge \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.clk )
\add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.sum_s1  <= _137_;
always @(posedge \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.clk )
\add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.carry_s1  <= _136_;
assign _135_ = \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.ce  ? \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.b [5:3] : \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.bin_s1 ;
assign _134_ = \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.ce  ? \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.a [5:3] : \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.ain_s1 ;
assign _136_ = \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.ce  ? \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.facout_s1  : \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.carry_s1 ;
assign _137_ = \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.ce  ? \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.fas_s1  : \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.sum_s1 ;
assign _138_ = \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.u1.a  + \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.u1.b ;
assign { \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.u1.cout , \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.u1.s  } = _138_ + \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.u1.cin ;
assign _139_ = \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.u2.a  + \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.u2.b ;
assign { \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.u2.cout , \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.u2.s  } = _139_ + \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.u2.cin ;
always @(posedge \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.clk )
\add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.bin_s1  <= _141_;
always @(posedge \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.clk )
\add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.ain_s1  <= _140_;
always @(posedge \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.clk )
\add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.sum_s1  <= _143_;
always @(posedge \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.clk )
\add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.carry_s1  <= _142_;
assign _141_ = \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.ce  ? \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.b [7:4] : \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.bin_s1 ;
assign _140_ = \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.ce  ? \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.a [7:4] : \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.ain_s1 ;
assign _142_ = \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.ce  ? \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.facout_s1  : \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.carry_s1 ;
assign _143_ = \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.ce  ? \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.fas_s1  : \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.sum_s1 ;
assign _144_ = \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.u1.a  + \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.u1.b ;
assign { \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.u1.cout , \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.u1.s  } = _144_ + \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.u1.cin ;
assign _145_ = \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.u2.a  + \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.u2.b ;
assign { \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.u2.cout , \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.u2.s  } = _145_ + \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.u2.cin ;
always @(posedge \ashr_32s_32s_32_7_1_U5.clk )
\ashr_32s_32s_32_7_1_U5.dout_array[5]  <= _157_;
always @(posedge \ashr_32s_32s_32_7_1_U5.clk )
\ashr_32s_32s_32_7_1_U5.din1_cast_array[5]  <= _151_;
always @(posedge \ashr_32s_32s_32_7_1_U5.clk )
\ashr_32s_32s_32_7_1_U5.dout_array[4]  <= _156_;
always @(posedge \ashr_32s_32s_32_7_1_U5.clk )
\ashr_32s_32s_32_7_1_U5.din1_cast_array[4]  <= _150_;
always @(posedge \ashr_32s_32s_32_7_1_U5.clk )
\ashr_32s_32s_32_7_1_U5.dout_array[3]  <= _155_;
always @(posedge \ashr_32s_32s_32_7_1_U5.clk )
\ashr_32s_32s_32_7_1_U5.din1_cast_array[3]  <= _149_;
always @(posedge \ashr_32s_32s_32_7_1_U5.clk )
\ashr_32s_32s_32_7_1_U5.dout_array[2]  <= _154_;
always @(posedge \ashr_32s_32s_32_7_1_U5.clk )
\ashr_32s_32s_32_7_1_U5.din1_cast_array[2]  <= _148_;
always @(posedge \ashr_32s_32s_32_7_1_U5.clk )
\ashr_32s_32s_32_7_1_U5.dout_array[1]  <= _153_;
always @(posedge \ashr_32s_32s_32_7_1_U5.clk )
\ashr_32s_32s_32_7_1_U5.din1_cast_array[1]  <= _147_;
always @(posedge \ashr_32s_32s_32_7_1_U5.clk )
\ashr_32s_32s_32_7_1_U5.dout_array[0]  <= _152_;
always @(posedge \ashr_32s_32s_32_7_1_U5.clk )
\ashr_32s_32s_32_7_1_U5.din1_cast_array[0]  <= _146_;
assign _158_ = \ashr_32s_32s_32_7_1_U5.ce  ? \ashr_32s_32s_32_7_1_U5.din1_cast_array[4]  : \ashr_32s_32s_32_7_1_U5.din1_cast_array[5] ;
assign _151_ = \ashr_32s_32s_32_7_1_U5.reset  ? 32'd0 : _158_;
assign _159_ = \ashr_32s_32s_32_7_1_U5.ce  ? _175_ : \ashr_32s_32s_32_7_1_U5.dout_array[5] ;
assign _157_ = \ashr_32s_32s_32_7_1_U5.reset  ? 32'd0 : _159_;
assign _160_ = \ashr_32s_32s_32_7_1_U5.ce  ? \ashr_32s_32s_32_7_1_U5.din1_cast_array[3]  : \ashr_32s_32s_32_7_1_U5.din1_cast_array[4] ;
assign _150_ = \ashr_32s_32s_32_7_1_U5.reset  ? 32'd0 : _160_;
assign _161_ = \ashr_32s_32s_32_7_1_U5.ce  ? _174_ : \ashr_32s_32s_32_7_1_U5.dout_array[4] ;
assign _156_ = \ashr_32s_32s_32_7_1_U5.reset  ? 32'd0 : _161_;
assign _162_ = \ashr_32s_32s_32_7_1_U5.ce  ? \ashr_32s_32s_32_7_1_U5.din1_cast_array[2]  : \ashr_32s_32s_32_7_1_U5.din1_cast_array[3] ;
assign _149_ = \ashr_32s_32s_32_7_1_U5.reset  ? 32'd0 : _162_;
assign _163_ = \ashr_32s_32s_32_7_1_U5.ce  ? _173_ : \ashr_32s_32s_32_7_1_U5.dout_array[3] ;
assign _155_ = \ashr_32s_32s_32_7_1_U5.reset  ? 32'd0 : _163_;
assign _164_ = \ashr_32s_32s_32_7_1_U5.ce  ? \ashr_32s_32s_32_7_1_U5.din1_cast_array[1]  : \ashr_32s_32s_32_7_1_U5.din1_cast_array[2] ;
assign _148_ = \ashr_32s_32s_32_7_1_U5.reset  ? 32'd0 : _164_;
assign _165_ = \ashr_32s_32s_32_7_1_U5.ce  ? _172_ : \ashr_32s_32s_32_7_1_U5.dout_array[2] ;
assign _154_ = \ashr_32s_32s_32_7_1_U5.reset  ? 32'd0 : _165_;
assign _166_ = \ashr_32s_32s_32_7_1_U5.ce  ? \ashr_32s_32s_32_7_1_U5.din1_cast_array[0]  : \ashr_32s_32s_32_7_1_U5.din1_cast_array[1] ;
assign _147_ = \ashr_32s_32s_32_7_1_U5.reset  ? 32'd0 : _166_;
assign _167_ = \ashr_32s_32s_32_7_1_U5.ce  ? _171_ : \ashr_32s_32s_32_7_1_U5.dout_array[1] ;
assign _153_ = \ashr_32s_32s_32_7_1_U5.reset  ? 32'd0 : _167_;
assign _168_ = \ashr_32s_32s_32_7_1_U5.ce  ? \ashr_32s_32s_32_7_1_U5.din1  : \ashr_32s_32s_32_7_1_U5.din1_cast_array[0] ;
assign _146_ = \ashr_32s_32s_32_7_1_U5.reset  ? 32'd0 : _168_;
assign _169_ = \ashr_32s_32s_32_7_1_U5.ce  ? _170_ : \ashr_32s_32s_32_7_1_U5.dout_array[0] ;
assign _152_ = \ashr_32s_32s_32_7_1_U5.reset  ? 32'd0 : _169_;
assign _170_ = $signed(\ashr_32s_32s_32_7_1_U5.din0 ) >>> { \ashr_32s_32s_32_7_1_U5.din1 [31:30], 30'h00000000 };
assign _171_ = $signed(\ashr_32s_32s_32_7_1_U5.dout_array[0] ) >>> { \ashr_32s_32s_32_7_1_U5.din1_cast_array[0] [29:25], 25'h0000000 };
assign _172_ = $signed(\ashr_32s_32s_32_7_1_U5.dout_array[1] ) >>> { \ashr_32s_32s_32_7_1_U5.din1_cast_array[1] [24:20], 20'h00000 };
assign _173_ = $signed(\ashr_32s_32s_32_7_1_U5.dout_array[2] ) >>> { \ashr_32s_32s_32_7_1_U5.din1_cast_array[2] [19:15], 15'h0000 };
assign _174_ = $signed(\ashr_32s_32s_32_7_1_U5.dout_array[3] ) >>> { \ashr_32s_32s_32_7_1_U5.din1_cast_array[3] [14:10], 10'h000 };
assign _175_ = $signed(\ashr_32s_32s_32_7_1_U5.dout_array[4] ) >>> { \ashr_32s_32s_32_7_1_U5.din1_cast_array[4] [9:5], 5'h00 };
assign \ashr_32s_32s_32_7_1_U5.dout  = $signed(\ashr_32s_32s_32_7_1_U5.dout_array[5] ) >>> \ashr_32s_32s_32_7_1_U5.din1_cast_array[5] [4:0];
assign \mul_4s_4s_4_7_1_U2.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.tmp_product  = $signed(\mul_4s_4s_4_7_1_U2.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.a_reg0 ) * $signed(\mul_4s_4s_4_7_1_U2.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.b_reg0 );
always @(posedge \mul_4s_4s_4_7_1_U2.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.clk )
\mul_4s_4s_4_7_1_U2.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.a_reg0  <= _176_;
always @(posedge \mul_4s_4s_4_7_1_U2.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.clk )
\mul_4s_4s_4_7_1_U2.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.b_reg0  <= _177_;
always @(posedge \mul_4s_4s_4_7_1_U2.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.clk )
\mul_4s_4s_4_7_1_U2.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.buff0  <= _178_;
always @(posedge \mul_4s_4s_4_7_1_U2.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.clk )
\mul_4s_4s_4_7_1_U2.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.buff1  <= _179_;
always @(posedge \mul_4s_4s_4_7_1_U2.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.clk )
\mul_4s_4s_4_7_1_U2.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.buff2  <= _180_;
always @(posedge \mul_4s_4s_4_7_1_U2.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.clk )
\mul_4s_4s_4_7_1_U2.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.buff3  <= _181_;
always @(posedge \mul_4s_4s_4_7_1_U2.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.clk )
\mul_4s_4s_4_7_1_U2.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.buff4  <= _182_;
assign _182_ = \mul_4s_4s_4_7_1_U2.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.ce  ? \mul_4s_4s_4_7_1_U2.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.buff3  : \mul_4s_4s_4_7_1_U2.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.buff4 ;
assign _181_ = \mul_4s_4s_4_7_1_U2.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.ce  ? \mul_4s_4s_4_7_1_U2.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.buff2  : \mul_4s_4s_4_7_1_U2.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.buff3 ;
assign _180_ = \mul_4s_4s_4_7_1_U2.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.ce  ? \mul_4s_4s_4_7_1_U2.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.buff1  : \mul_4s_4s_4_7_1_U2.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.buff2 ;
assign _179_ = \mul_4s_4s_4_7_1_U2.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.ce  ? \mul_4s_4s_4_7_1_U2.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.buff0  : \mul_4s_4s_4_7_1_U2.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.buff1 ;
assign _178_ = \mul_4s_4s_4_7_1_U2.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.ce  ? \mul_4s_4s_4_7_1_U2.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.tmp_product  : \mul_4s_4s_4_7_1_U2.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.buff0 ;
assign _177_ = \mul_4s_4s_4_7_1_U2.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.ce  ? \mul_4s_4s_4_7_1_U2.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.b  : \mul_4s_4s_4_7_1_U2.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.b_reg0 ;
assign _176_ = \mul_4s_4s_4_7_1_U2.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.ce  ? \mul_4s_4s_4_7_1_U2.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.a  : \mul_4s_4s_4_7_1_U2.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.a_reg0 ;
always @(posedge \shl_32s_32s_32_7_1_U6.clk )
\shl_32s_32s_32_7_1_U6.dout_array[5]  <= _194_;
always @(posedge \shl_32s_32s_32_7_1_U6.clk )
\shl_32s_32s_32_7_1_U6.din1_cast_array[5]  <= _188_;
always @(posedge \shl_32s_32s_32_7_1_U6.clk )
\shl_32s_32s_32_7_1_U6.dout_array[4]  <= _193_;
always @(posedge \shl_32s_32s_32_7_1_U6.clk )
\shl_32s_32s_32_7_1_U6.din1_cast_array[4]  <= _187_;
always @(posedge \shl_32s_32s_32_7_1_U6.clk )
\shl_32s_32s_32_7_1_U6.dout_array[3]  <= _192_;
always @(posedge \shl_32s_32s_32_7_1_U6.clk )
\shl_32s_32s_32_7_1_U6.din1_cast_array[3]  <= _186_;
always @(posedge \shl_32s_32s_32_7_1_U6.clk )
\shl_32s_32s_32_7_1_U6.dout_array[2]  <= _191_;
always @(posedge \shl_32s_32s_32_7_1_U6.clk )
\shl_32s_32s_32_7_1_U6.din1_cast_array[2]  <= _185_;
always @(posedge \shl_32s_32s_32_7_1_U6.clk )
\shl_32s_32s_32_7_1_U6.dout_array[1]  <= _190_;
always @(posedge \shl_32s_32s_32_7_1_U6.clk )
\shl_32s_32s_32_7_1_U6.din1_cast_array[1]  <= _184_;
always @(posedge \shl_32s_32s_32_7_1_U6.clk )
\shl_32s_32s_32_7_1_U6.dout_array[0]  <= _189_;
always @(posedge \shl_32s_32s_32_7_1_U6.clk )
\shl_32s_32s_32_7_1_U6.din1_cast_array[0]  <= _183_;
assign _195_ = \shl_32s_32s_32_7_1_U6.ce  ? \shl_32s_32s_32_7_1_U6.din1_cast_array[4]  : \shl_32s_32s_32_7_1_U6.din1_cast_array[5] ;
assign _188_ = \shl_32s_32s_32_7_1_U6.reset  ? 32'd0 : _195_;
assign _196_ = \shl_32s_32s_32_7_1_U6.ce  ? _212_ : \shl_32s_32s_32_7_1_U6.dout_array[5] ;
assign _194_ = \shl_32s_32s_32_7_1_U6.reset  ? 32'd0 : _196_;
assign _197_ = \shl_32s_32s_32_7_1_U6.ce  ? \shl_32s_32s_32_7_1_U6.din1_cast_array[3]  : \shl_32s_32s_32_7_1_U6.din1_cast_array[4] ;
assign _187_ = \shl_32s_32s_32_7_1_U6.reset  ? 32'd0 : _197_;
assign _198_ = \shl_32s_32s_32_7_1_U6.ce  ? _211_ : \shl_32s_32s_32_7_1_U6.dout_array[4] ;
assign _193_ = \shl_32s_32s_32_7_1_U6.reset  ? 32'd0 : _198_;
assign _199_ = \shl_32s_32s_32_7_1_U6.ce  ? \shl_32s_32s_32_7_1_U6.din1_cast_array[2]  : \shl_32s_32s_32_7_1_U6.din1_cast_array[3] ;
assign _186_ = \shl_32s_32s_32_7_1_U6.reset  ? 32'd0 : _199_;
assign _200_ = \shl_32s_32s_32_7_1_U6.ce  ? _210_ : \shl_32s_32s_32_7_1_U6.dout_array[3] ;
assign _192_ = \shl_32s_32s_32_7_1_U6.reset  ? 32'd0 : _200_;
assign _201_ = \shl_32s_32s_32_7_1_U6.ce  ? \shl_32s_32s_32_7_1_U6.din1_cast_array[1]  : \shl_32s_32s_32_7_1_U6.din1_cast_array[2] ;
assign _185_ = \shl_32s_32s_32_7_1_U6.reset  ? 32'd0 : _201_;
assign _202_ = \shl_32s_32s_32_7_1_U6.ce  ? _209_ : \shl_32s_32s_32_7_1_U6.dout_array[2] ;
assign _191_ = \shl_32s_32s_32_7_1_U6.reset  ? 32'd0 : _202_;
assign _203_ = \shl_32s_32s_32_7_1_U6.ce  ? \shl_32s_32s_32_7_1_U6.din1_cast_array[0]  : \shl_32s_32s_32_7_1_U6.din1_cast_array[1] ;
assign _184_ = \shl_32s_32s_32_7_1_U6.reset  ? 32'd0 : _203_;
assign _204_ = \shl_32s_32s_32_7_1_U6.ce  ? _208_ : \shl_32s_32s_32_7_1_U6.dout_array[1] ;
assign _190_ = \shl_32s_32s_32_7_1_U6.reset  ? 32'd0 : _204_;
assign _205_ = \shl_32s_32s_32_7_1_U6.ce  ? \shl_32s_32s_32_7_1_U6.din1  : \shl_32s_32s_32_7_1_U6.din1_cast_array[0] ;
assign _183_ = \shl_32s_32s_32_7_1_U6.reset  ? 32'd0 : _205_;
assign _206_ = \shl_32s_32s_32_7_1_U6.ce  ? _207_ : \shl_32s_32s_32_7_1_U6.dout_array[0] ;
assign _189_ = \shl_32s_32s_32_7_1_U6.reset  ? 32'd0 : _206_;
assign _207_ = \shl_32s_32s_32_7_1_U6.din0  << { \shl_32s_32s_32_7_1_U6.din1 [31:30], 30'h00000000 };
assign _208_ = \shl_32s_32s_32_7_1_U6.dout_array[0]  << { \shl_32s_32s_32_7_1_U6.din1_cast_array[0] [29:25], 25'h0000000 };
assign _209_ = \shl_32s_32s_32_7_1_U6.dout_array[1]  << { \shl_32s_32s_32_7_1_U6.din1_cast_array[1] [24:20], 20'h00000 };
assign _210_ = \shl_32s_32s_32_7_1_U6.dout_array[2]  << { \shl_32s_32s_32_7_1_U6.din1_cast_array[2] [19:15], 15'h0000 };
assign _211_ = \shl_32s_32s_32_7_1_U6.dout_array[3]  << { \shl_32s_32s_32_7_1_U6.din1_cast_array[3] [14:10], 10'h000 };
assign _212_ = \shl_32s_32s_32_7_1_U6.dout_array[4]  << { \shl_32s_32s_32_7_1_U6.din1_cast_array[4] [9:5], 5'h00 };
assign \shl_32s_32s_32_7_1_U6.dout  = \shl_32s_32s_32_7_1_U6.dout_array[5]  << \shl_32s_32s_32_7_1_U6.din1_cast_array[5] [4:0];
assign \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.bin_s0  = ~ \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.b ;
always @(posedge \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.clk )
\sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.bin_s1  <= _214_;
always @(posedge \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.clk )
\sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.ain_s1  <= _213_;
always @(posedge \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.clk )
\sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.sum_s1  <= _216_;
always @(posedge \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.clk )
\sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.carry_s1  <= _215_;
assign _214_ = \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.ce  ? \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.bin_s0 [1] : \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.bin_s1 ;
assign _213_ = \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.ce  ? \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.a [1] : \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.ain_s1 ;
assign _215_ = \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.ce  ? \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.facout_s1  : \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.carry_s1 ;
assign _216_ = \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.ce  ? \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.fas_s1  : \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.sum_s1 ;
assign _217_ = \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.u1.a  + \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.u1.b ;
assign { \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.u1.cout , \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.u1.s  } = _217_ + \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.u1.cin ;
assign _218_ = \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.u2.a  + \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.u2.b ;
assign { \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.u2.cout , \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.u2.s  } = _218_ + \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.u2.cin ;
assign \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.bin_s0  = ~ \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.b ;
always @(posedge \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.clk )
\sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.bin_s1  <= _220_;
always @(posedge \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.clk )
\sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.ain_s1  <= _219_;
always @(posedge \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.clk )
\sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.sum_s1  <= _222_;
always @(posedge \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.clk )
\sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.carry_s1  <= _221_;
assign _220_ = \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.ce  ? \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.bin_s0 [4:2] : \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.bin_s1 ;
assign _219_ = \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.ce  ? \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.a [4:2] : \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.ain_s1 ;
assign _221_ = \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.ce  ? \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.facout_s1  : \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.carry_s1 ;
assign _222_ = \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.ce  ? \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.fas_s1  : \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.sum_s1 ;
assign _223_ = \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.u1.a  + \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.u1.b ;
assign { \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.u1.cout , \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.u1.s  } = _223_ + \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.u1.cin ;
assign _224_ = \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.u2.a  + \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.u2.b ;
assign { \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.u2.cout , \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.u2.s  } = _224_ + \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.u2.cin ;
assign _225_ = $signed(op_5) < $signed(ret_V_3_reg_768);
assign _226_ = | tmp_1_reg_924;
assign _227_ = | op_10[2:0];
assign _228_ = op_3_V_reg_793 != op_5;
assign or_ln384_fu_502_p2 = p_Result_8_reg_918 | overflow_reg_951;
assign or_ln785_fu_473_p2 = p_Result_9_reg_912 | icmp_ln768_reg_939;
assign ret_V_6_fu_577_p2 = op_6 | op_3_V_reg_793;
always @(posedge ap_clk)
trunc_ln1497_reg_887 <= _045_;
always @(posedge ap_clk)
trunc_ln1497_1_reg_892 <= _044_;
always @(posedge ap_clk)
sext_ln703_3_reg_782 <= _035_;
always @(posedge ap_clk)
tmp_reg_788 <= _042_;
always @(posedge ap_clk)
select_ln850_3_reg_882 <= _034_;
always @(posedge ap_clk)
ret_V_9_reg_877 <= _030_;
always @(posedge ap_clk)
ret_V_3_reg_768 <= _027_;
always @(posedge ap_clk)
ret_V_2_reg_763 <= _026_;
always @(posedge ap_clk)
ret_V_19_reg_983 <= _024_;
always @(posedge ap_clk)
ret_V_21_cast_reg_988 <= _025_;
always @(posedge ap_clk)
ret_V_17_reg_855 <= _022_;
always @(posedge ap_clk)
ret_V_7_reg_860 <= _029_;
always @(posedge ap_clk)
trunc_ln851_1_reg_867 <= _046_;
always @(posedge ap_clk)
ret_V_16_reg_840 <= _021_;
always @(posedge ap_clk)
ret_V_15_reg_1000 <= _020_;
always @(posedge ap_clk)
ret_V_6_reg_1005 <= _028_;
always @(posedge ap_clk)
select_ln353_1_reg_1010 <= _032_;
always @(posedge ap_clk)
ret_V_14_reg_750 <= _019_;
always @(posedge ap_clk)
ret_V_reg_756 <= _031_;
always @(posedge ap_clk)
p_Result_9_reg_912 <= _018_;
always @(posedge ap_clk)
p_Result_8_reg_918 <= _017_;
always @(posedge ap_clk)
tmp_1_reg_924 <= _039_;
always @(posedge ap_clk)
ret_V_18_reg_929 <= _023_;
always @(posedge ap_clk)
tmp_2_reg_934 <= _040_;
always @(posedge ap_clk)
overflow_reg_951 <= _016_;
always @(posedge ap_clk)
op_3_V_reg_793 <= _015_;
always @(posedge ap_clk)
sub_ln1497_reg_799 <= _038_;
always @(posedge ap_clk)
trunc_ln1347_reg_804 <= _043_;
always @(posedge ap_clk)
tmp_V_reg_1050 <= _041_;
always @(posedge ap_clk)
op_25_V_reg_1055 <= _013_;
always @(posedge ap_clk)
op_17_V_reg_1075 <= _011_;
always @(posedge ap_clk)
op_26_V_reg_1080 <= _014_;
always @(posedge ap_clk)
op_12_V_reg_962 <= _010_;
always @(posedge ap_clk)
select_ln353_reg_968 <= _033_;
always @(posedge ap_clk)
icmp_ln890_reg_820 <= _009_;
always @(posedge ap_clk)
signbit_reg_835 <= _037_;
always @(posedge ap_clk)
icmp_ln851_reg_872 <= _008_;
always @(posedge ap_clk)
icmp_ln851_1_reg_907 <= _007_;
always @(posedge ap_clk)
icmp_ln768_reg_939 <= _006_;
always @(posedge ap_clk)
sext_ln850_reg_944 <= _036_;
always @(posedge ap_clk)
op_23_V_reg_1035 <= _012_;
always @(posedge ap_clk)
add_ln69_reg_1040 <= _004_;
always @(posedge ap_clk)
add_ln69_2_reg_1100 <= _002_;
always @(posedge ap_clk)
add_ln69_3_reg_1105 <= _003_;
always @(posedge ap_clk)
add_ln691_reg_957 <= _001_;
always @(posedge ap_clk)
add_ln691_1_reg_995 <= _000_;
always @(posedge ap_clk)
ap_CS_fsm <= _005_;
assign _047_ = _052_ ? 2'h2 : 2'h1;
assign _229_ = ap_CS_fsm == 1'h1;
function [36:0] _641_;
input [36:0] a;
input [1368:0] b;
input [36:0] s;
case (s)
37'b0000000000000000000000000000000000001:
_641_ = b[36:0];
37'b0000000000000000000000000000000000010:
_641_ = b[73:37];
37'b0000000000000000000000000000000000100:
_641_ = b[110:74];
37'b0000000000000000000000000000000001000:
_641_ = b[147:111];
37'b0000000000000000000000000000000010000:
_641_ = b[184:148];
37'b0000000000000000000000000000000100000:
_641_ = b[221:185];
37'b0000000000000000000000000000001000000:
_641_ = b[258:222];
37'b0000000000000000000000000000010000000:
_641_ = b[295:259];
37'b0000000000000000000000000000100000000:
_641_ = b[332:296];
37'b0000000000000000000000000001000000000:
_641_ = b[369:333];
37'b0000000000000000000000000010000000000:
_641_ = b[406:370];
37'b0000000000000000000000000100000000000:
_641_ = b[443:407];
37'b0000000000000000000000001000000000000:
_641_ = b[480:444];
37'b0000000000000000000000010000000000000:
_641_ = b[517:481];
37'b0000000000000000000000100000000000000:
_641_ = b[554:518];
37'b0000000000000000000001000000000000000:
_641_ = b[591:555];
37'b0000000000000000000010000000000000000:
_641_ = b[628:592];
37'b0000000000000000000100000000000000000:
_641_ = b[665:629];
37'b0000000000000000001000000000000000000:
_641_ = b[702:666];
37'b0000000000000000010000000000000000000:
_641_ = b[739:703];
37'b0000000000000000100000000000000000000:
_641_ = b[776:740];
37'b0000000000000001000000000000000000000:
_641_ = b[813:777];
37'b0000000000000010000000000000000000000:
_641_ = b[850:814];
37'b0000000000000100000000000000000000000:
_641_ = b[887:851];
37'b0000000000001000000000000000000000000:
_641_ = b[924:888];
37'b0000000000010000000000000000000000000:
_641_ = b[961:925];
37'b0000000000100000000000000000000000000:
_641_ = b[998:962];
37'b0000000001000000000000000000000000000:
_641_ = b[1035:999];
37'b0000000010000000000000000000000000000:
_641_ = b[1072:1036];
37'b0000000100000000000000000000000000000:
_641_ = b[1109:1073];
37'b0000001000000000000000000000000000000:
_641_ = b[1146:1110];
37'b0000010000000000000000000000000000000:
_641_ = b[1183:1147];
37'b0000100000000000000000000000000000000:
_641_ = b[1220:1184];
37'b0001000000000000000000000000000000000:
_641_ = b[1257:1221];
37'b0010000000000000000000000000000000000:
_641_ = b[1294:1258];
37'b0100000000000000000000000000000000000:
_641_ = b[1331:1295];
37'b1000000000000000000000000000000000000:
_641_ = b[1368:1332];
37'b0000000000000000000000000000000000000:
_641_ = a;
default:
_641_ = 37'bx;
endcase
endfunction
assign ap_NS_fsm = _641_(37'hxxxxxxxxxx, { 35'h000000000, _047_, 1332'h000000002000000002000000002000000002000000002000000002000000002000000002000000002000000002000000002000000002000000002000000002000000002000000002000000002000000002000000002000000002000000002000000002000000002000000002000000002000000002000000002000000002000000002000000002000000002000000002000000002000000002000000002000000000000000001 }, { _229_, _265_, _264_, _263_, _262_, _261_, _260_, _259_, _258_, _257_, _256_, _255_, _254_, _253_, _252_, _251_, _250_, _249_, _248_, _247_, _246_, _245_, _244_, _243_, _242_, _241_, _240_, _239_, _238_, _237_, _236_, _235_, _234_, _233_, _232_, _231_, _230_ });
assign _230_ = ap_CS_fsm == 37'h1000000000;
assign _231_ = ap_CS_fsm == 36'h800000000;
assign _232_ = ap_CS_fsm == 35'h400000000;
assign _233_ = ap_CS_fsm == 34'h200000000;
assign _234_ = ap_CS_fsm == 33'h100000000;
assign _235_ = ap_CS_fsm == 32'd2147483648;
assign _236_ = ap_CS_fsm == 31'h40000000;
assign _237_ = ap_CS_fsm == 30'h20000000;
assign _238_ = ap_CS_fsm == 29'h10000000;
assign _239_ = ap_CS_fsm == 28'h8000000;
assign _240_ = ap_CS_fsm == 27'h4000000;
assign _241_ = ap_CS_fsm == 26'h2000000;
assign _242_ = ap_CS_fsm == 25'h1000000;
assign _243_ = ap_CS_fsm == 24'h800000;
assign _244_ = ap_CS_fsm == 23'h400000;
assign _245_ = ap_CS_fsm == 22'h200000;
assign _246_ = ap_CS_fsm == 21'h100000;
assign _247_ = ap_CS_fsm == 20'h80000;
assign _248_ = ap_CS_fsm == 19'h40000;
assign _249_ = ap_CS_fsm == 18'h20000;
assign _250_ = ap_CS_fsm == 17'h10000;
assign _251_ = ap_CS_fsm == 16'h8000;
assign _252_ = ap_CS_fsm == 15'h4000;
assign _253_ = ap_CS_fsm == 14'h2000;
assign _254_ = ap_CS_fsm == 13'h1000;
assign _255_ = ap_CS_fsm == 12'h800;
assign _256_ = ap_CS_fsm == 11'h400;
assign _257_ = ap_CS_fsm == 10'h200;
assign _258_ = ap_CS_fsm == 9'h100;
assign _259_ = ap_CS_fsm == 8'h80;
assign _260_ = ap_CS_fsm == 7'h40;
assign _261_ = ap_CS_fsm == 6'h20;
assign _262_ = ap_CS_fsm == 5'h10;
assign _263_ = ap_CS_fsm == 4'h8;
assign _264_ = ap_CS_fsm == 3'h4;
assign _265_ = ap_CS_fsm == 2'h2;
assign op_29_ap_vld = ap_CS_fsm[36] ? 1'h1 : 1'h0;
assign ap_idle = _051_ ? 1'h1 : 1'h0;
assign _045_ = _050_ ? grp_fu_295_p2[3:0] : trunc_ln1497_reg_887;
assign _044_ = _049_ ? grp_fu_304_p2[11:0] : trunc_ln1497_1_reg_892;
assign _042_ = ap_CS_fsm[9] ? op_6[3] : tmp_reg_788;
assign _035_ = ap_CS_fsm[9] ? { op_6[3], op_6 } : sext_ln703_3_reg_782;
assign _034_ = ap_CS_fsm[16] ? select_ln850_3_fu_372_p3 : select_ln850_3_reg_882;
assign _030_ = ap_CS_fsm[15] ? grp_fu_355_p2 : ret_V_9_reg_877;
assign _027_ = ap_CS_fsm[3] ? ret_V_3_fu_242_p3 : ret_V_3_reg_768;
assign _026_ = ap_CS_fsm[2] ? grp_fu_221_p2 : ret_V_2_reg_763;
assign _025_ = ap_CS_fsm[23] ? grp_fu_547_p2[32:1] : ret_V_21_cast_reg_988;
assign _024_ = ap_CS_fsm[23] ? grp_fu_547_p2 : ret_V_19_reg_983;
assign _046_ = ap_CS_fsm[13] ? grp_fu_330_p2[12:0] : trunc_ln851_1_reg_867;
assign _029_ = ap_CS_fsm[13] ? grp_fu_330_p2[16:13] : ret_V_7_reg_860;
assign _022_ = ap_CS_fsm[13] ? grp_fu_330_p2 : ret_V_17_reg_855;
assign _021_ = ap_CS_fsm[12] ? grp_fu_279_p2 : ret_V_16_reg_840;
assign _032_ = ap_CS_fsm[26] ? select_ln353_1_fu_597_p3 : select_ln353_1_reg_1010;
assign _028_ = ap_CS_fsm[26] ? ret_V_6_fu_577_p2 : ret_V_6_reg_1005;
assign _020_ = ap_CS_fsm[26] ? ret_V_15_fu_572_p2 : ret_V_15_reg_1000;
assign _031_ = ap_CS_fsm[0] ? ret_V_14_fu_205_p2[4:1] : ret_V_reg_756;
assign _019_ = ap_CS_fsm[0] ? ret_V_14_fu_205_p2 : ret_V_14_reg_750;
assign _040_ = ap_CS_fsm[18] ? grp_fu_402_p2[7:3] : tmp_2_reg_934;
assign _023_ = ap_CS_fsm[18] ? grp_fu_402_p2 : ret_V_18_reg_929;
assign _039_ = ap_CS_fsm[18] ? r_fu_421_p3[11:1] : tmp_1_reg_924;
assign _017_ = ap_CS_fsm[18] ? r_fu_421_p3[11] : p_Result_8_reg_918;
assign _018_ = ap_CS_fsm[18] ? r_fu_421_p3[0] : p_Result_9_reg_912;
assign _016_ = ap_CS_fsm[20] ? overflow_fu_482_p2 : overflow_reg_951;
assign _043_ = ap_CS_fsm[10] ? grp_fu_249_p2[1:0] : trunc_ln1347_reg_804;
assign _038_ = ap_CS_fsm[10] ? grp_fu_265_p2 : sub_ln1497_reg_799;
assign _015_ = ap_CS_fsm[10] ? grp_fu_249_p2 : op_3_V_reg_793;
assign _013_ = ap_CS_fsm[30] ? grp_fu_661_p2 : op_25_V_reg_1055;
assign _041_ = ap_CS_fsm[30] ? tmp_V_fu_666_p2 : tmp_V_reg_1050;
assign _014_ = ap_CS_fsm[32] ? grp_fu_698_p2[35:4] : op_26_V_reg_1080;
assign _011_ = ap_CS_fsm[32] ? grp_fu_675_p2 : op_17_V_reg_1075;
assign _033_ = ap_CS_fsm[21] ? select_ln353_fu_526_p3 : select_ln353_reg_968;
assign _010_ = ap_CS_fsm[21] ? op_12_V_fu_506_p3 : op_12_V_reg_962;
assign _037_ = ap_CS_fsm[11] ? signbit_fu_310_p2 : signbit_reg_835;
assign _009_ = ap_CS_fsm[11] ? icmp_ln890_fu_287_p2 : icmp_ln890_reg_820;
assign _008_ = ap_CS_fsm[14] ? icmp_ln851_fu_350_p2 : icmp_ln851_reg_872;
assign _007_ = ap_CS_fsm[17] ? icmp_ln851_1_fu_412_p2 : icmp_ln851_1_reg_907;
assign _036_ = ap_CS_fsm[19] ? { tmp_2_reg_934[4], tmp_2_reg_934 } : sext_ln850_reg_944;
assign _006_ = ap_CS_fsm[19] ? icmp_ln768_fu_459_p2 : icmp_ln768_reg_939;
assign _004_ = ap_CS_fsm[28] ? grp_fu_642_p2 : add_ln69_reg_1040;
assign _012_ = ap_CS_fsm[28] ? grp_fu_622_p2[35:4] : op_23_V_reg_1035;
assign _003_ = ap_CS_fsm[34] ? grp_fu_730_p2 : add_ln69_3_reg_1105;
assign _002_ = ap_CS_fsm[34] ? grp_fu_725_p2 : add_ln69_2_reg_1100;
assign _001_ = _048_ ? grp_fu_467_p2 : add_ln691_reg_957;
assign _000_ = ap_CS_fsm[25] ? grp_fu_563_p2 : add_ln691_1_reg_995;
assign _005_ = ap_rst ? 37'h0000000001 : ap_NS_fsm;
assign icmp_ln768_fu_459_p2 = _226_ ? 1'h1 : 1'h0;
assign icmp_ln851_1_fu_412_p2 = _227_ ? 1'h1 : 1'h0;
assign icmp_ln851_fu_350_p2 = _055_ ? 1'h1 : 1'h0;
assign icmp_ln890_fu_287_p2 = _225_ ? 1'h1 : 1'h0;
assign op_12_V_fu_506_p3 = or_ln384_fu_502_p2 ? select_ln384_fu_495_p3 : { p_Result_9_reg_912, 1'h0 };
assign r_fu_421_p3 = tmp_reg_788 ? trunc_ln1497_1_reg_892 : { trunc_ln1497_reg_887[3], trunc_ln1497_reg_887[3], trunc_ln1497_reg_887[3], trunc_ln1497_reg_887[3], trunc_ln1497_reg_887[3], trunc_ln1497_reg_887[3], trunc_ln1497_reg_887[3], trunc_ln1497_reg_887[3], trunc_ln1497_reg_887 };
assign ret_V_3_fu_242_p3 = ret_V_14_reg_750[4] ? select_ln850_fu_236_p3 : ret_V_reg_756;
assign select_ln353_1_fu_597_p3 = ret_V_19_reg_983[33] ? select_ln850_5_fu_591_p3 : ret_V_21_cast_reg_988;
assign select_ln353_fu_526_p3 = ret_V_18_reg_929[7] ? select_ln850_4_fu_521_p3 : sext_ln850_reg_944;
assign select_ln384_fu_495_p3 = overflow_reg_951 ? 2'h1 : 2'h3;
assign select_ln850_2_fu_367_p3 = icmp_ln851_reg_872 ? ret_V_7_reg_860 : ret_V_9_reg_877;
assign select_ln850_3_fu_372_p3 = ret_V_17_reg_855[16] ? select_ln850_2_fu_367_p3 : ret_V_7_reg_860;
assign select_ln850_4_fu_521_p3 = icmp_ln851_1_reg_907 ? add_ln691_reg_957 : sext_ln850_reg_944;
assign select_ln850_5_fu_591_p3 = op_12_V_reg_962[0] ? add_ln691_1_reg_995 : ret_V_21_cast_reg_988;
assign select_ln850_fu_236_p3 = ret_V_14_reg_750[0] ? ret_V_2_reg_763 : ret_V_reg_756;
assign signbit_fu_310_p2 = _228_ ? 1'h1 : 1'h0;
assign ret_V_14_fu_205_p2 = { op_0[3], op_0 } ^ { op_1, 1'h0 };
assign ap_CS_fsm_state1 = ap_CS_fsm[0];
assign ap_CS_fsm_state10 = ap_CS_fsm[9];
assign ap_CS_fsm_state11 = ap_CS_fsm[10];
assign ap_CS_fsm_state12 = ap_CS_fsm[11];
assign ap_CS_fsm_state13 = ap_CS_fsm[12];
assign ap_CS_fsm_state14 = ap_CS_fsm[13];
assign ap_CS_fsm_state15 = ap_CS_fsm[14];
assign ap_CS_fsm_state16 = ap_CS_fsm[15];
assign ap_CS_fsm_state17 = ap_CS_fsm[16];
assign ap_CS_fsm_state18 = ap_CS_fsm[17];
assign ap_CS_fsm_state19 = ap_CS_fsm[18];
assign ap_CS_fsm_state2 = ap_CS_fsm[1];
assign ap_CS_fsm_state20 = ap_CS_fsm[19];
assign ap_CS_fsm_state21 = ap_CS_fsm[20];
assign ap_CS_fsm_state22 = ap_CS_fsm[21];
assign ap_CS_fsm_state23 = ap_CS_fsm[22];
assign ap_CS_fsm_state24 = ap_CS_fsm[23];
assign ap_CS_fsm_state25 = ap_CS_fsm[24];
assign ap_CS_fsm_state26 = ap_CS_fsm[25];
assign ap_CS_fsm_state27 = ap_CS_fsm[26];
assign ap_CS_fsm_state28 = ap_CS_fsm[27];
assign ap_CS_fsm_state29 = ap_CS_fsm[28];
assign ap_CS_fsm_state3 = ap_CS_fsm[2];
assign ap_CS_fsm_state30 = ap_CS_fsm[29];
assign ap_CS_fsm_state31 = ap_CS_fsm[30];
assign ap_CS_fsm_state32 = ap_CS_fsm[31];
assign ap_CS_fsm_state33 = ap_CS_fsm[32];
assign ap_CS_fsm_state34 = ap_CS_fsm[33];
assign ap_CS_fsm_state35 = ap_CS_fsm[34];
assign ap_CS_fsm_state36 = ap_CS_fsm[35];
assign ap_CS_fsm_state37 = ap_CS_fsm[36];
assign ap_CS_fsm_state4 = ap_CS_fsm[3];
assign ap_CS_fsm_state5 = ap_CS_fsm[4];
assign ap_done = op_29_ap_vld;
assign ap_ready = op_29_ap_vld;
assign grp_fu_265_p1 = { op_6[3], op_6 };
assign grp_fu_279_p1 = { op_5[3], op_5 };
assign grp_fu_295_p1 = { op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6 };
assign grp_fu_304_p1 = { sub_ln1497_reg_799[4], sub_ln1497_reg_799[4], sub_ln1497_reg_799[4], sub_ln1497_reg_799[4], sub_ln1497_reg_799[4], sub_ln1497_reg_799[4], sub_ln1497_reg_799[4], sub_ln1497_reg_799[4], sub_ln1497_reg_799[4], sub_ln1497_reg_799[4], sub_ln1497_reg_799[4], sub_ln1497_reg_799[4], sub_ln1497_reg_799[4], sub_ln1497_reg_799[4], sub_ln1497_reg_799[4], sub_ln1497_reg_799[4], sub_ln1497_reg_799[4], sub_ln1497_reg_799[4], sub_ln1497_reg_799[4], sub_ln1497_reg_799[4], sub_ln1497_reg_799[4], sub_ln1497_reg_799[4], sub_ln1497_reg_799[4], sub_ln1497_reg_799[4], sub_ln1497_reg_799[4], sub_ln1497_reg_799[4], sub_ln1497_reg_799[4], sub_ln1497_reg_799 };
assign grp_fu_330_p0 = { 3'h0, signbit_reg_835, 13'h0000 };
assign grp_fu_330_p1 = { op_7[15], op_7 };
assign grp_fu_402_p0 = { select_ln850_3_reg_882[3], select_ln850_3_reg_882, 3'h0 };
assign grp_fu_402_p1 = { op_10[3], op_10[3], op_10[3], op_10[3], op_10 };
assign grp_fu_467_p0 = { tmp_2_reg_934[4], tmp_2_reg_934 };
assign grp_fu_547_p0 = { select_ln353_reg_968[5], select_ln353_reg_968[5], select_ln353_reg_968[5], select_ln353_reg_968[5], select_ln353_reg_968[5], select_ln353_reg_968[5], select_ln353_reg_968[5], select_ln353_reg_968[5], select_ln353_reg_968[5], select_ln353_reg_968[5], select_ln353_reg_968[5], select_ln353_reg_968[5], select_ln353_reg_968[5], select_ln353_reg_968[5], select_ln353_reg_968[5], select_ln353_reg_968[5], select_ln353_reg_968[5], select_ln353_reg_968[5], select_ln353_reg_968[5], select_ln353_reg_968[5], select_ln353_reg_968[5], select_ln353_reg_968[5], select_ln353_reg_968[5], select_ln353_reg_968[5], select_ln353_reg_968[5], select_ln353_reg_968[5], select_ln353_reg_968[5], select_ln353_reg_968, 1'h0 };
assign grp_fu_547_p1 = { op_12_V_reg_962[1], op_12_V_reg_962[1], op_12_V_reg_962[1], op_12_V_reg_962[1], op_12_V_reg_962[1], op_12_V_reg_962[1], op_12_V_reg_962[1], op_12_V_reg_962[1], op_12_V_reg_962[1], op_12_V_reg_962[1], op_12_V_reg_962[1], op_12_V_reg_962[1], op_12_V_reg_962[1], op_12_V_reg_962[1], op_12_V_reg_962[1], op_12_V_reg_962[1], op_12_V_reg_962[1], op_12_V_reg_962[1], op_12_V_reg_962[1], op_12_V_reg_962[1], op_12_V_reg_962[1], op_12_V_reg_962[1], op_12_V_reg_962[1], op_12_V_reg_962[1], op_12_V_reg_962[1], op_12_V_reg_962[1], op_12_V_reg_962[1], op_12_V_reg_962[1], op_12_V_reg_962[1], op_12_V_reg_962[1], op_12_V_reg_962[1], op_12_V_reg_962[1], op_12_V_reg_962 };
assign grp_fu_622_p0 = { select_ln353_1_reg_1010, 4'h0 };
assign grp_fu_622_p1 = { ret_V_6_reg_1005[3], ret_V_6_reg_1005[3], ret_V_6_reg_1005[3], ret_V_6_reg_1005[3], ret_V_6_reg_1005[3], ret_V_6_reg_1005[3], ret_V_6_reg_1005[3], ret_V_6_reg_1005[3], ret_V_6_reg_1005[3], ret_V_6_reg_1005[3], ret_V_6_reg_1005[3], ret_V_6_reg_1005[3], ret_V_6_reg_1005[3], ret_V_6_reg_1005[3], ret_V_6_reg_1005[3], ret_V_6_reg_1005[3], ret_V_6_reg_1005[3], ret_V_6_reg_1005[3], ret_V_6_reg_1005[3], ret_V_6_reg_1005[3], ret_V_6_reg_1005[3], ret_V_6_reg_1005[3], ret_V_6_reg_1005[3], ret_V_6_reg_1005[3], ret_V_6_reg_1005[3], ret_V_6_reg_1005[3], ret_V_6_reg_1005[3], ret_V_6_reg_1005[3], ret_V_6_reg_1005, 4'h0 };
assign grp_fu_642_p0 = { 1'h0, ret_V_15_reg_1000[3], ret_V_15_reg_1000[3], ret_V_15_reg_1000[3], ret_V_15_reg_1000[3], ret_V_15_reg_1000[3], ret_V_15_reg_1000[3], ret_V_15_reg_1000[3], ret_V_15_reg_1000[3], ret_V_15_reg_1000[3], ret_V_15_reg_1000[3], ret_V_15_reg_1000[3], ret_V_15_reg_1000[3], ret_V_15_reg_1000 };
assign grp_fu_642_p1 = { 9'h000, ret_V_16_reg_840[4], ret_V_16_reg_840[4], ret_V_16_reg_840[4], ret_V_16_reg_840 };
assign grp_fu_661_p0 = { 15'h0000, add_ln69_reg_1040 };
assign grp_fu_675_p1 = op_11[1:0];
assign grp_fu_698_p0 = { op_25_V_reg_1055, 4'h0 };
assign grp_fu_698_p1 = { 31'h00000000, tmp_V_reg_1050, 4'h0 };
assign grp_fu_725_p1 = { op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19 };
assign grp_fu_730_p0 = { 2'h0, op_18 };
assign grp_fu_730_p1 = { op_17_V_reg_1075[1], op_17_V_reg_1075[1], op_17_V_reg_1075 };
assign grp_fu_739_p0 = { add_ln69_3_reg_1105[3], add_ln69_3_reg_1105[3], add_ln69_3_reg_1105[3], add_ln69_3_reg_1105[3], add_ln69_3_reg_1105[3], add_ln69_3_reg_1105[3], add_ln69_3_reg_1105[3], add_ln69_3_reg_1105[3], add_ln69_3_reg_1105[3], add_ln69_3_reg_1105[3], add_ln69_3_reg_1105[3], add_ln69_3_reg_1105[3], add_ln69_3_reg_1105[3], add_ln69_3_reg_1105[3], add_ln69_3_reg_1105[3], add_ln69_3_reg_1105[3], add_ln69_3_reg_1105[3], add_ln69_3_reg_1105[3], add_ln69_3_reg_1105[3], add_ln69_3_reg_1105[3], add_ln69_3_reg_1105[3], add_ln69_3_reg_1105[3], add_ln69_3_reg_1105[3], add_ln69_3_reg_1105[3], add_ln69_3_reg_1105[3], add_ln69_3_reg_1105[3], add_ln69_3_reg_1105[3], add_ln69_3_reg_1105[3], add_ln69_3_reg_1105 };
assign icmp_ln890_fu_287_p0 = op_5;
assign op_13_V_fu_604_p3 = { ret_V_6_reg_1005, 4'h0 };
assign op_29 = grp_fu_739_p2;
assign p_Result_5_fu_360_p3 = ret_V_17_reg_855[16];
assign p_Result_6_fu_514_p3 = ret_V_18_reg_929[7];
assign p_Result_7_fu_581_p3 = ret_V_19_reg_983[33];
assign p_Result_9_fu_427_p1 = r_fu_421_p3[0];
assign p_Result_s_fu_226_p3 = ret_V_14_reg_750[4];
assign p_Val2_4_fu_488_p3 = { p_Result_9_reg_912, 1'h0 };
assign p_Val2_s_fu_680_p3 = { tmp_V_reg_1050, 4'h0 };
assign ret_V_15_fu_572_p1 = op_6;
assign ret_V_6_fu_577_p1 = op_6;
assign rhs_1_fu_319_p3 = { signbit_reg_835, 13'h0000 };
assign rhs_2_fu_391_p3 = { select_ln850_3_reg_882, 3'h0 };
assign rhs_fu_197_p1 = op_1;
assign rhs_fu_197_p3 = { op_1, 1'h0 };
assign sext_ln1192_fu_387_p0 = op_10;
assign sext_ln1497_fu_418_p1 = { trunc_ln1497_reg_887[3], trunc_ln1497_reg_887[3], trunc_ln1497_reg_887[3], trunc_ln1497_reg_887[3], trunc_ln1497_reg_887[3], trunc_ln1497_reg_887[3], trunc_ln1497_reg_887[3], trunc_ln1497_reg_887[3], trunc_ln1497_reg_887 };
assign sext_ln545_fu_292_p0 = op_6;
assign sext_ln69_2_fu_635_p1 = { ret_V_16_reg_840[4], ret_V_16_reg_840[4], ret_V_16_reg_840[4], ret_V_16_reg_840 };
assign sext_ln69_fu_628_p1 = { ret_V_15_reg_1000[3], ret_V_15_reg_1000[3], ret_V_15_reg_1000[3], ret_V_15_reg_1000[3], ret_V_15_reg_1000[3], ret_V_15_reg_1000[3], ret_V_15_reg_1000[3], ret_V_15_reg_1000[3], ret_V_15_reg_1000[3], ret_V_15_reg_1000[3], ret_V_15_reg_1000[3], ret_V_15_reg_1000[3], ret_V_15_reg_1000 };
assign sext_ln703_1_fu_568_p1 = { op_4[1], op_4[1], op_4 };
assign sext_ln703_2_fu_275_p0 = op_5;
assign sext_ln703_3_fu_253_p0 = op_6;
assign sext_ln703_3_fu_253_p1 = { op_6[3], op_6 };
assign sext_ln703_fu_193_p1 = { op_0[3], op_0 };
assign sext_ln850_fu_464_p1 = { tmp_2_reg_934[4], tmp_2_reg_934 };
assign sext_ln890_fu_284_p1 = { ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768 };
assign signbit_fu_310_p1 = op_5;
assign tmp_6_fu_536_p3 = { select_ln353_reg_968, 1'h0 };
assign tmp_fu_257_p1 = op_6;
assign trunc_ln1347_fu_271_p1 = grp_fu_249_p2[1:0];
assign trunc_ln1497_1_fu_383_p1 = grp_fu_304_p2[11:0];
assign trunc_ln1497_fu_379_p1 = grp_fu_295_p2[3:0];
assign trunc_ln851_1_fu_346_p1 = grp_fu_330_p2[12:0];
assign trunc_ln851_2_fu_408_p0 = op_10;
assign trunc_ln851_2_fu_408_p1 = op_10[2:0];
assign trunc_ln851_3_fu_588_p1 = op_12_V_reg_962[0];
assign trunc_ln851_fu_233_p1 = ret_V_14_reg_750[0];
assign \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.ain_s0  = \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.a ;
assign \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.s  = { \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.fas_s2 , \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.sum_s1  };
assign \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.u2.a  = \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.ain_s1 ;
assign \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.u2.b  = \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.bin_s1 ;
assign \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.u2.cin  = \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.carry_s1 ;
assign \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.facout_s2  = \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.u2.cout ;
assign \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.fas_s2  = \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.u2.s ;
assign \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.u1.a  = \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.a [1:0];
assign \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.u1.b  = \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.bin_s0 [1:0];
assign \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.u1.cin  = 1'h1;
assign \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.facout_s1  = \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.u1.cout ;
assign \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.fas_s1  = \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.u1.s ;
assign \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.a  = \sub_5ns_5s_5_2_1_U3.din0 ;
assign \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.b  = \sub_5ns_5s_5_2_1_U3.din1 ;
assign \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.ce  = \sub_5ns_5s_5_2_1_U3.ce ;
assign \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.clk  = \sub_5ns_5s_5_2_1_U3.clk ;
assign \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.reset  = \sub_5ns_5s_5_2_1_U3.reset ;
assign \sub_5ns_5s_5_2_1_U3.dout  = \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.s ;
assign \sub_5ns_5s_5_2_1_U3.ce  = 1'h1;
assign \sub_5ns_5s_5_2_1_U3.clk  = ap_clk;
assign \sub_5ns_5s_5_2_1_U3.din0  = 5'h00;
assign \sub_5ns_5s_5_2_1_U3.din1  = { op_6[3], op_6 };
assign grp_fu_265_p2 = \sub_5ns_5s_5_2_1_U3.dout ;
assign \sub_5ns_5s_5_2_1_U3.reset  = ap_rst;
assign \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.ain_s0  = \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.a ;
assign \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.s  = { \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.fas_s2 , \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.sum_s1  };
assign \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.u2.a  = \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.ain_s1 ;
assign \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.u2.b  = \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.bin_s1 ;
assign \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.u2.cin  = \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.carry_s1 ;
assign \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.facout_s2  = \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.u2.cout ;
assign \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.fas_s2  = \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.u2.s ;
assign \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.u1.a  = \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.a [0];
assign \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.u1.b  = \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.bin_s0 [0];
assign \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.u1.cin  = 1'h1;
assign \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.facout_s1  = \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.u1.cout ;
assign \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.fas_s1  = \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.u1.s ;
assign \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.a  = \sub_2ns_2ns_2_2_1_U16.din0 ;
assign \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.b  = \sub_2ns_2ns_2_2_1_U16.din1 ;
assign \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.ce  = \sub_2ns_2ns_2_2_1_U16.ce ;
assign \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.clk  = \sub_2ns_2ns_2_2_1_U16.clk ;
assign \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.reset  = \sub_2ns_2ns_2_2_1_U16.reset ;
assign \sub_2ns_2ns_2_2_1_U16.dout  = \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.s ;
assign \sub_2ns_2ns_2_2_1_U16.ce  = 1'h1;
assign \sub_2ns_2ns_2_2_1_U16.clk  = ap_clk;
assign \sub_2ns_2ns_2_2_1_U16.din0  = trunc_ln1347_reg_804;
assign \sub_2ns_2ns_2_2_1_U16.din1  = op_11[1:0];
assign grp_fu_675_p2 = \sub_2ns_2ns_2_2_1_U16.dout ;
assign \sub_2ns_2ns_2_2_1_U16.reset  = ap_rst;
assign \shl_32s_32s_32_7_1_U6.din1_cast  = \shl_32s_32s_32_7_1_U6.din1 ;
assign \shl_32s_32s_32_7_1_U6.din1_mask  = 32'd31;
assign \shl_32s_32s_32_7_1_U6.ce  = 1'h1;
assign \shl_32s_32s_32_7_1_U6.clk  = ap_clk;
assign \shl_32s_32s_32_7_1_U6.din0  = { ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768 };
assign \shl_32s_32s_32_7_1_U6.din1  = { sub_ln1497_reg_799[4], sub_ln1497_reg_799[4], sub_ln1497_reg_799[4], sub_ln1497_reg_799[4], sub_ln1497_reg_799[4], sub_ln1497_reg_799[4], sub_ln1497_reg_799[4], sub_ln1497_reg_799[4], sub_ln1497_reg_799[4], sub_ln1497_reg_799[4], sub_ln1497_reg_799[4], sub_ln1497_reg_799[4], sub_ln1497_reg_799[4], sub_ln1497_reg_799[4], sub_ln1497_reg_799[4], sub_ln1497_reg_799[4], sub_ln1497_reg_799[4], sub_ln1497_reg_799[4], sub_ln1497_reg_799[4], sub_ln1497_reg_799[4], sub_ln1497_reg_799[4], sub_ln1497_reg_799[4], sub_ln1497_reg_799[4], sub_ln1497_reg_799[4], sub_ln1497_reg_799[4], sub_ln1497_reg_799[4], sub_ln1497_reg_799[4], sub_ln1497_reg_799 };
assign grp_fu_304_p2 = \shl_32s_32s_32_7_1_U6.dout ;
assign \shl_32s_32s_32_7_1_U6.reset  = ap_rst;
assign \mul_4s_4s_4_7_1_U2.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.p  = \mul_4s_4s_4_7_1_U2.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.buff4 ;
assign \mul_4s_4s_4_7_1_U2.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.a  = \mul_4s_4s_4_7_1_U2.din0 ;
assign \mul_4s_4s_4_7_1_U2.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.b  = \mul_4s_4s_4_7_1_U2.din1 ;
assign \mul_4s_4s_4_7_1_U2.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.ce  = \mul_4s_4s_4_7_1_U2.ce ;
assign \mul_4s_4s_4_7_1_U2.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.clk  = \mul_4s_4s_4_7_1_U2.clk ;
assign \mul_4s_4s_4_7_1_U2.dout  = \mul_4s_4s_4_7_1_U2.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.p ;
assign \mul_4s_4s_4_7_1_U2.ce  = 1'h1;
assign \mul_4s_4s_4_7_1_U2.clk  = ap_clk;
assign \mul_4s_4s_4_7_1_U2.din0  = ret_V_3_reg_768;
assign \mul_4s_4s_4_7_1_U2.din1  = op_1;
assign grp_fu_249_p2 = \mul_4s_4s_4_7_1_U2.dout ;
assign \mul_4s_4s_4_7_1_U2.reset  = ap_rst;
assign \ashr_32s_32s_32_7_1_U5.din1_cast  = \ashr_32s_32s_32_7_1_U5.din1 ;
assign \ashr_32s_32s_32_7_1_U5.din1_mask  = 32'd31;
assign \ashr_32s_32s_32_7_1_U5.ce  = 1'h1;
assign \ashr_32s_32s_32_7_1_U5.clk  = ap_clk;
assign \ashr_32s_32s_32_7_1_U5.din0  = { ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768 };
assign \ashr_32s_32s_32_7_1_U5.din1  = { op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6 };
assign grp_fu_295_p2 = \ashr_32s_32s_32_7_1_U5.dout ;
assign \ashr_32s_32s_32_7_1_U5.reset  = ap_rst;
assign \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.ain_s0  = \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.a ;
assign \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.bin_s0  = \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.b ;
assign \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.s  = { \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.fas_s2 , \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.sum_s1  };
assign \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.u2.a  = \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.ain_s1 ;
assign \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.u2.b  = \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.bin_s1 ;
assign \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.u2.cin  = \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.carry_s1 ;
assign \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.facout_s2  = \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.u2.cout ;
assign \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.fas_s2  = \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.u2.s ;
assign \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.u1.a  = \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.a [3:0];
assign \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.u1.b  = \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.b [3:0];
assign \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.u1.cin  = 1'h0;
assign \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.facout_s1  = \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.u1.cout ;
assign \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.fas_s1  = \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.u1.s ;
assign \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.a  = \add_8s_8s_8_2_1_U9.din0 ;
assign \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.b  = \add_8s_8s_8_2_1_U9.din1 ;
assign \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.ce  = \add_8s_8s_8_2_1_U9.ce ;
assign \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.clk  = \add_8s_8s_8_2_1_U9.clk ;
assign \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.reset  = \add_8s_8s_8_2_1_U9.reset ;
assign \add_8s_8s_8_2_1_U9.dout  = \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.s ;
assign \add_8s_8s_8_2_1_U9.ce  = 1'h1;
assign \add_8s_8s_8_2_1_U9.clk  = ap_clk;
assign \add_8s_8s_8_2_1_U9.din0  = { select_ln850_3_reg_882[3], select_ln850_3_reg_882, 3'h0 };
assign \add_8s_8s_8_2_1_U9.din1  = { op_10[3], op_10[3], op_10[3], op_10[3], op_10 };
assign grp_fu_402_p2 = \add_8s_8s_8_2_1_U9.dout ;
assign \add_8s_8s_8_2_1_U9.reset  = ap_rst;
assign \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.ain_s0  = \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.a ;
assign \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.bin_s0  = \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.b ;
assign \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.s  = { \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.fas_s2 , \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.sum_s1  };
assign \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.u2.a  = \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.ain_s1 ;
assign \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.u2.b  = \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.bin_s1 ;
assign \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.u2.cin  = \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.carry_s1 ;
assign \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.facout_s2  = \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.u2.cout ;
assign \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.fas_s2  = \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.u2.s ;
assign \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.u1.a  = \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.a [2:0];
assign \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.u1.b  = \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.b [2:0];
assign \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.u1.cin  = 1'h0;
assign \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.facout_s1  = \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.u1.cout ;
assign \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.fas_s1  = \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.u1.s ;
assign \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.a  = \add_6s_6ns_6_2_1_U10.din0 ;
assign \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.b  = \add_6s_6ns_6_2_1_U10.din1 ;
assign \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.ce  = \add_6s_6ns_6_2_1_U10.ce ;
assign \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.clk  = \add_6s_6ns_6_2_1_U10.clk ;
assign \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.reset  = \add_6s_6ns_6_2_1_U10.reset ;
assign \add_6s_6ns_6_2_1_U10.dout  = \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.s ;
assign \add_6s_6ns_6_2_1_U10.ce  = 1'h1;
assign \add_6s_6ns_6_2_1_U10.clk  = ap_clk;
assign \add_6s_6ns_6_2_1_U10.din0  = { tmp_2_reg_934[4], tmp_2_reg_934 };
assign \add_6s_6ns_6_2_1_U10.din1  = 6'h01;
assign grp_fu_467_p2 = \add_6s_6ns_6_2_1_U10.dout ;
assign \add_6s_6ns_6_2_1_U10.reset  = ap_rst;
assign \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.ain_s0  = \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.a ;
assign \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.bin_s0  = \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.b ;
assign \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.s  = { \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.fas_s2 , \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.sum_s1  };
assign \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.u2.a  = \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.ain_s1 ;
assign \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.u2.b  = \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.bin_s1 ;
assign \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.u2.cin  = \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.carry_s1 ;
assign \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.facout_s2  = \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.u2.cout ;
assign \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.fas_s2  = \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.u2.s ;
assign \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.u1.a  = \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.a [1:0];
assign \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.u1.b  = \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.b [1:0];
assign \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.u1.cin  = 1'h0;
assign \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.facout_s1  = \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.u1.cout ;
assign \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.fas_s1  = \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.u1.s ;
assign \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.a  = \add_5s_5s_5_2_1_U4.din0 ;
assign \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.b  = \add_5s_5s_5_2_1_U4.din1 ;
assign \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.ce  = \add_5s_5s_5_2_1_U4.ce ;
assign \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.clk  = \add_5s_5s_5_2_1_U4.clk ;
assign \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.reset  = \add_5s_5s_5_2_1_U4.reset ;
assign \add_5s_5s_5_2_1_U4.dout  = \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.s ;
assign \add_5s_5s_5_2_1_U4.ce  = 1'h1;
assign \add_5s_5s_5_2_1_U4.clk  = ap_clk;
assign \add_5s_5s_5_2_1_U4.din0  = sext_ln703_3_reg_782;
assign \add_5s_5s_5_2_1_U4.din1  = { op_5[3], op_5 };
assign grp_fu_279_p2 = \add_5s_5s_5_2_1_U4.dout ;
assign \add_5s_5s_5_2_1_U4.reset  = ap_rst;
assign \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.ain_s0  = \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.a ;
assign \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.bin_s0  = \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.b ;
assign \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.s  = { \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.fas_s2 , \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.sum_s1  };
assign \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.u2.a  = \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.ain_s1 ;
assign \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.u2.b  = \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.bin_s1 ;
assign \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.u2.cin  = \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.carry_s1 ;
assign \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.facout_s2  = \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.u2.cout ;
assign \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.fas_s2  = \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.u2.s ;
assign \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.u1.a  = \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.a [1:0];
assign \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.u1.b  = \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.b [1:0];
assign \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.u1.cin  = 1'h0;
assign \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.facout_s1  = \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.u1.cout ;
assign \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.fas_s1  = \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.u1.s ;
assign \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.a  = \add_4ns_4s_4_2_1_U19.din0 ;
assign \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.b  = \add_4ns_4s_4_2_1_U19.din1 ;
assign \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.ce  = \add_4ns_4s_4_2_1_U19.ce ;
assign \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.clk  = \add_4ns_4s_4_2_1_U19.clk ;
assign \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.reset  = \add_4ns_4s_4_2_1_U19.reset ;
assign \add_4ns_4s_4_2_1_U19.dout  = \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.s ;
assign \add_4ns_4s_4_2_1_U19.ce  = 1'h1;
assign \add_4ns_4s_4_2_1_U19.clk  = ap_clk;
assign \add_4ns_4s_4_2_1_U19.din0  = { 2'h0, op_18 };
assign \add_4ns_4s_4_2_1_U19.din1  = { op_17_V_reg_1075[1], op_17_V_reg_1075[1], op_17_V_reg_1075 };
assign grp_fu_730_p2 = \add_4ns_4s_4_2_1_U19.dout ;
assign \add_4ns_4s_4_2_1_U19.reset  = ap_rst;
assign \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.ain_s0  = \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.a ;
assign \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.bin_s0  = \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.b ;
assign \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.s  = { \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.fas_s2 , \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.sum_s1  };
assign \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.u2.a  = \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.ain_s1 ;
assign \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.u2.b  = \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.bin_s1 ;
assign \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.u2.cin  = \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.carry_s1 ;
assign \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.facout_s2  = \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.u2.cout ;
assign \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.fas_s2  = \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.u2.s ;
assign \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.u1.a  = \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.a [1:0];
assign \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.u1.b  = \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.b [1:0];
assign \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.u1.cin  = 1'h0;
assign \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.facout_s1  = \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.u1.cout ;
assign \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.fas_s1  = \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.u1.s ;
assign \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.a  = \add_4ns_4ns_4_2_1_U8.din0 ;
assign \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.b  = \add_4ns_4ns_4_2_1_U8.din1 ;
assign \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.ce  = \add_4ns_4ns_4_2_1_U8.ce ;
assign \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.clk  = \add_4ns_4ns_4_2_1_U8.clk ;
assign \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.reset  = \add_4ns_4ns_4_2_1_U8.reset ;
assign \add_4ns_4ns_4_2_1_U8.dout  = \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.s ;
assign \add_4ns_4ns_4_2_1_U8.ce  = 1'h1;
assign \add_4ns_4ns_4_2_1_U8.clk  = ap_clk;
assign \add_4ns_4ns_4_2_1_U8.din0  = ret_V_7_reg_860;
assign \add_4ns_4ns_4_2_1_U8.din1  = 4'h1;
assign grp_fu_355_p2 = \add_4ns_4ns_4_2_1_U8.dout ;
assign \add_4ns_4ns_4_2_1_U8.reset  = ap_rst;
assign \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.ain_s0  = \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.a ;
assign \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.bin_s0  = \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.b ;
assign \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.s  = { \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.fas_s2 , \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.sum_s1  };
assign \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.u2.a  = \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.ain_s1 ;
assign \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.u2.b  = \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.bin_s1 ;
assign \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.u2.cin  = \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.carry_s1 ;
assign \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.facout_s2  = \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.u2.cout ;
assign \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.fas_s2  = \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.u2.s ;
assign \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.u1.a  = \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.a [1:0];
assign \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.u1.b  = \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.b [1:0];
assign \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.u1.cin  = 1'h0;
assign \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.facout_s1  = \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.u1.cout ;
assign \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.fas_s1  = \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.u1.s ;
assign \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.a  = \add_4ns_4ns_4_2_1_U1.din0 ;
assign \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.b  = \add_4ns_4ns_4_2_1_U1.din1 ;
assign \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.ce  = \add_4ns_4ns_4_2_1_U1.ce ;
assign \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.clk  = \add_4ns_4ns_4_2_1_U1.clk ;
assign \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.reset  = \add_4ns_4ns_4_2_1_U1.reset ;
assign \add_4ns_4ns_4_2_1_U1.dout  = \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.s ;
assign \add_4ns_4ns_4_2_1_U1.ce  = 1'h1;
assign \add_4ns_4ns_4_2_1_U1.clk  = ap_clk;
assign \add_4ns_4ns_4_2_1_U1.din0  = ret_V_reg_756;
assign \add_4ns_4ns_4_2_1_U1.din1  = 4'h1;
assign grp_fu_221_p2 = \add_4ns_4ns_4_2_1_U1.dout ;
assign \add_4ns_4ns_4_2_1_U1.reset  = ap_rst;
assign \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.ain_s0  = \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.a ;
assign \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.bin_s0  = \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.b ;
assign \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.s  = { \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.fas_s2 , \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.sum_s1  };
assign \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.u2.a  = \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.ain_s1 ;
assign \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.u2.b  = \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.bin_s1 ;
assign \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.u2.cin  = \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.carry_s1 ;
assign \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.facout_s2  = \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.u2.cout ;
assign \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.fas_s2  = \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.u2.s ;
assign \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.u1.a  = \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.a [17:0];
assign \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.u1.b  = \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.b [17:0];
assign \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.u1.cin  = 1'h0;
assign \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.facout_s1  = \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.u1.cout ;
assign \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.fas_s1  = \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.u1.s ;
assign \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.a  = \add_36ns_36s_36_2_1_U13.din0 ;
assign \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.b  = \add_36ns_36s_36_2_1_U13.din1 ;
assign \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.ce  = \add_36ns_36s_36_2_1_U13.ce ;
assign \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.clk  = \add_36ns_36s_36_2_1_U13.clk ;
assign \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.reset  = \add_36ns_36s_36_2_1_U13.reset ;
assign \add_36ns_36s_36_2_1_U13.dout  = \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.s ;
assign \add_36ns_36s_36_2_1_U13.ce  = 1'h1;
assign \add_36ns_36s_36_2_1_U13.clk  = ap_clk;
assign \add_36ns_36s_36_2_1_U13.din0  = { select_ln353_1_reg_1010, 4'h0 };
assign \add_36ns_36s_36_2_1_U13.din1  = { ret_V_6_reg_1005[3], ret_V_6_reg_1005[3], ret_V_6_reg_1005[3], ret_V_6_reg_1005[3], ret_V_6_reg_1005[3], ret_V_6_reg_1005[3], ret_V_6_reg_1005[3], ret_V_6_reg_1005[3], ret_V_6_reg_1005[3], ret_V_6_reg_1005[3], ret_V_6_reg_1005[3], ret_V_6_reg_1005[3], ret_V_6_reg_1005[3], ret_V_6_reg_1005[3], ret_V_6_reg_1005[3], ret_V_6_reg_1005[3], ret_V_6_reg_1005[3], ret_V_6_reg_1005[3], ret_V_6_reg_1005[3], ret_V_6_reg_1005[3], ret_V_6_reg_1005[3], ret_V_6_reg_1005[3], ret_V_6_reg_1005[3], ret_V_6_reg_1005[3], ret_V_6_reg_1005[3], ret_V_6_reg_1005[3], ret_V_6_reg_1005[3], ret_V_6_reg_1005[3], ret_V_6_reg_1005, 4'h0 };
assign grp_fu_622_p2 = \add_36ns_36s_36_2_1_U13.dout ;
assign \add_36ns_36s_36_2_1_U13.reset  = ap_rst;
assign \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.ain_s0  = \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.a ;
assign \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.bin_s0  = \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.b ;
assign \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.s  = { \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.fas_s2 , \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.sum_s1  };
assign \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.u2.a  = \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.ain_s1 ;
assign \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.u2.b  = \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.bin_s1 ;
assign \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.u2.cin  = \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.carry_s1 ;
assign \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.facout_s2  = \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.u2.cout ;
assign \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.fas_s2  = \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.u2.s ;
assign \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.u1.a  = \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.a [17:0];
assign \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.u1.b  = \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.b [17:0];
assign \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.u1.cin  = 1'h0;
assign \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.facout_s1  = \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.u1.cout ;
assign \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.fas_s1  = \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.u1.s ;
assign \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.a  = \add_36ns_36ns_36_2_1_U17.din0 ;
assign \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.b  = \add_36ns_36ns_36_2_1_U17.din1 ;
assign \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.ce  = \add_36ns_36ns_36_2_1_U17.ce ;
assign \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.clk  = \add_36ns_36ns_36_2_1_U17.clk ;
assign \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.reset  = \add_36ns_36ns_36_2_1_U17.reset ;
assign \add_36ns_36ns_36_2_1_U17.dout  = \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.s ;
assign \add_36ns_36ns_36_2_1_U17.ce  = 1'h1;
assign \add_36ns_36ns_36_2_1_U17.clk  = ap_clk;
assign \add_36ns_36ns_36_2_1_U17.din0  = { op_25_V_reg_1055, 4'h0 };
assign \add_36ns_36ns_36_2_1_U17.din1  = { 31'h00000000, tmp_V_reg_1050, 4'h0 };
assign grp_fu_698_p2 = \add_36ns_36ns_36_2_1_U17.dout ;
assign \add_36ns_36ns_36_2_1_U17.reset  = ap_rst;
assign \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.ain_s0  = \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.a ;
assign \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.bin_s0  = \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.b ;
assign \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.s  = { \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.fas_s2 , \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.sum_s1  };
assign \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.u2.a  = \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.ain_s1 ;
assign \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.u2.b  = \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.bin_s1 ;
assign \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.u2.cin  = \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.carry_s1 ;
assign \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.facout_s2  = \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.u2.cout ;
assign \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.fas_s2  = \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.u2.s ;
assign \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.u1.a  = \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.a [16:0];
assign \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.u1.b  = \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.b [16:0];
assign \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.u1.cin  = 1'h0;
assign \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.facout_s1  = \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.u1.cout ;
assign \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.fas_s1  = \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.u1.s ;
assign \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.a  = \add_34s_34s_34_2_1_U11.din0 ;
assign \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.b  = \add_34s_34s_34_2_1_U11.din1 ;
assign \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.ce  = \add_34s_34s_34_2_1_U11.ce ;
assign \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.clk  = \add_34s_34s_34_2_1_U11.clk ;
assign \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.reset  = \add_34s_34s_34_2_1_U11.reset ;
assign \add_34s_34s_34_2_1_U11.dout  = \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.s ;
assign \add_34s_34s_34_2_1_U11.ce  = 1'h1;
assign \add_34s_34s_34_2_1_U11.clk  = ap_clk;
assign \add_34s_34s_34_2_1_U11.din0  = { select_ln353_reg_968[5], select_ln353_reg_968[5], select_ln353_reg_968[5], select_ln353_reg_968[5], select_ln353_reg_968[5], select_ln353_reg_968[5], select_ln353_reg_968[5], select_ln353_reg_968[5], select_ln353_reg_968[5], select_ln353_reg_968[5], select_ln353_reg_968[5], select_ln353_reg_968[5], select_ln353_reg_968[5], select_ln353_reg_968[5], select_ln353_reg_968[5], select_ln353_reg_968[5], select_ln353_reg_968[5], select_ln353_reg_968[5], select_ln353_reg_968[5], select_ln353_reg_968[5], select_ln353_reg_968[5], select_ln353_reg_968[5], select_ln353_reg_968[5], select_ln353_reg_968[5], select_ln353_reg_968[5], select_ln353_reg_968[5], select_ln353_reg_968[5], select_ln353_reg_968, 1'h0 };
assign \add_34s_34s_34_2_1_U11.din1  = { op_12_V_reg_962[1], op_12_V_reg_962[1], op_12_V_reg_962[1], op_12_V_reg_962[1], op_12_V_reg_962[1], op_12_V_reg_962[1], op_12_V_reg_962[1], op_12_V_reg_962[1], op_12_V_reg_962[1], op_12_V_reg_962[1], op_12_V_reg_962[1], op_12_V_reg_962[1], op_12_V_reg_962[1], op_12_V_reg_962[1], op_12_V_reg_962[1], op_12_V_reg_962[1], op_12_V_reg_962[1], op_12_V_reg_962[1], op_12_V_reg_962[1], op_12_V_reg_962[1], op_12_V_reg_962[1], op_12_V_reg_962[1], op_12_V_reg_962[1], op_12_V_reg_962[1], op_12_V_reg_962[1], op_12_V_reg_962[1], op_12_V_reg_962[1], op_12_V_reg_962[1], op_12_V_reg_962[1], op_12_V_reg_962[1], op_12_V_reg_962[1], op_12_V_reg_962[1], op_12_V_reg_962 };
assign grp_fu_547_p2 = \add_34s_34s_34_2_1_U11.dout ;
assign \add_34s_34s_34_2_1_U11.reset  = ap_rst;
assign \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.ain_s0  = \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.a ;
assign \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.bin_s0  = \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.b ;
assign \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.s  = { \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.fas_s2 , \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.sum_s1  };
assign \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.u2.a  = \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.ain_s1 ;
assign \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.u2.b  = \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.bin_s1 ;
assign \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.u2.cin  = \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.carry_s1 ;
assign \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.facout_s2  = \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.u2.cout ;
assign \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.fas_s2  = \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.u2.s ;
assign \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.u1.a  = \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.a [15:0];
assign \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.u1.b  = \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.b [15:0];
assign \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.u1.cin  = 1'h0;
assign \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.facout_s1  = \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.u1.cout ;
assign \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.fas_s1  = \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.u1.s ;
assign \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.a  = \add_32s_32ns_32_2_1_U20.din0 ;
assign \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.b  = \add_32s_32ns_32_2_1_U20.din1 ;
assign \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.ce  = \add_32s_32ns_32_2_1_U20.ce ;
assign \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.clk  = \add_32s_32ns_32_2_1_U20.clk ;
assign \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.reset  = \add_32s_32ns_32_2_1_U20.reset ;
assign \add_32s_32ns_32_2_1_U20.dout  = \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.s ;
assign \add_32s_32ns_32_2_1_U20.ce  = 1'h1;
assign \add_32s_32ns_32_2_1_U20.clk  = ap_clk;
assign \add_32s_32ns_32_2_1_U20.din0  = { add_ln69_3_reg_1105[3], add_ln69_3_reg_1105[3], add_ln69_3_reg_1105[3], add_ln69_3_reg_1105[3], add_ln69_3_reg_1105[3], add_ln69_3_reg_1105[3], add_ln69_3_reg_1105[3], add_ln69_3_reg_1105[3], add_ln69_3_reg_1105[3], add_ln69_3_reg_1105[3], add_ln69_3_reg_1105[3], add_ln69_3_reg_1105[3], add_ln69_3_reg_1105[3], add_ln69_3_reg_1105[3], add_ln69_3_reg_1105[3], add_ln69_3_reg_1105[3], add_ln69_3_reg_1105[3], add_ln69_3_reg_1105[3], add_ln69_3_reg_1105[3], add_ln69_3_reg_1105[3], add_ln69_3_reg_1105[3], add_ln69_3_reg_1105[3], add_ln69_3_reg_1105[3], add_ln69_3_reg_1105[3], add_ln69_3_reg_1105[3], add_ln69_3_reg_1105[3], add_ln69_3_reg_1105[3], add_ln69_3_reg_1105[3], add_ln69_3_reg_1105 };
assign \add_32s_32ns_32_2_1_U20.din1  = add_ln69_2_reg_1100;
assign grp_fu_739_p2 = \add_32s_32ns_32_2_1_U20.dout ;
assign \add_32s_32ns_32_2_1_U20.reset  = ap_rst;
assign \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.ain_s0  = \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.a ;
assign \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.bin_s0  = \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.b ;
assign \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.s  = { \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.fas_s2 , \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.sum_s1  };
assign \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.u2.a  = \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.ain_s1 ;
assign \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.u2.b  = \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.bin_s1 ;
assign \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.u2.cin  = \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.carry_s1 ;
assign \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.facout_s2  = \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.u2.cout ;
assign \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.fas_s2  = \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.u2.s ;
assign \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.u1.a  = \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.a [15:0];
assign \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.u1.b  = \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.b [15:0];
assign \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.u1.cin  = 1'h0;
assign \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.facout_s1  = \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.u1.cout ;
assign \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.fas_s1  = \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.u1.s ;
assign \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.a  = \add_32ns_32s_32_2_1_U18.din0 ;
assign \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.b  = \add_32ns_32s_32_2_1_U18.din1 ;
assign \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.ce  = \add_32ns_32s_32_2_1_U18.ce ;
assign \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.clk  = \add_32ns_32s_32_2_1_U18.clk ;
assign \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.reset  = \add_32ns_32s_32_2_1_U18.reset ;
assign \add_32ns_32s_32_2_1_U18.dout  = \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.s ;
assign \add_32ns_32s_32_2_1_U18.ce  = 1'h1;
assign \add_32ns_32s_32_2_1_U18.clk  = ap_clk;
assign \add_32ns_32s_32_2_1_U18.din0  = op_26_V_reg_1080;
assign \add_32ns_32s_32_2_1_U18.din1  = { op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19 };
assign grp_fu_725_p2 = \add_32ns_32s_32_2_1_U18.dout ;
assign \add_32ns_32s_32_2_1_U18.reset  = ap_rst;
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s0  = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.a ;
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s0  = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.b ;
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.s  = { \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s2 , \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.sum_s1  };
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.a  = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s1 ;
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.b  = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s1 ;
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cin  = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.carry_s1 ;
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.facout_s2  = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cout ;
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s2  = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.s ;
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.a  = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.a [15:0];
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.b  = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.b [15:0];
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cin  = 1'h0;
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.facout_s1  = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cout ;
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s1  = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.s ;
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.a  = \add_32ns_32ns_32_2_1_U15.din0 ;
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.b  = \add_32ns_32ns_32_2_1_U15.din1 ;
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.ce  = \add_32ns_32ns_32_2_1_U15.ce ;
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.clk  = \add_32ns_32ns_32_2_1_U15.clk ;
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.reset  = \add_32ns_32ns_32_2_1_U15.reset ;
assign \add_32ns_32ns_32_2_1_U15.dout  = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.s ;
assign \add_32ns_32ns_32_2_1_U15.ce  = 1'h1;
assign \add_32ns_32ns_32_2_1_U15.clk  = ap_clk;
assign \add_32ns_32ns_32_2_1_U15.din0  = { 15'h0000, add_ln69_reg_1040 };
assign \add_32ns_32ns_32_2_1_U15.din1  = op_23_V_reg_1035;
assign grp_fu_661_p2 = \add_32ns_32ns_32_2_1_U15.dout ;
assign \add_32ns_32ns_32_2_1_U15.reset  = ap_rst;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s0  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.a ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s0  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.b ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.s  = { \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s2 , \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.sum_s1  };
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.a  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s1 ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.b  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s1 ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cin  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.carry_s1 ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.facout_s2  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cout ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s2  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.s ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.a  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.a [15:0];
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.b  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.b [15:0];
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cin  = 1'h0;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.facout_s1  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cout ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s1  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.s ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.a  = \add_32ns_32ns_32_2_1_U12.din0 ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.b  = \add_32ns_32ns_32_2_1_U12.din1 ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.ce  = \add_32ns_32ns_32_2_1_U12.ce ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.clk  = \add_32ns_32ns_32_2_1_U12.clk ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.reset  = \add_32ns_32ns_32_2_1_U12.reset ;
assign \add_32ns_32ns_32_2_1_U12.dout  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.s ;
assign \add_32ns_32ns_32_2_1_U12.ce  = 1'h1;
assign \add_32ns_32ns_32_2_1_U12.clk  = ap_clk;
assign \add_32ns_32ns_32_2_1_U12.din0  = ret_V_21_cast_reg_988;
assign \add_32ns_32ns_32_2_1_U12.din1  = 32'd1;
assign grp_fu_563_p2 = \add_32ns_32ns_32_2_1_U12.dout ;
assign \add_32ns_32ns_32_2_1_U12.reset  = ap_rst;
assign \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.ain_s0  = \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.a ;
assign \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.bin_s0  = \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.b ;
assign \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.s  = { \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.fas_s2 , \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.sum_s1  };
assign \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.u2.a  = \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.ain_s1 ;
assign \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.u2.b  = \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.bin_s1 ;
assign \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.u2.cin  = \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.carry_s1 ;
assign \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.facout_s2  = \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.u2.cout ;
assign \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.fas_s2  = \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.u2.s ;
assign \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.u1.a  = \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.a [7:0];
assign \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.u1.b  = \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.b [7:0];
assign \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.u1.cin  = 1'h0;
assign \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.facout_s1  = \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.u1.cout ;
assign \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.fas_s1  = \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.u1.s ;
assign \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.a  = \add_17ns_17s_17_2_1_U7.din0 ;
assign \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.b  = \add_17ns_17s_17_2_1_U7.din1 ;
assign \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.ce  = \add_17ns_17s_17_2_1_U7.ce ;
assign \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.clk  = \add_17ns_17s_17_2_1_U7.clk ;
assign \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.reset  = \add_17ns_17s_17_2_1_U7.reset ;
assign \add_17ns_17s_17_2_1_U7.dout  = \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.s ;
assign \add_17ns_17s_17_2_1_U7.ce  = 1'h1;
assign \add_17ns_17s_17_2_1_U7.clk  = ap_clk;
assign \add_17ns_17s_17_2_1_U7.din0  = { 3'h0, signbit_reg_835, 13'h0000 };
assign \add_17ns_17s_17_2_1_U7.din1  = { op_7[15], op_7 };
assign grp_fu_330_p2 = \add_17ns_17s_17_2_1_U7.dout ;
assign \add_17ns_17s_17_2_1_U7.reset  = ap_rst;
assign \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.ain_s0  = \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.a ;
assign \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.bin_s0  = \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.b ;
assign \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.s  = { \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.fas_s2 , \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.sum_s1  };
assign \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.u2.a  = \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.ain_s1 ;
assign \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.u2.b  = \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.bin_s1 ;
assign \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.u2.cin  = \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.carry_s1 ;
assign \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.facout_s2  = \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.u2.cout ;
assign \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.fas_s2  = \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.u2.s ;
assign \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.u1.a  = \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.a [7:0];
assign \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.u1.b  = \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.b [7:0];
assign \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.u1.cin  = 1'h0;
assign \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.facout_s1  = \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.u1.cout ;
assign \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.fas_s1  = \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.u1.s ;
assign \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.a  = \add_17ns_17ns_17_2_1_U14.din0 ;
assign \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.b  = \add_17ns_17ns_17_2_1_U14.din1 ;
assign \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.ce  = \add_17ns_17ns_17_2_1_U14.ce ;
assign \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.clk  = \add_17ns_17ns_17_2_1_U14.clk ;
assign \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.reset  = \add_17ns_17ns_17_2_1_U14.reset ;
assign \add_17ns_17ns_17_2_1_U14.dout  = \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.s ;
assign \add_17ns_17ns_17_2_1_U14.ce  = 1'h1;
assign \add_17ns_17ns_17_2_1_U14.clk  = ap_clk;
assign \add_17ns_17ns_17_2_1_U14.din0  = { 1'h0, ret_V_15_reg_1000[3], ret_V_15_reg_1000[3], ret_V_15_reg_1000[3], ret_V_15_reg_1000[3], ret_V_15_reg_1000[3], ret_V_15_reg_1000[3], ret_V_15_reg_1000[3], ret_V_15_reg_1000[3], ret_V_15_reg_1000[3], ret_V_15_reg_1000[3], ret_V_15_reg_1000[3], ret_V_15_reg_1000[3], ret_V_15_reg_1000 };
assign \add_17ns_17ns_17_2_1_U14.din1  = { 9'h000, ret_V_16_reg_840[4], ret_V_16_reg_840[4], ret_V_16_reg_840[4], ret_V_16_reg_840 };
assign grp_fu_642_p2 = \add_17ns_17ns_17_2_1_U14.dout ;
assign \add_17ns_17ns_17_2_1_U14.reset  = ap_rst;
endmodule


// Machine B:
// Processed by function `add_clk_enable_signal` in `verilog_tricks.py`.
// Processed by function `remove_reset_signal` in `verilog_tricks.py`.
module top_B (
  ap_clk,
  ap_start,
  ap_done,
  ap_idle,
  ap_ready,
  op_0,
  op_1,
  op_4,
  op_5,
  op_6,
  op_7,
  op_10,
  op_11,
  op_18,
  op_19,
  op_29,
  op_29_ap_vld,
clk_enable
);
input clk_enable;


input ap_clk;
wire ap_rst;
assign ap_rst = op_29_ap_vld;
input ap_start;
input [3:0] op_0;
input [3:0] op_1;
input [3:0] op_10;
input [3:0] op_11;
input [1:0] op_18;
input [3:0] op_19;
input [1:0] op_4;
input [3:0] op_5;
input [3:0] op_6;
input [15:0] op_7;
output ap_done;
output ap_idle;
output ap_ready;
output [31:0] op_29;
output op_29_ap_vld;


reg [8:0] \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.ain_s1 ;
reg [8:0] \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.bin_s1 ;
reg \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.carry_s1 ;
reg [7:0] \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.sum_s1 ;
reg [8:0] \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.ain_s1 ;
reg [8:0] \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.bin_s1 ;
reg \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.carry_s1 ;
reg [7:0] \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.sum_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s1 ;
reg \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.carry_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.sum_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s1 ;
reg \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.carry_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.sum_s1 ;
reg [15:0] \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.ain_s1 ;
reg [15:0] \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.bin_s1 ;
reg \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.carry_s1 ;
reg [15:0] \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.sum_s1 ;
reg [15:0] \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.ain_s1 ;
reg [15:0] \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.bin_s1 ;
reg \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.carry_s1 ;
reg [15:0] \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.sum_s1 ;
reg [16:0] \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.ain_s1 ;
reg [16:0] \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.bin_s1 ;
reg \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.carry_s1 ;
reg [16:0] \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.sum_s1 ;
reg [17:0] \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.ain_s1 ;
reg [17:0] \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.bin_s1 ;
reg \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.carry_s1 ;
reg [17:0] \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.sum_s1 ;
reg [17:0] \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.ain_s1 ;
reg [17:0] \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.bin_s1 ;
reg \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.carry_s1 ;
reg [17:0] \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.sum_s1 ;
reg [1:0] \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.ain_s1 ;
reg [1:0] \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.bin_s1 ;
reg \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.carry_s1 ;
reg [1:0] \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.sum_s1 ;
reg [1:0] \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.ain_s1 ;
reg [1:0] \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.bin_s1 ;
reg \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.carry_s1 ;
reg [1:0] \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.sum_s1 ;
reg [1:0] \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.ain_s1 ;
reg [1:0] \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.bin_s1 ;
reg \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.carry_s1 ;
reg [1:0] \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.sum_s1 ;
reg [2:0] \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.ain_s1 ;
reg [2:0] \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.bin_s1 ;
reg \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.carry_s1 ;
reg [1:0] \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.sum_s1 ;
reg [2:0] \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.ain_s1 ;
reg [2:0] \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.bin_s1 ;
reg \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.carry_s1 ;
reg [2:0] \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.sum_s1 ;
reg [3:0] \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.ain_s1 ;
reg [3:0] \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.bin_s1 ;
reg \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.carry_s1 ;
reg [3:0] \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.sum_s1 ;
reg [31:0] add_ln691_1_reg_995;
reg [5:0] add_ln691_reg_957;
reg [31:0] add_ln69_2_reg_1100;
reg [3:0] add_ln69_3_reg_1105;
reg [16:0] add_ln69_reg_1040;
reg [36:0] ap_CS_fsm = 37'h0000000001;
reg [31:0] \ashr_32s_32s_32_7_1_U5.din1_cast_array[0] ;
reg [31:0] \ashr_32s_32s_32_7_1_U5.din1_cast_array[1] ;
reg [31:0] \ashr_32s_32s_32_7_1_U5.din1_cast_array[2] ;
reg [31:0] \ashr_32s_32s_32_7_1_U5.din1_cast_array[3] ;
reg [31:0] \ashr_32s_32s_32_7_1_U5.din1_cast_array[4] ;
reg [31:0] \ashr_32s_32s_32_7_1_U5.din1_cast_array[5] ;
reg [31:0] \ashr_32s_32s_32_7_1_U5.dout_array[0] ;
reg [31:0] \ashr_32s_32s_32_7_1_U5.dout_array[1] ;
reg [31:0] \ashr_32s_32s_32_7_1_U5.dout_array[2] ;
reg [31:0] \ashr_32s_32s_32_7_1_U5.dout_array[3] ;
reg [31:0] \ashr_32s_32s_32_7_1_U5.dout_array[4] ;
reg [31:0] \ashr_32s_32s_32_7_1_U5.dout_array[5] ;
reg icmp_ln768_reg_939;
reg icmp_ln851_1_reg_907;
reg icmp_ln851_reg_872;
reg icmp_ln890_reg_820;
reg [3:0] \mul_4s_4s_4_7_1_U2.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.a_reg0 ;
reg [3:0] \mul_4s_4s_4_7_1_U2.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.b_reg0 ;
reg [3:0] \mul_4s_4s_4_7_1_U2.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.buff0 ;
reg [3:0] \mul_4s_4s_4_7_1_U2.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.buff1 ;
reg [3:0] \mul_4s_4s_4_7_1_U2.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.buff2 ;
reg [3:0] \mul_4s_4s_4_7_1_U2.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.buff3 ;
reg [3:0] \mul_4s_4s_4_7_1_U2.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.buff4 ;
reg [1:0] op_12_V_reg_962;
reg [1:0] op_17_V_reg_1075;
reg [31:0] op_23_V_reg_1035;
reg [31:0] op_25_V_reg_1055;
reg [31:0] op_26_V_reg_1080;
reg [3:0] op_3_V_reg_793;
reg overflow_reg_951;
reg p_Result_8_reg_918;
reg p_Result_9_reg_912;
reg [4:0] ret_V_14_reg_750;
reg [3:0] ret_V_15_reg_1000;
reg [4:0] ret_V_16_reg_840;
reg [16:0] ret_V_17_reg_855;
reg [7:0] ret_V_18_reg_929;
reg [33:0] ret_V_19_reg_983;
reg [31:0] ret_V_21_cast_reg_988;
reg [3:0] ret_V_2_reg_763;
reg [3:0] ret_V_3_reg_768;
reg [3:0] ret_V_6_reg_1005;
reg [3:0] ret_V_7_reg_860;
reg [3:0] ret_V_9_reg_877;
reg [3:0] ret_V_reg_756;
reg [31:0] select_ln353_1_reg_1010;
reg [5:0] select_ln353_reg_968;
reg [3:0] select_ln850_3_reg_882;
reg [4:0] sext_ln703_3_reg_782;
reg [5:0] sext_ln850_reg_944;
reg [31:0] \shl_32s_32s_32_7_1_U6.din1_cast_array[0] ;
reg [31:0] \shl_32s_32s_32_7_1_U6.din1_cast_array[1] ;
reg [31:0] \shl_32s_32s_32_7_1_U6.din1_cast_array[2] ;
reg [31:0] \shl_32s_32s_32_7_1_U6.din1_cast_array[3] ;
reg [31:0] \shl_32s_32s_32_7_1_U6.din1_cast_array[4] ;
reg [31:0] \shl_32s_32s_32_7_1_U6.din1_cast_array[5] ;
reg [31:0] \shl_32s_32s_32_7_1_U6.dout_array[0] ;
reg [31:0] \shl_32s_32s_32_7_1_U6.dout_array[1] ;
reg [31:0] \shl_32s_32s_32_7_1_U6.dout_array[2] ;
reg [31:0] \shl_32s_32s_32_7_1_U6.dout_array[3] ;
reg [31:0] \shl_32s_32s_32_7_1_U6.dout_array[4] ;
reg [31:0] \shl_32s_32s_32_7_1_U6.dout_array[5] ;
reg signbit_reg_835;
reg \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.ain_s1 ;
reg \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.bin_s1 ;
reg \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.carry_s1 ;
reg \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.sum_s1 ;
reg [2:0] \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.ain_s1 ;
reg [2:0] \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.bin_s1 ;
reg \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.carry_s1 ;
reg [1:0] \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.sum_s1 ;
reg [4:0] sub_ln1497_reg_799;
reg [10:0] tmp_1_reg_924;
reg [4:0] tmp_2_reg_934;
reg tmp_V_reg_1050;
reg tmp_reg_788;
reg [1:0] trunc_ln1347_reg_804;
reg [11:0] trunc_ln1497_1_reg_892;
reg [3:0] trunc_ln1497_reg_887;
reg [12:0] trunc_ln851_1_reg_867;
wire [31:0] _000_;
wire [5:0] _001_;
wire [31:0] _002_;
wire [3:0] _003_;
wire [16:0] _004_;
wire [36:0] _005_;
wire _006_;
wire _007_;
wire _008_;
wire _009_;
wire [1:0] _010_;
wire [1:0] _011_;
wire [31:0] _012_;
wire [31:0] _013_;
wire [31:0] _014_;
wire [3:0] _015_;
wire _016_;
wire _017_;
wire _018_;
wire [4:0] _019_;
wire [3:0] _020_;
wire [4:0] _021_;
wire [16:0] _022_;
wire [7:0] _023_;
wire [33:0] _024_;
wire [31:0] _025_;
wire [3:0] _026_;
wire [3:0] _027_;
wire [3:0] _028_;
wire [3:0] _029_;
wire [3:0] _030_;
wire [3:0] _031_;
wire [31:0] _032_;
wire [5:0] _033_;
wire [3:0] _034_;
wire [4:0] _035_;
wire [5:0] _036_;
wire _037_;
wire [4:0] _038_;
wire [10:0] _039_;
wire [4:0] _040_;
wire _041_;
wire _042_;
wire [1:0] _043_;
wire [11:0] _044_;
wire [3:0] _045_;
wire [12:0] _046_;
wire [1:0] _047_;
wire _048_;
wire _049_;
wire _050_;
wire _051_;
wire _052_;
wire _053_;
wire _054_;
wire _055_;
wire [8:0] _056_;
wire [8:0] _057_;
wire _058_;
wire [7:0] _059_;
wire [8:0] _060_;
wire [9:0] _061_;
wire [8:0] _062_;
wire [8:0] _063_;
wire _064_;
wire [7:0] _065_;
wire [8:0] _066_;
wire [9:0] _067_;
wire [15:0] _068_;
wire [15:0] _069_;
wire _070_;
wire [15:0] _071_;
wire [16:0] _072_;
wire [16:0] _073_;
wire [15:0] _074_;
wire [15:0] _075_;
wire _076_;
wire [15:0] _077_;
wire [16:0] _078_;
wire [16:0] _079_;
wire [15:0] _080_;
wire [15:0] _081_;
wire _082_;
wire [15:0] _083_;
wire [16:0] _084_;
wire [16:0] _085_;
wire [15:0] _086_;
wire [15:0] _087_;
wire _088_;
wire [15:0] _089_;
wire [16:0] _090_;
wire [16:0] _091_;
wire [16:0] _092_;
wire [16:0] _093_;
wire _094_;
wire [16:0] _095_;
wire [17:0] _096_;
wire [17:0] _097_;
wire [17:0] _098_;
wire [17:0] _099_;
wire _100_;
wire [17:0] _101_;
wire [18:0] _102_;
wire [18:0] _103_;
wire [17:0] _104_;
wire [17:0] _105_;
wire _106_;
wire [17:0] _107_;
wire [18:0] _108_;
wire [18:0] _109_;
wire [1:0] _110_;
wire [1:0] _111_;
wire _112_;
wire [1:0] _113_;
wire [2:0] _114_;
wire [2:0] _115_;
wire [1:0] _116_;
wire [1:0] _117_;
wire _118_;
wire [1:0] _119_;
wire [2:0] _120_;
wire [2:0] _121_;
wire [1:0] _122_;
wire [1:0] _123_;
wire _124_;
wire [1:0] _125_;
wire [2:0] _126_;
wire [2:0] _127_;
wire [2:0] _128_;
wire [2:0] _129_;
wire _130_;
wire [1:0] _131_;
wire [2:0] _132_;
wire [3:0] _133_;
wire [2:0] _134_;
wire [2:0] _135_;
wire _136_;
wire [2:0] _137_;
wire [3:0] _138_;
wire [3:0] _139_;
wire [3:0] _140_;
wire [3:0] _141_;
wire _142_;
wire [3:0] _143_;
wire [4:0] _144_;
wire [4:0] _145_;
wire [31:0] _146_;
wire [31:0] _147_;
wire [31:0] _148_;
wire [31:0] _149_;
wire [31:0] _150_;
wire [31:0] _151_;
wire [31:0] _152_;
wire [31:0] _153_;
wire [31:0] _154_;
wire [31:0] _155_;
wire [31:0] _156_;
wire [31:0] _157_;
wire [31:0] _158_;
wire [31:0] _159_;
wire [31:0] _160_;
wire [31:0] _161_;
wire [31:0] _162_;
wire [31:0] _163_;
wire [31:0] _164_;
wire [31:0] _165_;
wire [31:0] _166_;
wire [31:0] _167_;
wire [31:0] _168_;
wire [31:0] _169_;
wire [31:0] _170_;
wire [31:0] _171_;
wire [31:0] _172_;
wire [31:0] _173_;
wire [31:0] _174_;
wire [31:0] _175_;
wire [3:0] _176_;
wire [3:0] _177_;
wire [3:0] _178_;
wire [3:0] _179_;
wire [3:0] _180_;
wire [3:0] _181_;
wire [3:0] _182_;
wire [31:0] _183_;
wire [31:0] _184_;
wire [31:0] _185_;
wire [31:0] _186_;
wire [31:0] _187_;
wire [31:0] _188_;
wire [31:0] _189_;
wire [31:0] _190_;
wire [31:0] _191_;
wire [31:0] _192_;
wire [31:0] _193_;
wire [31:0] _194_;
wire [31:0] _195_;
wire [31:0] _196_;
wire [31:0] _197_;
wire [31:0] _198_;
wire [31:0] _199_;
wire [31:0] _200_;
wire [31:0] _201_;
wire [31:0] _202_;
wire [31:0] _203_;
wire [31:0] _204_;
wire [31:0] _205_;
wire [31:0] _206_;
wire [31:0] _207_;
wire [31:0] _208_;
wire [31:0] _209_;
wire [31:0] _210_;
wire [31:0] _211_;
wire [31:0] _212_;
wire _213_;
wire _214_;
wire _215_;
wire _216_;
wire [1:0] _217_;
wire [1:0] _218_;
wire [2:0] _219_;
wire [2:0] _220_;
wire _221_;
wire [1:0] _222_;
wire [2:0] _223_;
wire [3:0] _224_;
wire _225_;
wire _226_;
wire _227_;
wire _228_;
wire _229_;
wire _230_;
wire _231_;
wire _232_;
wire _233_;
wire _234_;
wire _235_;
wire _236_;
wire _237_;
wire _238_;
wire _239_;
wire _240_;
wire _241_;
wire _242_;
wire _243_;
wire _244_;
wire _245_;
wire _246_;
wire _247_;
wire _248_;
wire _249_;
wire _250_;
wire _251_;
wire _252_;
wire _253_;
wire _254_;
wire _255_;
wire _256_;
wire _257_;
wire _258_;
wire _259_;
wire _260_;
wire _261_;
wire _262_;
wire _263_;
wire _264_;
wire _265_;
wire \add_17ns_17ns_17_2_1_U14.ce ;
wire \add_17ns_17ns_17_2_1_U14.clk ;
wire [16:0] \add_17ns_17ns_17_2_1_U14.din0 ;
wire [16:0] \add_17ns_17ns_17_2_1_U14.din1 ;
wire [16:0] \add_17ns_17ns_17_2_1_U14.dout ;
wire \add_17ns_17ns_17_2_1_U14.reset ;
wire [16:0] \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.a ;
wire [16:0] \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.ain_s0 ;
wire [16:0] \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.b ;
wire [16:0] \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.bin_s0 ;
wire \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.ce ;
wire \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.clk ;
wire \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.facout_s1 ;
wire \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.facout_s2 ;
wire [7:0] \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.fas_s1 ;
wire [8:0] \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.fas_s2 ;
wire \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.reset ;
wire [16:0] \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.s ;
wire [7:0] \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.u1.a ;
wire [7:0] \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.u1.b ;
wire \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.u1.cin ;
wire \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.u1.cout ;
wire [7:0] \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.u1.s ;
wire [8:0] \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.u2.a ;
wire [8:0] \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.u2.b ;
wire \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.u2.cin ;
wire \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.u2.cout ;
wire [8:0] \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.u2.s ;
wire \add_17ns_17s_17_2_1_U7.ce ;
wire \add_17ns_17s_17_2_1_U7.clk ;
wire [16:0] \add_17ns_17s_17_2_1_U7.din0 ;
wire [16:0] \add_17ns_17s_17_2_1_U7.din1 ;
wire [16:0] \add_17ns_17s_17_2_1_U7.dout ;
wire \add_17ns_17s_17_2_1_U7.reset ;
wire [16:0] \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.a ;
wire [16:0] \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.ain_s0 ;
wire [16:0] \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.b ;
wire [16:0] \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.bin_s0 ;
wire \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.ce ;
wire \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.clk ;
wire \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.facout_s1 ;
wire \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.facout_s2 ;
wire [7:0] \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.fas_s1 ;
wire [8:0] \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.fas_s2 ;
wire \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.reset ;
wire [16:0] \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.s ;
wire [7:0] \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.u1.a ;
wire [7:0] \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.u1.b ;
wire \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.u1.cin ;
wire \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.u1.cout ;
wire [7:0] \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.u1.s ;
wire [8:0] \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.u2.a ;
wire [8:0] \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.u2.b ;
wire \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.u2.cin ;
wire \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.u2.cout ;
wire [8:0] \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.u2.s ;
wire \add_32ns_32ns_32_2_1_U12.ce ;
wire \add_32ns_32ns_32_2_1_U12.clk ;
wire [31:0] \add_32ns_32ns_32_2_1_U12.din0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U12.din1 ;
wire [31:0] \add_32ns_32ns_32_2_1_U12.dout ;
wire \add_32ns_32ns_32_2_1_U12.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.a ;
wire [31:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.b ;
wire [31:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s0 ;
wire \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.ce ;
wire \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.clk ;
wire \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.facout_s1 ;
wire \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.facout_s2 ;
wire [15:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s1 ;
wire [15:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s2 ;
wire \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.b ;
wire \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cin ;
wire \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.b ;
wire \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cin ;
wire \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.s ;
wire \add_32ns_32ns_32_2_1_U15.ce ;
wire \add_32ns_32ns_32_2_1_U15.clk ;
wire [31:0] \add_32ns_32ns_32_2_1_U15.din0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U15.din1 ;
wire [31:0] \add_32ns_32ns_32_2_1_U15.dout ;
wire \add_32ns_32ns_32_2_1_U15.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.a ;
wire [31:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.b ;
wire [31:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s0 ;
wire \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.ce ;
wire \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.clk ;
wire \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.facout_s1 ;
wire \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.facout_s2 ;
wire [15:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s1 ;
wire [15:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s2 ;
wire \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.b ;
wire \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cin ;
wire \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.b ;
wire \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cin ;
wire \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.s ;
wire \add_32ns_32s_32_2_1_U18.ce ;
wire \add_32ns_32s_32_2_1_U18.clk ;
wire [31:0] \add_32ns_32s_32_2_1_U18.din0 ;
wire [31:0] \add_32ns_32s_32_2_1_U18.din1 ;
wire [31:0] \add_32ns_32s_32_2_1_U18.dout ;
wire \add_32ns_32s_32_2_1_U18.reset ;
wire [31:0] \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.a ;
wire [31:0] \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.ain_s0 ;
wire [31:0] \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.b ;
wire [31:0] \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.bin_s0 ;
wire \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.ce ;
wire \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.clk ;
wire \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.facout_s1 ;
wire \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.facout_s2 ;
wire [15:0] \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.fas_s1 ;
wire [15:0] \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.fas_s2 ;
wire \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.reset ;
wire [31:0] \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.s ;
wire [15:0] \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.u1.a ;
wire [15:0] \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.u1.b ;
wire \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.u1.cin ;
wire \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.u1.cout ;
wire [15:0] \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.u1.s ;
wire [15:0] \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.u2.a ;
wire [15:0] \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.u2.b ;
wire \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.u2.cin ;
wire \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.u2.cout ;
wire [15:0] \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.u2.s ;
wire \add_32s_32ns_32_2_1_U20.ce ;
wire \add_32s_32ns_32_2_1_U20.clk ;
wire [31:0] \add_32s_32ns_32_2_1_U20.din0 ;
wire [31:0] \add_32s_32ns_32_2_1_U20.din1 ;
wire [31:0] \add_32s_32ns_32_2_1_U20.dout ;
wire \add_32s_32ns_32_2_1_U20.reset ;
wire [31:0] \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.a ;
wire [31:0] \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.ain_s0 ;
wire [31:0] \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.b ;
wire [31:0] \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.bin_s0 ;
wire \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.ce ;
wire \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.clk ;
wire \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.facout_s1 ;
wire \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.facout_s2 ;
wire [15:0] \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.fas_s1 ;
wire [15:0] \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.fas_s2 ;
wire \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.reset ;
wire [31:0] \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.s ;
wire [15:0] \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.u1.a ;
wire [15:0] \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.u1.b ;
wire \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.u1.cin ;
wire \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.u1.cout ;
wire [15:0] \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.u1.s ;
wire [15:0] \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.u2.a ;
wire [15:0] \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.u2.b ;
wire \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.u2.cin ;
wire \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.u2.cout ;
wire [15:0] \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.u2.s ;
wire \add_34s_34s_34_2_1_U11.ce ;
wire \add_34s_34s_34_2_1_U11.clk ;
wire [33:0] \add_34s_34s_34_2_1_U11.din0 ;
wire [33:0] \add_34s_34s_34_2_1_U11.din1 ;
wire [33:0] \add_34s_34s_34_2_1_U11.dout ;
wire \add_34s_34s_34_2_1_U11.reset ;
wire [33:0] \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.a ;
wire [33:0] \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.ain_s0 ;
wire [33:0] \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.b ;
wire [33:0] \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.bin_s0 ;
wire \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.ce ;
wire \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.clk ;
wire \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.facout_s1 ;
wire \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.facout_s2 ;
wire [16:0] \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.fas_s1 ;
wire [16:0] \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.fas_s2 ;
wire \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.reset ;
wire [33:0] \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.s ;
wire [16:0] \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.u1.a ;
wire [16:0] \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.u1.b ;
wire \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.u1.cin ;
wire \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.u1.cout ;
wire [16:0] \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.u1.s ;
wire [16:0] \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.u2.a ;
wire [16:0] \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.u2.b ;
wire \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.u2.cin ;
wire \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.u2.cout ;
wire [16:0] \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.u2.s ;
wire \add_36ns_36ns_36_2_1_U17.ce ;
wire \add_36ns_36ns_36_2_1_U17.clk ;
wire [35:0] \add_36ns_36ns_36_2_1_U17.din0 ;
wire [35:0] \add_36ns_36ns_36_2_1_U17.din1 ;
wire [35:0] \add_36ns_36ns_36_2_1_U17.dout ;
wire \add_36ns_36ns_36_2_1_U17.reset ;
wire [35:0] \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.a ;
wire [35:0] \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.ain_s0 ;
wire [35:0] \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.b ;
wire [35:0] \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.bin_s0 ;
wire \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.ce ;
wire \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.clk ;
wire \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.facout_s1 ;
wire \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.facout_s2 ;
wire [17:0] \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.fas_s1 ;
wire [17:0] \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.fas_s2 ;
wire \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.reset ;
wire [35:0] \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.s ;
wire [17:0] \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.u1.a ;
wire [17:0] \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.u1.b ;
wire \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.u1.cin ;
wire \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.u1.cout ;
wire [17:0] \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.u1.s ;
wire [17:0] \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.u2.a ;
wire [17:0] \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.u2.b ;
wire \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.u2.cin ;
wire \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.u2.cout ;
wire [17:0] \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.u2.s ;
wire \add_36ns_36s_36_2_1_U13.ce ;
wire \add_36ns_36s_36_2_1_U13.clk ;
wire [35:0] \add_36ns_36s_36_2_1_U13.din0 ;
wire [35:0] \add_36ns_36s_36_2_1_U13.din1 ;
wire [35:0] \add_36ns_36s_36_2_1_U13.dout ;
wire \add_36ns_36s_36_2_1_U13.reset ;
wire [35:0] \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.a ;
wire [35:0] \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.ain_s0 ;
wire [35:0] \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.b ;
wire [35:0] \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.bin_s0 ;
wire \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.ce ;
wire \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.clk ;
wire \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.facout_s1 ;
wire \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.facout_s2 ;
wire [17:0] \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.fas_s1 ;
wire [17:0] \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.fas_s2 ;
wire \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.reset ;
wire [35:0] \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.s ;
wire [17:0] \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.u1.a ;
wire [17:0] \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.u1.b ;
wire \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.u1.cin ;
wire \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.u1.cout ;
wire [17:0] \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.u1.s ;
wire [17:0] \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.u2.a ;
wire [17:0] \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.u2.b ;
wire \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.u2.cin ;
wire \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.u2.cout ;
wire [17:0] \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.u2.s ;
wire \add_4ns_4ns_4_2_1_U1.ce ;
wire \add_4ns_4ns_4_2_1_U1.clk ;
wire [3:0] \add_4ns_4ns_4_2_1_U1.din0 ;
wire [3:0] \add_4ns_4ns_4_2_1_U1.din1 ;
wire [3:0] \add_4ns_4ns_4_2_1_U1.dout ;
wire \add_4ns_4ns_4_2_1_U1.reset ;
wire [3:0] \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.a ;
wire [3:0] \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.ain_s0 ;
wire [3:0] \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.b ;
wire [3:0] \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.bin_s0 ;
wire \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.ce ;
wire \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.clk ;
wire \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.facout_s1 ;
wire \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.facout_s2 ;
wire [1:0] \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.fas_s1 ;
wire [1:0] \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.fas_s2 ;
wire \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.reset ;
wire [3:0] \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.s ;
wire [1:0] \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.u1.a ;
wire [1:0] \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.u1.b ;
wire \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.u1.cin ;
wire \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.u1.cout ;
wire [1:0] \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.u1.s ;
wire [1:0] \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.u2.a ;
wire [1:0] \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.u2.b ;
wire \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.u2.cin ;
wire \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.u2.cout ;
wire [1:0] \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.u2.s ;
wire \add_4ns_4ns_4_2_1_U8.ce ;
wire \add_4ns_4ns_4_2_1_U8.clk ;
wire [3:0] \add_4ns_4ns_4_2_1_U8.din0 ;
wire [3:0] \add_4ns_4ns_4_2_1_U8.din1 ;
wire [3:0] \add_4ns_4ns_4_2_1_U8.dout ;
wire \add_4ns_4ns_4_2_1_U8.reset ;
wire [3:0] \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.a ;
wire [3:0] \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.ain_s0 ;
wire [3:0] \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.b ;
wire [3:0] \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.bin_s0 ;
wire \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.ce ;
wire \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.clk ;
wire \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.facout_s1 ;
wire \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.facout_s2 ;
wire [1:0] \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.fas_s1 ;
wire [1:0] \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.fas_s2 ;
wire \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.reset ;
wire [3:0] \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.s ;
wire [1:0] \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.u1.a ;
wire [1:0] \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.u1.b ;
wire \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.u1.cin ;
wire \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.u1.cout ;
wire [1:0] \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.u1.s ;
wire [1:0] \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.u2.a ;
wire [1:0] \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.u2.b ;
wire \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.u2.cin ;
wire \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.u2.cout ;
wire [1:0] \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.u2.s ;
wire \add_4ns_4s_4_2_1_U19.ce ;
wire \add_4ns_4s_4_2_1_U19.clk ;
wire [3:0] \add_4ns_4s_4_2_1_U19.din0 ;
wire [3:0] \add_4ns_4s_4_2_1_U19.din1 ;
wire [3:0] \add_4ns_4s_4_2_1_U19.dout ;
wire \add_4ns_4s_4_2_1_U19.reset ;
wire [3:0] \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.a ;
wire [3:0] \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.ain_s0 ;
wire [3:0] \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.b ;
wire [3:0] \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.bin_s0 ;
wire \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.ce ;
wire \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.clk ;
wire \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.facout_s1 ;
wire \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.facout_s2 ;
wire [1:0] \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.fas_s1 ;
wire [1:0] \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.fas_s2 ;
wire \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.reset ;
wire [3:0] \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.s ;
wire [1:0] \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.u1.a ;
wire [1:0] \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.u1.b ;
wire \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.u1.cin ;
wire \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.u1.cout ;
wire [1:0] \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.u1.s ;
wire [1:0] \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.u2.a ;
wire [1:0] \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.u2.b ;
wire \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.u2.cin ;
wire \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.u2.cout ;
wire [1:0] \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.u2.s ;
wire \add_5s_5s_5_2_1_U4.ce ;
wire \add_5s_5s_5_2_1_U4.clk ;
wire [4:0] \add_5s_5s_5_2_1_U4.din0 ;
wire [4:0] \add_5s_5s_5_2_1_U4.din1 ;
wire [4:0] \add_5s_5s_5_2_1_U4.dout ;
wire \add_5s_5s_5_2_1_U4.reset ;
wire [4:0] \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.a ;
wire [4:0] \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.ain_s0 ;
wire [4:0] \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.b ;
wire [4:0] \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.bin_s0 ;
wire \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.ce ;
wire \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.clk ;
wire \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.facout_s1 ;
wire \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.facout_s2 ;
wire [1:0] \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.fas_s1 ;
wire [2:0] \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.fas_s2 ;
wire \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.reset ;
wire [4:0] \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.s ;
wire [1:0] \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.u1.a ;
wire [1:0] \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.u1.b ;
wire \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.u1.cin ;
wire \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.u1.cout ;
wire [1:0] \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.u1.s ;
wire [2:0] \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.u2.a ;
wire [2:0] \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.u2.b ;
wire \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.u2.cin ;
wire \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.u2.cout ;
wire [2:0] \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.u2.s ;
wire \add_6s_6ns_6_2_1_U10.ce ;
wire \add_6s_6ns_6_2_1_U10.clk ;
wire [5:0] \add_6s_6ns_6_2_1_U10.din0 ;
wire [5:0] \add_6s_6ns_6_2_1_U10.din1 ;
wire [5:0] \add_6s_6ns_6_2_1_U10.dout ;
wire \add_6s_6ns_6_2_1_U10.reset ;
wire [5:0] \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.a ;
wire [5:0] \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.ain_s0 ;
wire [5:0] \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.b ;
wire [5:0] \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.bin_s0 ;
wire \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.ce ;
wire \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.clk ;
wire \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.facout_s1 ;
wire \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.facout_s2 ;
wire [2:0] \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.fas_s1 ;
wire [2:0] \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.fas_s2 ;
wire \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.reset ;
wire [5:0] \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.s ;
wire [2:0] \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.u1.a ;
wire [2:0] \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.u1.b ;
wire \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.u1.cin ;
wire \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.u1.cout ;
wire [2:0] \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.u1.s ;
wire [2:0] \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.u2.a ;
wire [2:0] \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.u2.b ;
wire \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.u2.cin ;
wire \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.u2.cout ;
wire [2:0] \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.u2.s ;
wire \add_8s_8s_8_2_1_U9.ce ;
wire \add_8s_8s_8_2_1_U9.clk ;
wire [7:0] \add_8s_8s_8_2_1_U9.din0 ;
wire [7:0] \add_8s_8s_8_2_1_U9.din1 ;
wire [7:0] \add_8s_8s_8_2_1_U9.dout ;
wire \add_8s_8s_8_2_1_U9.reset ;
wire [7:0] \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.a ;
wire [7:0] \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.ain_s0 ;
wire [7:0] \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.b ;
wire [7:0] \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.bin_s0 ;
wire \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.ce ;
wire \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.clk ;
wire \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.facout_s1 ;
wire \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.facout_s2 ;
wire [3:0] \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.fas_s1 ;
wire [3:0] \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.fas_s2 ;
wire \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.reset ;
wire [7:0] \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.s ;
wire [3:0] \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.u1.a ;
wire [3:0] \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.u1.b ;
wire \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.u1.cin ;
wire \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.u1.cout ;
wire [3:0] \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.u1.s ;
wire [3:0] \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.u2.a ;
wire [3:0] \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.u2.b ;
wire \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.u2.cin ;
wire \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.u2.cout ;
wire [3:0] \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.u2.s ;
wire ap_CS_fsm_state1;
wire ap_CS_fsm_state10;
wire ap_CS_fsm_state11;
wire ap_CS_fsm_state12;
wire ap_CS_fsm_state13;
wire ap_CS_fsm_state14;
wire ap_CS_fsm_state15;
wire ap_CS_fsm_state16;
wire ap_CS_fsm_state17;
wire ap_CS_fsm_state18;
wire ap_CS_fsm_state19;
wire ap_CS_fsm_state2;
wire ap_CS_fsm_state20;
wire ap_CS_fsm_state21;
wire ap_CS_fsm_state22;
wire ap_CS_fsm_state23;
wire ap_CS_fsm_state24;
wire ap_CS_fsm_state25;
wire ap_CS_fsm_state26;
wire ap_CS_fsm_state27;
wire ap_CS_fsm_state28;
wire ap_CS_fsm_state29;
wire ap_CS_fsm_state3;
wire ap_CS_fsm_state30;
wire ap_CS_fsm_state31;
wire ap_CS_fsm_state32;
wire ap_CS_fsm_state33;
wire ap_CS_fsm_state34;
wire ap_CS_fsm_state35;
wire ap_CS_fsm_state36;
wire ap_CS_fsm_state37;
wire ap_CS_fsm_state4;
wire ap_CS_fsm_state5;
wire [36:0] ap_NS_fsm;
wire ap_clk;
wire ap_done;
wire ap_idle;
wire ap_ready;
wire ap_rst;
wire ap_start;
wire \ashr_32s_32s_32_7_1_U5.ce ;
wire \ashr_32s_32s_32_7_1_U5.clk ;
wire [31:0] \ashr_32s_32s_32_7_1_U5.din0 ;
wire [31:0] \ashr_32s_32s_32_7_1_U5.din1 ;
wire [31:0] \ashr_32s_32s_32_7_1_U5.din1_cast ;
wire [31:0] \ashr_32s_32s_32_7_1_U5.din1_mask ;
wire [31:0] \ashr_32s_32s_32_7_1_U5.dout ;
wire \ashr_32s_32s_32_7_1_U5.reset ;
wire [3:0] grp_fu_221_p2;
wire [3:0] grp_fu_249_p2;
wire [4:0] grp_fu_265_p1;
wire [4:0] grp_fu_265_p2;
wire [4:0] grp_fu_279_p1;
wire [4:0] grp_fu_279_p2;
wire [31:0] grp_fu_295_p1;
wire [31:0] grp_fu_295_p2;
wire [31:0] grp_fu_304_p1;
wire [31:0] grp_fu_304_p2;
wire [16:0] grp_fu_330_p0;
wire [16:0] grp_fu_330_p1;
wire [16:0] grp_fu_330_p2;
wire [3:0] grp_fu_355_p2;
wire [7:0] grp_fu_402_p0;
wire [7:0] grp_fu_402_p1;
wire [7:0] grp_fu_402_p2;
wire [5:0] grp_fu_467_p0;
wire [5:0] grp_fu_467_p2;
wire [33:0] grp_fu_547_p0;
wire [33:0] grp_fu_547_p1;
wire [33:0] grp_fu_547_p2;
wire [31:0] grp_fu_563_p2;
wire [35:0] grp_fu_622_p0;
wire [35:0] grp_fu_622_p1;
wire [35:0] grp_fu_622_p2;
wire [16:0] grp_fu_642_p0;
wire [16:0] grp_fu_642_p1;
wire [16:0] grp_fu_642_p2;
wire [31:0] grp_fu_661_p0;
wire [31:0] grp_fu_661_p2;
wire [1:0] grp_fu_675_p1;
wire [1:0] grp_fu_675_p2;
wire [35:0] grp_fu_698_p0;
wire [35:0] grp_fu_698_p1;
wire [35:0] grp_fu_698_p2;
wire [31:0] grp_fu_725_p1;
wire [31:0] grp_fu_725_p2;
wire [3:0] grp_fu_730_p0;
wire [3:0] grp_fu_730_p1;
wire [3:0] grp_fu_730_p2;
wire [31:0] grp_fu_739_p0;
wire [31:0] grp_fu_739_p2;
wire icmp_ln768_fu_459_p2;
wire icmp_ln851_1_fu_412_p2;
wire icmp_ln851_fu_350_p2;
wire [3:0] icmp_ln890_fu_287_p0;
wire icmp_ln890_fu_287_p2;
wire \mul_4s_4s_4_7_1_U2.ce ;
wire \mul_4s_4s_4_7_1_U2.clk ;
wire [3:0] \mul_4s_4s_4_7_1_U2.din0 ;
wire [3:0] \mul_4s_4s_4_7_1_U2.din1 ;
wire [3:0] \mul_4s_4s_4_7_1_U2.dout ;
wire \mul_4s_4s_4_7_1_U2.reset ;
wire [3:0] \mul_4s_4s_4_7_1_U2.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.a ;
wire [3:0] \mul_4s_4s_4_7_1_U2.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.b ;
wire \mul_4s_4s_4_7_1_U2.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.ce ;
wire \mul_4s_4s_4_7_1_U2.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.clk ;
wire [3:0] \mul_4s_4s_4_7_1_U2.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.p ;
wire [3:0] \mul_4s_4s_4_7_1_U2.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.tmp_product ;
wire [3:0] op_0;
wire [3:0] op_1;
wire [3:0] op_10;
wire [3:0] op_11;
wire [1:0] op_12_V_fu_506_p3;
wire [7:0] op_13_V_fu_604_p3;
wire [1:0] op_18;
wire [3:0] op_19;
wire [31:0] op_29;
wire op_29_ap_vld;
wire [1:0] op_4;
wire [3:0] op_5;
wire [3:0] op_6;
wire [15:0] op_7;
wire or_ln384_fu_502_p2;
wire or_ln785_fu_473_p2;
wire overflow_fu_482_p2;
wire p_Result_5_fu_360_p3;
wire p_Result_6_fu_514_p3;
wire p_Result_7_fu_581_p3;
wire p_Result_9_fu_427_p1;
wire p_Result_s_fu_226_p3;
wire [1:0] p_Val2_4_fu_488_p3;
wire [4:0] p_Val2_s_fu_680_p3;
wire [11:0] r_fu_421_p3;
wire [4:0] ret_V_14_fu_205_p2;
wire [3:0] ret_V_15_fu_572_p1;
wire [3:0] ret_V_15_fu_572_p2;
wire [3:0] ret_V_3_fu_242_p3;
wire [3:0] ret_V_6_fu_577_p1;
wire [3:0] ret_V_6_fu_577_p2;
wire [13:0] rhs_1_fu_319_p3;
wire [6:0] rhs_2_fu_391_p3;
wire [3:0] rhs_fu_197_p1;
wire [4:0] rhs_fu_197_p3;
wire [31:0] select_ln353_1_fu_597_p3;
wire [5:0] select_ln353_fu_526_p3;
wire [1:0] select_ln384_fu_495_p3;
wire [3:0] select_ln850_2_fu_367_p3;
wire [3:0] select_ln850_3_fu_372_p3;
wire [5:0] select_ln850_4_fu_521_p3;
wire [31:0] select_ln850_5_fu_591_p3;
wire [3:0] select_ln850_fu_236_p3;
wire [3:0] sext_ln1192_fu_387_p0;
wire [11:0] sext_ln1497_fu_418_p1;
wire [3:0] sext_ln545_fu_292_p0;
wire [7:0] sext_ln69_2_fu_635_p1;
wire [15:0] sext_ln69_fu_628_p1;
wire [3:0] sext_ln703_1_fu_568_p1;
wire [3:0] sext_ln703_2_fu_275_p0;
wire [3:0] sext_ln703_3_fu_253_p0;
wire [4:0] sext_ln703_3_fu_253_p1;
wire [4:0] sext_ln703_fu_193_p1;
wire [5:0] sext_ln850_fu_464_p1;
wire [31:0] sext_ln890_fu_284_p1;
wire \shl_32s_32s_32_7_1_U6.ce ;
wire \shl_32s_32s_32_7_1_U6.clk ;
wire [31:0] \shl_32s_32s_32_7_1_U6.din0 ;
wire [31:0] \shl_32s_32s_32_7_1_U6.din1 ;
wire [31:0] \shl_32s_32s_32_7_1_U6.din1_cast ;
wire [31:0] \shl_32s_32s_32_7_1_U6.din1_mask ;
wire [31:0] \shl_32s_32s_32_7_1_U6.dout ;
wire \shl_32s_32s_32_7_1_U6.reset ;
wire [3:0] signbit_fu_310_p1;
wire signbit_fu_310_p2;
wire \sub_2ns_2ns_2_2_1_U16.ce ;
wire \sub_2ns_2ns_2_2_1_U16.clk ;
wire [1:0] \sub_2ns_2ns_2_2_1_U16.din0 ;
wire [1:0] \sub_2ns_2ns_2_2_1_U16.din1 ;
wire [1:0] \sub_2ns_2ns_2_2_1_U16.dout ;
wire \sub_2ns_2ns_2_2_1_U16.reset ;
wire [1:0] \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.a ;
wire [1:0] \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.ain_s0 ;
wire [1:0] \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.b ;
wire [1:0] \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.bin_s0 ;
wire \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.ce ;
wire \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.clk ;
wire \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.facout_s1 ;
wire \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.facout_s2 ;
wire \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.fas_s1 ;
wire \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.fas_s2 ;
wire \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.reset ;
wire [1:0] \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.s ;
wire \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.u1.a ;
wire \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.u1.b ;
wire \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.u1.cin ;
wire \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.u1.cout ;
wire \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.u1.s ;
wire \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.u2.a ;
wire \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.u2.b ;
wire \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.u2.cin ;
wire \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.u2.cout ;
wire \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.u2.s ;
wire \sub_5ns_5s_5_2_1_U3.ce ;
wire \sub_5ns_5s_5_2_1_U3.clk ;
wire [4:0] \sub_5ns_5s_5_2_1_U3.din0 ;
wire [4:0] \sub_5ns_5s_5_2_1_U3.din1 ;
wire [4:0] \sub_5ns_5s_5_2_1_U3.dout ;
wire \sub_5ns_5s_5_2_1_U3.reset ;
wire [4:0] \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.a ;
wire [4:0] \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.ain_s0 ;
wire [4:0] \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.b ;
wire [4:0] \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.bin_s0 ;
wire \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.ce ;
wire \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.clk ;
wire \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.facout_s1 ;
wire \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.facout_s2 ;
wire [1:0] \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.fas_s1 ;
wire [2:0] \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.fas_s2 ;
wire \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.reset ;
wire [4:0] \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.s ;
wire [1:0] \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.u1.a ;
wire [1:0] \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.u1.b ;
wire \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.u1.cin ;
wire \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.u1.cout ;
wire [1:0] \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.u1.s ;
wire [2:0] \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.u2.a ;
wire [2:0] \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.u2.b ;
wire \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.u2.cin ;
wire \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.u2.cout ;
wire [2:0] \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.u2.s ;
wire [6:0] tmp_6_fu_536_p3;
wire tmp_V_fu_666_p2;
wire [3:0] tmp_fu_257_p1;
wire [1:0] trunc_ln1347_fu_271_p1;
wire [11:0] trunc_ln1497_1_fu_383_p1;
wire [3:0] trunc_ln1497_fu_379_p1;
wire [12:0] trunc_ln851_1_fu_346_p1;
wire [3:0] trunc_ln851_2_fu_408_p0;
wire [2:0] trunc_ln851_2_fu_408_p1;
wire trunc_ln851_3_fu_588_p1;
wire trunc_ln851_fu_233_p1;
wire xor_ln785_fu_477_p2;


assign _048_ = ap_CS_fsm[20] & icmp_ln851_1_reg_907;
assign _049_ = tmp_reg_788 & ap_CS_fsm[17];
assign _050_ = _053_ & ap_CS_fsm[17];
assign _051_ = _054_ & ap_CS_fsm[0];
assign _052_ = ap_start & ap_CS_fsm[0];
assign overflow_fu_482_p2 = xor_ln785_fu_477_p2 & or_ln785_fu_473_p2;
assign ret_V_15_fu_572_p2 = $signed(op_4) & $signed(op_6);
assign xor_ln785_fu_477_p2 = ~ p_Result_8_reg_918;
assign tmp_V_fu_666_p2 = ~ icmp_ln890_reg_820;
assign _053_ = ~ tmp_reg_788;
assign _054_ = ~ ap_start;
assign _055_ = ! trunc_ln851_1_reg_867;
always @(posedge \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.clk )
\add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.bin_s1  <= _057_;
always @(posedge \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.clk )
\add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.ain_s1  <= _056_;
always @(posedge \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.clk )
\add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.sum_s1  <= _059_;
always @(posedge \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.clk )
\add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.carry_s1  <= _058_;
assign _057_ = \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.ce  ? \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.b [16:8] : \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.bin_s1 ;
assign _056_ = \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.ce  ? \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.a [16:8] : \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.ain_s1 ;
assign _058_ = \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.ce  ? \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.facout_s1  : \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.carry_s1 ;
assign _059_ = \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.ce  ? \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.fas_s1  : \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.sum_s1 ;
assign _060_ = \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.u1.a  + \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.u1.b ;
assign { \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.u1.cout , \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.u1.s  } = _060_ + \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.u1.cin ;
assign _061_ = \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.u2.a  + \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.u2.b ;
assign { \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.u2.cout , \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.u2.s  } = _061_ + \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.u2.cin ;
always @(posedge \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.clk )
\add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.bin_s1  <= _063_;
always @(posedge \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.clk )
\add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.ain_s1  <= _062_;
always @(posedge \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.clk )
\add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.sum_s1  <= _065_;
always @(posedge \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.clk )
\add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.carry_s1  <= _064_;
assign _063_ = \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.ce  ? \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.b [16:8] : \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.bin_s1 ;
assign _062_ = \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.ce  ? \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.a [16:8] : \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.ain_s1 ;
assign _064_ = \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.ce  ? \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.facout_s1  : \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.carry_s1 ;
assign _065_ = \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.ce  ? \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.fas_s1  : \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.sum_s1 ;
assign _066_ = \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.u1.a  + \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.u1.b ;
assign { \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.u1.cout , \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.u1.s  } = _066_ + \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.u1.cin ;
assign _067_ = \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.u2.a  + \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.u2.b ;
assign { \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.u2.cout , \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.u2.s  } = _067_ + \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.u2.cin ;
always @(posedge \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.clk )
\add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s1  <= _069_;
always @(posedge \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.clk )
\add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s1  <= _068_;
always @(posedge \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.clk )
\add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.sum_s1  <= _071_;
always @(posedge \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.clk )
\add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.carry_s1  <= _070_;
assign _069_ = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.ce  ? \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.b [31:16] : \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s1 ;
assign _068_ = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.ce  ? \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.a [31:16] : \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s1 ;
assign _070_ = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.ce  ? \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.facout_s1  : \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.carry_s1 ;
assign _071_ = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.ce  ? \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s1  : \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.sum_s1 ;
assign _072_ = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.a  + \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.b ;
assign { \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cout , \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.s  } = _072_ + \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cin ;
assign _073_ = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.a  + \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.b ;
assign { \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cout , \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.s  } = _073_ + \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cin ;
always @(posedge \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.clk )
\add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s1  <= _075_;
always @(posedge \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.clk )
\add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s1  <= _074_;
always @(posedge \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.clk )
\add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.sum_s1  <= _077_;
always @(posedge \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.clk )
\add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.carry_s1  <= _076_;
assign _075_ = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.ce  ? \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.b [31:16] : \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s1 ;
assign _074_ = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.ce  ? \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.a [31:16] : \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s1 ;
assign _076_ = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.ce  ? \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.facout_s1  : \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.carry_s1 ;
assign _077_ = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.ce  ? \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s1  : \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.sum_s1 ;
assign _078_ = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.a  + \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.b ;
assign { \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cout , \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.s  } = _078_ + \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cin ;
assign _079_ = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.a  + \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.b ;
assign { \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cout , \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.s  } = _079_ + \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cin ;
always @(posedge \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.clk )
\add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.bin_s1  <= _081_;
always @(posedge \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.clk )
\add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.ain_s1  <= _080_;
always @(posedge \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.clk )
\add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.sum_s1  <= _083_;
always @(posedge \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.clk )
\add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.carry_s1  <= _082_;
assign _081_ = \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.ce  ? \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.b [31:16] : \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.bin_s1 ;
assign _080_ = \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.ce  ? \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.a [31:16] : \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.ain_s1 ;
assign _082_ = \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.ce  ? \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.facout_s1  : \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.carry_s1 ;
assign _083_ = \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.ce  ? \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.fas_s1  : \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.sum_s1 ;
assign _084_ = \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.u1.a  + \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.u1.b ;
assign { \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.u1.cout , \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.u1.s  } = _084_ + \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.u1.cin ;
assign _085_ = \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.u2.a  + \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.u2.b ;
assign { \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.u2.cout , \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.u2.s  } = _085_ + \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.u2.cin ;
always @(posedge \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.clk )
\add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.bin_s1  <= _087_;
always @(posedge \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.clk )
\add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.ain_s1  <= _086_;
always @(posedge \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.clk )
\add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.sum_s1  <= _089_;
always @(posedge \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.clk )
\add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.carry_s1  <= _088_;
assign _087_ = \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.ce  ? \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.b [31:16] : \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.bin_s1 ;
assign _086_ = \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.ce  ? \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.a [31:16] : \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.ain_s1 ;
assign _088_ = \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.ce  ? \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.facout_s1  : \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.carry_s1 ;
assign _089_ = \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.ce  ? \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.fas_s1  : \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.sum_s1 ;
assign _090_ = \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.u1.a  + \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.u1.b ;
assign { \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.u1.cout , \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.u1.s  } = _090_ + \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.u1.cin ;
assign _091_ = \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.u2.a  + \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.u2.b ;
assign { \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.u2.cout , \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.u2.s  } = _091_ + \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.u2.cin ;
always @(posedge \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.clk )
\add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.bin_s1  <= _093_;
always @(posedge \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.clk )
\add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.ain_s1  <= _092_;
always @(posedge \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.clk )
\add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.sum_s1  <= _095_;
always @(posedge \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.clk )
\add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.carry_s1  <= _094_;
assign _093_ = \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.ce  ? \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.b [33:17] : \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.bin_s1 ;
assign _092_ = \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.ce  ? \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.a [33:17] : \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.ain_s1 ;
assign _094_ = \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.ce  ? \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.facout_s1  : \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.carry_s1 ;
assign _095_ = \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.ce  ? \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.fas_s1  : \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.sum_s1 ;
assign _096_ = \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.u1.a  + \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.u1.b ;
assign { \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.u1.cout , \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.u1.s  } = _096_ + \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.u1.cin ;
assign _097_ = \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.u2.a  + \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.u2.b ;
assign { \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.u2.cout , \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.u2.s  } = _097_ + \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.u2.cin ;
always @(posedge \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.clk )
\add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.bin_s1  <= _099_;
always @(posedge \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.clk )
\add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.ain_s1  <= _098_;
always @(posedge \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.clk )
\add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.sum_s1  <= _101_;
always @(posedge \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.clk )
\add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.carry_s1  <= _100_;
assign _099_ = \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.ce  ? \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.b [35:18] : \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.bin_s1 ;
assign _098_ = \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.ce  ? \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.a [35:18] : \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.ain_s1 ;
assign _100_ = \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.ce  ? \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.facout_s1  : \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.carry_s1 ;
assign _101_ = \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.ce  ? \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.fas_s1  : \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.sum_s1 ;
assign _102_ = \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.u1.a  + \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.u1.b ;
assign { \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.u1.cout , \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.u1.s  } = _102_ + \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.u1.cin ;
assign _103_ = \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.u2.a  + \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.u2.b ;
assign { \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.u2.cout , \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.u2.s  } = _103_ + \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.u2.cin ;
always @(posedge \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.clk )
\add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.bin_s1  <= _105_;
always @(posedge \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.clk )
\add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.ain_s1  <= _104_;
always @(posedge \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.clk )
\add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.sum_s1  <= _107_;
always @(posedge \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.clk )
\add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.carry_s1  <= _106_;
assign _105_ = \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.ce  ? \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.b [35:18] : \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.bin_s1 ;
assign _104_ = \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.ce  ? \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.a [35:18] : \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.ain_s1 ;
assign _106_ = \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.ce  ? \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.facout_s1  : \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.carry_s1 ;
assign _107_ = \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.ce  ? \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.fas_s1  : \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.sum_s1 ;
assign _108_ = \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.u1.a  + \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.u1.b ;
assign { \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.u1.cout , \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.u1.s  } = _108_ + \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.u1.cin ;
assign _109_ = \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.u2.a  + \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.u2.b ;
assign { \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.u2.cout , \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.u2.s  } = _109_ + \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.u2.cin ;
always @(posedge \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.clk )
\add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.bin_s1  <= _111_;
always @(posedge \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.clk )
\add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.ain_s1  <= _110_;
always @(posedge \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.clk )
\add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.sum_s1  <= _113_;
always @(posedge \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.clk )
\add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.carry_s1  <= _112_;
assign _111_ = \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.ce  ? \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.b [3:2] : \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.bin_s1 ;
assign _110_ = \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.ce  ? \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.a [3:2] : \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.ain_s1 ;
assign _112_ = \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.ce  ? \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.facout_s1  : \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.carry_s1 ;
assign _113_ = \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.ce  ? \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.fas_s1  : \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.sum_s1 ;
assign _114_ = \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.u1.a  + \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.u1.b ;
assign { \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.u1.cout , \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.u1.s  } = _114_ + \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.u1.cin ;
assign _115_ = \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.u2.a  + \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.u2.b ;
assign { \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.u2.cout , \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.u2.s  } = _115_ + \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.u2.cin ;
always @(posedge \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.clk )
\add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.bin_s1  <= _117_;
always @(posedge \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.clk )
\add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.ain_s1  <= _116_;
always @(posedge \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.clk )
\add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.sum_s1  <= _119_;
always @(posedge \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.clk )
\add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.carry_s1  <= _118_;
assign _117_ = \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.ce  ? \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.b [3:2] : \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.bin_s1 ;
assign _116_ = \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.ce  ? \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.a [3:2] : \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.ain_s1 ;
assign _118_ = \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.ce  ? \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.facout_s1  : \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.carry_s1 ;
assign _119_ = \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.ce  ? \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.fas_s1  : \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.sum_s1 ;
assign _120_ = \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.u1.a  + \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.u1.b ;
assign { \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.u1.cout , \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.u1.s  } = _120_ + \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.u1.cin ;
assign _121_ = \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.u2.a  + \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.u2.b ;
assign { \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.u2.cout , \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.u2.s  } = _121_ + \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.u2.cin ;
always @(posedge \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.clk )
\add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.bin_s1  <= _123_;
always @(posedge \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.clk )
\add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.ain_s1  <= _122_;
always @(posedge \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.clk )
\add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.sum_s1  <= _125_;
always @(posedge \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.clk )
\add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.carry_s1  <= _124_;
assign _123_ = \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.ce  ? \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.b [3:2] : \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.bin_s1 ;
assign _122_ = \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.ce  ? \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.a [3:2] : \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.ain_s1 ;
assign _124_ = \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.ce  ? \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.facout_s1  : \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.carry_s1 ;
assign _125_ = \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.ce  ? \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.fas_s1  : \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.sum_s1 ;
assign _126_ = \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.u1.a  + \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.u1.b ;
assign { \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.u1.cout , \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.u1.s  } = _126_ + \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.u1.cin ;
assign _127_ = \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.u2.a  + \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.u2.b ;
assign { \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.u2.cout , \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.u2.s  } = _127_ + \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.u2.cin ;
always @(posedge \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.clk )
\add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.bin_s1  <= _129_;
always @(posedge \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.clk )
\add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.ain_s1  <= _128_;
always @(posedge \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.clk )
\add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.sum_s1  <= _131_;
always @(posedge \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.clk )
\add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.carry_s1  <= _130_;
assign _129_ = \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.ce  ? \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.b [4:2] : \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.bin_s1 ;
assign _128_ = \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.ce  ? \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.a [4:2] : \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.ain_s1 ;
assign _130_ = \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.ce  ? \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.facout_s1  : \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.carry_s1 ;
assign _131_ = \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.ce  ? \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.fas_s1  : \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.sum_s1 ;
assign _132_ = \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.u1.a  + \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.u1.b ;
assign { \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.u1.cout , \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.u1.s  } = _132_ + \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.u1.cin ;
assign _133_ = \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.u2.a  + \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.u2.b ;
assign { \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.u2.cout , \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.u2.s  } = _133_ + \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.u2.cin ;
always @(posedge \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.clk )
\add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.bin_s1  <= _135_;
always @(posedge \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.clk )
\add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.ain_s1  <= _134_;
always @(posedge \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.clk )
\add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.sum_s1  <= _137_;
always @(posedge \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.clk )
\add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.carry_s1  <= _136_;
assign _135_ = \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.ce  ? \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.b [5:3] : \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.bin_s1 ;
assign _134_ = \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.ce  ? \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.a [5:3] : \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.ain_s1 ;
assign _136_ = \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.ce  ? \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.facout_s1  : \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.carry_s1 ;
assign _137_ = \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.ce  ? \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.fas_s1  : \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.sum_s1 ;
assign _138_ = \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.u1.a  + \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.u1.b ;
assign { \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.u1.cout , \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.u1.s  } = _138_ + \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.u1.cin ;
assign _139_ = \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.u2.a  + \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.u2.b ;
assign { \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.u2.cout , \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.u2.s  } = _139_ + \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.u2.cin ;
always @(posedge \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.clk )
\add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.bin_s1  <= _141_;
always @(posedge \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.clk )
\add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.ain_s1  <= _140_;
always @(posedge \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.clk )
\add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.sum_s1  <= _143_;
always @(posedge \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.clk )
\add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.carry_s1  <= _142_;
assign _141_ = \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.ce  ? \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.b [7:4] : \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.bin_s1 ;
assign _140_ = \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.ce  ? \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.a [7:4] : \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.ain_s1 ;
assign _142_ = \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.ce  ? \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.facout_s1  : \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.carry_s1 ;
assign _143_ = \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.ce  ? \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.fas_s1  : \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.sum_s1 ;
assign _144_ = \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.u1.a  + \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.u1.b ;
assign { \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.u1.cout , \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.u1.s  } = _144_ + \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.u1.cin ;
assign _145_ = \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.u2.a  + \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.u2.b ;
assign { \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.u2.cout , \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.u2.s  } = _145_ + \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.u2.cin ;
always @(posedge \ashr_32s_32s_32_7_1_U5.clk )
\ashr_32s_32s_32_7_1_U5.dout_array[5]  <= _157_;
always @(posedge \ashr_32s_32s_32_7_1_U5.clk )
\ashr_32s_32s_32_7_1_U5.din1_cast_array[5]  <= _151_;
always @(posedge \ashr_32s_32s_32_7_1_U5.clk )
\ashr_32s_32s_32_7_1_U5.dout_array[4]  <= _156_;
always @(posedge \ashr_32s_32s_32_7_1_U5.clk )
\ashr_32s_32s_32_7_1_U5.din1_cast_array[4]  <= _150_;
always @(posedge \ashr_32s_32s_32_7_1_U5.clk )
\ashr_32s_32s_32_7_1_U5.dout_array[3]  <= _155_;
always @(posedge \ashr_32s_32s_32_7_1_U5.clk )
\ashr_32s_32s_32_7_1_U5.din1_cast_array[3]  <= _149_;
always @(posedge \ashr_32s_32s_32_7_1_U5.clk )
\ashr_32s_32s_32_7_1_U5.dout_array[2]  <= _154_;
always @(posedge \ashr_32s_32s_32_7_1_U5.clk )
\ashr_32s_32s_32_7_1_U5.din1_cast_array[2]  <= _148_;
always @(posedge \ashr_32s_32s_32_7_1_U5.clk )
\ashr_32s_32s_32_7_1_U5.dout_array[1]  <= _153_;
always @(posedge \ashr_32s_32s_32_7_1_U5.clk )
\ashr_32s_32s_32_7_1_U5.din1_cast_array[1]  <= _147_;
always @(posedge \ashr_32s_32s_32_7_1_U5.clk )
\ashr_32s_32s_32_7_1_U5.dout_array[0]  <= _152_;
always @(posedge \ashr_32s_32s_32_7_1_U5.clk )
\ashr_32s_32s_32_7_1_U5.din1_cast_array[0]  <= _146_;
assign _158_ = \ashr_32s_32s_32_7_1_U5.ce  ? \ashr_32s_32s_32_7_1_U5.din1_cast_array[4]  : \ashr_32s_32s_32_7_1_U5.din1_cast_array[5] ;
assign _151_ = \ashr_32s_32s_32_7_1_U5.reset  ? 32'd0 : _158_;
assign _159_ = \ashr_32s_32s_32_7_1_U5.ce  ? _175_ : \ashr_32s_32s_32_7_1_U5.dout_array[5] ;
assign _157_ = \ashr_32s_32s_32_7_1_U5.reset  ? 32'd0 : _159_;
assign _160_ = \ashr_32s_32s_32_7_1_U5.ce  ? \ashr_32s_32s_32_7_1_U5.din1_cast_array[3]  : \ashr_32s_32s_32_7_1_U5.din1_cast_array[4] ;
assign _150_ = \ashr_32s_32s_32_7_1_U5.reset  ? 32'd0 : _160_;
assign _161_ = \ashr_32s_32s_32_7_1_U5.ce  ? _174_ : \ashr_32s_32s_32_7_1_U5.dout_array[4] ;
assign _156_ = \ashr_32s_32s_32_7_1_U5.reset  ? 32'd0 : _161_;
assign _162_ = \ashr_32s_32s_32_7_1_U5.ce  ? \ashr_32s_32s_32_7_1_U5.din1_cast_array[2]  : \ashr_32s_32s_32_7_1_U5.din1_cast_array[3] ;
assign _149_ = \ashr_32s_32s_32_7_1_U5.reset  ? 32'd0 : _162_;
assign _163_ = \ashr_32s_32s_32_7_1_U5.ce  ? _173_ : \ashr_32s_32s_32_7_1_U5.dout_array[3] ;
assign _155_ = \ashr_32s_32s_32_7_1_U5.reset  ? 32'd0 : _163_;
assign _164_ = \ashr_32s_32s_32_7_1_U5.ce  ? \ashr_32s_32s_32_7_1_U5.din1_cast_array[1]  : \ashr_32s_32s_32_7_1_U5.din1_cast_array[2] ;
assign _148_ = \ashr_32s_32s_32_7_1_U5.reset  ? 32'd0 : _164_;
assign _165_ = \ashr_32s_32s_32_7_1_U5.ce  ? _172_ : \ashr_32s_32s_32_7_1_U5.dout_array[2] ;
assign _154_ = \ashr_32s_32s_32_7_1_U5.reset  ? 32'd0 : _165_;
assign _166_ = \ashr_32s_32s_32_7_1_U5.ce  ? \ashr_32s_32s_32_7_1_U5.din1_cast_array[0]  : \ashr_32s_32s_32_7_1_U5.din1_cast_array[1] ;
assign _147_ = \ashr_32s_32s_32_7_1_U5.reset  ? 32'd0 : _166_;
assign _167_ = \ashr_32s_32s_32_7_1_U5.ce  ? _171_ : \ashr_32s_32s_32_7_1_U5.dout_array[1] ;
assign _153_ = \ashr_32s_32s_32_7_1_U5.reset  ? 32'd0 : _167_;
assign _168_ = \ashr_32s_32s_32_7_1_U5.ce  ? \ashr_32s_32s_32_7_1_U5.din1  : \ashr_32s_32s_32_7_1_U5.din1_cast_array[0] ;
assign _146_ = \ashr_32s_32s_32_7_1_U5.reset  ? 32'd0 : _168_;
assign _169_ = \ashr_32s_32s_32_7_1_U5.ce  ? _170_ : \ashr_32s_32s_32_7_1_U5.dout_array[0] ;
assign _152_ = \ashr_32s_32s_32_7_1_U5.reset  ? 32'd0 : _169_;
assign _170_ = $signed(\ashr_32s_32s_32_7_1_U5.din0 ) >>> { \ashr_32s_32s_32_7_1_U5.din1 [31:30], 30'h00000000 };
assign _171_ = $signed(\ashr_32s_32s_32_7_1_U5.dout_array[0] ) >>> { \ashr_32s_32s_32_7_1_U5.din1_cast_array[0] [29:25], 25'h0000000 };
assign _172_ = $signed(\ashr_32s_32s_32_7_1_U5.dout_array[1] ) >>> { \ashr_32s_32s_32_7_1_U5.din1_cast_array[1] [24:20], 20'h00000 };
assign _173_ = $signed(\ashr_32s_32s_32_7_1_U5.dout_array[2] ) >>> { \ashr_32s_32s_32_7_1_U5.din1_cast_array[2] [19:15], 15'h0000 };
assign _174_ = $signed(\ashr_32s_32s_32_7_1_U5.dout_array[3] ) >>> { \ashr_32s_32s_32_7_1_U5.din1_cast_array[3] [14:10], 10'h000 };
assign _175_ = $signed(\ashr_32s_32s_32_7_1_U5.dout_array[4] ) >>> { \ashr_32s_32s_32_7_1_U5.din1_cast_array[4] [9:5], 5'h00 };
assign \ashr_32s_32s_32_7_1_U5.dout  = $signed(\ashr_32s_32s_32_7_1_U5.dout_array[5] ) >>> \ashr_32s_32s_32_7_1_U5.din1_cast_array[5] [4:0];
assign \mul_4s_4s_4_7_1_U2.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.tmp_product  = $signed(\mul_4s_4s_4_7_1_U2.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.a_reg0 ) * $signed(\mul_4s_4s_4_7_1_U2.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.b_reg0 );
always @(posedge \mul_4s_4s_4_7_1_U2.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.clk )
\mul_4s_4s_4_7_1_U2.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.a_reg0  <= _176_;
always @(posedge \mul_4s_4s_4_7_1_U2.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.clk )
\mul_4s_4s_4_7_1_U2.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.b_reg0  <= _177_;
always @(posedge \mul_4s_4s_4_7_1_U2.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.clk )
\mul_4s_4s_4_7_1_U2.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.buff0  <= _178_;
always @(posedge \mul_4s_4s_4_7_1_U2.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.clk )
\mul_4s_4s_4_7_1_U2.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.buff1  <= _179_;
always @(posedge \mul_4s_4s_4_7_1_U2.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.clk )
\mul_4s_4s_4_7_1_U2.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.buff2  <= _180_;
always @(posedge \mul_4s_4s_4_7_1_U2.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.clk )
\mul_4s_4s_4_7_1_U2.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.buff3  <= _181_;
always @(posedge \mul_4s_4s_4_7_1_U2.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.clk )
\mul_4s_4s_4_7_1_U2.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.buff4  <= _182_;
assign _182_ = \mul_4s_4s_4_7_1_U2.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.ce  ? \mul_4s_4s_4_7_1_U2.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.buff3  : \mul_4s_4s_4_7_1_U2.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.buff4 ;
assign _181_ = \mul_4s_4s_4_7_1_U2.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.ce  ? \mul_4s_4s_4_7_1_U2.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.buff2  : \mul_4s_4s_4_7_1_U2.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.buff3 ;
assign _180_ = \mul_4s_4s_4_7_1_U2.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.ce  ? \mul_4s_4s_4_7_1_U2.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.buff1  : \mul_4s_4s_4_7_1_U2.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.buff2 ;
assign _179_ = \mul_4s_4s_4_7_1_U2.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.ce  ? \mul_4s_4s_4_7_1_U2.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.buff0  : \mul_4s_4s_4_7_1_U2.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.buff1 ;
assign _178_ = \mul_4s_4s_4_7_1_U2.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.ce  ? \mul_4s_4s_4_7_1_U2.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.tmp_product  : \mul_4s_4s_4_7_1_U2.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.buff0 ;
assign _177_ = \mul_4s_4s_4_7_1_U2.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.ce  ? \mul_4s_4s_4_7_1_U2.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.b  : \mul_4s_4s_4_7_1_U2.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.b_reg0 ;
assign _176_ = \mul_4s_4s_4_7_1_U2.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.ce  ? \mul_4s_4s_4_7_1_U2.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.a  : \mul_4s_4s_4_7_1_U2.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.a_reg0 ;
always @(posedge \shl_32s_32s_32_7_1_U6.clk )
\shl_32s_32s_32_7_1_U6.dout_array[5]  <= _194_;
always @(posedge \shl_32s_32s_32_7_1_U6.clk )
\shl_32s_32s_32_7_1_U6.din1_cast_array[5]  <= _188_;
always @(posedge \shl_32s_32s_32_7_1_U6.clk )
\shl_32s_32s_32_7_1_U6.dout_array[4]  <= _193_;
always @(posedge \shl_32s_32s_32_7_1_U6.clk )
\shl_32s_32s_32_7_1_U6.din1_cast_array[4]  <= _187_;
always @(posedge \shl_32s_32s_32_7_1_U6.clk )
\shl_32s_32s_32_7_1_U6.dout_array[3]  <= _192_;
always @(posedge \shl_32s_32s_32_7_1_U6.clk )
\shl_32s_32s_32_7_1_U6.din1_cast_array[3]  <= _186_;
always @(posedge \shl_32s_32s_32_7_1_U6.clk )
\shl_32s_32s_32_7_1_U6.dout_array[2]  <= _191_;
always @(posedge \shl_32s_32s_32_7_1_U6.clk )
\shl_32s_32s_32_7_1_U6.din1_cast_array[2]  <= _185_;
always @(posedge \shl_32s_32s_32_7_1_U6.clk )
\shl_32s_32s_32_7_1_U6.dout_array[1]  <= _190_;
always @(posedge \shl_32s_32s_32_7_1_U6.clk )
\shl_32s_32s_32_7_1_U6.din1_cast_array[1]  <= _184_;
always @(posedge \shl_32s_32s_32_7_1_U6.clk )
\shl_32s_32s_32_7_1_U6.dout_array[0]  <= _189_;
always @(posedge \shl_32s_32s_32_7_1_U6.clk )
\shl_32s_32s_32_7_1_U6.din1_cast_array[0]  <= _183_;
assign _195_ = \shl_32s_32s_32_7_1_U6.ce  ? \shl_32s_32s_32_7_1_U6.din1_cast_array[4]  : \shl_32s_32s_32_7_1_U6.din1_cast_array[5] ;
assign _188_ = \shl_32s_32s_32_7_1_U6.reset  ? 32'd0 : _195_;
assign _196_ = \shl_32s_32s_32_7_1_U6.ce  ? _212_ : \shl_32s_32s_32_7_1_U6.dout_array[5] ;
assign _194_ = \shl_32s_32s_32_7_1_U6.reset  ? 32'd0 : _196_;
assign _197_ = \shl_32s_32s_32_7_1_U6.ce  ? \shl_32s_32s_32_7_1_U6.din1_cast_array[3]  : \shl_32s_32s_32_7_1_U6.din1_cast_array[4] ;
assign _187_ = \shl_32s_32s_32_7_1_U6.reset  ? 32'd0 : _197_;
assign _198_ = \shl_32s_32s_32_7_1_U6.ce  ? _211_ : \shl_32s_32s_32_7_1_U6.dout_array[4] ;
assign _193_ = \shl_32s_32s_32_7_1_U6.reset  ? 32'd0 : _198_;
assign _199_ = \shl_32s_32s_32_7_1_U6.ce  ? \shl_32s_32s_32_7_1_U6.din1_cast_array[2]  : \shl_32s_32s_32_7_1_U6.din1_cast_array[3] ;
assign _186_ = \shl_32s_32s_32_7_1_U6.reset  ? 32'd0 : _199_;
assign _200_ = \shl_32s_32s_32_7_1_U6.ce  ? _210_ : \shl_32s_32s_32_7_1_U6.dout_array[3] ;
assign _192_ = \shl_32s_32s_32_7_1_U6.reset  ? 32'd0 : _200_;
assign _201_ = \shl_32s_32s_32_7_1_U6.ce  ? \shl_32s_32s_32_7_1_U6.din1_cast_array[1]  : \shl_32s_32s_32_7_1_U6.din1_cast_array[2] ;
assign _185_ = \shl_32s_32s_32_7_1_U6.reset  ? 32'd0 : _201_;
assign _202_ = \shl_32s_32s_32_7_1_U6.ce  ? _209_ : \shl_32s_32s_32_7_1_U6.dout_array[2] ;
assign _191_ = \shl_32s_32s_32_7_1_U6.reset  ? 32'd0 : _202_;
assign _203_ = \shl_32s_32s_32_7_1_U6.ce  ? \shl_32s_32s_32_7_1_U6.din1_cast_array[0]  : \shl_32s_32s_32_7_1_U6.din1_cast_array[1] ;
assign _184_ = \shl_32s_32s_32_7_1_U6.reset  ? 32'd0 : _203_;
assign _204_ = \shl_32s_32s_32_7_1_U6.ce  ? _208_ : \shl_32s_32s_32_7_1_U6.dout_array[1] ;
assign _190_ = \shl_32s_32s_32_7_1_U6.reset  ? 32'd0 : _204_;
assign _205_ = \shl_32s_32s_32_7_1_U6.ce  ? \shl_32s_32s_32_7_1_U6.din1  : \shl_32s_32s_32_7_1_U6.din1_cast_array[0] ;
assign _183_ = \shl_32s_32s_32_7_1_U6.reset  ? 32'd0 : _205_;
assign _206_ = \shl_32s_32s_32_7_1_U6.ce  ? _207_ : \shl_32s_32s_32_7_1_U6.dout_array[0] ;
assign _189_ = \shl_32s_32s_32_7_1_U6.reset  ? 32'd0 : _206_;
assign _207_ = \shl_32s_32s_32_7_1_U6.din0  << { \shl_32s_32s_32_7_1_U6.din1 [31:30], 30'h00000000 };
assign _208_ = \shl_32s_32s_32_7_1_U6.dout_array[0]  << { \shl_32s_32s_32_7_1_U6.din1_cast_array[0] [29:25], 25'h0000000 };
assign _209_ = \shl_32s_32s_32_7_1_U6.dout_array[1]  << { \shl_32s_32s_32_7_1_U6.din1_cast_array[1] [24:20], 20'h00000 };
assign _210_ = \shl_32s_32s_32_7_1_U6.dout_array[2]  << { \shl_32s_32s_32_7_1_U6.din1_cast_array[2] [19:15], 15'h0000 };
assign _211_ = \shl_32s_32s_32_7_1_U6.dout_array[3]  << { \shl_32s_32s_32_7_1_U6.din1_cast_array[3] [14:10], 10'h000 };
assign _212_ = \shl_32s_32s_32_7_1_U6.dout_array[4]  << { \shl_32s_32s_32_7_1_U6.din1_cast_array[4] [9:5], 5'h00 };
assign \shl_32s_32s_32_7_1_U6.dout  = \shl_32s_32s_32_7_1_U6.dout_array[5]  << \shl_32s_32s_32_7_1_U6.din1_cast_array[5] [4:0];
assign \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.bin_s0  = ~ \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.b ;
always @(posedge \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.clk )
\sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.bin_s1  <= _214_;
always @(posedge \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.clk )
\sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.ain_s1  <= _213_;
always @(posedge \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.clk )
\sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.sum_s1  <= _216_;
always @(posedge \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.clk )
\sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.carry_s1  <= _215_;
assign _214_ = \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.ce  ? \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.bin_s0 [1] : \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.bin_s1 ;
assign _213_ = \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.ce  ? \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.a [1] : \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.ain_s1 ;
assign _215_ = \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.ce  ? \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.facout_s1  : \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.carry_s1 ;
assign _216_ = \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.ce  ? \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.fas_s1  : \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.sum_s1 ;
assign _217_ = \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.u1.a  + \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.u1.b ;
assign { \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.u1.cout , \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.u1.s  } = _217_ + \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.u1.cin ;
assign _218_ = \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.u2.a  + \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.u2.b ;
assign { \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.u2.cout , \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.u2.s  } = _218_ + \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.u2.cin ;
assign \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.bin_s0  = ~ \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.b ;
always @(posedge \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.clk )
\sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.bin_s1  <= _220_;
always @(posedge \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.clk )
\sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.ain_s1  <= _219_;
always @(posedge \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.clk )
\sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.sum_s1  <= _222_;
always @(posedge \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.clk )
\sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.carry_s1  <= _221_;
assign _220_ = \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.ce  ? \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.bin_s0 [4:2] : \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.bin_s1 ;
assign _219_ = \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.ce  ? \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.a [4:2] : \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.ain_s1 ;
assign _221_ = \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.ce  ? \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.facout_s1  : \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.carry_s1 ;
assign _222_ = \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.ce  ? \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.fas_s1  : \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.sum_s1 ;
assign _223_ = \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.u1.a  + \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.u1.b ;
assign { \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.u1.cout , \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.u1.s  } = _223_ + \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.u1.cin ;
assign _224_ = \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.u2.a  + \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.u2.b ;
assign { \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.u2.cout , \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.u2.s  } = _224_ + \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.u2.cin ;
assign _225_ = $signed(op_5) < $signed(ret_V_3_reg_768);
assign _226_ = | tmp_1_reg_924;
assign _227_ = | op_10[2:0];
assign _228_ = op_3_V_reg_793 != op_5;
assign or_ln384_fu_502_p2 = p_Result_8_reg_918 | overflow_reg_951;
assign or_ln785_fu_473_p2 = p_Result_9_reg_912 | icmp_ln768_reg_939;
assign ret_V_6_fu_577_p2 = op_6 | op_3_V_reg_793;
always @(posedge ap_clk)
trunc_ln1497_reg_887 <= _045_;
always @(posedge ap_clk)
trunc_ln1497_1_reg_892 <= _044_;
always @(posedge ap_clk)
sext_ln703_3_reg_782 <= _035_;
always @(posedge ap_clk)
tmp_reg_788 <= _042_;
always @(posedge ap_clk)
select_ln850_3_reg_882 <= _034_;
always @(posedge ap_clk)
ret_V_9_reg_877 <= _030_;
always @(posedge ap_clk)
ret_V_3_reg_768 <= _027_;
always @(posedge ap_clk)
ret_V_2_reg_763 <= _026_;
always @(posedge ap_clk)
ret_V_19_reg_983 <= _024_;
always @(posedge ap_clk)
ret_V_21_cast_reg_988 <= _025_;
always @(posedge ap_clk)
ret_V_17_reg_855 <= _022_;
always @(posedge ap_clk)
ret_V_7_reg_860 <= _029_;
always @(posedge ap_clk)
trunc_ln851_1_reg_867 <= _046_;
always @(posedge ap_clk)
ret_V_16_reg_840 <= _021_;
always @(posedge ap_clk)
ret_V_15_reg_1000 <= _020_;
always @(posedge ap_clk)
ret_V_6_reg_1005 <= _028_;
always @(posedge ap_clk)
select_ln353_1_reg_1010 <= _032_;
always @(posedge ap_clk)
ret_V_14_reg_750 <= _019_;
always @(posedge ap_clk)
ret_V_reg_756 <= _031_;
always @(posedge ap_clk)
p_Result_9_reg_912 <= _018_;
always @(posedge ap_clk)
p_Result_8_reg_918 <= _017_;
always @(posedge ap_clk)
tmp_1_reg_924 <= _039_;
always @(posedge ap_clk)
ret_V_18_reg_929 <= _023_;
always @(posedge ap_clk)
tmp_2_reg_934 <= _040_;
always @(posedge ap_clk)
overflow_reg_951 <= _016_;
always @(posedge ap_clk)
op_3_V_reg_793 <= _015_;
always @(posedge ap_clk)
sub_ln1497_reg_799 <= _038_;
always @(posedge ap_clk)
trunc_ln1347_reg_804 <= _043_;
always @(posedge ap_clk)
tmp_V_reg_1050 <= _041_;
always @(posedge ap_clk)
op_25_V_reg_1055 <= _013_;
always @(posedge ap_clk)
op_17_V_reg_1075 <= _011_;
always @(posedge ap_clk)
op_26_V_reg_1080 <= _014_;
always @(posedge ap_clk)
op_12_V_reg_962 <= _010_;
always @(posedge ap_clk)
select_ln353_reg_968 <= _033_;
always @(posedge ap_clk)
icmp_ln890_reg_820 <= _009_;
always @(posedge ap_clk)
signbit_reg_835 <= _037_;
always @(posedge ap_clk)
icmp_ln851_reg_872 <= _008_;
always @(posedge ap_clk)
icmp_ln851_1_reg_907 <= _007_;
always @(posedge ap_clk)
icmp_ln768_reg_939 <= _006_;
always @(posedge ap_clk)
sext_ln850_reg_944 <= _036_;
always @(posedge ap_clk)
op_23_V_reg_1035 <= _012_;
always @(posedge ap_clk)
add_ln69_reg_1040 <= _004_;
always @(posedge ap_clk)
add_ln69_2_reg_1100 <= _002_;
always @(posedge ap_clk)
add_ln69_3_reg_1105 <= _003_;
always @(posedge ap_clk)
add_ln691_reg_957 <= _001_;
always @(posedge ap_clk)
add_ln691_1_reg_995 <= _000_;
always @(posedge ap_clk)
ap_CS_fsm <= _005_;
assign _047_ = _052_ ? 2'h2 : 2'h1;
assign _229_ = ap_CS_fsm == 1'h1;
function [36:0] _641_;
input [36:0] a;
input [1368:0] b;
input [36:0] s;
case (s)
37'b0000000000000000000000000000000000001:
_641_ = b[36:0];
37'b0000000000000000000000000000000000010:
_641_ = b[73:37];
37'b0000000000000000000000000000000000100:
_641_ = b[110:74];
37'b0000000000000000000000000000000001000:
_641_ = b[147:111];
37'b0000000000000000000000000000000010000:
_641_ = b[184:148];
37'b0000000000000000000000000000000100000:
_641_ = b[221:185];
37'b0000000000000000000000000000001000000:
_641_ = b[258:222];
37'b0000000000000000000000000000010000000:
_641_ = b[295:259];
37'b0000000000000000000000000000100000000:
_641_ = b[332:296];
37'b0000000000000000000000000001000000000:
_641_ = b[369:333];
37'b0000000000000000000000000010000000000:
_641_ = b[406:370];
37'b0000000000000000000000000100000000000:
_641_ = b[443:407];
37'b0000000000000000000000001000000000000:
_641_ = b[480:444];
37'b0000000000000000000000010000000000000:
_641_ = b[517:481];
37'b0000000000000000000000100000000000000:
_641_ = b[554:518];
37'b0000000000000000000001000000000000000:
_641_ = b[591:555];
37'b0000000000000000000010000000000000000:
_641_ = b[628:592];
37'b0000000000000000000100000000000000000:
_641_ = b[665:629];
37'b0000000000000000001000000000000000000:
_641_ = b[702:666];
37'b0000000000000000010000000000000000000:
_641_ = b[739:703];
37'b0000000000000000100000000000000000000:
_641_ = b[776:740];
37'b0000000000000001000000000000000000000:
_641_ = b[813:777];
37'b0000000000000010000000000000000000000:
_641_ = b[850:814];
37'b0000000000000100000000000000000000000:
_641_ = b[887:851];
37'b0000000000001000000000000000000000000:
_641_ = b[924:888];
37'b0000000000010000000000000000000000000:
_641_ = b[961:925];
37'b0000000000100000000000000000000000000:
_641_ = b[998:962];
37'b0000000001000000000000000000000000000:
_641_ = b[1035:999];
37'b0000000010000000000000000000000000000:
_641_ = b[1072:1036];
37'b0000000100000000000000000000000000000:
_641_ = b[1109:1073];
37'b0000001000000000000000000000000000000:
_641_ = b[1146:1110];
37'b0000010000000000000000000000000000000:
_641_ = b[1183:1147];
37'b0000100000000000000000000000000000000:
_641_ = b[1220:1184];
37'b0001000000000000000000000000000000000:
_641_ = b[1257:1221];
37'b0010000000000000000000000000000000000:
_641_ = b[1294:1258];
37'b0100000000000000000000000000000000000:
_641_ = b[1331:1295];
37'b1000000000000000000000000000000000000:
_641_ = b[1368:1332];
37'b0000000000000000000000000000000000000:
_641_ = a;
default:
_641_ = 37'bx;
endcase
endfunction
assign ap_NS_fsm = _641_(37'hxxxxxxxxxx, { 35'h000000000, _047_, 1332'h000000002000000002000000002000000002000000002000000002000000002000000002000000002000000002000000002000000002000000002000000002000000002000000002000000002000000002000000002000000002000000002000000002000000002000000002000000002000000002000000002000000002000000002000000002000000002000000002000000002000000002000000002000000000000000001 }, { _229_, _265_, _264_, _263_, _262_, _261_, _260_, _259_, _258_, _257_, _256_, _255_, _254_, _253_, _252_, _251_, _250_, _249_, _248_, _247_, _246_, _245_, _244_, _243_, _242_, _241_, _240_, _239_, _238_, _237_, _236_, _235_, _234_, _233_, _232_, _231_, _230_ });
assign _230_ = ap_CS_fsm == 37'h1000000000;
assign _231_ = ap_CS_fsm == 36'h800000000;
assign _232_ = ap_CS_fsm == 35'h400000000;
assign _233_ = ap_CS_fsm == 34'h200000000;
assign _234_ = ap_CS_fsm == 33'h100000000;
assign _235_ = ap_CS_fsm == 32'd2147483648;
assign _236_ = ap_CS_fsm == 31'h40000000;
assign _237_ = ap_CS_fsm == 30'h20000000;
assign _238_ = ap_CS_fsm == 29'h10000000;
assign _239_ = ap_CS_fsm == 28'h8000000;
assign _240_ = ap_CS_fsm == 27'h4000000;
assign _241_ = ap_CS_fsm == 26'h2000000;
assign _242_ = ap_CS_fsm == 25'h1000000;
assign _243_ = ap_CS_fsm == 24'h800000;
assign _244_ = ap_CS_fsm == 23'h400000;
assign _245_ = ap_CS_fsm == 22'h200000;
assign _246_ = ap_CS_fsm == 21'h100000;
assign _247_ = ap_CS_fsm == 20'h80000;
assign _248_ = ap_CS_fsm == 19'h40000;
assign _249_ = ap_CS_fsm == 18'h20000;
assign _250_ = ap_CS_fsm == 17'h10000;
assign _251_ = ap_CS_fsm == 16'h8000;
assign _252_ = ap_CS_fsm == 15'h4000;
assign _253_ = ap_CS_fsm == 14'h2000;
assign _254_ = ap_CS_fsm == 13'h1000;
assign _255_ = ap_CS_fsm == 12'h800;
assign _256_ = ap_CS_fsm == 11'h400;
assign _257_ = ap_CS_fsm == 10'h200;
assign _258_ = ap_CS_fsm == 9'h100;
assign _259_ = ap_CS_fsm == 8'h80;
assign _260_ = ap_CS_fsm == 7'h40;
assign _261_ = ap_CS_fsm == 6'h20;
assign _262_ = ap_CS_fsm == 5'h10;
assign _263_ = ap_CS_fsm == 4'h8;
assign _264_ = ap_CS_fsm == 3'h4;
assign _265_ = ap_CS_fsm == 2'h2;
assign op_29_ap_vld = ap_CS_fsm[36] ? 1'h1 : 1'h0;
assign ap_idle = _051_ ? 1'h1 : 1'h0;
assign _045_ = _050_ ? grp_fu_295_p2[3:0] : trunc_ln1497_reg_887;
assign _044_ = _049_ ? grp_fu_304_p2[11:0] : trunc_ln1497_1_reg_892;
assign _042_ = ap_CS_fsm[9] ? op_6[3] : tmp_reg_788;
assign _035_ = ap_CS_fsm[9] ? { op_6[3], op_6 } : sext_ln703_3_reg_782;
assign _034_ = ap_CS_fsm[16] ? select_ln850_3_fu_372_p3 : select_ln850_3_reg_882;
assign _030_ = ap_CS_fsm[15] ? grp_fu_355_p2 : ret_V_9_reg_877;
assign _027_ = ap_CS_fsm[3] ? ret_V_3_fu_242_p3 : ret_V_3_reg_768;
assign _026_ = ap_CS_fsm[2] ? grp_fu_221_p2 : ret_V_2_reg_763;
assign _025_ = ap_CS_fsm[23] ? grp_fu_547_p2[32:1] : ret_V_21_cast_reg_988;
assign _024_ = ap_CS_fsm[23] ? grp_fu_547_p2 : ret_V_19_reg_983;
assign _046_ = ap_CS_fsm[13] ? grp_fu_330_p2[12:0] : trunc_ln851_1_reg_867;
assign _029_ = ap_CS_fsm[13] ? grp_fu_330_p2[16:13] : ret_V_7_reg_860;
assign _022_ = ap_CS_fsm[13] ? grp_fu_330_p2 : ret_V_17_reg_855;
assign _021_ = ap_CS_fsm[12] ? grp_fu_279_p2 : ret_V_16_reg_840;
assign _032_ = ap_CS_fsm[26] ? select_ln353_1_fu_597_p3 : select_ln353_1_reg_1010;
assign _028_ = ap_CS_fsm[26] ? ret_V_6_fu_577_p2 : ret_V_6_reg_1005;
assign _020_ = ap_CS_fsm[26] ? ret_V_15_fu_572_p2 : ret_V_15_reg_1000;
assign _031_ = ap_CS_fsm[0] ? ret_V_14_fu_205_p2[4:1] : ret_V_reg_756;
assign _019_ = ap_CS_fsm[0] ? ret_V_14_fu_205_p2 : ret_V_14_reg_750;
assign _040_ = ap_CS_fsm[18] ? grp_fu_402_p2[7:3] : tmp_2_reg_934;
assign _023_ = ap_CS_fsm[18] ? grp_fu_402_p2 : ret_V_18_reg_929;
assign _039_ = ap_CS_fsm[18] ? r_fu_421_p3[11:1] : tmp_1_reg_924;
assign _017_ = ap_CS_fsm[18] ? r_fu_421_p3[11] : p_Result_8_reg_918;
assign _018_ = ap_CS_fsm[18] ? r_fu_421_p3[0] : p_Result_9_reg_912;
assign _016_ = ap_CS_fsm[20] ? overflow_fu_482_p2 : overflow_reg_951;
assign _043_ = ap_CS_fsm[10] ? grp_fu_249_p2[1:0] : trunc_ln1347_reg_804;
assign _038_ = ap_CS_fsm[10] ? grp_fu_265_p2 : sub_ln1497_reg_799;
assign _015_ = ap_CS_fsm[10] ? grp_fu_249_p2 : op_3_V_reg_793;
assign _013_ = ap_CS_fsm[30] ? grp_fu_661_p2 : op_25_V_reg_1055;
assign _041_ = ap_CS_fsm[30] ? tmp_V_fu_666_p2 : tmp_V_reg_1050;
assign _014_ = ap_CS_fsm[32] ? grp_fu_698_p2[35:4] : op_26_V_reg_1080;
assign _011_ = ap_CS_fsm[32] ? grp_fu_675_p2 : op_17_V_reg_1075;
assign _033_ = ap_CS_fsm[21] ? select_ln353_fu_526_p3 : select_ln353_reg_968;
assign _010_ = ap_CS_fsm[21] ? op_12_V_fu_506_p3 : op_12_V_reg_962;
assign _037_ = ap_CS_fsm[11] ? signbit_fu_310_p2 : signbit_reg_835;
assign _009_ = ap_CS_fsm[11] ? icmp_ln890_fu_287_p2 : icmp_ln890_reg_820;
assign _008_ = ap_CS_fsm[14] ? icmp_ln851_fu_350_p2 : icmp_ln851_reg_872;
assign _007_ = ap_CS_fsm[17] ? icmp_ln851_1_fu_412_p2 : icmp_ln851_1_reg_907;
assign _036_ = ap_CS_fsm[19] ? { tmp_2_reg_934[4], tmp_2_reg_934 } : sext_ln850_reg_944;
assign _006_ = ap_CS_fsm[19] ? icmp_ln768_fu_459_p2 : icmp_ln768_reg_939;
assign _004_ = ap_CS_fsm[28] ? grp_fu_642_p2 : add_ln69_reg_1040;
assign _012_ = ap_CS_fsm[28] ? grp_fu_622_p2[35:4] : op_23_V_reg_1035;
assign _003_ = ap_CS_fsm[34] ? grp_fu_730_p2 : add_ln69_3_reg_1105;
assign _002_ = ap_CS_fsm[34] ? grp_fu_725_p2 : add_ln69_2_reg_1100;
assign _001_ = _048_ ? grp_fu_467_p2 : add_ln691_reg_957;
assign _000_ = ap_CS_fsm[25] ? grp_fu_563_p2 : add_ln691_1_reg_995;
assign _005_ = ap_rst ? 37'h0000000001 : ap_NS_fsm;
assign icmp_ln768_fu_459_p2 = _226_ ? 1'h1 : 1'h0;
assign icmp_ln851_1_fu_412_p2 = _227_ ? 1'h1 : 1'h0;
assign icmp_ln851_fu_350_p2 = _055_ ? 1'h1 : 1'h0;
assign icmp_ln890_fu_287_p2 = _225_ ? 1'h1 : 1'h0;
assign op_12_V_fu_506_p3 = or_ln384_fu_502_p2 ? select_ln384_fu_495_p3 : { p_Result_9_reg_912, 1'h0 };
assign r_fu_421_p3 = tmp_reg_788 ? trunc_ln1497_1_reg_892 : { trunc_ln1497_reg_887[3], trunc_ln1497_reg_887[3], trunc_ln1497_reg_887[3], trunc_ln1497_reg_887[3], trunc_ln1497_reg_887[3], trunc_ln1497_reg_887[3], trunc_ln1497_reg_887[3], trunc_ln1497_reg_887[3], trunc_ln1497_reg_887 };
assign ret_V_3_fu_242_p3 = ret_V_14_reg_750[4] ? select_ln850_fu_236_p3 : ret_V_reg_756;
assign select_ln353_1_fu_597_p3 = ret_V_19_reg_983[33] ? select_ln850_5_fu_591_p3 : ret_V_21_cast_reg_988;
assign select_ln353_fu_526_p3 = ret_V_18_reg_929[7] ? select_ln850_4_fu_521_p3 : sext_ln850_reg_944;
assign select_ln384_fu_495_p3 = overflow_reg_951 ? 2'h1 : 2'h3;
assign select_ln850_2_fu_367_p3 = icmp_ln851_reg_872 ? ret_V_7_reg_860 : ret_V_9_reg_877;
assign select_ln850_3_fu_372_p3 = ret_V_17_reg_855[16] ? select_ln850_2_fu_367_p3 : ret_V_7_reg_860;
assign select_ln850_4_fu_521_p3 = icmp_ln851_1_reg_907 ? add_ln691_reg_957 : sext_ln850_reg_944;
assign select_ln850_5_fu_591_p3 = op_12_V_reg_962[0] ? add_ln691_1_reg_995 : ret_V_21_cast_reg_988;
assign select_ln850_fu_236_p3 = ret_V_14_reg_750[0] ? ret_V_2_reg_763 : ret_V_reg_756;
assign signbit_fu_310_p2 = _228_ ? 1'h1 : 1'h0;
assign ret_V_14_fu_205_p2 = { op_0[3], op_0 } ^ { op_1, 1'h0 };
assign ap_CS_fsm_state1 = ap_CS_fsm[0];
assign ap_CS_fsm_state10 = ap_CS_fsm[9];
assign ap_CS_fsm_state11 = ap_CS_fsm[10];
assign ap_CS_fsm_state12 = ap_CS_fsm[11];
assign ap_CS_fsm_state13 = ap_CS_fsm[12];
assign ap_CS_fsm_state14 = ap_CS_fsm[13];
assign ap_CS_fsm_state15 = ap_CS_fsm[14];
assign ap_CS_fsm_state16 = ap_CS_fsm[15];
assign ap_CS_fsm_state17 = ap_CS_fsm[16];
assign ap_CS_fsm_state18 = ap_CS_fsm[17];
assign ap_CS_fsm_state19 = ap_CS_fsm[18];
assign ap_CS_fsm_state2 = ap_CS_fsm[1];
assign ap_CS_fsm_state20 = ap_CS_fsm[19];
assign ap_CS_fsm_state21 = ap_CS_fsm[20];
assign ap_CS_fsm_state22 = ap_CS_fsm[21];
assign ap_CS_fsm_state23 = ap_CS_fsm[22];
assign ap_CS_fsm_state24 = ap_CS_fsm[23];
assign ap_CS_fsm_state25 = ap_CS_fsm[24];
assign ap_CS_fsm_state26 = ap_CS_fsm[25];
assign ap_CS_fsm_state27 = ap_CS_fsm[26];
assign ap_CS_fsm_state28 = ap_CS_fsm[27];
assign ap_CS_fsm_state29 = ap_CS_fsm[28];
assign ap_CS_fsm_state3 = ap_CS_fsm[2];
assign ap_CS_fsm_state30 = ap_CS_fsm[29];
assign ap_CS_fsm_state31 = ap_CS_fsm[30];
assign ap_CS_fsm_state32 = ap_CS_fsm[31];
assign ap_CS_fsm_state33 = ap_CS_fsm[32];
assign ap_CS_fsm_state34 = ap_CS_fsm[33];
assign ap_CS_fsm_state35 = ap_CS_fsm[34];
assign ap_CS_fsm_state36 = ap_CS_fsm[35];
assign ap_CS_fsm_state37 = ap_CS_fsm[36];
assign ap_CS_fsm_state4 = ap_CS_fsm[3];
assign ap_CS_fsm_state5 = ap_CS_fsm[4];
assign ap_done = op_29_ap_vld;
assign ap_ready = op_29_ap_vld;
assign grp_fu_265_p1 = { op_6[3], op_6 };
assign grp_fu_279_p1 = { op_5[3], op_5 };
assign grp_fu_295_p1 = { op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6 };
assign grp_fu_304_p1 = { sub_ln1497_reg_799[4], sub_ln1497_reg_799[4], sub_ln1497_reg_799[4], sub_ln1497_reg_799[4], sub_ln1497_reg_799[4], sub_ln1497_reg_799[4], sub_ln1497_reg_799[4], sub_ln1497_reg_799[4], sub_ln1497_reg_799[4], sub_ln1497_reg_799[4], sub_ln1497_reg_799[4], sub_ln1497_reg_799[4], sub_ln1497_reg_799[4], sub_ln1497_reg_799[4], sub_ln1497_reg_799[4], sub_ln1497_reg_799[4], sub_ln1497_reg_799[4], sub_ln1497_reg_799[4], sub_ln1497_reg_799[4], sub_ln1497_reg_799[4], sub_ln1497_reg_799[4], sub_ln1497_reg_799[4], sub_ln1497_reg_799[4], sub_ln1497_reg_799[4], sub_ln1497_reg_799[4], sub_ln1497_reg_799[4], sub_ln1497_reg_799[4], sub_ln1497_reg_799 };
assign grp_fu_330_p0 = { 3'h0, signbit_reg_835, 13'h0000 };
assign grp_fu_330_p1 = { op_7[15], op_7 };
assign grp_fu_402_p0 = { select_ln850_3_reg_882[3], select_ln850_3_reg_882, 3'h0 };
assign grp_fu_402_p1 = { op_10[3], op_10[3], op_10[3], op_10[3], op_10 };
assign grp_fu_467_p0 = { tmp_2_reg_934[4], tmp_2_reg_934 };
assign grp_fu_547_p0 = { select_ln353_reg_968[5], select_ln353_reg_968[5], select_ln353_reg_968[5], select_ln353_reg_968[5], select_ln353_reg_968[5], select_ln353_reg_968[5], select_ln353_reg_968[5], select_ln353_reg_968[5], select_ln353_reg_968[5], select_ln353_reg_968[5], select_ln353_reg_968[5], select_ln353_reg_968[5], select_ln353_reg_968[5], select_ln353_reg_968[5], select_ln353_reg_968[5], select_ln353_reg_968[5], select_ln353_reg_968[5], select_ln353_reg_968[5], select_ln353_reg_968[5], select_ln353_reg_968[5], select_ln353_reg_968[5], select_ln353_reg_968[5], select_ln353_reg_968[5], select_ln353_reg_968[5], select_ln353_reg_968[5], select_ln353_reg_968[5], select_ln353_reg_968[5], select_ln353_reg_968, 1'h0 };
assign grp_fu_547_p1 = { op_12_V_reg_962[1], op_12_V_reg_962[1], op_12_V_reg_962[1], op_12_V_reg_962[1], op_12_V_reg_962[1], op_12_V_reg_962[1], op_12_V_reg_962[1], op_12_V_reg_962[1], op_12_V_reg_962[1], op_12_V_reg_962[1], op_12_V_reg_962[1], op_12_V_reg_962[1], op_12_V_reg_962[1], op_12_V_reg_962[1], op_12_V_reg_962[1], op_12_V_reg_962[1], op_12_V_reg_962[1], op_12_V_reg_962[1], op_12_V_reg_962[1], op_12_V_reg_962[1], op_12_V_reg_962[1], op_12_V_reg_962[1], op_12_V_reg_962[1], op_12_V_reg_962[1], op_12_V_reg_962[1], op_12_V_reg_962[1], op_12_V_reg_962[1], op_12_V_reg_962[1], op_12_V_reg_962[1], op_12_V_reg_962[1], op_12_V_reg_962[1], op_12_V_reg_962[1], op_12_V_reg_962 };
assign grp_fu_622_p0 = { select_ln353_1_reg_1010, 4'h0 };
assign grp_fu_622_p1 = { ret_V_6_reg_1005[3], ret_V_6_reg_1005[3], ret_V_6_reg_1005[3], ret_V_6_reg_1005[3], ret_V_6_reg_1005[3], ret_V_6_reg_1005[3], ret_V_6_reg_1005[3], ret_V_6_reg_1005[3], ret_V_6_reg_1005[3], ret_V_6_reg_1005[3], ret_V_6_reg_1005[3], ret_V_6_reg_1005[3], ret_V_6_reg_1005[3], ret_V_6_reg_1005[3], ret_V_6_reg_1005[3], ret_V_6_reg_1005[3], ret_V_6_reg_1005[3], ret_V_6_reg_1005[3], ret_V_6_reg_1005[3], ret_V_6_reg_1005[3], ret_V_6_reg_1005[3], ret_V_6_reg_1005[3], ret_V_6_reg_1005[3], ret_V_6_reg_1005[3], ret_V_6_reg_1005[3], ret_V_6_reg_1005[3], ret_V_6_reg_1005[3], ret_V_6_reg_1005[3], ret_V_6_reg_1005, 4'h0 };
assign grp_fu_642_p0 = { 1'h0, ret_V_15_reg_1000[3], ret_V_15_reg_1000[3], ret_V_15_reg_1000[3], ret_V_15_reg_1000[3], ret_V_15_reg_1000[3], ret_V_15_reg_1000[3], ret_V_15_reg_1000[3], ret_V_15_reg_1000[3], ret_V_15_reg_1000[3], ret_V_15_reg_1000[3], ret_V_15_reg_1000[3], ret_V_15_reg_1000[3], ret_V_15_reg_1000 };
assign grp_fu_642_p1 = { 9'h000, ret_V_16_reg_840[4], ret_V_16_reg_840[4], ret_V_16_reg_840[4], ret_V_16_reg_840 };
assign grp_fu_661_p0 = { 15'h0000, add_ln69_reg_1040 };
assign grp_fu_675_p1 = op_11[1:0];
assign grp_fu_698_p0 = { op_25_V_reg_1055, 4'h0 };
assign grp_fu_698_p1 = { 31'h00000000, tmp_V_reg_1050, 4'h0 };
assign grp_fu_725_p1 = { op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19 };
assign grp_fu_730_p0 = { 2'h0, op_18 };
assign grp_fu_730_p1 = { op_17_V_reg_1075[1], op_17_V_reg_1075[1], op_17_V_reg_1075 };
assign grp_fu_739_p0 = { add_ln69_3_reg_1105[3], add_ln69_3_reg_1105[3], add_ln69_3_reg_1105[3], add_ln69_3_reg_1105[3], add_ln69_3_reg_1105[3], add_ln69_3_reg_1105[3], add_ln69_3_reg_1105[3], add_ln69_3_reg_1105[3], add_ln69_3_reg_1105[3], add_ln69_3_reg_1105[3], add_ln69_3_reg_1105[3], add_ln69_3_reg_1105[3], add_ln69_3_reg_1105[3], add_ln69_3_reg_1105[3], add_ln69_3_reg_1105[3], add_ln69_3_reg_1105[3], add_ln69_3_reg_1105[3], add_ln69_3_reg_1105[3], add_ln69_3_reg_1105[3], add_ln69_3_reg_1105[3], add_ln69_3_reg_1105[3], add_ln69_3_reg_1105[3], add_ln69_3_reg_1105[3], add_ln69_3_reg_1105[3], add_ln69_3_reg_1105[3], add_ln69_3_reg_1105[3], add_ln69_3_reg_1105[3], add_ln69_3_reg_1105[3], add_ln69_3_reg_1105 };
assign icmp_ln890_fu_287_p0 = op_5;
assign op_13_V_fu_604_p3 = { ret_V_6_reg_1005, 4'h0 };
assign op_29 = grp_fu_739_p2;
assign p_Result_5_fu_360_p3 = ret_V_17_reg_855[16];
assign p_Result_6_fu_514_p3 = ret_V_18_reg_929[7];
assign p_Result_7_fu_581_p3 = ret_V_19_reg_983[33];
assign p_Result_9_fu_427_p1 = r_fu_421_p3[0];
assign p_Result_s_fu_226_p3 = ret_V_14_reg_750[4];
assign p_Val2_4_fu_488_p3 = { p_Result_9_reg_912, 1'h0 };
assign p_Val2_s_fu_680_p3 = { tmp_V_reg_1050, 4'h0 };
assign ret_V_15_fu_572_p1 = op_6;
assign ret_V_6_fu_577_p1 = op_6;
assign rhs_1_fu_319_p3 = { signbit_reg_835, 13'h0000 };
assign rhs_2_fu_391_p3 = { select_ln850_3_reg_882, 3'h0 };
assign rhs_fu_197_p1 = op_1;
assign rhs_fu_197_p3 = { op_1, 1'h0 };
assign sext_ln1192_fu_387_p0 = op_10;
assign sext_ln1497_fu_418_p1 = { trunc_ln1497_reg_887[3], trunc_ln1497_reg_887[3], trunc_ln1497_reg_887[3], trunc_ln1497_reg_887[3], trunc_ln1497_reg_887[3], trunc_ln1497_reg_887[3], trunc_ln1497_reg_887[3], trunc_ln1497_reg_887[3], trunc_ln1497_reg_887 };
assign sext_ln545_fu_292_p0 = op_6;
assign sext_ln69_2_fu_635_p1 = { ret_V_16_reg_840[4], ret_V_16_reg_840[4], ret_V_16_reg_840[4], ret_V_16_reg_840 };
assign sext_ln69_fu_628_p1 = { ret_V_15_reg_1000[3], ret_V_15_reg_1000[3], ret_V_15_reg_1000[3], ret_V_15_reg_1000[3], ret_V_15_reg_1000[3], ret_V_15_reg_1000[3], ret_V_15_reg_1000[3], ret_V_15_reg_1000[3], ret_V_15_reg_1000[3], ret_V_15_reg_1000[3], ret_V_15_reg_1000[3], ret_V_15_reg_1000[3], ret_V_15_reg_1000 };
assign sext_ln703_1_fu_568_p1 = { op_4[1], op_4[1], op_4 };
assign sext_ln703_2_fu_275_p0 = op_5;
assign sext_ln703_3_fu_253_p0 = op_6;
assign sext_ln703_3_fu_253_p1 = { op_6[3], op_6 };
assign sext_ln703_fu_193_p1 = { op_0[3], op_0 };
assign sext_ln850_fu_464_p1 = { tmp_2_reg_934[4], tmp_2_reg_934 };
assign sext_ln890_fu_284_p1 = { ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768 };
assign signbit_fu_310_p1 = op_5;
assign tmp_6_fu_536_p3 = { select_ln353_reg_968, 1'h0 };
assign tmp_fu_257_p1 = op_6;
assign trunc_ln1347_fu_271_p1 = grp_fu_249_p2[1:0];
assign trunc_ln1497_1_fu_383_p1 = grp_fu_304_p2[11:0];
assign trunc_ln1497_fu_379_p1 = grp_fu_295_p2[3:0];
assign trunc_ln851_1_fu_346_p1 = grp_fu_330_p2[12:0];
assign trunc_ln851_2_fu_408_p0 = op_10;
assign trunc_ln851_2_fu_408_p1 = op_10[2:0];
assign trunc_ln851_3_fu_588_p1 = op_12_V_reg_962[0];
assign trunc_ln851_fu_233_p1 = ret_V_14_reg_750[0];
assign \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.ain_s0  = \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.a ;
assign \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.s  = { \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.fas_s2 , \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.sum_s1  };
assign \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.u2.a  = \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.ain_s1 ;
assign \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.u2.b  = \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.bin_s1 ;
assign \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.u2.cin  = \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.carry_s1 ;
assign \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.facout_s2  = \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.u2.cout ;
assign \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.fas_s2  = \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.u2.s ;
assign \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.u1.a  = \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.a [1:0];
assign \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.u1.b  = \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.bin_s0 [1:0];
assign \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.u1.cin  = 1'h1;
assign \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.facout_s1  = \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.u1.cout ;
assign \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.fas_s1  = \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.u1.s ;
assign \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.a  = \sub_5ns_5s_5_2_1_U3.din0 ;
assign \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.b  = \sub_5ns_5s_5_2_1_U3.din1 ;
assign \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.ce  = \sub_5ns_5s_5_2_1_U3.ce ;
assign \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.clk  = \sub_5ns_5s_5_2_1_U3.clk ;
assign \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.reset  = \sub_5ns_5s_5_2_1_U3.reset ;
assign \sub_5ns_5s_5_2_1_U3.dout  = \sub_5ns_5s_5_2_1_U3.top_sub_5ns_5s_5_2_1_Adder_1_U.s ;
assign \sub_5ns_5s_5_2_1_U3.ce  = 1'h1;
assign \sub_5ns_5s_5_2_1_U3.clk  = ap_clk;
assign \sub_5ns_5s_5_2_1_U3.din0  = 5'h00;
assign \sub_5ns_5s_5_2_1_U3.din1  = { op_6[3], op_6 };
assign grp_fu_265_p2 = \sub_5ns_5s_5_2_1_U3.dout ;
assign \sub_5ns_5s_5_2_1_U3.reset  = ap_rst;
assign \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.ain_s0  = \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.a ;
assign \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.s  = { \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.fas_s2 , \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.sum_s1  };
assign \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.u2.a  = \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.ain_s1 ;
assign \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.u2.b  = \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.bin_s1 ;
assign \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.u2.cin  = \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.carry_s1 ;
assign \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.facout_s2  = \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.u2.cout ;
assign \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.fas_s2  = \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.u2.s ;
assign \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.u1.a  = \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.a [0];
assign \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.u1.b  = \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.bin_s0 [0];
assign \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.u1.cin  = 1'h1;
assign \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.facout_s1  = \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.u1.cout ;
assign \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.fas_s1  = \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.u1.s ;
assign \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.a  = \sub_2ns_2ns_2_2_1_U16.din0 ;
assign \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.b  = \sub_2ns_2ns_2_2_1_U16.din1 ;
assign \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.ce  = \sub_2ns_2ns_2_2_1_U16.ce ;
assign \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.clk  = \sub_2ns_2ns_2_2_1_U16.clk ;
assign \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.reset  = \sub_2ns_2ns_2_2_1_U16.reset ;
assign \sub_2ns_2ns_2_2_1_U16.dout  = \sub_2ns_2ns_2_2_1_U16.top_sub_2ns_2ns_2_2_1_Adder_10_U.s ;
assign \sub_2ns_2ns_2_2_1_U16.ce  = 1'h1;
assign \sub_2ns_2ns_2_2_1_U16.clk  = ap_clk;
assign \sub_2ns_2ns_2_2_1_U16.din0  = trunc_ln1347_reg_804;
assign \sub_2ns_2ns_2_2_1_U16.din1  = op_11[1:0];
assign grp_fu_675_p2 = \sub_2ns_2ns_2_2_1_U16.dout ;
assign \sub_2ns_2ns_2_2_1_U16.reset  = ap_rst;
assign \shl_32s_32s_32_7_1_U6.din1_cast  = \shl_32s_32s_32_7_1_U6.din1 ;
assign \shl_32s_32s_32_7_1_U6.din1_mask  = 32'd31;
assign \shl_32s_32s_32_7_1_U6.ce  = 1'h1;
assign \shl_32s_32s_32_7_1_U6.clk  = ap_clk;
assign \shl_32s_32s_32_7_1_U6.din0  = { ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768 };
assign \shl_32s_32s_32_7_1_U6.din1  = { sub_ln1497_reg_799[4], sub_ln1497_reg_799[4], sub_ln1497_reg_799[4], sub_ln1497_reg_799[4], sub_ln1497_reg_799[4], sub_ln1497_reg_799[4], sub_ln1497_reg_799[4], sub_ln1497_reg_799[4], sub_ln1497_reg_799[4], sub_ln1497_reg_799[4], sub_ln1497_reg_799[4], sub_ln1497_reg_799[4], sub_ln1497_reg_799[4], sub_ln1497_reg_799[4], sub_ln1497_reg_799[4], sub_ln1497_reg_799[4], sub_ln1497_reg_799[4], sub_ln1497_reg_799[4], sub_ln1497_reg_799[4], sub_ln1497_reg_799[4], sub_ln1497_reg_799[4], sub_ln1497_reg_799[4], sub_ln1497_reg_799[4], sub_ln1497_reg_799[4], sub_ln1497_reg_799[4], sub_ln1497_reg_799[4], sub_ln1497_reg_799[4], sub_ln1497_reg_799 };
assign grp_fu_304_p2 = \shl_32s_32s_32_7_1_U6.dout ;
assign \shl_32s_32s_32_7_1_U6.reset  = ap_rst;
assign \mul_4s_4s_4_7_1_U2.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.p  = \mul_4s_4s_4_7_1_U2.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.buff4 ;
assign \mul_4s_4s_4_7_1_U2.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.a  = \mul_4s_4s_4_7_1_U2.din0 ;
assign \mul_4s_4s_4_7_1_U2.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.b  = \mul_4s_4s_4_7_1_U2.din1 ;
assign \mul_4s_4s_4_7_1_U2.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.ce  = \mul_4s_4s_4_7_1_U2.ce ;
assign \mul_4s_4s_4_7_1_U2.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.clk  = \mul_4s_4s_4_7_1_U2.clk ;
assign \mul_4s_4s_4_7_1_U2.dout  = \mul_4s_4s_4_7_1_U2.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.p ;
assign \mul_4s_4s_4_7_1_U2.ce  = 1'h1;
assign \mul_4s_4s_4_7_1_U2.clk  = ap_clk;
assign \mul_4s_4s_4_7_1_U2.din0  = ret_V_3_reg_768;
assign \mul_4s_4s_4_7_1_U2.din1  = op_1;
assign grp_fu_249_p2 = \mul_4s_4s_4_7_1_U2.dout ;
assign \mul_4s_4s_4_7_1_U2.reset  = ap_rst;
assign \ashr_32s_32s_32_7_1_U5.din1_cast  = \ashr_32s_32s_32_7_1_U5.din1 ;
assign \ashr_32s_32s_32_7_1_U5.din1_mask  = 32'd31;
assign \ashr_32s_32s_32_7_1_U5.ce  = 1'h1;
assign \ashr_32s_32s_32_7_1_U5.clk  = ap_clk;
assign \ashr_32s_32s_32_7_1_U5.din0  = { ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768[3], ret_V_3_reg_768 };
assign \ashr_32s_32s_32_7_1_U5.din1  = { op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6 };
assign grp_fu_295_p2 = \ashr_32s_32s_32_7_1_U5.dout ;
assign \ashr_32s_32s_32_7_1_U5.reset  = ap_rst;
assign \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.ain_s0  = \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.a ;
assign \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.bin_s0  = \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.b ;
assign \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.s  = { \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.fas_s2 , \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.sum_s1  };
assign \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.u2.a  = \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.ain_s1 ;
assign \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.u2.b  = \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.bin_s1 ;
assign \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.u2.cin  = \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.carry_s1 ;
assign \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.facout_s2  = \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.u2.cout ;
assign \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.fas_s2  = \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.u2.s ;
assign \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.u1.a  = \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.a [3:0];
assign \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.u1.b  = \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.b [3:0];
assign \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.u1.cin  = 1'h0;
assign \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.facout_s1  = \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.u1.cout ;
assign \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.fas_s1  = \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.u1.s ;
assign \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.a  = \add_8s_8s_8_2_1_U9.din0 ;
assign \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.b  = \add_8s_8s_8_2_1_U9.din1 ;
assign \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.ce  = \add_8s_8s_8_2_1_U9.ce ;
assign \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.clk  = \add_8s_8s_8_2_1_U9.clk ;
assign \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.reset  = \add_8s_8s_8_2_1_U9.reset ;
assign \add_8s_8s_8_2_1_U9.dout  = \add_8s_8s_8_2_1_U9.top_add_8s_8s_8_2_1_Adder_4_U.s ;
assign \add_8s_8s_8_2_1_U9.ce  = 1'h1;
assign \add_8s_8s_8_2_1_U9.clk  = ap_clk;
assign \add_8s_8s_8_2_1_U9.din0  = { select_ln850_3_reg_882[3], select_ln850_3_reg_882, 3'h0 };
assign \add_8s_8s_8_2_1_U9.din1  = { op_10[3], op_10[3], op_10[3], op_10[3], op_10 };
assign grp_fu_402_p2 = \add_8s_8s_8_2_1_U9.dout ;
assign \add_8s_8s_8_2_1_U9.reset  = ap_rst;
assign \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.ain_s0  = \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.a ;
assign \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.bin_s0  = \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.b ;
assign \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.s  = { \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.fas_s2 , \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.sum_s1  };
assign \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.u2.a  = \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.ain_s1 ;
assign \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.u2.b  = \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.bin_s1 ;
assign \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.u2.cin  = \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.carry_s1 ;
assign \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.facout_s2  = \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.u2.cout ;
assign \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.fas_s2  = \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.u2.s ;
assign \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.u1.a  = \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.a [2:0];
assign \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.u1.b  = \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.b [2:0];
assign \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.u1.cin  = 1'h0;
assign \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.facout_s1  = \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.u1.cout ;
assign \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.fas_s1  = \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.u1.s ;
assign \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.a  = \add_6s_6ns_6_2_1_U10.din0 ;
assign \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.b  = \add_6s_6ns_6_2_1_U10.din1 ;
assign \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.ce  = \add_6s_6ns_6_2_1_U10.ce ;
assign \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.clk  = \add_6s_6ns_6_2_1_U10.clk ;
assign \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.reset  = \add_6s_6ns_6_2_1_U10.reset ;
assign \add_6s_6ns_6_2_1_U10.dout  = \add_6s_6ns_6_2_1_U10.top_add_6s_6ns_6_2_1_Adder_5_U.s ;
assign \add_6s_6ns_6_2_1_U10.ce  = 1'h1;
assign \add_6s_6ns_6_2_1_U10.clk  = ap_clk;
assign \add_6s_6ns_6_2_1_U10.din0  = { tmp_2_reg_934[4], tmp_2_reg_934 };
assign \add_6s_6ns_6_2_1_U10.din1  = 6'h01;
assign grp_fu_467_p2 = \add_6s_6ns_6_2_1_U10.dout ;
assign \add_6s_6ns_6_2_1_U10.reset  = ap_rst;
assign \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.ain_s0  = \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.a ;
assign \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.bin_s0  = \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.b ;
assign \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.s  = { \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.fas_s2 , \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.sum_s1  };
assign \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.u2.a  = \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.ain_s1 ;
assign \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.u2.b  = \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.bin_s1 ;
assign \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.u2.cin  = \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.carry_s1 ;
assign \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.facout_s2  = \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.u2.cout ;
assign \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.fas_s2  = \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.u2.s ;
assign \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.u1.a  = \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.a [1:0];
assign \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.u1.b  = \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.b [1:0];
assign \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.u1.cin  = 1'h0;
assign \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.facout_s1  = \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.u1.cout ;
assign \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.fas_s1  = \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.u1.s ;
assign \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.a  = \add_5s_5s_5_2_1_U4.din0 ;
assign \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.b  = \add_5s_5s_5_2_1_U4.din1 ;
assign \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.ce  = \add_5s_5s_5_2_1_U4.ce ;
assign \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.clk  = \add_5s_5s_5_2_1_U4.clk ;
assign \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.reset  = \add_5s_5s_5_2_1_U4.reset ;
assign \add_5s_5s_5_2_1_U4.dout  = \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_2_U.s ;
assign \add_5s_5s_5_2_1_U4.ce  = 1'h1;
assign \add_5s_5s_5_2_1_U4.clk  = ap_clk;
assign \add_5s_5s_5_2_1_U4.din0  = sext_ln703_3_reg_782;
assign \add_5s_5s_5_2_1_U4.din1  = { op_5[3], op_5 };
assign grp_fu_279_p2 = \add_5s_5s_5_2_1_U4.dout ;
assign \add_5s_5s_5_2_1_U4.reset  = ap_rst;
assign \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.ain_s0  = \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.a ;
assign \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.bin_s0  = \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.b ;
assign \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.s  = { \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.fas_s2 , \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.sum_s1  };
assign \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.u2.a  = \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.ain_s1 ;
assign \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.u2.b  = \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.bin_s1 ;
assign \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.u2.cin  = \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.carry_s1 ;
assign \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.facout_s2  = \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.u2.cout ;
assign \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.fas_s2  = \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.u2.s ;
assign \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.u1.a  = \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.a [1:0];
assign \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.u1.b  = \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.b [1:0];
assign \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.u1.cin  = 1'h0;
assign \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.facout_s1  = \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.u1.cout ;
assign \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.fas_s1  = \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.u1.s ;
assign \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.a  = \add_4ns_4s_4_2_1_U19.din0 ;
assign \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.b  = \add_4ns_4s_4_2_1_U19.din1 ;
assign \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.ce  = \add_4ns_4s_4_2_1_U19.ce ;
assign \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.clk  = \add_4ns_4s_4_2_1_U19.clk ;
assign \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.reset  = \add_4ns_4s_4_2_1_U19.reset ;
assign \add_4ns_4s_4_2_1_U19.dout  = \add_4ns_4s_4_2_1_U19.top_add_4ns_4s_4_2_1_Adder_13_U.s ;
assign \add_4ns_4s_4_2_1_U19.ce  = 1'h1;
assign \add_4ns_4s_4_2_1_U19.clk  = ap_clk;
assign \add_4ns_4s_4_2_1_U19.din0  = { 2'h0, op_18 };
assign \add_4ns_4s_4_2_1_U19.din1  = { op_17_V_reg_1075[1], op_17_V_reg_1075[1], op_17_V_reg_1075 };
assign grp_fu_730_p2 = \add_4ns_4s_4_2_1_U19.dout ;
assign \add_4ns_4s_4_2_1_U19.reset  = ap_rst;
assign \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.ain_s0  = \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.a ;
assign \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.bin_s0  = \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.b ;
assign \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.s  = { \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.fas_s2 , \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.sum_s1  };
assign \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.u2.a  = \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.ain_s1 ;
assign \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.u2.b  = \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.bin_s1 ;
assign \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.u2.cin  = \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.carry_s1 ;
assign \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.facout_s2  = \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.u2.cout ;
assign \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.fas_s2  = \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.u2.s ;
assign \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.u1.a  = \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.a [1:0];
assign \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.u1.b  = \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.b [1:0];
assign \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.u1.cin  = 1'h0;
assign \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.facout_s1  = \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.u1.cout ;
assign \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.fas_s1  = \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.u1.s ;
assign \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.a  = \add_4ns_4ns_4_2_1_U8.din0 ;
assign \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.b  = \add_4ns_4ns_4_2_1_U8.din1 ;
assign \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.ce  = \add_4ns_4ns_4_2_1_U8.ce ;
assign \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.clk  = \add_4ns_4ns_4_2_1_U8.clk ;
assign \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.reset  = \add_4ns_4ns_4_2_1_U8.reset ;
assign \add_4ns_4ns_4_2_1_U8.dout  = \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_0_U.s ;
assign \add_4ns_4ns_4_2_1_U8.ce  = 1'h1;
assign \add_4ns_4ns_4_2_1_U8.clk  = ap_clk;
assign \add_4ns_4ns_4_2_1_U8.din0  = ret_V_7_reg_860;
assign \add_4ns_4ns_4_2_1_U8.din1  = 4'h1;
assign grp_fu_355_p2 = \add_4ns_4ns_4_2_1_U8.dout ;
assign \add_4ns_4ns_4_2_1_U8.reset  = ap_rst;
assign \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.ain_s0  = \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.a ;
assign \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.bin_s0  = \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.b ;
assign \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.s  = { \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.fas_s2 , \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.sum_s1  };
assign \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.u2.a  = \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.ain_s1 ;
assign \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.u2.b  = \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.bin_s1 ;
assign \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.u2.cin  = \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.carry_s1 ;
assign \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.facout_s2  = \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.u2.cout ;
assign \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.fas_s2  = \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.u2.s ;
assign \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.u1.a  = \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.a [1:0];
assign \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.u1.b  = \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.b [1:0];
assign \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.u1.cin  = 1'h0;
assign \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.facout_s1  = \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.u1.cout ;
assign \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.fas_s1  = \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.u1.s ;
assign \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.a  = \add_4ns_4ns_4_2_1_U1.din0 ;
assign \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.b  = \add_4ns_4ns_4_2_1_U1.din1 ;
assign \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.ce  = \add_4ns_4ns_4_2_1_U1.ce ;
assign \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.clk  = \add_4ns_4ns_4_2_1_U1.clk ;
assign \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.reset  = \add_4ns_4ns_4_2_1_U1.reset ;
assign \add_4ns_4ns_4_2_1_U1.dout  = \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.s ;
assign \add_4ns_4ns_4_2_1_U1.ce  = 1'h1;
assign \add_4ns_4ns_4_2_1_U1.clk  = ap_clk;
assign \add_4ns_4ns_4_2_1_U1.din0  = ret_V_reg_756;
assign \add_4ns_4ns_4_2_1_U1.din1  = 4'h1;
assign grp_fu_221_p2 = \add_4ns_4ns_4_2_1_U1.dout ;
assign \add_4ns_4ns_4_2_1_U1.reset  = ap_rst;
assign \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.ain_s0  = \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.a ;
assign \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.bin_s0  = \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.b ;
assign \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.s  = { \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.fas_s2 , \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.sum_s1  };
assign \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.u2.a  = \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.ain_s1 ;
assign \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.u2.b  = \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.bin_s1 ;
assign \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.u2.cin  = \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.carry_s1 ;
assign \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.facout_s2  = \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.u2.cout ;
assign \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.fas_s2  = \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.u2.s ;
assign \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.u1.a  = \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.a [17:0];
assign \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.u1.b  = \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.b [17:0];
assign \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.u1.cin  = 1'h0;
assign \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.facout_s1  = \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.u1.cout ;
assign \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.fas_s1  = \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.u1.s ;
assign \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.a  = \add_36ns_36s_36_2_1_U13.din0 ;
assign \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.b  = \add_36ns_36s_36_2_1_U13.din1 ;
assign \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.ce  = \add_36ns_36s_36_2_1_U13.ce ;
assign \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.clk  = \add_36ns_36s_36_2_1_U13.clk ;
assign \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.reset  = \add_36ns_36s_36_2_1_U13.reset ;
assign \add_36ns_36s_36_2_1_U13.dout  = \add_36ns_36s_36_2_1_U13.top_add_36ns_36s_36_2_1_Adder_8_U.s ;
assign \add_36ns_36s_36_2_1_U13.ce  = 1'h1;
assign \add_36ns_36s_36_2_1_U13.clk  = ap_clk;
assign \add_36ns_36s_36_2_1_U13.din0  = { select_ln353_1_reg_1010, 4'h0 };
assign \add_36ns_36s_36_2_1_U13.din1  = { ret_V_6_reg_1005[3], ret_V_6_reg_1005[3], ret_V_6_reg_1005[3], ret_V_6_reg_1005[3], ret_V_6_reg_1005[3], ret_V_6_reg_1005[3], ret_V_6_reg_1005[3], ret_V_6_reg_1005[3], ret_V_6_reg_1005[3], ret_V_6_reg_1005[3], ret_V_6_reg_1005[3], ret_V_6_reg_1005[3], ret_V_6_reg_1005[3], ret_V_6_reg_1005[3], ret_V_6_reg_1005[3], ret_V_6_reg_1005[3], ret_V_6_reg_1005[3], ret_V_6_reg_1005[3], ret_V_6_reg_1005[3], ret_V_6_reg_1005[3], ret_V_6_reg_1005[3], ret_V_6_reg_1005[3], ret_V_6_reg_1005[3], ret_V_6_reg_1005[3], ret_V_6_reg_1005[3], ret_V_6_reg_1005[3], ret_V_6_reg_1005[3], ret_V_6_reg_1005[3], ret_V_6_reg_1005, 4'h0 };
assign grp_fu_622_p2 = \add_36ns_36s_36_2_1_U13.dout ;
assign \add_36ns_36s_36_2_1_U13.reset  = ap_rst;
assign \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.ain_s0  = \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.a ;
assign \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.bin_s0  = \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.b ;
assign \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.s  = { \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.fas_s2 , \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.sum_s1  };
assign \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.u2.a  = \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.ain_s1 ;
assign \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.u2.b  = \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.bin_s1 ;
assign \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.u2.cin  = \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.carry_s1 ;
assign \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.facout_s2  = \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.u2.cout ;
assign \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.fas_s2  = \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.u2.s ;
assign \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.u1.a  = \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.a [17:0];
assign \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.u1.b  = \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.b [17:0];
assign \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.u1.cin  = 1'h0;
assign \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.facout_s1  = \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.u1.cout ;
assign \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.fas_s1  = \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.u1.s ;
assign \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.a  = \add_36ns_36ns_36_2_1_U17.din0 ;
assign \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.b  = \add_36ns_36ns_36_2_1_U17.din1 ;
assign \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.ce  = \add_36ns_36ns_36_2_1_U17.ce ;
assign \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.clk  = \add_36ns_36ns_36_2_1_U17.clk ;
assign \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.reset  = \add_36ns_36ns_36_2_1_U17.reset ;
assign \add_36ns_36ns_36_2_1_U17.dout  = \add_36ns_36ns_36_2_1_U17.top_add_36ns_36ns_36_2_1_Adder_11_U.s ;
assign \add_36ns_36ns_36_2_1_U17.ce  = 1'h1;
assign \add_36ns_36ns_36_2_1_U17.clk  = ap_clk;
assign \add_36ns_36ns_36_2_1_U17.din0  = { op_25_V_reg_1055, 4'h0 };
assign \add_36ns_36ns_36_2_1_U17.din1  = { 31'h00000000, tmp_V_reg_1050, 4'h0 };
assign grp_fu_698_p2 = \add_36ns_36ns_36_2_1_U17.dout ;
assign \add_36ns_36ns_36_2_1_U17.reset  = ap_rst;
assign \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.ain_s0  = \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.a ;
assign \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.bin_s0  = \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.b ;
assign \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.s  = { \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.fas_s2 , \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.sum_s1  };
assign \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.u2.a  = \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.ain_s1 ;
assign \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.u2.b  = \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.bin_s1 ;
assign \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.u2.cin  = \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.carry_s1 ;
assign \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.facout_s2  = \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.u2.cout ;
assign \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.fas_s2  = \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.u2.s ;
assign \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.u1.a  = \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.a [16:0];
assign \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.u1.b  = \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.b [16:0];
assign \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.u1.cin  = 1'h0;
assign \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.facout_s1  = \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.u1.cout ;
assign \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.fas_s1  = \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.u1.s ;
assign \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.a  = \add_34s_34s_34_2_1_U11.din0 ;
assign \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.b  = \add_34s_34s_34_2_1_U11.din1 ;
assign \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.ce  = \add_34s_34s_34_2_1_U11.ce ;
assign \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.clk  = \add_34s_34s_34_2_1_U11.clk ;
assign \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.reset  = \add_34s_34s_34_2_1_U11.reset ;
assign \add_34s_34s_34_2_1_U11.dout  = \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_6_U.s ;
assign \add_34s_34s_34_2_1_U11.ce  = 1'h1;
assign \add_34s_34s_34_2_1_U11.clk  = ap_clk;
assign \add_34s_34s_34_2_1_U11.din0  = { select_ln353_reg_968[5], select_ln353_reg_968[5], select_ln353_reg_968[5], select_ln353_reg_968[5], select_ln353_reg_968[5], select_ln353_reg_968[5], select_ln353_reg_968[5], select_ln353_reg_968[5], select_ln353_reg_968[5], select_ln353_reg_968[5], select_ln353_reg_968[5], select_ln353_reg_968[5], select_ln353_reg_968[5], select_ln353_reg_968[5], select_ln353_reg_968[5], select_ln353_reg_968[5], select_ln353_reg_968[5], select_ln353_reg_968[5], select_ln353_reg_968[5], select_ln353_reg_968[5], select_ln353_reg_968[5], select_ln353_reg_968[5], select_ln353_reg_968[5], select_ln353_reg_968[5], select_ln353_reg_968[5], select_ln353_reg_968[5], select_ln353_reg_968[5], select_ln353_reg_968, 1'h0 };
assign \add_34s_34s_34_2_1_U11.din1  = { op_12_V_reg_962[1], op_12_V_reg_962[1], op_12_V_reg_962[1], op_12_V_reg_962[1], op_12_V_reg_962[1], op_12_V_reg_962[1], op_12_V_reg_962[1], op_12_V_reg_962[1], op_12_V_reg_962[1], op_12_V_reg_962[1], op_12_V_reg_962[1], op_12_V_reg_962[1], op_12_V_reg_962[1], op_12_V_reg_962[1], op_12_V_reg_962[1], op_12_V_reg_962[1], op_12_V_reg_962[1], op_12_V_reg_962[1], op_12_V_reg_962[1], op_12_V_reg_962[1], op_12_V_reg_962[1], op_12_V_reg_962[1], op_12_V_reg_962[1], op_12_V_reg_962[1], op_12_V_reg_962[1], op_12_V_reg_962[1], op_12_V_reg_962[1], op_12_V_reg_962[1], op_12_V_reg_962[1], op_12_V_reg_962[1], op_12_V_reg_962[1], op_12_V_reg_962[1], op_12_V_reg_962 };
assign grp_fu_547_p2 = \add_34s_34s_34_2_1_U11.dout ;
assign \add_34s_34s_34_2_1_U11.reset  = ap_rst;
assign \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.ain_s0  = \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.a ;
assign \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.bin_s0  = \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.b ;
assign \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.s  = { \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.fas_s2 , \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.sum_s1  };
assign \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.u2.a  = \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.ain_s1 ;
assign \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.u2.b  = \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.bin_s1 ;
assign \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.u2.cin  = \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.carry_s1 ;
assign \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.facout_s2  = \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.u2.cout ;
assign \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.fas_s2  = \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.u2.s ;
assign \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.u1.a  = \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.a [15:0];
assign \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.u1.b  = \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.b [15:0];
assign \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.u1.cin  = 1'h0;
assign \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.facout_s1  = \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.u1.cout ;
assign \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.fas_s1  = \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.u1.s ;
assign \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.a  = \add_32s_32ns_32_2_1_U20.din0 ;
assign \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.b  = \add_32s_32ns_32_2_1_U20.din1 ;
assign \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.ce  = \add_32s_32ns_32_2_1_U20.ce ;
assign \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.clk  = \add_32s_32ns_32_2_1_U20.clk ;
assign \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.reset  = \add_32s_32ns_32_2_1_U20.reset ;
assign \add_32s_32ns_32_2_1_U20.dout  = \add_32s_32ns_32_2_1_U20.top_add_32s_32ns_32_2_1_Adder_14_U.s ;
assign \add_32s_32ns_32_2_1_U20.ce  = 1'h1;
assign \add_32s_32ns_32_2_1_U20.clk  = ap_clk;
assign \add_32s_32ns_32_2_1_U20.din0  = { add_ln69_3_reg_1105[3], add_ln69_3_reg_1105[3], add_ln69_3_reg_1105[3], add_ln69_3_reg_1105[3], add_ln69_3_reg_1105[3], add_ln69_3_reg_1105[3], add_ln69_3_reg_1105[3], add_ln69_3_reg_1105[3], add_ln69_3_reg_1105[3], add_ln69_3_reg_1105[3], add_ln69_3_reg_1105[3], add_ln69_3_reg_1105[3], add_ln69_3_reg_1105[3], add_ln69_3_reg_1105[3], add_ln69_3_reg_1105[3], add_ln69_3_reg_1105[3], add_ln69_3_reg_1105[3], add_ln69_3_reg_1105[3], add_ln69_3_reg_1105[3], add_ln69_3_reg_1105[3], add_ln69_3_reg_1105[3], add_ln69_3_reg_1105[3], add_ln69_3_reg_1105[3], add_ln69_3_reg_1105[3], add_ln69_3_reg_1105[3], add_ln69_3_reg_1105[3], add_ln69_3_reg_1105[3], add_ln69_3_reg_1105[3], add_ln69_3_reg_1105 };
assign \add_32s_32ns_32_2_1_U20.din1  = add_ln69_2_reg_1100;
assign grp_fu_739_p2 = \add_32s_32ns_32_2_1_U20.dout ;
assign \add_32s_32ns_32_2_1_U20.reset  = ap_rst;
assign \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.ain_s0  = \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.a ;
assign \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.bin_s0  = \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.b ;
assign \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.s  = { \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.fas_s2 , \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.sum_s1  };
assign \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.u2.a  = \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.ain_s1 ;
assign \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.u2.b  = \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.bin_s1 ;
assign \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.u2.cin  = \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.carry_s1 ;
assign \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.facout_s2  = \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.u2.cout ;
assign \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.fas_s2  = \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.u2.s ;
assign \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.u1.a  = \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.a [15:0];
assign \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.u1.b  = \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.b [15:0];
assign \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.u1.cin  = 1'h0;
assign \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.facout_s1  = \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.u1.cout ;
assign \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.fas_s1  = \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.u1.s ;
assign \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.a  = \add_32ns_32s_32_2_1_U18.din0 ;
assign \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.b  = \add_32ns_32s_32_2_1_U18.din1 ;
assign \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.ce  = \add_32ns_32s_32_2_1_U18.ce ;
assign \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.clk  = \add_32ns_32s_32_2_1_U18.clk ;
assign \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.reset  = \add_32ns_32s_32_2_1_U18.reset ;
assign \add_32ns_32s_32_2_1_U18.dout  = \add_32ns_32s_32_2_1_U18.top_add_32ns_32s_32_2_1_Adder_12_U.s ;
assign \add_32ns_32s_32_2_1_U18.ce  = 1'h1;
assign \add_32ns_32s_32_2_1_U18.clk  = ap_clk;
assign \add_32ns_32s_32_2_1_U18.din0  = op_26_V_reg_1080;
assign \add_32ns_32s_32_2_1_U18.din1  = { op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19 };
assign grp_fu_725_p2 = \add_32ns_32s_32_2_1_U18.dout ;
assign \add_32ns_32s_32_2_1_U18.reset  = ap_rst;
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s0  = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.a ;
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s0  = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.b ;
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.s  = { \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s2 , \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.sum_s1  };
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.a  = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s1 ;
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.b  = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s1 ;
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cin  = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.carry_s1 ;
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.facout_s2  = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cout ;
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s2  = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.s ;
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.a  = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.a [15:0];
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.b  = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.b [15:0];
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cin  = 1'h0;
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.facout_s1  = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cout ;
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s1  = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.s ;
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.a  = \add_32ns_32ns_32_2_1_U15.din0 ;
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.b  = \add_32ns_32ns_32_2_1_U15.din1 ;
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.ce  = \add_32ns_32ns_32_2_1_U15.ce ;
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.clk  = \add_32ns_32ns_32_2_1_U15.clk ;
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.reset  = \add_32ns_32ns_32_2_1_U15.reset ;
assign \add_32ns_32ns_32_2_1_U15.dout  = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_7_U.s ;
assign \add_32ns_32ns_32_2_1_U15.ce  = 1'h1;
assign \add_32ns_32ns_32_2_1_U15.clk  = ap_clk;
assign \add_32ns_32ns_32_2_1_U15.din0  = { 15'h0000, add_ln69_reg_1040 };
assign \add_32ns_32ns_32_2_1_U15.din1  = op_23_V_reg_1035;
assign grp_fu_661_p2 = \add_32ns_32ns_32_2_1_U15.dout ;
assign \add_32ns_32ns_32_2_1_U15.reset  = ap_rst;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s0  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.a ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s0  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.b ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.s  = { \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s2 , \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.sum_s1  };
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.a  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s1 ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.b  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s1 ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cin  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.carry_s1 ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.facout_s2  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cout ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s2  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.s ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.a  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.a [15:0];
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.b  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.b [15:0];
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cin  = 1'h0;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.facout_s1  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cout ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s1  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.s ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.a  = \add_32ns_32ns_32_2_1_U12.din0 ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.b  = \add_32ns_32ns_32_2_1_U12.din1 ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.ce  = \add_32ns_32ns_32_2_1_U12.ce ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.clk  = \add_32ns_32ns_32_2_1_U12.clk ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.reset  = \add_32ns_32ns_32_2_1_U12.reset ;
assign \add_32ns_32ns_32_2_1_U12.dout  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.s ;
assign \add_32ns_32ns_32_2_1_U12.ce  = 1'h1;
assign \add_32ns_32ns_32_2_1_U12.clk  = ap_clk;
assign \add_32ns_32ns_32_2_1_U12.din0  = ret_V_21_cast_reg_988;
assign \add_32ns_32ns_32_2_1_U12.din1  = 32'd1;
assign grp_fu_563_p2 = \add_32ns_32ns_32_2_1_U12.dout ;
assign \add_32ns_32ns_32_2_1_U12.reset  = ap_rst;
assign \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.ain_s0  = \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.a ;
assign \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.bin_s0  = \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.b ;
assign \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.s  = { \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.fas_s2 , \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.sum_s1  };
assign \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.u2.a  = \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.ain_s1 ;
assign \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.u2.b  = \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.bin_s1 ;
assign \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.u2.cin  = \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.carry_s1 ;
assign \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.facout_s2  = \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.u2.cout ;
assign \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.fas_s2  = \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.u2.s ;
assign \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.u1.a  = \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.a [7:0];
assign \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.u1.b  = \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.b [7:0];
assign \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.u1.cin  = 1'h0;
assign \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.facout_s1  = \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.u1.cout ;
assign \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.fas_s1  = \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.u1.s ;
assign \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.a  = \add_17ns_17s_17_2_1_U7.din0 ;
assign \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.b  = \add_17ns_17s_17_2_1_U7.din1 ;
assign \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.ce  = \add_17ns_17s_17_2_1_U7.ce ;
assign \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.clk  = \add_17ns_17s_17_2_1_U7.clk ;
assign \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.reset  = \add_17ns_17s_17_2_1_U7.reset ;
assign \add_17ns_17s_17_2_1_U7.dout  = \add_17ns_17s_17_2_1_U7.top_add_17ns_17s_17_2_1_Adder_3_U.s ;
assign \add_17ns_17s_17_2_1_U7.ce  = 1'h1;
assign \add_17ns_17s_17_2_1_U7.clk  = ap_clk;
assign \add_17ns_17s_17_2_1_U7.din0  = { 3'h0, signbit_reg_835, 13'h0000 };
assign \add_17ns_17s_17_2_1_U7.din1  = { op_7[15], op_7 };
assign grp_fu_330_p2 = \add_17ns_17s_17_2_1_U7.dout ;
assign \add_17ns_17s_17_2_1_U7.reset  = ap_rst;
assign \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.ain_s0  = \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.a ;
assign \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.bin_s0  = \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.b ;
assign \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.s  = { \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.fas_s2 , \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.sum_s1  };
assign \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.u2.a  = \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.ain_s1 ;
assign \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.u2.b  = \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.bin_s1 ;
assign \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.u2.cin  = \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.carry_s1 ;
assign \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.facout_s2  = \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.u2.cout ;
assign \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.fas_s2  = \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.u2.s ;
assign \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.u1.a  = \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.a [7:0];
assign \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.u1.b  = \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.b [7:0];
assign \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.u1.cin  = 1'h0;
assign \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.facout_s1  = \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.u1.cout ;
assign \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.fas_s1  = \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.u1.s ;
assign \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.a  = \add_17ns_17ns_17_2_1_U14.din0 ;
assign \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.b  = \add_17ns_17ns_17_2_1_U14.din1 ;
assign \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.ce  = \add_17ns_17ns_17_2_1_U14.ce ;
assign \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.clk  = \add_17ns_17ns_17_2_1_U14.clk ;
assign \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.reset  = \add_17ns_17ns_17_2_1_U14.reset ;
assign \add_17ns_17ns_17_2_1_U14.dout  = \add_17ns_17ns_17_2_1_U14.top_add_17ns_17ns_17_2_1_Adder_9_U.s ;
assign \add_17ns_17ns_17_2_1_U14.ce  = 1'h1;
assign \add_17ns_17ns_17_2_1_U14.clk  = ap_clk;
assign \add_17ns_17ns_17_2_1_U14.din0  = { 1'h0, ret_V_15_reg_1000[3], ret_V_15_reg_1000[3], ret_V_15_reg_1000[3], ret_V_15_reg_1000[3], ret_V_15_reg_1000[3], ret_V_15_reg_1000[3], ret_V_15_reg_1000[3], ret_V_15_reg_1000[3], ret_V_15_reg_1000[3], ret_V_15_reg_1000[3], ret_V_15_reg_1000[3], ret_V_15_reg_1000[3], ret_V_15_reg_1000 };
assign \add_17ns_17ns_17_2_1_U14.din1  = { 9'h000, ret_V_16_reg_840[4], ret_V_16_reg_840[4], ret_V_16_reg_840[4], ret_V_16_reg_840 };
assign grp_fu_642_p2 = \add_17ns_17ns_17_2_1_U14.dout ;
assign \add_17ns_17ns_17_2_1_U14.reset  = ap_rst;
endmodule


// Product machine:
module top_A_times_top_B (ap_start, op_0, op_1, op_10, op_11, op_18, op_19, op_4, op_5, op_6, op_7, ap_clk, unsafe_signal);
input ap_start;
input [3:0] op_0;
input [3:0] op_1;
input [3:0] op_10;
input [3:0] op_11;
input [1:0] op_18;
input [3:0] op_19;
input [1:0] op_4;
input [3:0] op_5;
input [3:0] op_6;
input [15:0] op_7;
input ap_clk;
output unsafe_signal;
reg _setup;
initial _setup = 1'b0;
always @ (posedge ap_clk) _setup <= 1'b1;
reg ap_start_internal;
always @ (posedge ap_clk) if (!_setup) ap_start_internal <= ap_start;
reg [3:0] op_0_internal;
always @ (posedge ap_clk) if (!_setup) op_0_internal <= op_0;
reg [3:0] op_1_internal;
always @ (posedge ap_clk) if (!_setup) op_1_internal <= op_1;
reg [3:0] op_10_internal;
always @ (posedge ap_clk) if (!_setup) op_10_internal <= op_10;
reg [3:0] op_11_internal;
always @ (posedge ap_clk) if (!_setup) op_11_internal <= op_11;
reg [1:0] op_18_internal;
always @ (posedge ap_clk) if (!_setup) op_18_internal <= op_18;
reg [3:0] op_19_internal;
always @ (posedge ap_clk) if (!_setup) op_19_internal <= op_19;
reg [1:0] op_4_internal;
always @ (posedge ap_clk) if (!_setup) op_4_internal <= op_4;
reg [3:0] op_5_internal;
always @ (posedge ap_clk) if (!_setup) op_5_internal <= op_5;
reg [3:0] op_6_internal;
always @ (posedge ap_clk) if (!_setup) op_6_internal <= op_6;
reg [15:0] op_7_internal;
always @ (posedge ap_clk) if (!_setup) op_7_internal <= op_7;
wire ap_done_A;
wire ap_done_B;
wire ap_done_eq;
assign ap_done_eq = ap_done_A == ap_done_B;
wire ap_idle_A;
wire ap_idle_B;
wire ap_idle_eq;
assign ap_idle_eq = ap_idle_A == ap_idle_B;
wire ap_ready_A;
wire ap_ready_B;
wire ap_ready_eq;
assign ap_ready_eq = ap_ready_A == ap_ready_B;
wire [31:0] op_29_A;
wire [31:0] op_29_B;
wire op_29_eq;
assign op_29_eq = op_29_A == op_29_B;
wire op_29_ap_vld_A;
wire op_29_ap_vld_B;
wire clk_enable_A;
wire clk_enable_B;
assign clk_enable_A = _setup & (~op_29_ap_vld_A | op_29_ap_vld_B);
assign clk_enable_B = _setup;
wire divergent;
assign divergent = ~(ap_done_eq & ap_idle_eq & ap_ready_eq & op_29_eq);
assign unsafe_signal = op_29_ap_vld_A & op_29_ap_vld_B & divergent;
top_A instance_A (
    .ap_clk(ap_clk),
    .clk_enable(clk_enable_A),
    .ap_start(ap_start_internal),
    .op_0(op_0_internal),
    .op_1(op_1_internal),
    .op_10(op_10_internal),
    .op_11(op_11_internal),
    .op_18(op_18_internal),
    .op_19(op_19_internal),
    .op_4(op_4_internal),
    .op_5(op_5_internal),
    .op_6(op_6_internal),
    .op_7(op_7_internal),
    .ap_done(ap_done_A),
    .ap_idle(ap_idle_A),
    .ap_ready(ap_ready_A),
    .op_29(op_29_A),
    .op_29_ap_vld(op_29_ap_vld_A)
);
top_B instance_B (
    .ap_clk(ap_clk),
    .clk_enable(clk_enable_B),
    .ap_start(ap_start_internal),
    .op_0(op_0_internal),
    .op_1(op_1_internal),
    .op_10(op_10_internal),
    .op_11(op_11_internal),
    .op_18(op_18_internal),
    .op_19(op_19_internal),
    .op_4(op_4_internal),
    .op_5(op_5_internal),
    .op_6(op_6_internal),
    .op_7(op_7_internal),
    .ap_done(ap_done_B),
    .ap_idle(ap_idle_B),
    .ap_ready(ap_ready_B),
    .op_29(op_29_B),
    .op_29_ap_vld(op_29_ap_vld_B)
);
endmodule
