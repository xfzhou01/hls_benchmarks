// Processed by function `construct_kairos` in `verilog_tricks.py`.
// Machine A:
// Processed by function `add_clk_enable_signal` in `verilog_tricks.py`.
// Processed by function `remove_reset_signal` in `verilog_tricks.py`.
module top_A (
  ap_clk,
  ap_start,
  ap_done,
  ap_idle,
  ap_ready,
  op_0,
  op_1,
  op_2,
  op_3,
  op_4,
  op_5,
  op_10,
  op_12,
  op_13,
  op_14,
  op_18,
  op_19,
  op_32,
  op_32_ap_vld,
clk_enable
);
input clk_enable;


input ap_clk;
wire ap_rst;
assign ap_rst = op_32_ap_vld;
input ap_start;
input [7:0] op_0;
input [3:0] op_1;
input [31:0] op_10;
input [1:0] op_12;
input op_13;
input [31:0] op_14;
input op_18;
input [3:0] op_19;
input [3:0] op_2;
input [1:0] op_3;
input [15:0] op_4;
input [1:0] op_5;
output ap_done;
output ap_idle;
output ap_ready;
output [31:0] op_32;
output op_32_ap_vld;


reg [2:0] add_ln69_1_reg_522;
reg [8:0] add_ln69_2_reg_527;
reg [31:0] add_ln69_4_reg_584;
reg [1:0] add_ln69_7_reg_579;
reg [2:0] add_ln69_8_reg_589;
reg [9:0] ap_CS_fsm = 10'h001;
reg icmp_ln851_reg_611;
reg icmp_ln890_reg_517;
reg [24:0] \mac_muladd_4ns_4s_32ns_32_4_1_U2.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.a_reg ;
reg [17:0] \mac_muladd_4ns_4s_32ns_32_4_1_U2.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.b_reg ;
reg [42:0] \mac_muladd_4ns_4s_32ns_32_4_1_U2.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.m_reg ;
reg [47:0] \mac_muladd_4ns_4s_32ns_32_4_1_U2.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.p_reg ;
reg [1:0] op_16_V_reg_552;
reg [31:0] op_24_V_reg_532;
reg [31:0] op_31_V_reg_594;
reg [3:0] r_reg_507;
reg [31:0] ret_V_3_cast_reg_604;
reg [33:0] ret_V_4_reg_557;
reg [31:0] ret_V_5_reg_569;
reg [35:0] ret_V_6_reg_599;
reg [31:0] ret_V_cast_reg_562;
reg [2:0] select_ln69_reg_574;
reg [1:0] zext_ln11_reg_512;
wire [2:0] _000_;
wire [8:0] _001_;
wire [31:0] _002_;
wire [1:0] _003_;
wire [2:0] _004_;
wire [9:0] _005_;
wire _006_;
wire _007_;
wire [1:0] _008_;
wire [31:0] _009_;
wire [31:0] _010_;
wire [3:0] _011_;
wire [31:0] _012_;
wire [33:0] _013_;
wire [31:0] _014_;
wire [35:0] _015_;
wire [31:0] _016_;
wire [2:0] _017_;
wire _018_;
wire [1:0] _019_;
wire _020_;
wire _021_;
wire _022_;
wire [24:0] _023_;
wire [17:0] _024_;
wire [42:0] _025_;
wire [47:0] _026_;
wire _027_;
wire _028_;
wire _029_;
wire _030_;
wire _031_;
wire _032_;
wire _033_;
wire _034_;
wire _035_;
wire _036_;
wire _037_;
wire _038_;
wire _039_;
wire [31:0] add_ln691_1_fu_476_p2;
wire [31:0] add_ln691_fu_347_p2;
wire [2:0] add_ln69_1_fu_233_p2;
wire [8:0] add_ln69_2_fu_256_p2;
wire [31:0] add_ln69_5_fu_414_p2;
wire [2:0] add_ln69_6_fu_400_p2;
wire [1:0] add_ln69_7_fu_391_p2;
wire [2:0] add_ln69_8_fu_408_p2;
wire [31:0] add_ln69_fu_266_p2;
wire ap_CS_fsm_state1;
wire ap_CS_fsm_state10;
wire ap_CS_fsm_state2;
wire ap_CS_fsm_state3;
wire ap_CS_fsm_state4;
wire ap_CS_fsm_state5;
wire ap_CS_fsm_state6;
wire ap_CS_fsm_state7;
wire ap_CS_fsm_state8;
wire ap_CS_fsm_state9;
wire [9:0] ap_NS_fsm;
wire ap_clk;
wire ap_done;
wire ap_idle;
wire ap_ready;
wire ap_rst;
wire ap_start;
wire [3:0] grp_fu_495_p0;
wire [7:0] grp_fu_495_p00;
wire [31:0] grp_fu_495_p3;
wire icmp_ln851_fu_463_p2;
wire icmp_ln890_fu_213_p2;
wire lhs_V_fu_189_p2;
wire \mac_muladd_4ns_4s_32ns_32_4_1_U2.ce ;
wire \mac_muladd_4ns_4s_32ns_32_4_1_U2.clk ;
wire [3:0] \mac_muladd_4ns_4s_32ns_32_4_1_U2.din0 ;
wire [3:0] \mac_muladd_4ns_4s_32ns_32_4_1_U2.din1 ;
wire [31:0] \mac_muladd_4ns_4s_32ns_32_4_1_U2.din2 ;
wire [31:0] \mac_muladd_4ns_4s_32ns_32_4_1_U2.dout ;
wire \mac_muladd_4ns_4s_32ns_32_4_1_U2.reset ;
wire [24:0] \mac_muladd_4ns_4s_32ns_32_4_1_U2.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.a ;
wire [17:0] \mac_muladd_4ns_4s_32ns_32_4_1_U2.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.b ;
wire [47:0] \mac_muladd_4ns_4s_32ns_32_4_1_U2.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.c ;
wire \mac_muladd_4ns_4s_32ns_32_4_1_U2.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.ce ;
wire \mac_muladd_4ns_4s_32ns_32_4_1_U2.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.clk ;
wire [31:0] \mac_muladd_4ns_4s_32ns_32_4_1_U2.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.dout ;
wire [3:0] \mac_muladd_4ns_4s_32ns_32_4_1_U2.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.in0 ;
wire [3:0] \mac_muladd_4ns_4s_32ns_32_4_1_U2.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.in1 ;
wire [31:0] \mac_muladd_4ns_4s_32ns_32_4_1_U2.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.in2 ;
wire [42:0] \mac_muladd_4ns_4s_32ns_32_4_1_U2.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.m ;
wire [47:0] \mac_muladd_4ns_4s_32ns_32_4_1_U2.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.p ;
wire \mac_muladd_4ns_4s_32ns_32_4_1_U2.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.rst ;
wire [1:0] \mul_2ns_2ns_4_1_1_U1.din0 ;
wire [1:0] \mul_2ns_2ns_4_1_1_U1.din1 ;
wire [3:0] \mul_2ns_2ns_4_1_1_U1.dout ;
wire [1:0] \mul_2ns_2ns_4_1_1_U1.top_mul_2ns_2ns_4_1_1_Multiplier_0_U.a ;
wire [1:0] \mul_2ns_2ns_4_1_1_U1.top_mul_2ns_2ns_4_1_1_Multiplier_0_U.b ;
wire [3:0] \mul_2ns_2ns_4_1_1_U1.top_mul_2ns_2ns_4_1_1_Multiplier_0_U.p ;
wire [7:0] op_0;
wire [3:0] op_1;
wire [31:0] op_10;
wire [1:0] op_12;
wire op_13;
wire [31:0] op_14;
wire [1:0] op_16_V_fu_301_p2;
wire op_18;
wire [3:0] op_19;
wire [3:0] op_2;
wire [31:0] op_24_V_fu_275_p2;
wire [1:0] op_3;
wire [31:0] op_31_V_fu_422_p2;
wire [31:0] op_32;
wire op_32_ap_vld;
wire [15:0] op_4;
wire [1:0] op_5;
wire op_9_V_fu_207_p2;
wire p_Result_1_fu_469_p3;
wire p_Result_s_fu_337_p3;
wire [1:0] r_1_fu_219_p2;
wire [3:0] r_fu_171_p2;
wire [1:0] ret_1_fu_284_p0;
wire [1:0] ret_1_fu_284_p1;
wire [3:0] ret_1_fu_284_p2;
wire [33:0] ret_V_4_fu_321_p2;
wire [31:0] ret_V_5_fu_359_p3;
wire [35:0] ret_V_6_fu_443_p2;
wire [8:0] ret_fu_247_p2;
wire [32:0] rhs_1_fu_310_p3;
wire [34:0] rhs_3_fu_432_p3;
wire [1:0] select_ln69_1_fu_383_p3;
wire [2:0] select_ln69_fu_371_p3;
wire [31:0] select_ln850_1_fu_481_p3;
wire [31:0] select_ln850_fu_352_p3;
wire [35:0] sext_ln1192_1_fu_439_p1;
wire [33:0] sext_ln1192_fu_317_p1;
wire [8:0] sext_ln215_1_fu_243_p1;
wire [8:0] sext_ln215_fu_239_p1;
wire [31:0] sext_ln69_1_fu_272_p1;
wire [2:0] sext_ln69_2_fu_397_p1;
wire [2:0] sext_ln69_4_fu_405_p1;
wire [31:0] sext_ln69_5_fu_419_p1;
wire [3:0] sext_ln703_1_fu_428_p0;
wire [35:0] sext_ln703_1_fu_428_p1;
wire [1:0] sext_ln703_fu_306_p0;
wire [33:0] sext_ln703_fu_306_p1;
wire [1:0] sext_ln874_1_fu_185_p0;
wire [2:0] sext_ln874_1_fu_185_p1;
wire [1:0] sext_ln874_fu_181_p0;
wire [3:0] sext_ln874_fu_181_p1;
wire [1:0] trunc_ln1350_fu_297_p1;
wire [1:0] trunc_ln213_1_fu_203_p0;
wire trunc_ln213_1_fu_203_p1;
wire trunc_ln213_fu_199_p1;
wire [3:0] trunc_ln851_1_fu_459_p0;
wire [2:0] trunc_ln851_1_fu_459_p1;
wire [1:0] trunc_ln851_fu_344_p0;
wire trunc_ln851_fu_344_p1;
wire xor_ln890_fu_366_p2;
wire [1:0] zext_ln11_fu_195_p1;
wire [3:0] zext_ln1345_fu_281_p1;
wire [2:0] zext_ln69_2_fu_225_p1;
wire [2:0] zext_ln69_3_fu_229_p1;
wire [8:0] zext_ln69_4_fu_253_p1;
wire [1:0] zext_ln69_5_fu_379_p1;
wire [31:0] zext_ln69_fu_262_p1;
wire [2:0] zext_ln874_fu_177_p1;


assign add_ln691_1_fu_476_p2 = ret_V_3_cast_reg_604 + 1'h1;
assign add_ln691_fu_347_p2 = ret_V_cast_reg_562 + 1'h1;
assign add_ln69_1_fu_233_p2 = r_1_fu_219_p2 + op_9_V_fu_207_p2;
assign add_ln69_2_fu_256_p2 = add_ln69_1_reg_522 + ret_fu_247_p2;
assign add_ln69_5_fu_414_p2 = $signed(add_ln69_4_reg_584) + $signed(op_14);
assign add_ln69_6_fu_400_p2 = $signed(op_16_V_reg_552) + $signed(select_ln69_reg_574);
assign add_ln69_7_fu_391_p2 = select_ln69_1_fu_383_p3 + xor_ln890_fu_366_p2;
assign add_ln69_8_fu_408_p2 = $signed(add_ln69_7_reg_579) + $signed(add_ln69_6_fu_400_p2);
assign add_ln69_fu_266_p2 = op_4 + op_10;
assign op_24_V_fu_275_p2 = $signed(add_ln69_2_reg_527) + $signed(add_ln69_fu_266_p2);
assign op_31_V_fu_422_p2 = $signed(add_ln69_8_reg_589) + $signed(add_ln69_5_fu_414_p2);
assign ret_V_4_fu_321_p2 = $signed({ op_24_V_reg_532, 1'h0 }) + $signed(op_12);
assign ret_V_6_fu_443_p2 = $signed({ op_31_V_reg_594, 3'h0 }) + $signed(op_19);
assign ret_fu_247_p2 = $signed(op_0) + $signed(op_1);
assign _020_ = ap_CS_fsm[0] & _022_;
assign _021_ = ap_CS_fsm[0] & ap_start;
assign xor_ln890_fu_366_p2 = ~ icmp_ln890_reg_517;
assign r_fu_171_p2 = ~ op_2;
assign _022_ = ~ ap_start;
assign { \mac_muladd_4ns_4s_32ns_32_4_1_U2.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.p [47], \mac_muladd_4ns_4s_32ns_32_4_1_U2.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.p [42:0] } = $signed(\mac_muladd_4ns_4s_32ns_32_4_1_U2.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.m_reg ) + $signed({ 1'h0, \mac_muladd_4ns_4s_32ns_32_4_1_U2.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.in2  });
assign \mac_muladd_4ns_4s_32ns_32_4_1_U2.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.m  = $signed(\mac_muladd_4ns_4s_32ns_32_4_1_U2.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.a_reg ) * $signed(\mac_muladd_4ns_4s_32ns_32_4_1_U2.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.b_reg );
always @(posedge \mac_muladd_4ns_4s_32ns_32_4_1_U2.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.clk )
\mac_muladd_4ns_4s_32ns_32_4_1_U2.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.m_reg  <= _025_;
always @(posedge \mac_muladd_4ns_4s_32ns_32_4_1_U2.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.clk )
\mac_muladd_4ns_4s_32ns_32_4_1_U2.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.a_reg  <= _023_;
always @(posedge \mac_muladd_4ns_4s_32ns_32_4_1_U2.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.clk )
\mac_muladd_4ns_4s_32ns_32_4_1_U2.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.b_reg  <= _024_;
always @(posedge \mac_muladd_4ns_4s_32ns_32_4_1_U2.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.clk )
\mac_muladd_4ns_4s_32ns_32_4_1_U2.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.p_reg  <= _026_;
assign _026_ = \mac_muladd_4ns_4s_32ns_32_4_1_U2.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.ce  ? { \mac_muladd_4ns_4s_32ns_32_4_1_U2.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.p [47], \mac_muladd_4ns_4s_32ns_32_4_1_U2.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.p [47], \mac_muladd_4ns_4s_32ns_32_4_1_U2.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.p [47], \mac_muladd_4ns_4s_32ns_32_4_1_U2.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.p [47], \mac_muladd_4ns_4s_32ns_32_4_1_U2.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.p [47], \mac_muladd_4ns_4s_32ns_32_4_1_U2.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.p [42:0] } : \mac_muladd_4ns_4s_32ns_32_4_1_U2.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.p_reg ;
assign _024_ = \mac_muladd_4ns_4s_32ns_32_4_1_U2.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.ce  ? { \mac_muladd_4ns_4s_32ns_32_4_1_U2.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.in1 [3], \mac_muladd_4ns_4s_32ns_32_4_1_U2.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.in1 [3], \mac_muladd_4ns_4s_32ns_32_4_1_U2.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.in1 [3], \mac_muladd_4ns_4s_32ns_32_4_1_U2.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.in1 [3], \mac_muladd_4ns_4s_32ns_32_4_1_U2.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.in1 [3], \mac_muladd_4ns_4s_32ns_32_4_1_U2.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.in1 [3], \mac_muladd_4ns_4s_32ns_32_4_1_U2.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.in1 [3], \mac_muladd_4ns_4s_32ns_32_4_1_U2.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.in1 [3], \mac_muladd_4ns_4s_32ns_32_4_1_U2.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.in1 [3], \mac_muladd_4ns_4s_32ns_32_4_1_U2.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.in1 [3], \mac_muladd_4ns_4s_32ns_32_4_1_U2.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.in1 [3], \mac_muladd_4ns_4s_32ns_32_4_1_U2.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.in1 [3], \mac_muladd_4ns_4s_32ns_32_4_1_U2.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.in1 [3], \mac_muladd_4ns_4s_32ns_32_4_1_U2.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.in1 [3], \mac_muladd_4ns_4s_32ns_32_4_1_U2.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.in1  } : \mac_muladd_4ns_4s_32ns_32_4_1_U2.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.b_reg ;
assign _023_ = \mac_muladd_4ns_4s_32ns_32_4_1_U2.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.ce  ? { 21'h000000, \mac_muladd_4ns_4s_32ns_32_4_1_U2.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.in0  } : \mac_muladd_4ns_4s_32ns_32_4_1_U2.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.a_reg ;
assign _025_ = \mac_muladd_4ns_4s_32ns_32_4_1_U2.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.ce  ? \mac_muladd_4ns_4s_32ns_32_4_1_U2.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.m  : \mac_muladd_4ns_4s_32ns_32_4_1_U2.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.m_reg ;
assign \mul_2ns_2ns_4_1_1_U1.top_mul_2ns_2ns_4_1_1_Multiplier_0_U.p  = \mul_2ns_2ns_4_1_1_U1.top_mul_2ns_2ns_4_1_1_Multiplier_0_U.a  * \mul_2ns_2ns_4_1_1_U1.top_mul_2ns_2ns_4_1_1_Multiplier_0_U.b ;
assign _027_ = $signed(r_fu_171_p2) < $signed(op_5);
assign _028_ = | op_19[2:0];
assign _029_ = op_3 != { op_5[1], op_5 };
always @(posedge ap_clk)
zext_ln11_reg_512[1] <= 1'h0;
always @(posedge ap_clk)
ret_V_5_reg_569 <= _014_;
always @(posedge ap_clk)
op_31_V_reg_594 <= _010_;
always @(posedge ap_clk)
op_24_V_reg_532 <= _009_;
always @(posedge ap_clk)
op_16_V_reg_552 <= _008_;
always @(posedge ap_clk)
ret_V_4_reg_557 <= _013_;
always @(posedge ap_clk)
ret_V_cast_reg_562 <= _016_;
always @(posedge ap_clk)
ret_V_6_reg_599 <= _015_;
always @(posedge ap_clk)
ret_V_3_cast_reg_604 <= _012_;
always @(posedge ap_clk)
icmp_ln851_reg_611 <= _006_;
always @(posedge ap_clk)
select_ln69_reg_574 <= _017_;
always @(posedge ap_clk)
add_ln69_7_reg_579 <= _003_;
always @(posedge ap_clk)
add_ln69_4_reg_584 <= _002_;
always @(posedge ap_clk)
add_ln69_8_reg_589 <= _004_;
always @(posedge ap_clk)
add_ln69_2_reg_527 <= _001_;
always @(posedge ap_clk)
r_reg_507 <= _011_;
always @(posedge ap_clk)
zext_ln11_reg_512[0] <= _018_;
always @(posedge ap_clk)
icmp_ln890_reg_517 <= _007_;
always @(posedge ap_clk)
add_ln69_1_reg_522 <= _000_;
always @(posedge ap_clk)
ap_CS_fsm <= _005_;
assign _030_ = ap_CS_fsm == 1'h1;
function [9:0] _094_;
input [9:0] a;
input [99:0] b;
input [9:0] s;
case (s)
10'b0000000001:
_094_ = b[9:0];
10'b0000000010:
_094_ = b[19:10];
10'b0000000100:
_094_ = b[29:20];
10'b0000001000:
_094_ = b[39:30];
10'b0000010000:
_094_ = b[49:40];
10'b0000100000:
_094_ = b[59:50];
10'b0001000000:
_094_ = b[69:60];
10'b0010000000:
_094_ = b[79:70];
10'b0100000000:
_094_ = b[89:80];
10'b1000000000:
_094_ = b[99:90];
10'b0000000000:
_094_ = a;
default:
_094_ = 10'bx;
endcase
endfunction
assign ap_NS_fsm = _094_(10'hxxx, { 8'h00, _019_, 90'h00402010080402010080001 }, { _030_, _039_, _038_, _037_, _036_, _035_, _034_, _033_, _032_, _031_ });
assign _031_ = ap_CS_fsm == 10'h200;
assign _032_ = ap_CS_fsm == 9'h100;
assign _033_ = ap_CS_fsm == 8'h80;
assign _034_ = ap_CS_fsm == 7'h40;
assign _035_ = ap_CS_fsm == 6'h20;
assign _036_ = ap_CS_fsm == 5'h10;
assign _037_ = ap_CS_fsm == 4'h8;
assign _038_ = ap_CS_fsm == 3'h4;
assign _039_ = ap_CS_fsm == 2'h2;
assign op_32_ap_vld = ap_CS_fsm[9] ? 1'h1 : 1'h0;
assign ap_idle = _020_ ? 1'h1 : 1'h0;
assign _014_ = ap_CS_fsm[4] ? ret_V_5_fu_359_p3 : ret_V_5_reg_569;
assign _010_ = ap_CS_fsm[7] ? op_31_V_fu_422_p2 : op_31_V_reg_594;
assign _009_ = ap_CS_fsm[2] ? op_24_V_fu_275_p2 : op_24_V_reg_532;
assign _016_ = ap_CS_fsm[3] ? ret_V_4_fu_321_p2[32:1] : ret_V_cast_reg_562;
assign _013_ = ap_CS_fsm[3] ? ret_V_4_fu_321_p2 : ret_V_4_reg_557;
assign _008_ = ap_CS_fsm[3] ? op_16_V_fu_301_p2 : op_16_V_reg_552;
assign _006_ = ap_CS_fsm[8] ? icmp_ln851_fu_463_p2 : icmp_ln851_reg_611;
assign _012_ = ap_CS_fsm[8] ? ret_V_6_fu_443_p2[34:3] : ret_V_3_cast_reg_604;
assign _015_ = ap_CS_fsm[8] ? ret_V_6_fu_443_p2 : ret_V_6_reg_599;
assign _003_ = ap_CS_fsm[5] ? add_ln69_7_fu_391_p2 : add_ln69_7_reg_579;
assign _017_ = ap_CS_fsm[5] ? select_ln69_fu_371_p3 : select_ln69_reg_574;
assign _004_ = ap_CS_fsm[6] ? add_ln69_8_fu_408_p2 : add_ln69_8_reg_589;
assign _002_ = ap_CS_fsm[6] ? grp_fu_495_p3 : add_ln69_4_reg_584;
assign _001_ = ap_CS_fsm[1] ? add_ln69_2_fu_256_p2 : add_ln69_2_reg_527;
assign _000_ = ap_CS_fsm[0] ? add_ln69_1_fu_233_p2 : add_ln69_1_reg_522;
assign _007_ = ap_CS_fsm[0] ? icmp_ln890_fu_213_p2 : icmp_ln890_reg_517;
assign _018_ = ap_CS_fsm[0] ? lhs_V_fu_189_p2 : zext_ln11_reg_512[0];
assign _011_ = ap_CS_fsm[0] ? r_fu_171_p2 : r_reg_507;
assign _005_ = ap_rst ? 10'h001 : ap_NS_fsm;
assign _019_ = _021_ ? 2'h2 : 2'h1;
assign r_1_fu_219_p2 = op_3 >> lhs_V_fu_189_p2;
assign icmp_ln851_fu_463_p2 = _028_ ? 1'h1 : 1'h0;
assign icmp_ln890_fu_213_p2 = _027_ ? 1'h1 : 1'h0;
assign lhs_V_fu_189_p2 = _029_ ? 1'h1 : 1'h0;
assign op_32 = ret_V_6_reg_599[35] ? select_ln850_1_fu_481_p3 : ret_V_3_cast_reg_604;
assign ret_V_5_fu_359_p3 = ret_V_4_reg_557[33] ? select_ln850_fu_352_p3 : ret_V_cast_reg_562;
assign select_ln69_1_fu_383_p3 = op_18 ? 2'h3 : 2'h0;
assign select_ln69_fu_371_p3 = op_13 ? 3'h7 : 3'h0;
assign select_ln850_1_fu_481_p3 = icmp_ln851_reg_611 ? add_ln691_1_fu_476_p2 : ret_V_3_cast_reg_604;
assign select_ln850_fu_352_p3 = op_12[0] ? add_ln691_fu_347_p2 : ret_V_cast_reg_562;
assign op_16_V_fu_301_p2 = zext_ln11_reg_512 ^ grp_fu_495_p0[1:0];
assign op_9_V_fu_207_p2 = op_2[0] ^ op_5[0];
assign ap_CS_fsm_state1 = ap_CS_fsm[0];
assign ap_CS_fsm_state10 = ap_CS_fsm[9];
assign ap_CS_fsm_state2 = ap_CS_fsm[1];
assign ap_CS_fsm_state3 = ap_CS_fsm[2];
assign ap_CS_fsm_state4 = ap_CS_fsm[3];
assign ap_CS_fsm_state5 = ap_CS_fsm[4];
assign ap_CS_fsm_state6 = ap_CS_fsm[5];
assign ap_CS_fsm_state7 = ap_CS_fsm[6];
assign ap_CS_fsm_state8 = ap_CS_fsm[7];
assign ap_CS_fsm_state9 = ap_CS_fsm[8];
assign ap_done = op_32_ap_vld;
assign ap_ready = op_32_ap_vld;
assign grp_fu_495_p00 = { 4'h0, grp_fu_495_p0 };
assign p_Result_1_fu_469_p3 = ret_V_6_reg_599[35];
assign p_Result_s_fu_337_p3 = ret_V_4_reg_557[33];
assign ret_1_fu_284_p0 = op_3;
assign ret_1_fu_284_p1 = op_3;
assign ret_1_fu_284_p2 = grp_fu_495_p0;
assign rhs_1_fu_310_p3 = { op_24_V_reg_532, 1'h0 };
assign rhs_3_fu_432_p3 = { op_31_V_reg_594, 3'h0 };
assign sext_ln1192_1_fu_439_p1 = { op_31_V_reg_594[31], op_31_V_reg_594, 3'h0 };
assign sext_ln1192_fu_317_p1 = { op_24_V_reg_532[31], op_24_V_reg_532, 1'h0 };
assign sext_ln215_1_fu_243_p1 = { op_1[3], op_1[3], op_1[3], op_1[3], op_1[3], op_1 };
assign sext_ln215_fu_239_p1 = { op_0[7], op_0 };
assign sext_ln69_1_fu_272_p1 = { add_ln69_2_reg_527[8], add_ln69_2_reg_527[8], add_ln69_2_reg_527[8], add_ln69_2_reg_527[8], add_ln69_2_reg_527[8], add_ln69_2_reg_527[8], add_ln69_2_reg_527[8], add_ln69_2_reg_527[8], add_ln69_2_reg_527[8], add_ln69_2_reg_527[8], add_ln69_2_reg_527[8], add_ln69_2_reg_527[8], add_ln69_2_reg_527[8], add_ln69_2_reg_527[8], add_ln69_2_reg_527[8], add_ln69_2_reg_527[8], add_ln69_2_reg_527[8], add_ln69_2_reg_527[8], add_ln69_2_reg_527[8], add_ln69_2_reg_527[8], add_ln69_2_reg_527[8], add_ln69_2_reg_527[8], add_ln69_2_reg_527[8], add_ln69_2_reg_527 };
assign sext_ln69_2_fu_397_p1 = { op_16_V_reg_552[1], op_16_V_reg_552 };
assign sext_ln69_4_fu_405_p1 = { add_ln69_7_reg_579[1], add_ln69_7_reg_579 };
assign sext_ln69_5_fu_419_p1 = { add_ln69_8_reg_589[2], add_ln69_8_reg_589[2], add_ln69_8_reg_589[2], add_ln69_8_reg_589[2], add_ln69_8_reg_589[2], add_ln69_8_reg_589[2], add_ln69_8_reg_589[2], add_ln69_8_reg_589[2], add_ln69_8_reg_589[2], add_ln69_8_reg_589[2], add_ln69_8_reg_589[2], add_ln69_8_reg_589[2], add_ln69_8_reg_589[2], add_ln69_8_reg_589[2], add_ln69_8_reg_589[2], add_ln69_8_reg_589[2], add_ln69_8_reg_589[2], add_ln69_8_reg_589[2], add_ln69_8_reg_589[2], add_ln69_8_reg_589[2], add_ln69_8_reg_589[2], add_ln69_8_reg_589[2], add_ln69_8_reg_589[2], add_ln69_8_reg_589[2], add_ln69_8_reg_589[2], add_ln69_8_reg_589[2], add_ln69_8_reg_589[2], add_ln69_8_reg_589[2], add_ln69_8_reg_589[2], add_ln69_8_reg_589 };
assign sext_ln703_1_fu_428_p0 = op_19;
assign sext_ln703_1_fu_428_p1 = { op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19 };
assign sext_ln703_fu_306_p0 = op_12;
assign sext_ln703_fu_306_p1 = { op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12 };
assign sext_ln874_1_fu_185_p0 = op_5;
assign sext_ln874_1_fu_185_p1 = { op_5[1], op_5 };
assign sext_ln874_fu_181_p0 = op_5;
assign sext_ln874_fu_181_p1 = { op_5[1], op_5[1], op_5 };
assign trunc_ln1350_fu_297_p1 = grp_fu_495_p0[1:0];
assign trunc_ln213_1_fu_203_p0 = op_5;
assign trunc_ln213_1_fu_203_p1 = op_5[0];
assign trunc_ln213_fu_199_p1 = op_2[0];
assign trunc_ln851_1_fu_459_p0 = op_19;
assign trunc_ln851_1_fu_459_p1 = op_19[2:0];
assign trunc_ln851_fu_344_p0 = op_12;
assign trunc_ln851_fu_344_p1 = op_12[0];
assign zext_ln11_fu_195_p1 = { 1'h0, lhs_V_fu_189_p2 };
assign zext_ln1345_fu_281_p1 = { 2'h0, op_3 };
assign zext_ln69_2_fu_225_p1 = { 2'h0, op_9_V_fu_207_p2 };
assign zext_ln69_3_fu_229_p1 = { 1'h0, r_1_fu_219_p2 };
assign zext_ln69_4_fu_253_p1 = { 6'h00, add_ln69_1_reg_522 };
assign zext_ln69_5_fu_379_p1 = { 1'h0, xor_ln890_fu_366_p2 };
assign zext_ln69_fu_262_p1 = { 16'h0000, op_4 };
assign zext_ln874_fu_177_p1 = { 1'h0, op_3 };
assign \mul_2ns_2ns_4_1_1_U1.top_mul_2ns_2ns_4_1_1_Multiplier_0_U.a  = \mul_2ns_2ns_4_1_1_U1.din0 ;
assign \mul_2ns_2ns_4_1_1_U1.top_mul_2ns_2ns_4_1_1_Multiplier_0_U.b  = \mul_2ns_2ns_4_1_1_U1.din1 ;
assign \mul_2ns_2ns_4_1_1_U1.dout  = \mul_2ns_2ns_4_1_1_U1.top_mul_2ns_2ns_4_1_1_Multiplier_0_U.p ;
assign \mul_2ns_2ns_4_1_1_U1.din0  = op_3;
assign \mul_2ns_2ns_4_1_1_U1.din1  = op_3;
assign grp_fu_495_p0 = \mul_2ns_2ns_4_1_1_U1.dout ;
assign \mac_muladd_4ns_4s_32ns_32_4_1_U2.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.a  = { 21'h000000, \mac_muladd_4ns_4s_32ns_32_4_1_U2.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.in0  };
assign \mac_muladd_4ns_4s_32ns_32_4_1_U2.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.b  = { \mac_muladd_4ns_4s_32ns_32_4_1_U2.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.in1 [3], \mac_muladd_4ns_4s_32ns_32_4_1_U2.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.in1 [3], \mac_muladd_4ns_4s_32ns_32_4_1_U2.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.in1 [3], \mac_muladd_4ns_4s_32ns_32_4_1_U2.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.in1 [3], \mac_muladd_4ns_4s_32ns_32_4_1_U2.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.in1 [3], \mac_muladd_4ns_4s_32ns_32_4_1_U2.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.in1 [3], \mac_muladd_4ns_4s_32ns_32_4_1_U2.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.in1 [3], \mac_muladd_4ns_4s_32ns_32_4_1_U2.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.in1 [3], \mac_muladd_4ns_4s_32ns_32_4_1_U2.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.in1 [3], \mac_muladd_4ns_4s_32ns_32_4_1_U2.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.in1 [3], \mac_muladd_4ns_4s_32ns_32_4_1_U2.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.in1 [3], \mac_muladd_4ns_4s_32ns_32_4_1_U2.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.in1 [3], \mac_muladd_4ns_4s_32ns_32_4_1_U2.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.in1 [3], \mac_muladd_4ns_4s_32ns_32_4_1_U2.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.in1 [3], \mac_muladd_4ns_4s_32ns_32_4_1_U2.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.in1  };
assign \mac_muladd_4ns_4s_32ns_32_4_1_U2.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.c  = { 16'h0000, \mac_muladd_4ns_4s_32ns_32_4_1_U2.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.in2  };
assign \mac_muladd_4ns_4s_32ns_32_4_1_U2.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.dout  = \mac_muladd_4ns_4s_32ns_32_4_1_U2.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.p_reg [31:0];
assign \mac_muladd_4ns_4s_32ns_32_4_1_U2.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.p [46:43] = { \mac_muladd_4ns_4s_32ns_32_4_1_U2.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.p [47], \mac_muladd_4ns_4s_32ns_32_4_1_U2.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.p [47], \mac_muladd_4ns_4s_32ns_32_4_1_U2.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.p [47], \mac_muladd_4ns_4s_32ns_32_4_1_U2.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.p [47] };
assign \mac_muladd_4ns_4s_32ns_32_4_1_U2.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.ce  = \mac_muladd_4ns_4s_32ns_32_4_1_U2.ce ;
assign \mac_muladd_4ns_4s_32ns_32_4_1_U2.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.clk  = \mac_muladd_4ns_4s_32ns_32_4_1_U2.clk ;
assign \mac_muladd_4ns_4s_32ns_32_4_1_U2.dout  = \mac_muladd_4ns_4s_32ns_32_4_1_U2.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.dout ;
assign \mac_muladd_4ns_4s_32ns_32_4_1_U2.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.in0  = \mac_muladd_4ns_4s_32ns_32_4_1_U2.din0 ;
assign \mac_muladd_4ns_4s_32ns_32_4_1_U2.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.in1  = \mac_muladd_4ns_4s_32ns_32_4_1_U2.din1 ;
assign \mac_muladd_4ns_4s_32ns_32_4_1_U2.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.in2  = \mac_muladd_4ns_4s_32ns_32_4_1_U2.din2 ;
assign \mac_muladd_4ns_4s_32ns_32_4_1_U2.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.rst  = \mac_muladd_4ns_4s_32ns_32_4_1_U2.reset ;
assign \mac_muladd_4ns_4s_32ns_32_4_1_U2.ce  = 1'h1;
assign \mac_muladd_4ns_4s_32ns_32_4_1_U2.clk  = ap_clk;
assign \mac_muladd_4ns_4s_32ns_32_4_1_U2.din0  = grp_fu_495_p0;
assign \mac_muladd_4ns_4s_32ns_32_4_1_U2.din1  = r_reg_507;
assign \mac_muladd_4ns_4s_32ns_32_4_1_U2.din2  = ret_V_5_reg_569;
assign grp_fu_495_p3 = \mac_muladd_4ns_4s_32ns_32_4_1_U2.dout ;
assign \mac_muladd_4ns_4s_32ns_32_4_1_U2.reset  = ap_rst;
endmodule


// Machine B:
// Processed by function `add_clk_enable_signal` in `verilog_tricks.py`.
// Processed by function `remove_reset_signal` in `verilog_tricks.py`.
module top_B (
  ap_clk,
  ap_start,
  ap_done,
  ap_idle,
  ap_ready,
  op_0,
  op_1,
  op_2,
  op_3,
  op_4,
  op_5,
  op_10,
  op_12,
  op_13,
  op_14,
  op_18,
  op_19,
  op_32,
  op_32_ap_vld,
clk_enable
);
input clk_enable;


input ap_clk;
wire ap_rst;
assign ap_rst = op_32_ap_vld;
input ap_start;
input [7:0] op_0;
input [3:0] op_1;
input [31:0] op_10;
input [1:0] op_12;
input op_13;
input [31:0] op_14;
input op_18;
input [3:0] op_19;
input [3:0] op_2;
input [1:0] op_3;
input [15:0] op_4;
input [1:0] op_5;
output ap_done;
output ap_idle;
output ap_ready;
output [31:0] op_32;
output op_32_ap_vld;


reg \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_7_U.ain_s1 ;
reg \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_7_U.bin_s1 ;
reg \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_7_U.carry_s1 ;
reg \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_7_U.sum_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_2_U.ain_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_2_U.bin_s1 ;
reg \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_2_U.carry_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_2_U.sum_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_2_U.ain_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_2_U.bin_s1 ;
reg \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_2_U.carry_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_2_U.sum_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_2_U.ain_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_2_U.bin_s1 ;
reg \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_2_U.carry_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_2_U.sum_s1 ;
reg [15:0] \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_4_U.ain_s1 ;
reg [15:0] \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_4_U.bin_s1 ;
reg \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_4_U.carry_s1 ;
reg [15:0] \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_4_U.sum_s1 ;
reg [15:0] \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_4_U.ain_s1 ;
reg [15:0] \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_4_U.bin_s1 ;
reg \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_4_U.carry_s1 ;
reg [15:0] \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_4_U.sum_s1 ;
reg [15:0] \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_4_U.ain_s1 ;
reg [15:0] \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_4_U.bin_s1 ;
reg \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_4_U.carry_s1 ;
reg [15:0] \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_4_U.sum_s1 ;
reg [16:0] \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_5_U.ain_s1 ;
reg [16:0] \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_5_U.bin_s1 ;
reg \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_5_U.carry_s1 ;
reg [16:0] \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_5_U.sum_s1 ;
reg [17:0] \add_36s_36s_36_2_1_U15.top_add_36s_36s_36_2_1_Adder_8_U.ain_s1 ;
reg [17:0] \add_36s_36s_36_2_1_U15.top_add_36s_36s_36_2_1_Adder_8_U.bin_s1 ;
reg \add_36s_36s_36_2_1_U15.top_add_36s_36s_36_2_1_Adder_8_U.carry_s1 ;
reg [17:0] \add_36s_36s_36_2_1_U15.top_add_36s_36s_36_2_1_Adder_8_U.sum_s1 ;
reg [1:0] \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_1_U.ain_s1 ;
reg [1:0] \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_1_U.bin_s1 ;
reg \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_1_U.carry_s1 ;
reg \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_1_U.sum_s1 ;
reg [1:0] \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.ain_s1 ;
reg [1:0] \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.bin_s1 ;
reg \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.carry_s1 ;
reg \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.sum_s1 ;
reg [1:0] \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_6_U.ain_s1 ;
reg [1:0] \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_6_U.bin_s1 ;
reg \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_6_U.carry_s1 ;
reg \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_6_U.sum_s1 ;
reg [4:0] \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_3_U.ain_s1 ;
reg [4:0] \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_3_U.bin_s1 ;
reg \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_3_U.carry_s1 ;
reg [3:0] \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_3_U.sum_s1 ;
reg [4:0] \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_0_U.ain_s1 ;
reg [4:0] \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_0_U.bin_s1 ;
reg \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_0_U.carry_s1 ;
reg [3:0] \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_0_U.sum_s1 ;
reg [31:0] add_ln691_1_reg_757;
reg [31:0] add_ln691_reg_650;
reg [2:0] add_ln69_1_reg_558;
reg [8:0] add_ln69_2_reg_583;
reg [31:0] add_ln69_4_reg_685;
reg [31:0] add_ln69_5_reg_710;
reg [2:0] add_ln69_6_reg_690;
reg [1:0] add_ln69_7_reg_695;
reg [2:0] add_ln69_8_reg_715;
reg [31:0] add_ln69_reg_578;
reg [29:0] ap_CS_fsm = 30'h00000001;
reg icmp_ln851_reg_740;
reg icmp_ln890_reg_538;
reg lhs_V_reg_496;
reg \lshr_2ns_1ns_2_7_1_U1.din1_cast_array[0] ;
reg \lshr_2ns_1ns_2_7_1_U1.din1_cast_array[1] ;
reg \lshr_2ns_1ns_2_7_1_U1.din1_cast_array[2] ;
reg \lshr_2ns_1ns_2_7_1_U1.din1_cast_array[3] ;
reg \lshr_2ns_1ns_2_7_1_U1.din1_cast_array[4] ;
reg \lshr_2ns_1ns_2_7_1_U1.din1_cast_array[5] ;
reg [1:0] \lshr_2ns_1ns_2_7_1_U1.dout_array[0] ;
reg [1:0] \lshr_2ns_1ns_2_7_1_U1.dout_array[1] ;
reg [1:0] \lshr_2ns_1ns_2_7_1_U1.dout_array[2] ;
reg [1:0] \lshr_2ns_1ns_2_7_1_U1.dout_array[3] ;
reg [1:0] \lshr_2ns_1ns_2_7_1_U1.dout_array[4] ;
reg [1:0] \lshr_2ns_1ns_2_7_1_U1.dout_array[5] ;
reg [24:0] \mac_muladd_4ns_4s_32ns_32_4_1_U17.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.a_reg ;
reg [17:0] \mac_muladd_4ns_4s_32ns_32_4_1_U17.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.b_reg ;
reg [42:0] \mac_muladd_4ns_4s_32ns_32_4_1_U17.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.m_reg ;
reg [47:0] \mac_muladd_4ns_4s_32ns_32_4_1_U17.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.p_reg ;
reg [1:0] op_16_V_reg_645;
reg [31:0] op_24_V_reg_593;
reg [31:0] op_31_V_reg_725;
reg op_9_V_reg_518;
reg [1:0] r_1_reg_523;
reg [3:0] r_reg_512;
reg [3:0] ret_1_reg_625;
reg [31:0] ret_V_3_cast_reg_750;
reg [33:0] ret_V_4_reg_613;
reg [31:0] ret_V_5_reg_660;
reg [35:0] ret_V_6_reg_745;
reg [31:0] ret_V_cast_reg_618;
reg [8:0] ret_reg_553;
reg [1:0] select_ln69_1_reg_670;
reg [2:0] select_ln69_reg_665;
reg [1:0] trunc_ln1350_reg_630;
reg trunc_ln213_1_reg_501;
reg xor_ln890_reg_655;
reg [1:0] zext_ln11_reg_506;
wire [31:0] _000_;
wire [31:0] _001_;
wire [2:0] _002_;
wire [8:0] _003_;
wire [31:0] _004_;
wire [31:0] _005_;
wire [2:0] _006_;
wire [1:0] _007_;
wire [2:0] _008_;
wire [31:0] _009_;
wire [29:0] _010_;
wire _011_;
wire _012_;
wire _013_;
wire [1:0] _014_;
wire [31:0] _015_;
wire [31:0] _016_;
wire _017_;
wire [1:0] _018_;
wire [3:0] _019_;
wire [3:0] _020_;
wire [31:0] _021_;
wire [33:0] _022_;
wire [31:0] _023_;
wire [35:0] _024_;
wire [31:0] _025_;
wire [8:0] _026_;
wire [1:0] _027_;
wire [2:0] _028_;
wire [1:0] _029_;
wire _030_;
wire _031_;
wire _032_;
wire [1:0] _033_;
wire _034_;
wire _035_;
wire _036_;
wire _037_;
wire _038_;
wire _039_;
wire _040_;
wire _041_;
wire [1:0] _042_;
wire [1:0] _043_;
wire [15:0] _044_;
wire [15:0] _045_;
wire _046_;
wire [15:0] _047_;
wire [16:0] _048_;
wire [16:0] _049_;
wire [15:0] _050_;
wire [15:0] _051_;
wire _052_;
wire [15:0] _053_;
wire [16:0] _054_;
wire [16:0] _055_;
wire [15:0] _056_;
wire [15:0] _057_;
wire _058_;
wire [15:0] _059_;
wire [16:0] _060_;
wire [16:0] _061_;
wire [15:0] _062_;
wire [15:0] _063_;
wire _064_;
wire [15:0] _065_;
wire [16:0] _066_;
wire [16:0] _067_;
wire [15:0] _068_;
wire [15:0] _069_;
wire _070_;
wire [15:0] _071_;
wire [16:0] _072_;
wire [16:0] _073_;
wire [15:0] _074_;
wire [15:0] _075_;
wire _076_;
wire [15:0] _077_;
wire [16:0] _078_;
wire [16:0] _079_;
wire [16:0] _080_;
wire [16:0] _081_;
wire _082_;
wire [16:0] _083_;
wire [17:0] _084_;
wire [17:0] _085_;
wire [17:0] _086_;
wire [17:0] _087_;
wire _088_;
wire [17:0] _089_;
wire [18:0] _090_;
wire [18:0] _091_;
wire [1:0] _092_;
wire [1:0] _093_;
wire _094_;
wire _095_;
wire [1:0] _096_;
wire [2:0] _097_;
wire [1:0] _098_;
wire [1:0] _099_;
wire _100_;
wire _101_;
wire [1:0] _102_;
wire [2:0] _103_;
wire [1:0] _104_;
wire [1:0] _105_;
wire _106_;
wire _107_;
wire [1:0] _108_;
wire [2:0] _109_;
wire [4:0] _110_;
wire [4:0] _111_;
wire _112_;
wire [3:0] _113_;
wire [4:0] _114_;
wire [5:0] _115_;
wire [4:0] _116_;
wire [4:0] _117_;
wire _118_;
wire [3:0] _119_;
wire [4:0] _120_;
wire [5:0] _121_;
wire _122_;
wire _123_;
wire _124_;
wire _125_;
wire _126_;
wire _127_;
wire [1:0] _128_;
wire [1:0] _129_;
wire [1:0] _130_;
wire [1:0] _131_;
wire [1:0] _132_;
wire [1:0] _133_;
wire _134_;
wire [1:0] _135_;
wire _136_;
wire [1:0] _137_;
wire _138_;
wire [1:0] _139_;
wire _140_;
wire [1:0] _141_;
wire _142_;
wire [1:0] _143_;
wire _144_;
wire [1:0] _145_;
wire [24:0] _146_;
wire [17:0] _147_;
wire [42:0] _148_;
wire [47:0] _149_;
wire _150_;
wire _151_;
wire _152_;
wire _153_;
wire _154_;
wire _155_;
wire _156_;
wire _157_;
wire _158_;
wire _159_;
wire _160_;
wire _161_;
wire _162_;
wire _163_;
wire _164_;
wire _165_;
wire _166_;
wire _167_;
wire _168_;
wire _169_;
wire _170_;
wire _171_;
wire _172_;
wire _173_;
wire _174_;
wire _175_;
wire _176_;
wire _177_;
wire _178_;
wire _179_;
wire _180_;
wire _181_;
wire _182_;
wire \add_2ns_2ns_2_2_1_U11.ce ;
wire \add_2ns_2ns_2_2_1_U11.clk ;
wire [1:0] \add_2ns_2ns_2_2_1_U11.din0 ;
wire [1:0] \add_2ns_2ns_2_2_1_U11.din1 ;
wire [1:0] \add_2ns_2ns_2_2_1_U11.dout ;
wire \add_2ns_2ns_2_2_1_U11.reset ;
wire [1:0] \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_7_U.a ;
wire [1:0] \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_7_U.ain_s0 ;
wire [1:0] \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_7_U.b ;
wire [1:0] \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_7_U.bin_s0 ;
wire \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_7_U.ce ;
wire \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_7_U.clk ;
wire \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_7_U.facout_s1 ;
wire \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_7_U.facout_s2 ;
wire \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_7_U.fas_s1 ;
wire \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_7_U.fas_s2 ;
wire \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_7_U.reset ;
wire [1:0] \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_7_U.s ;
wire \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_7_U.u1.a ;
wire \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_7_U.u1.b ;
wire \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_7_U.u1.cin ;
wire \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_7_U.u1.cout ;
wire \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_7_U.u1.s ;
wire \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_7_U.u2.a ;
wire \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_7_U.u2.b ;
wire \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_7_U.u2.cin ;
wire \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_7_U.u2.cout ;
wire \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_7_U.u2.s ;
wire \add_32ns_32ns_32_2_1_U16.ce ;
wire \add_32ns_32ns_32_2_1_U16.clk ;
wire [31:0] \add_32ns_32ns_32_2_1_U16.din0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U16.din1 ;
wire [31:0] \add_32ns_32ns_32_2_1_U16.dout ;
wire \add_32ns_32ns_32_2_1_U16.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_2_U.a ;
wire [31:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_2_U.ain_s0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_2_U.b ;
wire [31:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_2_U.bin_s0 ;
wire \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_2_U.ce ;
wire \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_2_U.clk ;
wire \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_2_U.facout_s1 ;
wire \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_2_U.facout_s2 ;
wire [15:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_2_U.fas_s1 ;
wire [15:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_2_U.fas_s2 ;
wire \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_2_U.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_2_U.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_2_U.u1.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_2_U.u1.b ;
wire \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_2_U.u1.cin ;
wire \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_2_U.u1.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_2_U.u1.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_2_U.u2.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_2_U.u2.b ;
wire \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_2_U.u2.cin ;
wire \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_2_U.u2.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_2_U.u2.s ;
wire \add_32ns_32ns_32_2_1_U4.ce ;
wire \add_32ns_32ns_32_2_1_U4.clk ;
wire [31:0] \add_32ns_32ns_32_2_1_U4.din0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U4.din1 ;
wire [31:0] \add_32ns_32ns_32_2_1_U4.dout ;
wire \add_32ns_32ns_32_2_1_U4.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_2_U.a ;
wire [31:0] \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_2_U.ain_s0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_2_U.b ;
wire [31:0] \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_2_U.bin_s0 ;
wire \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_2_U.ce ;
wire \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_2_U.clk ;
wire \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_2_U.facout_s1 ;
wire \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_2_U.facout_s2 ;
wire [15:0] \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_2_U.fas_s1 ;
wire [15:0] \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_2_U.fas_s2 ;
wire \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_2_U.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_2_U.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_2_U.u1.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_2_U.u1.b ;
wire \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_2_U.u1.cin ;
wire \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_2_U.u1.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_2_U.u1.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_2_U.u2.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_2_U.u2.b ;
wire \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_2_U.u2.cin ;
wire \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_2_U.u2.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_2_U.u2.s ;
wire \add_32ns_32ns_32_2_1_U9.ce ;
wire \add_32ns_32ns_32_2_1_U9.clk ;
wire [31:0] \add_32ns_32ns_32_2_1_U9.din0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U9.din1 ;
wire [31:0] \add_32ns_32ns_32_2_1_U9.dout ;
wire \add_32ns_32ns_32_2_1_U9.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_2_U.a ;
wire [31:0] \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_2_U.ain_s0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_2_U.b ;
wire [31:0] \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_2_U.bin_s0 ;
wire \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_2_U.ce ;
wire \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_2_U.clk ;
wire \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_2_U.facout_s1 ;
wire \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_2_U.facout_s2 ;
wire [15:0] \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_2_U.fas_s1 ;
wire [15:0] \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_2_U.fas_s2 ;
wire \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_2_U.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_2_U.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_2_U.u1.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_2_U.u1.b ;
wire \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_2_U.u1.cin ;
wire \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_2_U.u1.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_2_U.u1.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_2_U.u2.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_2_U.u2.b ;
wire \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_2_U.u2.cin ;
wire \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_2_U.u2.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_2_U.u2.s ;
wire \add_32s_32ns_32_2_1_U12.ce ;
wire \add_32s_32ns_32_2_1_U12.clk ;
wire [31:0] \add_32s_32ns_32_2_1_U12.din0 ;
wire [31:0] \add_32s_32ns_32_2_1_U12.din1 ;
wire [31:0] \add_32s_32ns_32_2_1_U12.dout ;
wire \add_32s_32ns_32_2_1_U12.reset ;
wire [31:0] \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_4_U.a ;
wire [31:0] \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_4_U.ain_s0 ;
wire [31:0] \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_4_U.b ;
wire [31:0] \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_4_U.bin_s0 ;
wire \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_4_U.ce ;
wire \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_4_U.clk ;
wire \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_4_U.facout_s1 ;
wire \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_4_U.facout_s2 ;
wire [15:0] \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_4_U.fas_s1 ;
wire [15:0] \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_4_U.fas_s2 ;
wire \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_4_U.reset ;
wire [31:0] \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_4_U.s ;
wire [15:0] \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_4_U.u1.a ;
wire [15:0] \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_4_U.u1.b ;
wire \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_4_U.u1.cin ;
wire \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_4_U.u1.cout ;
wire [15:0] \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_4_U.u1.s ;
wire [15:0] \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_4_U.u2.a ;
wire [15:0] \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_4_U.u2.b ;
wire \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_4_U.u2.cin ;
wire \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_4_U.u2.cout ;
wire [15:0] \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_4_U.u2.s ;
wire \add_32s_32ns_32_2_1_U14.ce ;
wire \add_32s_32ns_32_2_1_U14.clk ;
wire [31:0] \add_32s_32ns_32_2_1_U14.din0 ;
wire [31:0] \add_32s_32ns_32_2_1_U14.din1 ;
wire [31:0] \add_32s_32ns_32_2_1_U14.dout ;
wire \add_32s_32ns_32_2_1_U14.reset ;
wire [31:0] \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_4_U.a ;
wire [31:0] \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_4_U.ain_s0 ;
wire [31:0] \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_4_U.b ;
wire [31:0] \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_4_U.bin_s0 ;
wire \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_4_U.ce ;
wire \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_4_U.clk ;
wire \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_4_U.facout_s1 ;
wire \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_4_U.facout_s2 ;
wire [15:0] \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_4_U.fas_s1 ;
wire [15:0] \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_4_U.fas_s2 ;
wire \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_4_U.reset ;
wire [31:0] \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_4_U.s ;
wire [15:0] \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_4_U.u1.a ;
wire [15:0] \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_4_U.u1.b ;
wire \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_4_U.u1.cin ;
wire \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_4_U.u1.cout ;
wire [15:0] \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_4_U.u1.s ;
wire [15:0] \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_4_U.u2.a ;
wire [15:0] \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_4_U.u2.b ;
wire \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_4_U.u2.cin ;
wire \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_4_U.u2.cout ;
wire [15:0] \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_4_U.u2.s ;
wire \add_32s_32ns_32_2_1_U6.ce ;
wire \add_32s_32ns_32_2_1_U6.clk ;
wire [31:0] \add_32s_32ns_32_2_1_U6.din0 ;
wire [31:0] \add_32s_32ns_32_2_1_U6.din1 ;
wire [31:0] \add_32s_32ns_32_2_1_U6.dout ;
wire \add_32s_32ns_32_2_1_U6.reset ;
wire [31:0] \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_4_U.a ;
wire [31:0] \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_4_U.ain_s0 ;
wire [31:0] \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_4_U.b ;
wire [31:0] \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_4_U.bin_s0 ;
wire \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_4_U.ce ;
wire \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_4_U.clk ;
wire \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_4_U.facout_s1 ;
wire \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_4_U.facout_s2 ;
wire [15:0] \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_4_U.fas_s1 ;
wire [15:0] \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_4_U.fas_s2 ;
wire \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_4_U.reset ;
wire [31:0] \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_4_U.s ;
wire [15:0] \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_4_U.u1.a ;
wire [15:0] \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_4_U.u1.b ;
wire \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_4_U.u1.cin ;
wire \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_4_U.u1.cout ;
wire [15:0] \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_4_U.u1.s ;
wire [15:0] \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_4_U.u2.a ;
wire [15:0] \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_4_U.u2.b ;
wire \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_4_U.u2.cin ;
wire \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_4_U.u2.cout ;
wire [15:0] \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_4_U.u2.s ;
wire \add_34s_34s_34_2_1_U7.ce ;
wire \add_34s_34s_34_2_1_U7.clk ;
wire [33:0] \add_34s_34s_34_2_1_U7.din0 ;
wire [33:0] \add_34s_34s_34_2_1_U7.din1 ;
wire [33:0] \add_34s_34s_34_2_1_U7.dout ;
wire \add_34s_34s_34_2_1_U7.reset ;
wire [33:0] \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_5_U.a ;
wire [33:0] \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_5_U.ain_s0 ;
wire [33:0] \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_5_U.b ;
wire [33:0] \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_5_U.bin_s0 ;
wire \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_5_U.ce ;
wire \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_5_U.clk ;
wire \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_5_U.facout_s1 ;
wire \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_5_U.facout_s2 ;
wire [16:0] \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_5_U.fas_s1 ;
wire [16:0] \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_5_U.fas_s2 ;
wire \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_5_U.reset ;
wire [33:0] \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_5_U.s ;
wire [16:0] \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_5_U.u1.a ;
wire [16:0] \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_5_U.u1.b ;
wire \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_5_U.u1.cin ;
wire \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_5_U.u1.cout ;
wire [16:0] \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_5_U.u1.s ;
wire [16:0] \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_5_U.u2.a ;
wire [16:0] \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_5_U.u2.b ;
wire \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_5_U.u2.cin ;
wire \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_5_U.u2.cout ;
wire [16:0] \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_5_U.u2.s ;
wire \add_36s_36s_36_2_1_U15.ce ;
wire \add_36s_36s_36_2_1_U15.clk ;
wire [35:0] \add_36s_36s_36_2_1_U15.din0 ;
wire [35:0] \add_36s_36s_36_2_1_U15.din1 ;
wire [35:0] \add_36s_36s_36_2_1_U15.dout ;
wire \add_36s_36s_36_2_1_U15.reset ;
wire [35:0] \add_36s_36s_36_2_1_U15.top_add_36s_36s_36_2_1_Adder_8_U.a ;
wire [35:0] \add_36s_36s_36_2_1_U15.top_add_36s_36s_36_2_1_Adder_8_U.ain_s0 ;
wire [35:0] \add_36s_36s_36_2_1_U15.top_add_36s_36s_36_2_1_Adder_8_U.b ;
wire [35:0] \add_36s_36s_36_2_1_U15.top_add_36s_36s_36_2_1_Adder_8_U.bin_s0 ;
wire \add_36s_36s_36_2_1_U15.top_add_36s_36s_36_2_1_Adder_8_U.ce ;
wire \add_36s_36s_36_2_1_U15.top_add_36s_36s_36_2_1_Adder_8_U.clk ;
wire \add_36s_36s_36_2_1_U15.top_add_36s_36s_36_2_1_Adder_8_U.facout_s1 ;
wire \add_36s_36s_36_2_1_U15.top_add_36s_36s_36_2_1_Adder_8_U.facout_s2 ;
wire [17:0] \add_36s_36s_36_2_1_U15.top_add_36s_36s_36_2_1_Adder_8_U.fas_s1 ;
wire [17:0] \add_36s_36s_36_2_1_U15.top_add_36s_36s_36_2_1_Adder_8_U.fas_s2 ;
wire \add_36s_36s_36_2_1_U15.top_add_36s_36s_36_2_1_Adder_8_U.reset ;
wire [35:0] \add_36s_36s_36_2_1_U15.top_add_36s_36s_36_2_1_Adder_8_U.s ;
wire [17:0] \add_36s_36s_36_2_1_U15.top_add_36s_36s_36_2_1_Adder_8_U.u1.a ;
wire [17:0] \add_36s_36s_36_2_1_U15.top_add_36s_36s_36_2_1_Adder_8_U.u1.b ;
wire \add_36s_36s_36_2_1_U15.top_add_36s_36s_36_2_1_Adder_8_U.u1.cin ;
wire \add_36s_36s_36_2_1_U15.top_add_36s_36s_36_2_1_Adder_8_U.u1.cout ;
wire [17:0] \add_36s_36s_36_2_1_U15.top_add_36s_36s_36_2_1_Adder_8_U.u1.s ;
wire [17:0] \add_36s_36s_36_2_1_U15.top_add_36s_36s_36_2_1_Adder_8_U.u2.a ;
wire [17:0] \add_36s_36s_36_2_1_U15.top_add_36s_36s_36_2_1_Adder_8_U.u2.b ;
wire \add_36s_36s_36_2_1_U15.top_add_36s_36s_36_2_1_Adder_8_U.u2.cin ;
wire \add_36s_36s_36_2_1_U15.top_add_36s_36s_36_2_1_Adder_8_U.u2.cout ;
wire [17:0] \add_36s_36s_36_2_1_U15.top_add_36s_36s_36_2_1_Adder_8_U.u2.s ;
wire \add_3ns_3ns_3_2_1_U3.ce ;
wire \add_3ns_3ns_3_2_1_U3.clk ;
wire [2:0] \add_3ns_3ns_3_2_1_U3.din0 ;
wire [2:0] \add_3ns_3ns_3_2_1_U3.din1 ;
wire [2:0] \add_3ns_3ns_3_2_1_U3.dout ;
wire \add_3ns_3ns_3_2_1_U3.reset ;
wire [2:0] \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_1_U.a ;
wire [2:0] \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_1_U.ain_s0 ;
wire [2:0] \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_1_U.b ;
wire [2:0] \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_1_U.bin_s0 ;
wire \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_1_U.ce ;
wire \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_1_U.clk ;
wire \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_1_U.facout_s1 ;
wire \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_1_U.facout_s2 ;
wire \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_1_U.fas_s1 ;
wire [1:0] \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_1_U.fas_s2 ;
wire \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_1_U.reset ;
wire [2:0] \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_1_U.s ;
wire \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_1_U.u1.a ;
wire \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_1_U.u1.b ;
wire \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_1_U.u1.cin ;
wire \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_1_U.u1.cout ;
wire \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_1_U.u1.s ;
wire [1:0] \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_1_U.u2.a ;
wire [1:0] \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_1_U.u2.b ;
wire \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_1_U.u2.cin ;
wire \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_1_U.u2.cout ;
wire [1:0] \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_1_U.u2.s ;
wire \add_3s_3ns_3_2_1_U10.ce ;
wire \add_3s_3ns_3_2_1_U10.clk ;
wire [2:0] \add_3s_3ns_3_2_1_U10.din0 ;
wire [2:0] \add_3s_3ns_3_2_1_U10.din1 ;
wire [2:0] \add_3s_3ns_3_2_1_U10.dout ;
wire \add_3s_3ns_3_2_1_U10.reset ;
wire [2:0] \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.a ;
wire [2:0] \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.ain_s0 ;
wire [2:0] \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.b ;
wire [2:0] \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.bin_s0 ;
wire \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.ce ;
wire \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.clk ;
wire \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.facout_s1 ;
wire \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.facout_s2 ;
wire \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.fas_s1 ;
wire [1:0] \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.fas_s2 ;
wire \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.reset ;
wire [2:0] \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.s ;
wire \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.u1.a ;
wire \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.u1.b ;
wire \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.u1.cin ;
wire \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.u1.cout ;
wire \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.u1.s ;
wire [1:0] \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.u2.a ;
wire [1:0] \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.u2.b ;
wire \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.u2.cin ;
wire \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.u2.cout ;
wire [1:0] \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.u2.s ;
wire \add_3s_3ns_3_2_1_U13.ce ;
wire \add_3s_3ns_3_2_1_U13.clk ;
wire [2:0] \add_3s_3ns_3_2_1_U13.din0 ;
wire [2:0] \add_3s_3ns_3_2_1_U13.din1 ;
wire [2:0] \add_3s_3ns_3_2_1_U13.dout ;
wire \add_3s_3ns_3_2_1_U13.reset ;
wire [2:0] \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_6_U.a ;
wire [2:0] \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_6_U.ain_s0 ;
wire [2:0] \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_6_U.b ;
wire [2:0] \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_6_U.bin_s0 ;
wire \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_6_U.ce ;
wire \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_6_U.clk ;
wire \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_6_U.facout_s1 ;
wire \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_6_U.facout_s2 ;
wire \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_6_U.fas_s1 ;
wire [1:0] \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_6_U.fas_s2 ;
wire \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_6_U.reset ;
wire [2:0] \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_6_U.s ;
wire \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_6_U.u1.a ;
wire \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_6_U.u1.b ;
wire \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_6_U.u1.cin ;
wire \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_6_U.u1.cout ;
wire \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_6_U.u1.s ;
wire [1:0] \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_6_U.u2.a ;
wire [1:0] \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_6_U.u2.b ;
wire \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_6_U.u2.cin ;
wire \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_6_U.u2.cout ;
wire [1:0] \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_6_U.u2.s ;
wire \add_9ns_9ns_9_2_1_U5.ce ;
wire \add_9ns_9ns_9_2_1_U5.clk ;
wire [8:0] \add_9ns_9ns_9_2_1_U5.din0 ;
wire [8:0] \add_9ns_9ns_9_2_1_U5.din1 ;
wire [8:0] \add_9ns_9ns_9_2_1_U5.dout ;
wire \add_9ns_9ns_9_2_1_U5.reset ;
wire [8:0] \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_3_U.a ;
wire [8:0] \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_3_U.ain_s0 ;
wire [8:0] \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_3_U.b ;
wire [8:0] \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_3_U.bin_s0 ;
wire \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_3_U.ce ;
wire \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_3_U.clk ;
wire \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_3_U.facout_s1 ;
wire \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_3_U.facout_s2 ;
wire [3:0] \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_3_U.fas_s1 ;
wire [4:0] \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_3_U.fas_s2 ;
wire \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_3_U.reset ;
wire [8:0] \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_3_U.s ;
wire [3:0] \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_3_U.u1.a ;
wire [3:0] \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_3_U.u1.b ;
wire \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_3_U.u1.cin ;
wire \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_3_U.u1.cout ;
wire [3:0] \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_3_U.u1.s ;
wire [4:0] \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_3_U.u2.a ;
wire [4:0] \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_3_U.u2.b ;
wire \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_3_U.u2.cin ;
wire \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_3_U.u2.cout ;
wire [4:0] \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_3_U.u2.s ;
wire \add_9s_9s_9_2_1_U2.ce ;
wire \add_9s_9s_9_2_1_U2.clk ;
wire [8:0] \add_9s_9s_9_2_1_U2.din0 ;
wire [8:0] \add_9s_9s_9_2_1_U2.din1 ;
wire [8:0] \add_9s_9s_9_2_1_U2.dout ;
wire \add_9s_9s_9_2_1_U2.reset ;
wire [8:0] \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_0_U.a ;
wire [8:0] \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_0_U.ain_s0 ;
wire [8:0] \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_0_U.b ;
wire [8:0] \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_0_U.bin_s0 ;
wire \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_0_U.ce ;
wire \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_0_U.clk ;
wire \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_0_U.facout_s1 ;
wire \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_0_U.facout_s2 ;
wire [3:0] \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_0_U.fas_s1 ;
wire [4:0] \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_0_U.fas_s2 ;
wire \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_0_U.reset ;
wire [8:0] \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_0_U.s ;
wire [3:0] \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_0_U.u1.a ;
wire [3:0] \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_0_U.u1.b ;
wire \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_0_U.u1.cin ;
wire \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_0_U.u1.cout ;
wire [3:0] \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_0_U.u1.s ;
wire [4:0] \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_0_U.u2.a ;
wire [4:0] \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_0_U.u2.b ;
wire \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_0_U.u2.cin ;
wire \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_0_U.u2.cout ;
wire [4:0] \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_0_U.u2.s ;
wire ap_CS_fsm_state1;
wire ap_CS_fsm_state10;
wire ap_CS_fsm_state11;
wire ap_CS_fsm_state12;
wire ap_CS_fsm_state13;
wire ap_CS_fsm_state14;
wire ap_CS_fsm_state15;
wire ap_CS_fsm_state16;
wire ap_CS_fsm_state17;
wire ap_CS_fsm_state18;
wire ap_CS_fsm_state19;
wire ap_CS_fsm_state2;
wire ap_CS_fsm_state20;
wire ap_CS_fsm_state21;
wire ap_CS_fsm_state22;
wire ap_CS_fsm_state23;
wire ap_CS_fsm_state24;
wire ap_CS_fsm_state25;
wire ap_CS_fsm_state26;
wire ap_CS_fsm_state27;
wire ap_CS_fsm_state28;
wire ap_CS_fsm_state29;
wire ap_CS_fsm_state30;
wire ap_CS_fsm_state8;
wire ap_CS_fsm_state9;
wire [29:0] ap_NS_fsm;
wire ap_clk;
wire ap_done;
wire ap_idle;
wire ap_ready;
wire ap_rst;
wire ap_start;
wire [1:0] grp_fu_192_p1;
wire [1:0] grp_fu_192_p2;
wire [8:0] grp_fu_220_p0;
wire [8:0] grp_fu_220_p1;
wire [8:0] grp_fu_220_p2;
wire [2:0] grp_fu_240_p0;
wire [2:0] grp_fu_240_p1;
wire [2:0] grp_fu_240_p2;
wire [31:0] grp_fu_250_p0;
wire [31:0] grp_fu_250_p2;
wire [8:0] grp_fu_259_p0;
wire [8:0] grp_fu_259_p2;
wire [31:0] grp_fu_267_p0;
wire [31:0] grp_fu_267_p2;
wire [33:0] grp_fu_287_p0;
wire [33:0] grp_fu_287_p1;
wire [33:0] grp_fu_287_p2;
wire [31:0] grp_fu_316_p2;
wire [2:0] grp_fu_381_p0;
wire [2:0] grp_fu_381_p2;
wire [1:0] grp_fu_386_p1;
wire [1:0] grp_fu_386_p2;
wire [31:0] grp_fu_391_p2;
wire [2:0] grp_fu_399_p0;
wire [2:0] grp_fu_399_p2;
wire [31:0] grp_fu_407_p0;
wire [31:0] grp_fu_407_p2;
wire [35:0] grp_fu_427_p0;
wire [35:0] grp_fu_427_p1;
wire [35:0] grp_fu_427_p2;
wire [31:0] grp_fu_453_p2;
wire [3:0] grp_fu_478_p0;
wire [7:0] grp_fu_478_p00;
wire [31:0] grp_fu_478_p3;
wire icmp_ln851_fu_437_p2;
wire icmp_ln890_fu_229_p2;
wire lhs_V_fu_179_p2;
wire \lshr_2ns_1ns_2_7_1_U1.ce ;
wire \lshr_2ns_1ns_2_7_1_U1.clk ;
wire [1:0] \lshr_2ns_1ns_2_7_1_U1.din0 ;
wire [1:0] \lshr_2ns_1ns_2_7_1_U1.din1 ;
wire \lshr_2ns_1ns_2_7_1_U1.din1_cast ;
wire \lshr_2ns_1ns_2_7_1_U1.din1_mask ;
wire [1:0] \lshr_2ns_1ns_2_7_1_U1.dout ;
wire \lshr_2ns_1ns_2_7_1_U1.reset ;
wire \mac_muladd_4ns_4s_32ns_32_4_1_U17.ce ;
wire \mac_muladd_4ns_4s_32ns_32_4_1_U17.clk ;
wire [3:0] \mac_muladd_4ns_4s_32ns_32_4_1_U17.din0 ;
wire [3:0] \mac_muladd_4ns_4s_32ns_32_4_1_U17.din1 ;
wire [31:0] \mac_muladd_4ns_4s_32ns_32_4_1_U17.din2 ;
wire [31:0] \mac_muladd_4ns_4s_32ns_32_4_1_U17.dout ;
wire \mac_muladd_4ns_4s_32ns_32_4_1_U17.reset ;
wire [24:0] \mac_muladd_4ns_4s_32ns_32_4_1_U17.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.a ;
wire [17:0] \mac_muladd_4ns_4s_32ns_32_4_1_U17.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.b ;
wire [47:0] \mac_muladd_4ns_4s_32ns_32_4_1_U17.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.c ;
wire \mac_muladd_4ns_4s_32ns_32_4_1_U17.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.ce ;
wire \mac_muladd_4ns_4s_32ns_32_4_1_U17.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.clk ;
wire [31:0] \mac_muladd_4ns_4s_32ns_32_4_1_U17.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.dout ;
wire [3:0] \mac_muladd_4ns_4s_32ns_32_4_1_U17.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.in0 ;
wire [3:0] \mac_muladd_4ns_4s_32ns_32_4_1_U17.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.in1 ;
wire [31:0] \mac_muladd_4ns_4s_32ns_32_4_1_U17.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.in2 ;
wire [42:0] \mac_muladd_4ns_4s_32ns_32_4_1_U17.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.m ;
wire [47:0] \mac_muladd_4ns_4s_32ns_32_4_1_U17.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.p ;
wire \mac_muladd_4ns_4s_32ns_32_4_1_U17.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.rst ;
wire [1:0] \mul_2ns_2ns_4_1_1_U8.din0 ;
wire [1:0] \mul_2ns_2ns_4_1_1_U8.din1 ;
wire [3:0] \mul_2ns_2ns_4_1_1_U8.dout ;
wire [1:0] \mul_2ns_2ns_4_1_1_U8.top_mul_2ns_2ns_4_1_1_Multiplier_0_U.a ;
wire [1:0] \mul_2ns_2ns_4_1_1_U8.top_mul_2ns_2ns_4_1_1_Multiplier_0_U.b ;
wire [3:0] \mul_2ns_2ns_4_1_1_U8.top_mul_2ns_2ns_4_1_1_Multiplier_0_U.p ;
wire [7:0] op_0;
wire [3:0] op_1;
wire [31:0] op_10;
wire [1:0] op_12;
wire op_13;
wire [31:0] op_14;
wire [1:0] op_16_V_fu_327_p2;
wire op_18;
wire [3:0] op_19;
wire [3:0] op_2;
wire [1:0] op_3;
wire [31:0] op_32;
wire op_32_ap_vld;
wire [15:0] op_4;
wire [1:0] op_5;
wire op_9_V_fu_207_p2;
wire p_Result_1_fu_458_p3;
wire p_Result_s_fu_336_p3;
wire [3:0] r_fu_197_p2;
wire [1:0] ret_1_fu_306_p0;
wire [1:0] ret_1_fu_306_p1;
wire [3:0] ret_1_fu_306_p2;
wire [31:0] ret_V_5_fu_352_p3;
wire [32:0] rhs_1_fu_276_p3;
wire [34:0] rhs_3_fu_416_p3;
wire [1:0] select_ln69_1_fu_367_p3;
wire [2:0] select_ln69_fu_359_p3;
wire [31:0] select_ln850_1_fu_465_p3;
wire [31:0] select_ln850_fu_346_p3;
wire [3:0] sext_ln703_1_fu_412_p0;
wire [1:0] sext_ln703_fu_272_p0;
wire [1:0] sext_ln874_1_fu_175_p0;
wire [2:0] sext_ln874_1_fu_175_p1;
wire [1:0] sext_ln874_fu_226_p0;
wire [3:0] sext_ln874_fu_226_p1;
wire [1:0] trunc_ln1350_fu_312_p1;
wire [1:0] trunc_ln213_1_fu_185_p0;
wire trunc_ln213_1_fu_185_p1;
wire trunc_ln213_fu_203_p1;
wire [3:0] trunc_ln851_1_fu_433_p0;
wire [2:0] trunc_ln851_1_fu_433_p1;
wire [1:0] trunc_ln851_fu_343_p0;
wire trunc_ln851_fu_343_p1;
wire xor_ln890_fu_331_p2;
wire [1:0] zext_ln11_fu_189_p1;
wire [3:0] zext_ln1345_fu_303_p1;
wire [2:0] zext_ln874_fu_171_p1;


assign _034_ = icmp_ln851_reg_740 & ap_CS_fsm[28];
assign _035_ = _037_ & ap_CS_fsm[0];
assign _036_ = ap_start & ap_CS_fsm[0];
assign xor_ln890_fu_331_p2 = ~ icmp_ln890_reg_538;
assign r_fu_197_p2 = ~ op_2;
assign _037_ = ~ ap_start;
always @(posedge \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_7_U.clk )
\add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_7_U.bin_s1  <= _039_;
always @(posedge \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_7_U.clk )
\add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_7_U.ain_s1  <= _038_;
always @(posedge \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_7_U.clk )
\add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_7_U.sum_s1  <= _041_;
always @(posedge \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_7_U.clk )
\add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_7_U.carry_s1  <= _040_;
assign _039_ = \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_7_U.ce  ? \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_7_U.b [1] : \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_7_U.bin_s1 ;
assign _038_ = \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_7_U.ce  ? \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_7_U.a [1] : \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_7_U.ain_s1 ;
assign _040_ = \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_7_U.ce  ? \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_7_U.facout_s1  : \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_7_U.carry_s1 ;
assign _041_ = \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_7_U.ce  ? \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_7_U.fas_s1  : \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_7_U.sum_s1 ;
assign _042_ = \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_7_U.u1.a  + \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_7_U.u1.b ;
assign { \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_7_U.u1.cout , \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_7_U.u1.s  } = _042_ + \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_7_U.u1.cin ;
assign _043_ = \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_7_U.u2.a  + \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_7_U.u2.b ;
assign { \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_7_U.u2.cout , \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_7_U.u2.s  } = _043_ + \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_7_U.u2.cin ;
always @(posedge \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_2_U.clk )
\add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_2_U.bin_s1  <= _045_;
always @(posedge \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_2_U.clk )
\add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_2_U.ain_s1  <= _044_;
always @(posedge \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_2_U.clk )
\add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_2_U.sum_s1  <= _047_;
always @(posedge \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_2_U.clk )
\add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_2_U.carry_s1  <= _046_;
assign _045_ = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_2_U.ce  ? \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_2_U.b [31:16] : \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_2_U.bin_s1 ;
assign _044_ = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_2_U.ce  ? \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_2_U.a [31:16] : \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_2_U.ain_s1 ;
assign _046_ = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_2_U.ce  ? \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_2_U.facout_s1  : \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_2_U.carry_s1 ;
assign _047_ = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_2_U.ce  ? \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_2_U.fas_s1  : \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_2_U.sum_s1 ;
assign _048_ = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_2_U.u1.a  + \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_2_U.u1.b ;
assign { \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_2_U.u1.cout , \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_2_U.u1.s  } = _048_ + \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_2_U.u1.cin ;
assign _049_ = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_2_U.u2.a  + \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_2_U.u2.b ;
assign { \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_2_U.u2.cout , \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_2_U.u2.s  } = _049_ + \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_2_U.u2.cin ;
always @(posedge \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_2_U.clk )
\add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_2_U.bin_s1  <= _051_;
always @(posedge \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_2_U.clk )
\add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_2_U.ain_s1  <= _050_;
always @(posedge \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_2_U.clk )
\add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_2_U.sum_s1  <= _053_;
always @(posedge \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_2_U.clk )
\add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_2_U.carry_s1  <= _052_;
assign _051_ = \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_2_U.ce  ? \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_2_U.b [31:16] : \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_2_U.bin_s1 ;
assign _050_ = \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_2_U.ce  ? \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_2_U.a [31:16] : \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_2_U.ain_s1 ;
assign _052_ = \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_2_U.ce  ? \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_2_U.facout_s1  : \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_2_U.carry_s1 ;
assign _053_ = \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_2_U.ce  ? \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_2_U.fas_s1  : \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_2_U.sum_s1 ;
assign _054_ = \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_2_U.u1.a  + \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_2_U.u1.b ;
assign { \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_2_U.u1.cout , \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_2_U.u1.s  } = _054_ + \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_2_U.u1.cin ;
assign _055_ = \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_2_U.u2.a  + \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_2_U.u2.b ;
assign { \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_2_U.u2.cout , \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_2_U.u2.s  } = _055_ + \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_2_U.u2.cin ;
always @(posedge \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_2_U.clk )
\add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_2_U.bin_s1  <= _057_;
always @(posedge \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_2_U.clk )
\add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_2_U.ain_s1  <= _056_;
always @(posedge \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_2_U.clk )
\add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_2_U.sum_s1  <= _059_;
always @(posedge \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_2_U.clk )
\add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_2_U.carry_s1  <= _058_;
assign _057_ = \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_2_U.ce  ? \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_2_U.b [31:16] : \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_2_U.bin_s1 ;
assign _056_ = \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_2_U.ce  ? \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_2_U.a [31:16] : \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_2_U.ain_s1 ;
assign _058_ = \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_2_U.ce  ? \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_2_U.facout_s1  : \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_2_U.carry_s1 ;
assign _059_ = \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_2_U.ce  ? \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_2_U.fas_s1  : \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_2_U.sum_s1 ;
assign _060_ = \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_2_U.u1.a  + \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_2_U.u1.b ;
assign { \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_2_U.u1.cout , \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_2_U.u1.s  } = _060_ + \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_2_U.u1.cin ;
assign _061_ = \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_2_U.u2.a  + \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_2_U.u2.b ;
assign { \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_2_U.u2.cout , \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_2_U.u2.s  } = _061_ + \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_2_U.u2.cin ;
always @(posedge \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_4_U.clk )
\add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_4_U.bin_s1  <= _063_;
always @(posedge \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_4_U.clk )
\add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_4_U.ain_s1  <= _062_;
always @(posedge \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_4_U.clk )
\add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_4_U.sum_s1  <= _065_;
always @(posedge \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_4_U.clk )
\add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_4_U.carry_s1  <= _064_;
assign _063_ = \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_4_U.ce  ? \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_4_U.b [31:16] : \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_4_U.bin_s1 ;
assign _062_ = \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_4_U.ce  ? \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_4_U.a [31:16] : \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_4_U.ain_s1 ;
assign _064_ = \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_4_U.ce  ? \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_4_U.facout_s1  : \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_4_U.carry_s1 ;
assign _065_ = \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_4_U.ce  ? \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_4_U.fas_s1  : \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_4_U.sum_s1 ;
assign _066_ = \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_4_U.u1.a  + \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_4_U.u1.b ;
assign { \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_4_U.u1.cout , \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_4_U.u1.s  } = _066_ + \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_4_U.u1.cin ;
assign _067_ = \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_4_U.u2.a  + \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_4_U.u2.b ;
assign { \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_4_U.u2.cout , \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_4_U.u2.s  } = _067_ + \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_4_U.u2.cin ;
always @(posedge \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_4_U.clk )
\add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_4_U.bin_s1  <= _069_;
always @(posedge \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_4_U.clk )
\add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_4_U.ain_s1  <= _068_;
always @(posedge \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_4_U.clk )
\add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_4_U.sum_s1  <= _071_;
always @(posedge \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_4_U.clk )
\add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_4_U.carry_s1  <= _070_;
assign _069_ = \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_4_U.ce  ? \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_4_U.b [31:16] : \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_4_U.bin_s1 ;
assign _068_ = \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_4_U.ce  ? \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_4_U.a [31:16] : \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_4_U.ain_s1 ;
assign _070_ = \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_4_U.ce  ? \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_4_U.facout_s1  : \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_4_U.carry_s1 ;
assign _071_ = \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_4_U.ce  ? \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_4_U.fas_s1  : \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_4_U.sum_s1 ;
assign _072_ = \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_4_U.u1.a  + \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_4_U.u1.b ;
assign { \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_4_U.u1.cout , \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_4_U.u1.s  } = _072_ + \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_4_U.u1.cin ;
assign _073_ = \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_4_U.u2.a  + \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_4_U.u2.b ;
assign { \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_4_U.u2.cout , \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_4_U.u2.s  } = _073_ + \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_4_U.u2.cin ;
always @(posedge \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_4_U.clk )
\add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_4_U.bin_s1  <= _075_;
always @(posedge \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_4_U.clk )
\add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_4_U.ain_s1  <= _074_;
always @(posedge \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_4_U.clk )
\add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_4_U.sum_s1  <= _077_;
always @(posedge \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_4_U.clk )
\add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_4_U.carry_s1  <= _076_;
assign _075_ = \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_4_U.ce  ? \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_4_U.b [31:16] : \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_4_U.bin_s1 ;
assign _074_ = \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_4_U.ce  ? \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_4_U.a [31:16] : \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_4_U.ain_s1 ;
assign _076_ = \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_4_U.ce  ? \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_4_U.facout_s1  : \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_4_U.carry_s1 ;
assign _077_ = \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_4_U.ce  ? \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_4_U.fas_s1  : \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_4_U.sum_s1 ;
assign _078_ = \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_4_U.u1.a  + \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_4_U.u1.b ;
assign { \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_4_U.u1.cout , \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_4_U.u1.s  } = _078_ + \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_4_U.u1.cin ;
assign _079_ = \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_4_U.u2.a  + \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_4_U.u2.b ;
assign { \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_4_U.u2.cout , \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_4_U.u2.s  } = _079_ + \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_4_U.u2.cin ;
always @(posedge \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_5_U.clk )
\add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_5_U.bin_s1  <= _081_;
always @(posedge \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_5_U.clk )
\add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_5_U.ain_s1  <= _080_;
always @(posedge \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_5_U.clk )
\add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_5_U.sum_s1  <= _083_;
always @(posedge \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_5_U.clk )
\add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_5_U.carry_s1  <= _082_;
assign _081_ = \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_5_U.ce  ? \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_5_U.b [33:17] : \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_5_U.bin_s1 ;
assign _080_ = \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_5_U.ce  ? \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_5_U.a [33:17] : \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_5_U.ain_s1 ;
assign _082_ = \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_5_U.ce  ? \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_5_U.facout_s1  : \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_5_U.carry_s1 ;
assign _083_ = \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_5_U.ce  ? \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_5_U.fas_s1  : \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_5_U.sum_s1 ;
assign _084_ = \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_5_U.u1.a  + \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_5_U.u1.b ;
assign { \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_5_U.u1.cout , \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_5_U.u1.s  } = _084_ + \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_5_U.u1.cin ;
assign _085_ = \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_5_U.u2.a  + \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_5_U.u2.b ;
assign { \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_5_U.u2.cout , \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_5_U.u2.s  } = _085_ + \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_5_U.u2.cin ;
always @(posedge \add_36s_36s_36_2_1_U15.top_add_36s_36s_36_2_1_Adder_8_U.clk )
\add_36s_36s_36_2_1_U15.top_add_36s_36s_36_2_1_Adder_8_U.bin_s1  <= _087_;
always @(posedge \add_36s_36s_36_2_1_U15.top_add_36s_36s_36_2_1_Adder_8_U.clk )
\add_36s_36s_36_2_1_U15.top_add_36s_36s_36_2_1_Adder_8_U.ain_s1  <= _086_;
always @(posedge \add_36s_36s_36_2_1_U15.top_add_36s_36s_36_2_1_Adder_8_U.clk )
\add_36s_36s_36_2_1_U15.top_add_36s_36s_36_2_1_Adder_8_U.sum_s1  <= _089_;
always @(posedge \add_36s_36s_36_2_1_U15.top_add_36s_36s_36_2_1_Adder_8_U.clk )
\add_36s_36s_36_2_1_U15.top_add_36s_36s_36_2_1_Adder_8_U.carry_s1  <= _088_;
assign _087_ = \add_36s_36s_36_2_1_U15.top_add_36s_36s_36_2_1_Adder_8_U.ce  ? \add_36s_36s_36_2_1_U15.top_add_36s_36s_36_2_1_Adder_8_U.b [35:18] : \add_36s_36s_36_2_1_U15.top_add_36s_36s_36_2_1_Adder_8_U.bin_s1 ;
assign _086_ = \add_36s_36s_36_2_1_U15.top_add_36s_36s_36_2_1_Adder_8_U.ce  ? \add_36s_36s_36_2_1_U15.top_add_36s_36s_36_2_1_Adder_8_U.a [35:18] : \add_36s_36s_36_2_1_U15.top_add_36s_36s_36_2_1_Adder_8_U.ain_s1 ;
assign _088_ = \add_36s_36s_36_2_1_U15.top_add_36s_36s_36_2_1_Adder_8_U.ce  ? \add_36s_36s_36_2_1_U15.top_add_36s_36s_36_2_1_Adder_8_U.facout_s1  : \add_36s_36s_36_2_1_U15.top_add_36s_36s_36_2_1_Adder_8_U.carry_s1 ;
assign _089_ = \add_36s_36s_36_2_1_U15.top_add_36s_36s_36_2_1_Adder_8_U.ce  ? \add_36s_36s_36_2_1_U15.top_add_36s_36s_36_2_1_Adder_8_U.fas_s1  : \add_36s_36s_36_2_1_U15.top_add_36s_36s_36_2_1_Adder_8_U.sum_s1 ;
assign _090_ = \add_36s_36s_36_2_1_U15.top_add_36s_36s_36_2_1_Adder_8_U.u1.a  + \add_36s_36s_36_2_1_U15.top_add_36s_36s_36_2_1_Adder_8_U.u1.b ;
assign { \add_36s_36s_36_2_1_U15.top_add_36s_36s_36_2_1_Adder_8_U.u1.cout , \add_36s_36s_36_2_1_U15.top_add_36s_36s_36_2_1_Adder_8_U.u1.s  } = _090_ + \add_36s_36s_36_2_1_U15.top_add_36s_36s_36_2_1_Adder_8_U.u1.cin ;
assign _091_ = \add_36s_36s_36_2_1_U15.top_add_36s_36s_36_2_1_Adder_8_U.u2.a  + \add_36s_36s_36_2_1_U15.top_add_36s_36s_36_2_1_Adder_8_U.u2.b ;
assign { \add_36s_36s_36_2_1_U15.top_add_36s_36s_36_2_1_Adder_8_U.u2.cout , \add_36s_36s_36_2_1_U15.top_add_36s_36s_36_2_1_Adder_8_U.u2.s  } = _091_ + \add_36s_36s_36_2_1_U15.top_add_36s_36s_36_2_1_Adder_8_U.u2.cin ;
always @(posedge \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_1_U.clk )
\add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_1_U.bin_s1  <= _093_;
always @(posedge \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_1_U.clk )
\add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_1_U.ain_s1  <= _092_;
always @(posedge \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_1_U.clk )
\add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_1_U.sum_s1  <= _095_;
always @(posedge \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_1_U.clk )
\add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_1_U.carry_s1  <= _094_;
assign _093_ = \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_1_U.ce  ? \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_1_U.b [2:1] : \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_1_U.bin_s1 ;
assign _092_ = \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_1_U.ce  ? \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_1_U.a [2:1] : \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_1_U.ain_s1 ;
assign _094_ = \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_1_U.ce  ? \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_1_U.facout_s1  : \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_1_U.carry_s1 ;
assign _095_ = \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_1_U.ce  ? \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_1_U.fas_s1  : \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_1_U.sum_s1 ;
assign _096_ = \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_1_U.u1.a  + \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_1_U.u1.b ;
assign { \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_1_U.u1.cout , \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_1_U.u1.s  } = _096_ + \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_1_U.u1.cin ;
assign _097_ = \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_1_U.u2.a  + \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_1_U.u2.b ;
assign { \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_1_U.u2.cout , \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_1_U.u2.s  } = _097_ + \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_1_U.u2.cin ;
always @(posedge \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.clk )
\add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.bin_s1  <= _099_;
always @(posedge \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.clk )
\add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.ain_s1  <= _098_;
always @(posedge \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.clk )
\add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.sum_s1  <= _101_;
always @(posedge \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.clk )
\add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.carry_s1  <= _100_;
assign _099_ = \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.ce  ? \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.b [2:1] : \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.bin_s1 ;
assign _098_ = \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.ce  ? \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.a [2:1] : \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.ain_s1 ;
assign _100_ = \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.ce  ? \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.facout_s1  : \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.carry_s1 ;
assign _101_ = \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.ce  ? \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.fas_s1  : \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.sum_s1 ;
assign _102_ = \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.u1.a  + \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.u1.b ;
assign { \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.u1.cout , \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.u1.s  } = _102_ + \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.u1.cin ;
assign _103_ = \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.u2.a  + \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.u2.b ;
assign { \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.u2.cout , \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.u2.s  } = _103_ + \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.u2.cin ;
always @(posedge \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_6_U.clk )
\add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_6_U.bin_s1  <= _105_;
always @(posedge \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_6_U.clk )
\add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_6_U.ain_s1  <= _104_;
always @(posedge \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_6_U.clk )
\add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_6_U.sum_s1  <= _107_;
always @(posedge \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_6_U.clk )
\add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_6_U.carry_s1  <= _106_;
assign _105_ = \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_6_U.ce  ? \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_6_U.b [2:1] : \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_6_U.bin_s1 ;
assign _104_ = \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_6_U.ce  ? \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_6_U.a [2:1] : \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_6_U.ain_s1 ;
assign _106_ = \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_6_U.ce  ? \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_6_U.facout_s1  : \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_6_U.carry_s1 ;
assign _107_ = \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_6_U.ce  ? \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_6_U.fas_s1  : \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_6_U.sum_s1 ;
assign _108_ = \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_6_U.u1.a  + \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_6_U.u1.b ;
assign { \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_6_U.u1.cout , \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_6_U.u1.s  } = _108_ + \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_6_U.u1.cin ;
assign _109_ = \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_6_U.u2.a  + \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_6_U.u2.b ;
assign { \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_6_U.u2.cout , \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_6_U.u2.s  } = _109_ + \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_6_U.u2.cin ;
always @(posedge \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_3_U.clk )
\add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_3_U.bin_s1  <= _111_;
always @(posedge \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_3_U.clk )
\add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_3_U.ain_s1  <= _110_;
always @(posedge \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_3_U.clk )
\add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_3_U.sum_s1  <= _113_;
always @(posedge \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_3_U.clk )
\add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_3_U.carry_s1  <= _112_;
assign _111_ = \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_3_U.ce  ? \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_3_U.b [8:4] : \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_3_U.bin_s1 ;
assign _110_ = \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_3_U.ce  ? \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_3_U.a [8:4] : \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_3_U.ain_s1 ;
assign _112_ = \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_3_U.ce  ? \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_3_U.facout_s1  : \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_3_U.carry_s1 ;
assign _113_ = \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_3_U.ce  ? \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_3_U.fas_s1  : \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_3_U.sum_s1 ;
assign _114_ = \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_3_U.u1.a  + \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_3_U.u1.b ;
assign { \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_3_U.u1.cout , \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_3_U.u1.s  } = _114_ + \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_3_U.u1.cin ;
assign _115_ = \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_3_U.u2.a  + \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_3_U.u2.b ;
assign { \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_3_U.u2.cout , \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_3_U.u2.s  } = _115_ + \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_3_U.u2.cin ;
always @(posedge \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_0_U.clk )
\add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_0_U.bin_s1  <= _117_;
always @(posedge \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_0_U.clk )
\add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_0_U.ain_s1  <= _116_;
always @(posedge \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_0_U.clk )
\add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_0_U.sum_s1  <= _119_;
always @(posedge \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_0_U.clk )
\add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_0_U.carry_s1  <= _118_;
assign _117_ = \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_0_U.ce  ? \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_0_U.b [8:4] : \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_0_U.bin_s1 ;
assign _116_ = \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_0_U.ce  ? \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_0_U.a [8:4] : \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_0_U.ain_s1 ;
assign _118_ = \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_0_U.ce  ? \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_0_U.facout_s1  : \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_0_U.carry_s1 ;
assign _119_ = \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_0_U.ce  ? \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_0_U.fas_s1  : \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_0_U.sum_s1 ;
assign _120_ = \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_0_U.u1.a  + \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_0_U.u1.b ;
assign { \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_0_U.u1.cout , \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_0_U.u1.s  } = _120_ + \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_0_U.u1.cin ;
assign _121_ = \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_0_U.u2.a  + \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_0_U.u2.b ;
assign { \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_0_U.u2.cout , \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_0_U.u2.s  } = _121_ + \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_0_U.u2.cin ;
always @(posedge \lshr_2ns_1ns_2_7_1_U1.clk )
\lshr_2ns_1ns_2_7_1_U1.dout_array[5]  <= _133_;
always @(posedge \lshr_2ns_1ns_2_7_1_U1.clk )
\lshr_2ns_1ns_2_7_1_U1.din1_cast_array[5]  <= _127_;
always @(posedge \lshr_2ns_1ns_2_7_1_U1.clk )
\lshr_2ns_1ns_2_7_1_U1.dout_array[4]  <= _132_;
always @(posedge \lshr_2ns_1ns_2_7_1_U1.clk )
\lshr_2ns_1ns_2_7_1_U1.din1_cast_array[4]  <= _126_;
always @(posedge \lshr_2ns_1ns_2_7_1_U1.clk )
\lshr_2ns_1ns_2_7_1_U1.dout_array[3]  <= _131_;
always @(posedge \lshr_2ns_1ns_2_7_1_U1.clk )
\lshr_2ns_1ns_2_7_1_U1.din1_cast_array[3]  <= _125_;
always @(posedge \lshr_2ns_1ns_2_7_1_U1.clk )
\lshr_2ns_1ns_2_7_1_U1.dout_array[2]  <= _130_;
always @(posedge \lshr_2ns_1ns_2_7_1_U1.clk )
\lshr_2ns_1ns_2_7_1_U1.din1_cast_array[2]  <= _124_;
always @(posedge \lshr_2ns_1ns_2_7_1_U1.clk )
\lshr_2ns_1ns_2_7_1_U1.dout_array[1]  <= _129_;
always @(posedge \lshr_2ns_1ns_2_7_1_U1.clk )
\lshr_2ns_1ns_2_7_1_U1.din1_cast_array[1]  <= _123_;
always @(posedge \lshr_2ns_1ns_2_7_1_U1.clk )
\lshr_2ns_1ns_2_7_1_U1.dout_array[0]  <= _128_;
always @(posedge \lshr_2ns_1ns_2_7_1_U1.clk )
\lshr_2ns_1ns_2_7_1_U1.din1_cast_array[0]  <= _122_;
assign _134_ = \lshr_2ns_1ns_2_7_1_U1.ce  ? \lshr_2ns_1ns_2_7_1_U1.din1_cast_array[4]  : \lshr_2ns_1ns_2_7_1_U1.din1_cast_array[5] ;
assign _127_ = \lshr_2ns_1ns_2_7_1_U1.reset  ? 1'h0 : _134_;
assign _135_ = \lshr_2ns_1ns_2_7_1_U1.ce  ? \lshr_2ns_1ns_2_7_1_U1.dout_array[4]  : \lshr_2ns_1ns_2_7_1_U1.dout_array[5] ;
assign _133_ = \lshr_2ns_1ns_2_7_1_U1.reset  ? 2'h0 : _135_;
assign _136_ = \lshr_2ns_1ns_2_7_1_U1.ce  ? \lshr_2ns_1ns_2_7_1_U1.din1_cast_array[3]  : \lshr_2ns_1ns_2_7_1_U1.din1_cast_array[4] ;
assign _126_ = \lshr_2ns_1ns_2_7_1_U1.reset  ? 1'h0 : _136_;
assign _137_ = \lshr_2ns_1ns_2_7_1_U1.ce  ? \lshr_2ns_1ns_2_7_1_U1.dout_array[3]  : \lshr_2ns_1ns_2_7_1_U1.dout_array[4] ;
assign _132_ = \lshr_2ns_1ns_2_7_1_U1.reset  ? 2'h0 : _137_;
assign _138_ = \lshr_2ns_1ns_2_7_1_U1.ce  ? \lshr_2ns_1ns_2_7_1_U1.din1_cast_array[2]  : \lshr_2ns_1ns_2_7_1_U1.din1_cast_array[3] ;
assign _125_ = \lshr_2ns_1ns_2_7_1_U1.reset  ? 1'h0 : _138_;
assign _139_ = \lshr_2ns_1ns_2_7_1_U1.ce  ? \lshr_2ns_1ns_2_7_1_U1.dout_array[2]  : \lshr_2ns_1ns_2_7_1_U1.dout_array[3] ;
assign _131_ = \lshr_2ns_1ns_2_7_1_U1.reset  ? 2'h0 : _139_;
assign _140_ = \lshr_2ns_1ns_2_7_1_U1.ce  ? \lshr_2ns_1ns_2_7_1_U1.din1_cast_array[1]  : \lshr_2ns_1ns_2_7_1_U1.din1_cast_array[2] ;
assign _124_ = \lshr_2ns_1ns_2_7_1_U1.reset  ? 1'h0 : _140_;
assign _141_ = \lshr_2ns_1ns_2_7_1_U1.ce  ? \lshr_2ns_1ns_2_7_1_U1.dout_array[1]  : \lshr_2ns_1ns_2_7_1_U1.dout_array[2] ;
assign _130_ = \lshr_2ns_1ns_2_7_1_U1.reset  ? 2'h0 : _141_;
assign _142_ = \lshr_2ns_1ns_2_7_1_U1.ce  ? \lshr_2ns_1ns_2_7_1_U1.din1_cast_array[0]  : \lshr_2ns_1ns_2_7_1_U1.din1_cast_array[1] ;
assign _123_ = \lshr_2ns_1ns_2_7_1_U1.reset  ? 1'h0 : _142_;
assign _143_ = \lshr_2ns_1ns_2_7_1_U1.ce  ? \lshr_2ns_1ns_2_7_1_U1.dout_array[0]  : \lshr_2ns_1ns_2_7_1_U1.dout_array[1] ;
assign _129_ = \lshr_2ns_1ns_2_7_1_U1.reset  ? 2'h0 : _143_;
assign _144_ = \lshr_2ns_1ns_2_7_1_U1.ce  ? \lshr_2ns_1ns_2_7_1_U1.din1 [0] : \lshr_2ns_1ns_2_7_1_U1.din1_cast_array[0] ;
assign _122_ = \lshr_2ns_1ns_2_7_1_U1.reset  ? 1'h0 : _144_;
assign _145_ = \lshr_2ns_1ns_2_7_1_U1.ce  ? \lshr_2ns_1ns_2_7_1_U1.din0  : \lshr_2ns_1ns_2_7_1_U1.dout_array[0] ;
assign _128_ = \lshr_2ns_1ns_2_7_1_U1.reset  ? 2'h0 : _145_;
assign \lshr_2ns_1ns_2_7_1_U1.dout  = \lshr_2ns_1ns_2_7_1_U1.dout_array[5]  >> \lshr_2ns_1ns_2_7_1_U1.din1_cast_array[5] ;
assign { \mac_muladd_4ns_4s_32ns_32_4_1_U17.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.p [47], \mac_muladd_4ns_4s_32ns_32_4_1_U17.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.p [42:0] } = $signed(\mac_muladd_4ns_4s_32ns_32_4_1_U17.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.m_reg ) + $signed({ 1'h0, \mac_muladd_4ns_4s_32ns_32_4_1_U17.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.in2  });
assign \mac_muladd_4ns_4s_32ns_32_4_1_U17.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.m  = $signed(\mac_muladd_4ns_4s_32ns_32_4_1_U17.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.a_reg ) * $signed(\mac_muladd_4ns_4s_32ns_32_4_1_U17.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.b_reg );
always @(posedge \mac_muladd_4ns_4s_32ns_32_4_1_U17.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.clk )
\mac_muladd_4ns_4s_32ns_32_4_1_U17.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.m_reg  <= _148_;
always @(posedge \mac_muladd_4ns_4s_32ns_32_4_1_U17.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.clk )
\mac_muladd_4ns_4s_32ns_32_4_1_U17.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.a_reg  <= _146_;
always @(posedge \mac_muladd_4ns_4s_32ns_32_4_1_U17.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.clk )
\mac_muladd_4ns_4s_32ns_32_4_1_U17.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.b_reg  <= _147_;
always @(posedge \mac_muladd_4ns_4s_32ns_32_4_1_U17.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.clk )
\mac_muladd_4ns_4s_32ns_32_4_1_U17.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.p_reg  <= _149_;
assign _149_ = \mac_muladd_4ns_4s_32ns_32_4_1_U17.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.ce  ? { \mac_muladd_4ns_4s_32ns_32_4_1_U17.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.p [47], \mac_muladd_4ns_4s_32ns_32_4_1_U17.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.p [47], \mac_muladd_4ns_4s_32ns_32_4_1_U17.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.p [47], \mac_muladd_4ns_4s_32ns_32_4_1_U17.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.p [47], \mac_muladd_4ns_4s_32ns_32_4_1_U17.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.p [47], \mac_muladd_4ns_4s_32ns_32_4_1_U17.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.p [42:0] } : \mac_muladd_4ns_4s_32ns_32_4_1_U17.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.p_reg ;
assign _147_ = \mac_muladd_4ns_4s_32ns_32_4_1_U17.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.ce  ? { \mac_muladd_4ns_4s_32ns_32_4_1_U17.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.in1 [3], \mac_muladd_4ns_4s_32ns_32_4_1_U17.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.in1 [3], \mac_muladd_4ns_4s_32ns_32_4_1_U17.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.in1 [3], \mac_muladd_4ns_4s_32ns_32_4_1_U17.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.in1 [3], \mac_muladd_4ns_4s_32ns_32_4_1_U17.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.in1 [3], \mac_muladd_4ns_4s_32ns_32_4_1_U17.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.in1 [3], \mac_muladd_4ns_4s_32ns_32_4_1_U17.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.in1 [3], \mac_muladd_4ns_4s_32ns_32_4_1_U17.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.in1 [3], \mac_muladd_4ns_4s_32ns_32_4_1_U17.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.in1 [3], \mac_muladd_4ns_4s_32ns_32_4_1_U17.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.in1 [3], \mac_muladd_4ns_4s_32ns_32_4_1_U17.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.in1 [3], \mac_muladd_4ns_4s_32ns_32_4_1_U17.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.in1 [3], \mac_muladd_4ns_4s_32ns_32_4_1_U17.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.in1 [3], \mac_muladd_4ns_4s_32ns_32_4_1_U17.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.in1 [3], \mac_muladd_4ns_4s_32ns_32_4_1_U17.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.in1  } : \mac_muladd_4ns_4s_32ns_32_4_1_U17.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.b_reg ;
assign _146_ = \mac_muladd_4ns_4s_32ns_32_4_1_U17.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.ce  ? { 21'h000000, \mac_muladd_4ns_4s_32ns_32_4_1_U17.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.in0  } : \mac_muladd_4ns_4s_32ns_32_4_1_U17.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.a_reg ;
assign _148_ = \mac_muladd_4ns_4s_32ns_32_4_1_U17.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.ce  ? \mac_muladd_4ns_4s_32ns_32_4_1_U17.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.m  : \mac_muladd_4ns_4s_32ns_32_4_1_U17.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.m_reg ;
assign \mul_2ns_2ns_4_1_1_U8.top_mul_2ns_2ns_4_1_1_Multiplier_0_U.p  = \mul_2ns_2ns_4_1_1_U8.top_mul_2ns_2ns_4_1_1_Multiplier_0_U.a  * \mul_2ns_2ns_4_1_1_U8.top_mul_2ns_2ns_4_1_1_Multiplier_0_U.b ;
assign _150_ = $signed(r_reg_512) < $signed(op_5);
assign _151_ = | op_19[2:0];
assign _152_ = op_3 != { op_5[1], op_5 };
always @(posedge ap_clk)
zext_ln11_reg_506[1] <= 1'h0;
always @(posedge ap_clk)
zext_ln11_reg_506[0] <= _032_;
always @(posedge ap_clk)
xor_ln890_reg_655 <= _031_;
always @(posedge ap_clk)
ret_V_5_reg_660 <= _023_;
always @(posedge ap_clk)
select_ln69_reg_665 <= _028_;
always @(posedge ap_clk)
select_ln69_1_reg_670 <= _027_;
always @(posedge ap_clk)
ret_V_4_reg_613 <= _022_;
always @(posedge ap_clk)
ret_V_cast_reg_618 <= _025_;
always @(posedge ap_clk)
ret_V_6_reg_745 <= _024_;
always @(posedge ap_clk)
ret_V_3_cast_reg_750 <= _021_;
always @(posedge ap_clk)
ret_1_reg_625 <= _020_;
always @(posedge ap_clk)
trunc_ln1350_reg_630 <= _029_;
always @(posedge ap_clk)
r_reg_512 <= _019_;
always @(posedge ap_clk)
op_9_V_reg_518 <= _017_;
always @(posedge ap_clk)
r_1_reg_523 <= _018_;
always @(posedge ap_clk)
op_31_V_reg_725 <= _016_;
always @(posedge ap_clk)
op_24_V_reg_593 <= _015_;
always @(posedge ap_clk)
lhs_V_reg_496 <= _013_;
always @(posedge ap_clk)
trunc_ln213_1_reg_501 <= _030_;
always @(posedge ap_clk)
icmp_ln890_reg_538 <= _012_;
always @(posedge ap_clk)
icmp_ln851_reg_740 <= _011_;
always @(posedge ap_clk)
add_ln69_5_reg_710 <= _005_;
always @(posedge ap_clk)
add_ln69_8_reg_715 <= _008_;
always @(posedge ap_clk)
add_ln69_4_reg_685 <= _004_;
always @(posedge ap_clk)
add_ln69_6_reg_690 <= _006_;
always @(posedge ap_clk)
add_ln69_7_reg_695 <= _007_;
always @(posedge ap_clk)
add_ln69_reg_578 <= _009_;
always @(posedge ap_clk)
add_ln69_2_reg_583 <= _003_;
always @(posedge ap_clk)
ret_reg_553 <= _026_;
always @(posedge ap_clk)
add_ln69_1_reg_558 <= _002_;
always @(posedge ap_clk)
op_16_V_reg_645 <= _014_;
always @(posedge ap_clk)
add_ln691_reg_650 <= _001_;
always @(posedge ap_clk)
add_ln691_1_reg_757 <= _000_;
always @(posedge ap_clk)
ap_CS_fsm <= _010_;
assign _033_ = _036_ ? 2'h2 : 2'h1;
assign _153_ = ap_CS_fsm == 1'h1;
function [29:0] _444_;
input [29:0] a;
input [899:0] b;
input [29:0] s;
case (s)
30'b000000000000000000000000000001:
_444_ = b[29:0];
30'b000000000000000000000000000010:
_444_ = b[59:30];
30'b000000000000000000000000000100:
_444_ = b[89:60];
30'b000000000000000000000000001000:
_444_ = b[119:90];
30'b000000000000000000000000010000:
_444_ = b[149:120];
30'b000000000000000000000000100000:
_444_ = b[179:150];
30'b000000000000000000000001000000:
_444_ = b[209:180];
30'b000000000000000000000010000000:
_444_ = b[239:210];
30'b000000000000000000000100000000:
_444_ = b[269:240];
30'b000000000000000000001000000000:
_444_ = b[299:270];
30'b000000000000000000010000000000:
_444_ = b[329:300];
30'b000000000000000000100000000000:
_444_ = b[359:330];
30'b000000000000000001000000000000:
_444_ = b[389:360];
30'b000000000000000010000000000000:
_444_ = b[419:390];
30'b000000000000000100000000000000:
_444_ = b[449:420];
30'b000000000000001000000000000000:
_444_ = b[479:450];
30'b000000000000010000000000000000:
_444_ = b[509:480];
30'b000000000000100000000000000000:
_444_ = b[539:510];
30'b000000000001000000000000000000:
_444_ = b[569:540];
30'b000000000010000000000000000000:
_444_ = b[599:570];
30'b000000000100000000000000000000:
_444_ = b[629:600];
30'b000000001000000000000000000000:
_444_ = b[659:630];
30'b000000010000000000000000000000:
_444_ = b[689:660];
30'b000000100000000000000000000000:
_444_ = b[719:690];
30'b000001000000000000000000000000:
_444_ = b[749:720];
30'b000010000000000000000000000000:
_444_ = b[779:750];
30'b000100000000000000000000000000:
_444_ = b[809:780];
30'b001000000000000000000000000000:
_444_ = b[839:810];
30'b010000000000000000000000000000:
_444_ = b[869:840];
30'b100000000000000000000000000000:
_444_ = b[899:870];
30'b000000000000000000000000000000:
_444_ = a;
default:
_444_ = 30'bx;
endcase
endfunction
assign ap_NS_fsm = _444_(30'hxxxxxxxx, { 28'h0000000, _033_, 870'h00000004000000200000010000000800000040000002000000100000008000000400000020000001000000080000004000000200000010000000800000040000002000000100000008000000400000020000001000000080000004000000200000010000000800000000000001 }, { _153_, _182_, _181_, _180_, _179_, _178_, _177_, _176_, _175_, _174_, _173_, _172_, _171_, _170_, _169_, _168_, _167_, _166_, _165_, _164_, _163_, _162_, _161_, _160_, _159_, _158_, _157_, _156_, _155_, _154_ });
assign _154_ = ap_CS_fsm == 30'h20000000;
assign _155_ = ap_CS_fsm == 29'h10000000;
assign _156_ = ap_CS_fsm == 28'h8000000;
assign _157_ = ap_CS_fsm == 27'h4000000;
assign _158_ = ap_CS_fsm == 26'h2000000;
assign _159_ = ap_CS_fsm == 25'h1000000;
assign _160_ = ap_CS_fsm == 24'h800000;
assign _161_ = ap_CS_fsm == 23'h400000;
assign _162_ = ap_CS_fsm == 22'h200000;
assign _163_ = ap_CS_fsm == 21'h100000;
assign _164_ = ap_CS_fsm == 20'h80000;
assign _165_ = ap_CS_fsm == 19'h40000;
assign _166_ = ap_CS_fsm == 18'h20000;
assign _167_ = ap_CS_fsm == 17'h10000;
assign _168_ = ap_CS_fsm == 16'h8000;
assign _169_ = ap_CS_fsm == 15'h4000;
assign _170_ = ap_CS_fsm == 14'h2000;
assign _171_ = ap_CS_fsm == 13'h1000;
assign _172_ = ap_CS_fsm == 12'h800;
assign _173_ = ap_CS_fsm == 11'h400;
assign _174_ = ap_CS_fsm == 10'h200;
assign _175_ = ap_CS_fsm == 9'h100;
assign _176_ = ap_CS_fsm == 8'h80;
assign _177_ = ap_CS_fsm == 7'h40;
assign _178_ = ap_CS_fsm == 6'h20;
assign _179_ = ap_CS_fsm == 5'h10;
assign _180_ = ap_CS_fsm == 4'h8;
assign _181_ = ap_CS_fsm == 3'h4;
assign _182_ = ap_CS_fsm == 2'h2;
assign op_32_ap_vld = ap_CS_fsm[29] ? 1'h1 : 1'h0;
assign ap_idle = _035_ ? 1'h1 : 1'h0;
assign _032_ = ap_CS_fsm[1] ? lhs_V_reg_496 : zext_ln11_reg_506[0];
assign _027_ = ap_CS_fsm[18] ? select_ln69_1_fu_367_p3 : select_ln69_1_reg_670;
assign _028_ = ap_CS_fsm[18] ? select_ln69_fu_359_p3 : select_ln69_reg_665;
assign _023_ = ap_CS_fsm[18] ? ret_V_5_fu_352_p3 : ret_V_5_reg_660;
assign _031_ = ap_CS_fsm[18] ? xor_ln890_fu_331_p2 : xor_ln890_reg_655;
assign _025_ = ap_CS_fsm[15] ? grp_fu_287_p2[32:1] : ret_V_cast_reg_618;
assign _022_ = ap_CS_fsm[15] ? grp_fu_287_p2 : ret_V_4_reg_613;
assign _021_ = ap_CS_fsm[26] ? grp_fu_427_p2[34:3] : ret_V_3_cast_reg_750;
assign _024_ = ap_CS_fsm[26] ? grp_fu_427_p2 : ret_V_6_reg_745;
assign _029_ = ap_CS_fsm[16] ? ret_1_fu_306_p2[1:0] : trunc_ln1350_reg_630;
assign _020_ = ap_CS_fsm[16] ? ret_1_fu_306_p2 : ret_1_reg_625;
assign _018_ = ap_CS_fsm[7] ? grp_fu_192_p2 : r_1_reg_523;
assign _017_ = ap_CS_fsm[7] ? op_9_V_fu_207_p2 : op_9_V_reg_518;
assign _019_ = ap_CS_fsm[7] ? r_fu_197_p2 : r_reg_512;
assign _016_ = ap_CS_fsm[24] ? grp_fu_407_p2 : op_31_V_reg_725;
assign _015_ = ap_CS_fsm[13] ? grp_fu_267_p2 : op_24_V_reg_593;
assign _030_ = ap_CS_fsm[0] ? op_5[0] : trunc_ln213_1_reg_501;
assign _013_ = ap_CS_fsm[0] ? lhs_V_fu_179_p2 : lhs_V_reg_496;
assign _012_ = ap_CS_fsm[8] ? icmp_ln890_fu_229_p2 : icmp_ln890_reg_538;
assign _011_ = ap_CS_fsm[25] ? icmp_ln851_fu_437_p2 : icmp_ln851_reg_740;
assign _008_ = ap_CS_fsm[22] ? grp_fu_399_p2 : add_ln69_8_reg_715;
assign _005_ = ap_CS_fsm[22] ? grp_fu_391_p2 : add_ln69_5_reg_710;
assign _007_ = ap_CS_fsm[20] ? grp_fu_386_p2 : add_ln69_7_reg_695;
assign _006_ = ap_CS_fsm[20] ? grp_fu_381_p2 : add_ln69_6_reg_690;
assign _004_ = ap_CS_fsm[20] ? grp_fu_478_p3 : add_ln69_4_reg_685;
assign _003_ = ap_CS_fsm[11] ? grp_fu_259_p2 : add_ln69_2_reg_583;
assign _009_ = ap_CS_fsm[11] ? grp_fu_250_p2 : add_ln69_reg_578;
assign _002_ = ap_CS_fsm[9] ? grp_fu_240_p2 : add_ln69_1_reg_558;
assign _026_ = ap_CS_fsm[9] ? grp_fu_220_p2 : ret_reg_553;
assign _001_ = ap_CS_fsm[17] ? grp_fu_316_p2 : add_ln691_reg_650;
assign _014_ = ap_CS_fsm[17] ? op_16_V_fu_327_p2 : op_16_V_reg_645;
assign _000_ = _034_ ? grp_fu_453_p2 : add_ln691_1_reg_757;
assign _010_ = ap_rst ? 30'h00000001 : ap_NS_fsm;
assign icmp_ln851_fu_437_p2 = _151_ ? 1'h1 : 1'h0;
assign icmp_ln890_fu_229_p2 = _150_ ? 1'h1 : 1'h0;
assign lhs_V_fu_179_p2 = _152_ ? 1'h1 : 1'h0;
assign op_32 = ret_V_6_reg_745[35] ? select_ln850_1_fu_465_p3 : ret_V_3_cast_reg_750;
assign ret_V_5_fu_352_p3 = ret_V_4_reg_613[33] ? select_ln850_fu_346_p3 : ret_V_cast_reg_618;
assign select_ln69_1_fu_367_p3 = op_18 ? 2'h3 : 2'h0;
assign select_ln69_fu_359_p3 = op_13 ? 3'h7 : 3'h0;
assign select_ln850_1_fu_465_p3 = icmp_ln851_reg_740 ? add_ln691_1_reg_757 : ret_V_3_cast_reg_750;
assign select_ln850_fu_346_p3 = op_12[0] ? add_ln691_reg_650 : ret_V_cast_reg_618;
assign op_16_V_fu_327_p2 = zext_ln11_reg_506 ^ trunc_ln1350_reg_630;
assign op_9_V_fu_207_p2 = op_2[0] ^ trunc_ln213_1_reg_501;
assign ap_CS_fsm_state1 = ap_CS_fsm[0];
assign ap_CS_fsm_state10 = ap_CS_fsm[9];
assign ap_CS_fsm_state11 = ap_CS_fsm[10];
assign ap_CS_fsm_state12 = ap_CS_fsm[11];
assign ap_CS_fsm_state13 = ap_CS_fsm[12];
assign ap_CS_fsm_state14 = ap_CS_fsm[13];
assign ap_CS_fsm_state15 = ap_CS_fsm[14];
assign ap_CS_fsm_state16 = ap_CS_fsm[15];
assign ap_CS_fsm_state17 = ap_CS_fsm[16];
assign ap_CS_fsm_state18 = ap_CS_fsm[17];
assign ap_CS_fsm_state19 = ap_CS_fsm[18];
assign ap_CS_fsm_state2 = ap_CS_fsm[1];
assign ap_CS_fsm_state20 = ap_CS_fsm[19];
assign ap_CS_fsm_state21 = ap_CS_fsm[20];
assign ap_CS_fsm_state22 = ap_CS_fsm[21];
assign ap_CS_fsm_state23 = ap_CS_fsm[22];
assign ap_CS_fsm_state24 = ap_CS_fsm[23];
assign ap_CS_fsm_state25 = ap_CS_fsm[24];
assign ap_CS_fsm_state26 = ap_CS_fsm[25];
assign ap_CS_fsm_state27 = ap_CS_fsm[26];
assign ap_CS_fsm_state28 = ap_CS_fsm[27];
assign ap_CS_fsm_state29 = ap_CS_fsm[28];
assign ap_CS_fsm_state30 = ap_CS_fsm[29];
assign ap_CS_fsm_state8 = ap_CS_fsm[7];
assign ap_CS_fsm_state9 = ap_CS_fsm[8];
assign ap_done = op_32_ap_vld;
assign ap_ready = op_32_ap_vld;
assign grp_fu_192_p1 = { 1'h0, lhs_V_reg_496 };
assign grp_fu_220_p0 = { op_0[7], op_0 };
assign grp_fu_220_p1 = { op_1[3], op_1[3], op_1[3], op_1[3], op_1[3], op_1 };
assign grp_fu_240_p0 = { 1'h0, r_1_reg_523 };
assign grp_fu_240_p1 = { 2'h0, op_9_V_reg_518 };
assign grp_fu_250_p0 = { 16'h0000, op_4 };
assign grp_fu_259_p0 = { 6'h00, add_ln69_1_reg_558 };
assign grp_fu_267_p0 = { add_ln69_2_reg_583[8], add_ln69_2_reg_583[8], add_ln69_2_reg_583[8], add_ln69_2_reg_583[8], add_ln69_2_reg_583[8], add_ln69_2_reg_583[8], add_ln69_2_reg_583[8], add_ln69_2_reg_583[8], add_ln69_2_reg_583[8], add_ln69_2_reg_583[8], add_ln69_2_reg_583[8], add_ln69_2_reg_583[8], add_ln69_2_reg_583[8], add_ln69_2_reg_583[8], add_ln69_2_reg_583[8], add_ln69_2_reg_583[8], add_ln69_2_reg_583[8], add_ln69_2_reg_583[8], add_ln69_2_reg_583[8], add_ln69_2_reg_583[8], add_ln69_2_reg_583[8], add_ln69_2_reg_583[8], add_ln69_2_reg_583[8], add_ln69_2_reg_583 };
assign grp_fu_287_p0 = { op_24_V_reg_593[31], op_24_V_reg_593, 1'h0 };
assign grp_fu_287_p1 = { op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12 };
assign grp_fu_381_p0 = { op_16_V_reg_645[1], op_16_V_reg_645 };
assign grp_fu_386_p1 = { 1'h0, xor_ln890_reg_655 };
assign grp_fu_399_p0 = { add_ln69_7_reg_695[1], add_ln69_7_reg_695 };
assign grp_fu_407_p0 = { add_ln69_8_reg_715[2], add_ln69_8_reg_715[2], add_ln69_8_reg_715[2], add_ln69_8_reg_715[2], add_ln69_8_reg_715[2], add_ln69_8_reg_715[2], add_ln69_8_reg_715[2], add_ln69_8_reg_715[2], add_ln69_8_reg_715[2], add_ln69_8_reg_715[2], add_ln69_8_reg_715[2], add_ln69_8_reg_715[2], add_ln69_8_reg_715[2], add_ln69_8_reg_715[2], add_ln69_8_reg_715[2], add_ln69_8_reg_715[2], add_ln69_8_reg_715[2], add_ln69_8_reg_715[2], add_ln69_8_reg_715[2], add_ln69_8_reg_715[2], add_ln69_8_reg_715[2], add_ln69_8_reg_715[2], add_ln69_8_reg_715[2], add_ln69_8_reg_715[2], add_ln69_8_reg_715[2], add_ln69_8_reg_715[2], add_ln69_8_reg_715[2], add_ln69_8_reg_715[2], add_ln69_8_reg_715[2], add_ln69_8_reg_715 };
assign grp_fu_427_p0 = { op_31_V_reg_725[31], op_31_V_reg_725, 3'h0 };
assign grp_fu_427_p1 = { op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19 };
assign grp_fu_478_p0 = ret_1_reg_625;
assign grp_fu_478_p00 = { 4'h0, ret_1_reg_625 };
assign p_Result_1_fu_458_p3 = ret_V_6_reg_745[35];
assign p_Result_s_fu_336_p3 = ret_V_4_reg_613[33];
assign ret_1_fu_306_p0 = op_3;
assign ret_1_fu_306_p1 = op_3;
assign rhs_1_fu_276_p3 = { op_24_V_reg_593, 1'h0 };
assign rhs_3_fu_416_p3 = { op_31_V_reg_725, 3'h0 };
assign sext_ln703_1_fu_412_p0 = op_19;
assign sext_ln703_fu_272_p0 = op_12;
assign sext_ln874_1_fu_175_p0 = op_5;
assign sext_ln874_1_fu_175_p1 = { op_5[1], op_5 };
assign sext_ln874_fu_226_p0 = op_5;
assign sext_ln874_fu_226_p1 = { op_5[1], op_5[1], op_5 };
assign trunc_ln1350_fu_312_p1 = ret_1_fu_306_p2[1:0];
assign trunc_ln213_1_fu_185_p0 = op_5;
assign trunc_ln213_1_fu_185_p1 = op_5[0];
assign trunc_ln213_fu_203_p1 = op_2[0];
assign trunc_ln851_1_fu_433_p0 = op_19;
assign trunc_ln851_1_fu_433_p1 = op_19[2:0];
assign trunc_ln851_fu_343_p0 = op_12;
assign trunc_ln851_fu_343_p1 = op_12[0];
assign zext_ln11_fu_189_p1 = { 1'h0, lhs_V_reg_496 };
assign zext_ln1345_fu_303_p1 = { 2'h0, op_3 };
assign zext_ln874_fu_171_p1 = { 1'h0, op_3 };
assign \mul_2ns_2ns_4_1_1_U8.top_mul_2ns_2ns_4_1_1_Multiplier_0_U.a  = \mul_2ns_2ns_4_1_1_U8.din0 ;
assign \mul_2ns_2ns_4_1_1_U8.top_mul_2ns_2ns_4_1_1_Multiplier_0_U.b  = \mul_2ns_2ns_4_1_1_U8.din1 ;
assign \mul_2ns_2ns_4_1_1_U8.dout  = \mul_2ns_2ns_4_1_1_U8.top_mul_2ns_2ns_4_1_1_Multiplier_0_U.p ;
assign \mul_2ns_2ns_4_1_1_U8.din0  = op_3;
assign \mul_2ns_2ns_4_1_1_U8.din1  = op_3;
assign ret_1_fu_306_p2 = \mul_2ns_2ns_4_1_1_U8.dout ;
assign \mac_muladd_4ns_4s_32ns_32_4_1_U17.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.a  = { 21'h000000, \mac_muladd_4ns_4s_32ns_32_4_1_U17.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.in0  };
assign \mac_muladd_4ns_4s_32ns_32_4_1_U17.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.b  = { \mac_muladd_4ns_4s_32ns_32_4_1_U17.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.in1 [3], \mac_muladd_4ns_4s_32ns_32_4_1_U17.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.in1 [3], \mac_muladd_4ns_4s_32ns_32_4_1_U17.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.in1 [3], \mac_muladd_4ns_4s_32ns_32_4_1_U17.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.in1 [3], \mac_muladd_4ns_4s_32ns_32_4_1_U17.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.in1 [3], \mac_muladd_4ns_4s_32ns_32_4_1_U17.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.in1 [3], \mac_muladd_4ns_4s_32ns_32_4_1_U17.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.in1 [3], \mac_muladd_4ns_4s_32ns_32_4_1_U17.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.in1 [3], \mac_muladd_4ns_4s_32ns_32_4_1_U17.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.in1 [3], \mac_muladd_4ns_4s_32ns_32_4_1_U17.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.in1 [3], \mac_muladd_4ns_4s_32ns_32_4_1_U17.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.in1 [3], \mac_muladd_4ns_4s_32ns_32_4_1_U17.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.in1 [3], \mac_muladd_4ns_4s_32ns_32_4_1_U17.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.in1 [3], \mac_muladd_4ns_4s_32ns_32_4_1_U17.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.in1 [3], \mac_muladd_4ns_4s_32ns_32_4_1_U17.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.in1  };
assign \mac_muladd_4ns_4s_32ns_32_4_1_U17.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.c  = { 16'h0000, \mac_muladd_4ns_4s_32ns_32_4_1_U17.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.in2  };
assign \mac_muladd_4ns_4s_32ns_32_4_1_U17.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.dout  = \mac_muladd_4ns_4s_32ns_32_4_1_U17.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.p_reg [31:0];
assign \mac_muladd_4ns_4s_32ns_32_4_1_U17.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.p [46:43] = { \mac_muladd_4ns_4s_32ns_32_4_1_U17.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.p [47], \mac_muladd_4ns_4s_32ns_32_4_1_U17.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.p [47], \mac_muladd_4ns_4s_32ns_32_4_1_U17.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.p [47], \mac_muladd_4ns_4s_32ns_32_4_1_U17.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.p [47] };
assign \mac_muladd_4ns_4s_32ns_32_4_1_U17.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.ce  = \mac_muladd_4ns_4s_32ns_32_4_1_U17.ce ;
assign \mac_muladd_4ns_4s_32ns_32_4_1_U17.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.clk  = \mac_muladd_4ns_4s_32ns_32_4_1_U17.clk ;
assign \mac_muladd_4ns_4s_32ns_32_4_1_U17.dout  = \mac_muladd_4ns_4s_32ns_32_4_1_U17.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.dout ;
assign \mac_muladd_4ns_4s_32ns_32_4_1_U17.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.in0  = \mac_muladd_4ns_4s_32ns_32_4_1_U17.din0 ;
assign \mac_muladd_4ns_4s_32ns_32_4_1_U17.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.in1  = \mac_muladd_4ns_4s_32ns_32_4_1_U17.din1 ;
assign \mac_muladd_4ns_4s_32ns_32_4_1_U17.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.in2  = \mac_muladd_4ns_4s_32ns_32_4_1_U17.din2 ;
assign \mac_muladd_4ns_4s_32ns_32_4_1_U17.top_mac_muladd_4ns_4s_32ns_32_4_1_DSP48_0_U.rst  = \mac_muladd_4ns_4s_32ns_32_4_1_U17.reset ;
assign \mac_muladd_4ns_4s_32ns_32_4_1_U17.ce  = 1'h1;
assign \mac_muladd_4ns_4s_32ns_32_4_1_U17.clk  = ap_clk;
assign \mac_muladd_4ns_4s_32ns_32_4_1_U17.din0  = ret_1_reg_625;
assign \mac_muladd_4ns_4s_32ns_32_4_1_U17.din1  = r_reg_512;
assign \mac_muladd_4ns_4s_32ns_32_4_1_U17.din2  = ret_V_5_reg_660;
assign grp_fu_478_p3 = \mac_muladd_4ns_4s_32ns_32_4_1_U17.dout ;
assign \mac_muladd_4ns_4s_32ns_32_4_1_U17.reset  = ap_rst;
assign \lshr_2ns_1ns_2_7_1_U1.din1_cast  = \lshr_2ns_1ns_2_7_1_U1.din1 [0];
assign \lshr_2ns_1ns_2_7_1_U1.din1_mask  = 1'h1;
assign \lshr_2ns_1ns_2_7_1_U1.ce  = 1'h1;
assign \lshr_2ns_1ns_2_7_1_U1.clk  = ap_clk;
assign \lshr_2ns_1ns_2_7_1_U1.din0  = op_3;
assign \lshr_2ns_1ns_2_7_1_U1.din1  = { 1'h0, lhs_V_reg_496 };
assign grp_fu_192_p2 = \lshr_2ns_1ns_2_7_1_U1.dout ;
assign \lshr_2ns_1ns_2_7_1_U1.reset  = ap_rst;
assign \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_0_U.ain_s0  = \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_0_U.a ;
assign \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_0_U.bin_s0  = \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_0_U.b ;
assign \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_0_U.s  = { \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_0_U.fas_s2 , \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_0_U.sum_s1  };
assign \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_0_U.u2.a  = \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_0_U.ain_s1 ;
assign \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_0_U.u2.b  = \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_0_U.bin_s1 ;
assign \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_0_U.u2.cin  = \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_0_U.carry_s1 ;
assign \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_0_U.facout_s2  = \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_0_U.u2.cout ;
assign \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_0_U.fas_s2  = \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_0_U.u2.s ;
assign \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_0_U.u1.a  = \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_0_U.a [3:0];
assign \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_0_U.u1.b  = \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_0_U.b [3:0];
assign \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_0_U.u1.cin  = 1'h0;
assign \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_0_U.facout_s1  = \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_0_U.u1.cout ;
assign \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_0_U.fas_s1  = \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_0_U.u1.s ;
assign \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_0_U.a  = \add_9s_9s_9_2_1_U2.din0 ;
assign \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_0_U.b  = \add_9s_9s_9_2_1_U2.din1 ;
assign \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_0_U.ce  = \add_9s_9s_9_2_1_U2.ce ;
assign \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_0_U.clk  = \add_9s_9s_9_2_1_U2.clk ;
assign \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_0_U.reset  = \add_9s_9s_9_2_1_U2.reset ;
assign \add_9s_9s_9_2_1_U2.dout  = \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_0_U.s ;
assign \add_9s_9s_9_2_1_U2.ce  = 1'h1;
assign \add_9s_9s_9_2_1_U2.clk  = ap_clk;
assign \add_9s_9s_9_2_1_U2.din0  = { op_0[7], op_0 };
assign \add_9s_9s_9_2_1_U2.din1  = { op_1[3], op_1[3], op_1[3], op_1[3], op_1[3], op_1 };
assign grp_fu_220_p2 = \add_9s_9s_9_2_1_U2.dout ;
assign \add_9s_9s_9_2_1_U2.reset  = ap_rst;
assign \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_3_U.ain_s0  = \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_3_U.a ;
assign \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_3_U.bin_s0  = \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_3_U.b ;
assign \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_3_U.s  = { \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_3_U.fas_s2 , \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_3_U.sum_s1  };
assign \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_3_U.u2.a  = \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_3_U.ain_s1 ;
assign \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_3_U.u2.b  = \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_3_U.bin_s1 ;
assign \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_3_U.u2.cin  = \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_3_U.carry_s1 ;
assign \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_3_U.facout_s2  = \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_3_U.u2.cout ;
assign \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_3_U.fas_s2  = \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_3_U.u2.s ;
assign \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_3_U.u1.a  = \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_3_U.a [3:0];
assign \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_3_U.u1.b  = \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_3_U.b [3:0];
assign \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_3_U.u1.cin  = 1'h0;
assign \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_3_U.facout_s1  = \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_3_U.u1.cout ;
assign \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_3_U.fas_s1  = \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_3_U.u1.s ;
assign \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_3_U.a  = \add_9ns_9ns_9_2_1_U5.din0 ;
assign \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_3_U.b  = \add_9ns_9ns_9_2_1_U5.din1 ;
assign \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_3_U.ce  = \add_9ns_9ns_9_2_1_U5.ce ;
assign \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_3_U.clk  = \add_9ns_9ns_9_2_1_U5.clk ;
assign \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_3_U.reset  = \add_9ns_9ns_9_2_1_U5.reset ;
assign \add_9ns_9ns_9_2_1_U5.dout  = \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_3_U.s ;
assign \add_9ns_9ns_9_2_1_U5.ce  = 1'h1;
assign \add_9ns_9ns_9_2_1_U5.clk  = ap_clk;
assign \add_9ns_9ns_9_2_1_U5.din0  = { 6'h00, add_ln69_1_reg_558 };
assign \add_9ns_9ns_9_2_1_U5.din1  = ret_reg_553;
assign grp_fu_259_p2 = \add_9ns_9ns_9_2_1_U5.dout ;
assign \add_9ns_9ns_9_2_1_U5.reset  = ap_rst;
assign \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_6_U.ain_s0  = \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_6_U.a ;
assign \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_6_U.bin_s0  = \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_6_U.b ;
assign \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_6_U.s  = { \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_6_U.fas_s2 , \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_6_U.sum_s1  };
assign \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_6_U.u2.a  = \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_6_U.ain_s1 ;
assign \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_6_U.u2.b  = \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_6_U.bin_s1 ;
assign \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_6_U.u2.cin  = \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_6_U.carry_s1 ;
assign \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_6_U.facout_s2  = \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_6_U.u2.cout ;
assign \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_6_U.fas_s2  = \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_6_U.u2.s ;
assign \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_6_U.u1.a  = \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_6_U.a [0];
assign \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_6_U.u1.b  = \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_6_U.b [0];
assign \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_6_U.u1.cin  = 1'h0;
assign \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_6_U.facout_s1  = \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_6_U.u1.cout ;
assign \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_6_U.fas_s1  = \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_6_U.u1.s ;
assign \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_6_U.a  = \add_3s_3ns_3_2_1_U13.din0 ;
assign \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_6_U.b  = \add_3s_3ns_3_2_1_U13.din1 ;
assign \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_6_U.ce  = \add_3s_3ns_3_2_1_U13.ce ;
assign \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_6_U.clk  = \add_3s_3ns_3_2_1_U13.clk ;
assign \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_6_U.reset  = \add_3s_3ns_3_2_1_U13.reset ;
assign \add_3s_3ns_3_2_1_U13.dout  = \add_3s_3ns_3_2_1_U13.top_add_3s_3ns_3_2_1_Adder_6_U.s ;
assign \add_3s_3ns_3_2_1_U13.ce  = 1'h1;
assign \add_3s_3ns_3_2_1_U13.clk  = ap_clk;
assign \add_3s_3ns_3_2_1_U13.din0  = { add_ln69_7_reg_695[1], add_ln69_7_reg_695 };
assign \add_3s_3ns_3_2_1_U13.din1  = add_ln69_6_reg_690;
assign grp_fu_399_p2 = \add_3s_3ns_3_2_1_U13.dout ;
assign \add_3s_3ns_3_2_1_U13.reset  = ap_rst;
assign \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.ain_s0  = \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.a ;
assign \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.bin_s0  = \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.b ;
assign \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.s  = { \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.fas_s2 , \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.sum_s1  };
assign \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.u2.a  = \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.ain_s1 ;
assign \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.u2.b  = \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.bin_s1 ;
assign \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.u2.cin  = \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.carry_s1 ;
assign \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.facout_s2  = \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.u2.cout ;
assign \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.fas_s2  = \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.u2.s ;
assign \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.u1.a  = \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.a [0];
assign \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.u1.b  = \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.b [0];
assign \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.u1.cin  = 1'h0;
assign \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.facout_s1  = \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.u1.cout ;
assign \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.fas_s1  = \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.u1.s ;
assign \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.a  = \add_3s_3ns_3_2_1_U10.din0 ;
assign \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.b  = \add_3s_3ns_3_2_1_U10.din1 ;
assign \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.ce  = \add_3s_3ns_3_2_1_U10.ce ;
assign \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.clk  = \add_3s_3ns_3_2_1_U10.clk ;
assign \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.reset  = \add_3s_3ns_3_2_1_U10.reset ;
assign \add_3s_3ns_3_2_1_U10.dout  = \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.s ;
assign \add_3s_3ns_3_2_1_U10.ce  = 1'h1;
assign \add_3s_3ns_3_2_1_U10.clk  = ap_clk;
assign \add_3s_3ns_3_2_1_U10.din0  = { op_16_V_reg_645[1], op_16_V_reg_645 };
assign \add_3s_3ns_3_2_1_U10.din1  = select_ln69_reg_665;
assign grp_fu_381_p2 = \add_3s_3ns_3_2_1_U10.dout ;
assign \add_3s_3ns_3_2_1_U10.reset  = ap_rst;
assign \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_1_U.ain_s0  = \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_1_U.a ;
assign \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_1_U.bin_s0  = \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_1_U.b ;
assign \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_1_U.s  = { \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_1_U.fas_s2 , \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_1_U.sum_s1  };
assign \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_1_U.u2.a  = \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_1_U.ain_s1 ;
assign \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_1_U.u2.b  = \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_1_U.bin_s1 ;
assign \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_1_U.u2.cin  = \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_1_U.carry_s1 ;
assign \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_1_U.facout_s2  = \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_1_U.u2.cout ;
assign \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_1_U.fas_s2  = \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_1_U.u2.s ;
assign \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_1_U.u1.a  = \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_1_U.a [0];
assign \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_1_U.u1.b  = \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_1_U.b [0];
assign \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_1_U.u1.cin  = 1'h0;
assign \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_1_U.facout_s1  = \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_1_U.u1.cout ;
assign \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_1_U.fas_s1  = \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_1_U.u1.s ;
assign \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_1_U.a  = \add_3ns_3ns_3_2_1_U3.din0 ;
assign \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_1_U.b  = \add_3ns_3ns_3_2_1_U3.din1 ;
assign \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_1_U.ce  = \add_3ns_3ns_3_2_1_U3.ce ;
assign \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_1_U.clk  = \add_3ns_3ns_3_2_1_U3.clk ;
assign \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_1_U.reset  = \add_3ns_3ns_3_2_1_U3.reset ;
assign \add_3ns_3ns_3_2_1_U3.dout  = \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_1_U.s ;
assign \add_3ns_3ns_3_2_1_U3.ce  = 1'h1;
assign \add_3ns_3ns_3_2_1_U3.clk  = ap_clk;
assign \add_3ns_3ns_3_2_1_U3.din0  = { 1'h0, r_1_reg_523 };
assign \add_3ns_3ns_3_2_1_U3.din1  = { 2'h0, op_9_V_reg_518 };
assign grp_fu_240_p2 = \add_3ns_3ns_3_2_1_U3.dout ;
assign \add_3ns_3ns_3_2_1_U3.reset  = ap_rst;
assign \add_36s_36s_36_2_1_U15.top_add_36s_36s_36_2_1_Adder_8_U.ain_s0  = \add_36s_36s_36_2_1_U15.top_add_36s_36s_36_2_1_Adder_8_U.a ;
assign \add_36s_36s_36_2_1_U15.top_add_36s_36s_36_2_1_Adder_8_U.bin_s0  = \add_36s_36s_36_2_1_U15.top_add_36s_36s_36_2_1_Adder_8_U.b ;
assign \add_36s_36s_36_2_1_U15.top_add_36s_36s_36_2_1_Adder_8_U.s  = { \add_36s_36s_36_2_1_U15.top_add_36s_36s_36_2_1_Adder_8_U.fas_s2 , \add_36s_36s_36_2_1_U15.top_add_36s_36s_36_2_1_Adder_8_U.sum_s1  };
assign \add_36s_36s_36_2_1_U15.top_add_36s_36s_36_2_1_Adder_8_U.u2.a  = \add_36s_36s_36_2_1_U15.top_add_36s_36s_36_2_1_Adder_8_U.ain_s1 ;
assign \add_36s_36s_36_2_1_U15.top_add_36s_36s_36_2_1_Adder_8_U.u2.b  = \add_36s_36s_36_2_1_U15.top_add_36s_36s_36_2_1_Adder_8_U.bin_s1 ;
assign \add_36s_36s_36_2_1_U15.top_add_36s_36s_36_2_1_Adder_8_U.u2.cin  = \add_36s_36s_36_2_1_U15.top_add_36s_36s_36_2_1_Adder_8_U.carry_s1 ;
assign \add_36s_36s_36_2_1_U15.top_add_36s_36s_36_2_1_Adder_8_U.facout_s2  = \add_36s_36s_36_2_1_U15.top_add_36s_36s_36_2_1_Adder_8_U.u2.cout ;
assign \add_36s_36s_36_2_1_U15.top_add_36s_36s_36_2_1_Adder_8_U.fas_s2  = \add_36s_36s_36_2_1_U15.top_add_36s_36s_36_2_1_Adder_8_U.u2.s ;
assign \add_36s_36s_36_2_1_U15.top_add_36s_36s_36_2_1_Adder_8_U.u1.a  = \add_36s_36s_36_2_1_U15.top_add_36s_36s_36_2_1_Adder_8_U.a [17:0];
assign \add_36s_36s_36_2_1_U15.top_add_36s_36s_36_2_1_Adder_8_U.u1.b  = \add_36s_36s_36_2_1_U15.top_add_36s_36s_36_2_1_Adder_8_U.b [17:0];
assign \add_36s_36s_36_2_1_U15.top_add_36s_36s_36_2_1_Adder_8_U.u1.cin  = 1'h0;
assign \add_36s_36s_36_2_1_U15.top_add_36s_36s_36_2_1_Adder_8_U.facout_s1  = \add_36s_36s_36_2_1_U15.top_add_36s_36s_36_2_1_Adder_8_U.u1.cout ;
assign \add_36s_36s_36_2_1_U15.top_add_36s_36s_36_2_1_Adder_8_U.fas_s1  = \add_36s_36s_36_2_1_U15.top_add_36s_36s_36_2_1_Adder_8_U.u1.s ;
assign \add_36s_36s_36_2_1_U15.top_add_36s_36s_36_2_1_Adder_8_U.a  = \add_36s_36s_36_2_1_U15.din0 ;
assign \add_36s_36s_36_2_1_U15.top_add_36s_36s_36_2_1_Adder_8_U.b  = \add_36s_36s_36_2_1_U15.din1 ;
assign \add_36s_36s_36_2_1_U15.top_add_36s_36s_36_2_1_Adder_8_U.ce  = \add_36s_36s_36_2_1_U15.ce ;
assign \add_36s_36s_36_2_1_U15.top_add_36s_36s_36_2_1_Adder_8_U.clk  = \add_36s_36s_36_2_1_U15.clk ;
assign \add_36s_36s_36_2_1_U15.top_add_36s_36s_36_2_1_Adder_8_U.reset  = \add_36s_36s_36_2_1_U15.reset ;
assign \add_36s_36s_36_2_1_U15.dout  = \add_36s_36s_36_2_1_U15.top_add_36s_36s_36_2_1_Adder_8_U.s ;
assign \add_36s_36s_36_2_1_U15.ce  = 1'h1;
assign \add_36s_36s_36_2_1_U15.clk  = ap_clk;
assign \add_36s_36s_36_2_1_U15.din0  = { op_31_V_reg_725[31], op_31_V_reg_725, 3'h0 };
assign \add_36s_36s_36_2_1_U15.din1  = { op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19 };
assign grp_fu_427_p2 = \add_36s_36s_36_2_1_U15.dout ;
assign \add_36s_36s_36_2_1_U15.reset  = ap_rst;
assign \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_5_U.ain_s0  = \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_5_U.a ;
assign \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_5_U.bin_s0  = \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_5_U.b ;
assign \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_5_U.s  = { \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_5_U.fas_s2 , \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_5_U.sum_s1  };
assign \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_5_U.u2.a  = \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_5_U.ain_s1 ;
assign \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_5_U.u2.b  = \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_5_U.bin_s1 ;
assign \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_5_U.u2.cin  = \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_5_U.carry_s1 ;
assign \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_5_U.facout_s2  = \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_5_U.u2.cout ;
assign \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_5_U.fas_s2  = \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_5_U.u2.s ;
assign \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_5_U.u1.a  = \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_5_U.a [16:0];
assign \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_5_U.u1.b  = \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_5_U.b [16:0];
assign \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_5_U.u1.cin  = 1'h0;
assign \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_5_U.facout_s1  = \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_5_U.u1.cout ;
assign \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_5_U.fas_s1  = \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_5_U.u1.s ;
assign \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_5_U.a  = \add_34s_34s_34_2_1_U7.din0 ;
assign \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_5_U.b  = \add_34s_34s_34_2_1_U7.din1 ;
assign \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_5_U.ce  = \add_34s_34s_34_2_1_U7.ce ;
assign \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_5_U.clk  = \add_34s_34s_34_2_1_U7.clk ;
assign \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_5_U.reset  = \add_34s_34s_34_2_1_U7.reset ;
assign \add_34s_34s_34_2_1_U7.dout  = \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_5_U.s ;
assign \add_34s_34s_34_2_1_U7.ce  = 1'h1;
assign \add_34s_34s_34_2_1_U7.clk  = ap_clk;
assign \add_34s_34s_34_2_1_U7.din0  = { op_24_V_reg_593[31], op_24_V_reg_593, 1'h0 };
assign \add_34s_34s_34_2_1_U7.din1  = { op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12 };
assign grp_fu_287_p2 = \add_34s_34s_34_2_1_U7.dout ;
assign \add_34s_34s_34_2_1_U7.reset  = ap_rst;
assign \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_4_U.ain_s0  = \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_4_U.a ;
assign \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_4_U.bin_s0  = \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_4_U.b ;
assign \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_4_U.s  = { \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_4_U.fas_s2 , \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_4_U.sum_s1  };
assign \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_4_U.u2.a  = \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_4_U.ain_s1 ;
assign \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_4_U.u2.b  = \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_4_U.bin_s1 ;
assign \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_4_U.u2.cin  = \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_4_U.carry_s1 ;
assign \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_4_U.facout_s2  = \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_4_U.u2.cout ;
assign \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_4_U.fas_s2  = \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_4_U.u2.s ;
assign \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_4_U.u1.a  = \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_4_U.a [15:0];
assign \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_4_U.u1.b  = \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_4_U.b [15:0];
assign \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_4_U.u1.cin  = 1'h0;
assign \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_4_U.facout_s1  = \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_4_U.u1.cout ;
assign \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_4_U.fas_s1  = \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_4_U.u1.s ;
assign \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_4_U.a  = \add_32s_32ns_32_2_1_U6.din0 ;
assign \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_4_U.b  = \add_32s_32ns_32_2_1_U6.din1 ;
assign \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_4_U.ce  = \add_32s_32ns_32_2_1_U6.ce ;
assign \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_4_U.clk  = \add_32s_32ns_32_2_1_U6.clk ;
assign \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_4_U.reset  = \add_32s_32ns_32_2_1_U6.reset ;
assign \add_32s_32ns_32_2_1_U6.dout  = \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_4_U.s ;
assign \add_32s_32ns_32_2_1_U6.ce  = 1'h1;
assign \add_32s_32ns_32_2_1_U6.clk  = ap_clk;
assign \add_32s_32ns_32_2_1_U6.din0  = { add_ln69_2_reg_583[8], add_ln69_2_reg_583[8], add_ln69_2_reg_583[8], add_ln69_2_reg_583[8], add_ln69_2_reg_583[8], add_ln69_2_reg_583[8], add_ln69_2_reg_583[8], add_ln69_2_reg_583[8], add_ln69_2_reg_583[8], add_ln69_2_reg_583[8], add_ln69_2_reg_583[8], add_ln69_2_reg_583[8], add_ln69_2_reg_583[8], add_ln69_2_reg_583[8], add_ln69_2_reg_583[8], add_ln69_2_reg_583[8], add_ln69_2_reg_583[8], add_ln69_2_reg_583[8], add_ln69_2_reg_583[8], add_ln69_2_reg_583[8], add_ln69_2_reg_583[8], add_ln69_2_reg_583[8], add_ln69_2_reg_583[8], add_ln69_2_reg_583 };
assign \add_32s_32ns_32_2_1_U6.din1  = add_ln69_reg_578;
assign grp_fu_267_p2 = \add_32s_32ns_32_2_1_U6.dout ;
assign \add_32s_32ns_32_2_1_U6.reset  = ap_rst;
assign \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_4_U.ain_s0  = \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_4_U.a ;
assign \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_4_U.bin_s0  = \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_4_U.b ;
assign \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_4_U.s  = { \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_4_U.fas_s2 , \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_4_U.sum_s1  };
assign \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_4_U.u2.a  = \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_4_U.ain_s1 ;
assign \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_4_U.u2.b  = \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_4_U.bin_s1 ;
assign \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_4_U.u2.cin  = \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_4_U.carry_s1 ;
assign \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_4_U.facout_s2  = \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_4_U.u2.cout ;
assign \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_4_U.fas_s2  = \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_4_U.u2.s ;
assign \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_4_U.u1.a  = \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_4_U.a [15:0];
assign \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_4_U.u1.b  = \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_4_U.b [15:0];
assign \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_4_U.u1.cin  = 1'h0;
assign \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_4_U.facout_s1  = \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_4_U.u1.cout ;
assign \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_4_U.fas_s1  = \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_4_U.u1.s ;
assign \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_4_U.a  = \add_32s_32ns_32_2_1_U14.din0 ;
assign \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_4_U.b  = \add_32s_32ns_32_2_1_U14.din1 ;
assign \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_4_U.ce  = \add_32s_32ns_32_2_1_U14.ce ;
assign \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_4_U.clk  = \add_32s_32ns_32_2_1_U14.clk ;
assign \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_4_U.reset  = \add_32s_32ns_32_2_1_U14.reset ;
assign \add_32s_32ns_32_2_1_U14.dout  = \add_32s_32ns_32_2_1_U14.top_add_32s_32ns_32_2_1_Adder_4_U.s ;
assign \add_32s_32ns_32_2_1_U14.ce  = 1'h1;
assign \add_32s_32ns_32_2_1_U14.clk  = ap_clk;
assign \add_32s_32ns_32_2_1_U14.din0  = { add_ln69_8_reg_715[2], add_ln69_8_reg_715[2], add_ln69_8_reg_715[2], add_ln69_8_reg_715[2], add_ln69_8_reg_715[2], add_ln69_8_reg_715[2], add_ln69_8_reg_715[2], add_ln69_8_reg_715[2], add_ln69_8_reg_715[2], add_ln69_8_reg_715[2], add_ln69_8_reg_715[2], add_ln69_8_reg_715[2], add_ln69_8_reg_715[2], add_ln69_8_reg_715[2], add_ln69_8_reg_715[2], add_ln69_8_reg_715[2], add_ln69_8_reg_715[2], add_ln69_8_reg_715[2], add_ln69_8_reg_715[2], add_ln69_8_reg_715[2], add_ln69_8_reg_715[2], add_ln69_8_reg_715[2], add_ln69_8_reg_715[2], add_ln69_8_reg_715[2], add_ln69_8_reg_715[2], add_ln69_8_reg_715[2], add_ln69_8_reg_715[2], add_ln69_8_reg_715[2], add_ln69_8_reg_715[2], add_ln69_8_reg_715 };
assign \add_32s_32ns_32_2_1_U14.din1  = add_ln69_5_reg_710;
assign grp_fu_407_p2 = \add_32s_32ns_32_2_1_U14.dout ;
assign \add_32s_32ns_32_2_1_U14.reset  = ap_rst;
assign \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_4_U.ain_s0  = \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_4_U.a ;
assign \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_4_U.bin_s0  = \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_4_U.b ;
assign \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_4_U.s  = { \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_4_U.fas_s2 , \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_4_U.sum_s1  };
assign \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_4_U.u2.a  = \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_4_U.ain_s1 ;
assign \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_4_U.u2.b  = \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_4_U.bin_s1 ;
assign \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_4_U.u2.cin  = \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_4_U.carry_s1 ;
assign \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_4_U.facout_s2  = \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_4_U.u2.cout ;
assign \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_4_U.fas_s2  = \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_4_U.u2.s ;
assign \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_4_U.u1.a  = \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_4_U.a [15:0];
assign \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_4_U.u1.b  = \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_4_U.b [15:0];
assign \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_4_U.u1.cin  = 1'h0;
assign \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_4_U.facout_s1  = \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_4_U.u1.cout ;
assign \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_4_U.fas_s1  = \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_4_U.u1.s ;
assign \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_4_U.a  = \add_32s_32ns_32_2_1_U12.din0 ;
assign \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_4_U.b  = \add_32s_32ns_32_2_1_U12.din1 ;
assign \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_4_U.ce  = \add_32s_32ns_32_2_1_U12.ce ;
assign \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_4_U.clk  = \add_32s_32ns_32_2_1_U12.clk ;
assign \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_4_U.reset  = \add_32s_32ns_32_2_1_U12.reset ;
assign \add_32s_32ns_32_2_1_U12.dout  = \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_4_U.s ;
assign \add_32s_32ns_32_2_1_U12.ce  = 1'h1;
assign \add_32s_32ns_32_2_1_U12.clk  = ap_clk;
assign \add_32s_32ns_32_2_1_U12.din0  = add_ln69_4_reg_685;
assign \add_32s_32ns_32_2_1_U12.din1  = op_14;
assign grp_fu_391_p2 = \add_32s_32ns_32_2_1_U12.dout ;
assign \add_32s_32ns_32_2_1_U12.reset  = ap_rst;
assign \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_2_U.ain_s0  = \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_2_U.a ;
assign \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_2_U.bin_s0  = \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_2_U.b ;
assign \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_2_U.s  = { \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_2_U.fas_s2 , \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_2_U.sum_s1  };
assign \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_2_U.u2.a  = \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_2_U.ain_s1 ;
assign \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_2_U.u2.b  = \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_2_U.bin_s1 ;
assign \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_2_U.u2.cin  = \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_2_U.carry_s1 ;
assign \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_2_U.facout_s2  = \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_2_U.u2.cout ;
assign \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_2_U.fas_s2  = \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_2_U.u2.s ;
assign \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_2_U.u1.a  = \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_2_U.a [15:0];
assign \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_2_U.u1.b  = \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_2_U.b [15:0];
assign \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_2_U.u1.cin  = 1'h0;
assign \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_2_U.facout_s1  = \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_2_U.u1.cout ;
assign \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_2_U.fas_s1  = \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_2_U.u1.s ;
assign \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_2_U.a  = \add_32ns_32ns_32_2_1_U9.din0 ;
assign \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_2_U.b  = \add_32ns_32ns_32_2_1_U9.din1 ;
assign \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_2_U.ce  = \add_32ns_32ns_32_2_1_U9.ce ;
assign \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_2_U.clk  = \add_32ns_32ns_32_2_1_U9.clk ;
assign \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_2_U.reset  = \add_32ns_32ns_32_2_1_U9.reset ;
assign \add_32ns_32ns_32_2_1_U9.dout  = \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_2_U.s ;
assign \add_32ns_32ns_32_2_1_U9.ce  = 1'h1;
assign \add_32ns_32ns_32_2_1_U9.clk  = ap_clk;
assign \add_32ns_32ns_32_2_1_U9.din0  = ret_V_cast_reg_618;
assign \add_32ns_32ns_32_2_1_U9.din1  = 32'd1;
assign grp_fu_316_p2 = \add_32ns_32ns_32_2_1_U9.dout ;
assign \add_32ns_32ns_32_2_1_U9.reset  = ap_rst;
assign \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_2_U.ain_s0  = \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_2_U.a ;
assign \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_2_U.bin_s0  = \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_2_U.b ;
assign \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_2_U.s  = { \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_2_U.fas_s2 , \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_2_U.sum_s1  };
assign \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_2_U.u2.a  = \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_2_U.ain_s1 ;
assign \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_2_U.u2.b  = \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_2_U.bin_s1 ;
assign \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_2_U.u2.cin  = \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_2_U.carry_s1 ;
assign \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_2_U.facout_s2  = \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_2_U.u2.cout ;
assign \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_2_U.fas_s2  = \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_2_U.u2.s ;
assign \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_2_U.u1.a  = \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_2_U.a [15:0];
assign \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_2_U.u1.b  = \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_2_U.b [15:0];
assign \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_2_U.u1.cin  = 1'h0;
assign \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_2_U.facout_s1  = \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_2_U.u1.cout ;
assign \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_2_U.fas_s1  = \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_2_U.u1.s ;
assign \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_2_U.a  = \add_32ns_32ns_32_2_1_U4.din0 ;
assign \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_2_U.b  = \add_32ns_32ns_32_2_1_U4.din1 ;
assign \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_2_U.ce  = \add_32ns_32ns_32_2_1_U4.ce ;
assign \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_2_U.clk  = \add_32ns_32ns_32_2_1_U4.clk ;
assign \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_2_U.reset  = \add_32ns_32ns_32_2_1_U4.reset ;
assign \add_32ns_32ns_32_2_1_U4.dout  = \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_2_U.s ;
assign \add_32ns_32ns_32_2_1_U4.ce  = 1'h1;
assign \add_32ns_32ns_32_2_1_U4.clk  = ap_clk;
assign \add_32ns_32ns_32_2_1_U4.din0  = { 16'h0000, op_4 };
assign \add_32ns_32ns_32_2_1_U4.din1  = op_10;
assign grp_fu_250_p2 = \add_32ns_32ns_32_2_1_U4.dout ;
assign \add_32ns_32ns_32_2_1_U4.reset  = ap_rst;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_2_U.ain_s0  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_2_U.a ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_2_U.bin_s0  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_2_U.b ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_2_U.s  = { \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_2_U.fas_s2 , \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_2_U.sum_s1  };
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_2_U.u2.a  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_2_U.ain_s1 ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_2_U.u2.b  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_2_U.bin_s1 ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_2_U.u2.cin  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_2_U.carry_s1 ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_2_U.facout_s2  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_2_U.u2.cout ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_2_U.fas_s2  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_2_U.u2.s ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_2_U.u1.a  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_2_U.a [15:0];
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_2_U.u1.b  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_2_U.b [15:0];
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_2_U.u1.cin  = 1'h0;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_2_U.facout_s1  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_2_U.u1.cout ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_2_U.fas_s1  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_2_U.u1.s ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_2_U.a  = \add_32ns_32ns_32_2_1_U16.din0 ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_2_U.b  = \add_32ns_32ns_32_2_1_U16.din1 ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_2_U.ce  = \add_32ns_32ns_32_2_1_U16.ce ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_2_U.clk  = \add_32ns_32ns_32_2_1_U16.clk ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_2_U.reset  = \add_32ns_32ns_32_2_1_U16.reset ;
assign \add_32ns_32ns_32_2_1_U16.dout  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_2_U.s ;
assign \add_32ns_32ns_32_2_1_U16.ce  = 1'h1;
assign \add_32ns_32ns_32_2_1_U16.clk  = ap_clk;
assign \add_32ns_32ns_32_2_1_U16.din0  = ret_V_3_cast_reg_750;
assign \add_32ns_32ns_32_2_1_U16.din1  = 32'd1;
assign grp_fu_453_p2 = \add_32ns_32ns_32_2_1_U16.dout ;
assign \add_32ns_32ns_32_2_1_U16.reset  = ap_rst;
assign \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_7_U.ain_s0  = \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_7_U.a ;
assign \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_7_U.bin_s0  = \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_7_U.b ;
assign \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_7_U.s  = { \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_7_U.fas_s2 , \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_7_U.sum_s1  };
assign \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_7_U.u2.a  = \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_7_U.ain_s1 ;
assign \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_7_U.u2.b  = \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_7_U.bin_s1 ;
assign \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_7_U.u2.cin  = \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_7_U.carry_s1 ;
assign \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_7_U.facout_s2  = \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_7_U.u2.cout ;
assign \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_7_U.fas_s2  = \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_7_U.u2.s ;
assign \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_7_U.u1.a  = \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_7_U.a [0];
assign \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_7_U.u1.b  = \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_7_U.b [0];
assign \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_7_U.u1.cin  = 1'h0;
assign \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_7_U.facout_s1  = \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_7_U.u1.cout ;
assign \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_7_U.fas_s1  = \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_7_U.u1.s ;
assign \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_7_U.a  = \add_2ns_2ns_2_2_1_U11.din0 ;
assign \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_7_U.b  = \add_2ns_2ns_2_2_1_U11.din1 ;
assign \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_7_U.ce  = \add_2ns_2ns_2_2_1_U11.ce ;
assign \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_7_U.clk  = \add_2ns_2ns_2_2_1_U11.clk ;
assign \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_7_U.reset  = \add_2ns_2ns_2_2_1_U11.reset ;
assign \add_2ns_2ns_2_2_1_U11.dout  = \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_7_U.s ;
assign \add_2ns_2ns_2_2_1_U11.ce  = 1'h1;
assign \add_2ns_2ns_2_2_1_U11.clk  = ap_clk;
assign \add_2ns_2ns_2_2_1_U11.din0  = select_ln69_1_reg_670;
assign \add_2ns_2ns_2_2_1_U11.din1  = { 1'h0, xor_ln890_reg_655 };
assign grp_fu_386_p2 = \add_2ns_2ns_2_2_1_U11.dout ;
assign \add_2ns_2ns_2_2_1_U11.reset  = ap_rst;
endmodule


// Product machine:
module top_A_times_top_B (ap_start, op_0, op_1, op_10, op_12, op_13, op_14, op_18, op_19, op_2, op_3, op_4, op_5, ap_clk, unsafe_signal);
input ap_start;
input [7:0] op_0;
input [3:0] op_1;
input [31:0] op_10;
input [1:0] op_12;
input op_13;
input [31:0] op_14;
input op_18;
input [3:0] op_19;
input [3:0] op_2;
input [1:0] op_3;
input [15:0] op_4;
input [1:0] op_5;
input ap_clk;
output unsafe_signal;
reg _setup;
initial _setup = 1'b0;
always @ (posedge ap_clk) _setup <= 1'b1;
reg ap_start_internal;
always @ (posedge ap_clk) if (!_setup) ap_start_internal <= ap_start;
reg [7:0] op_0_internal;
always @ (posedge ap_clk) if (!_setup) op_0_internal <= op_0;
reg [3:0] op_1_internal;
always @ (posedge ap_clk) if (!_setup) op_1_internal <= op_1;
reg [31:0] op_10_internal;
always @ (posedge ap_clk) if (!_setup) op_10_internal <= op_10;
reg [1:0] op_12_internal;
always @ (posedge ap_clk) if (!_setup) op_12_internal <= op_12;
reg op_13_internal;
always @ (posedge ap_clk) if (!_setup) op_13_internal <= op_13;
reg [31:0] op_14_internal;
always @ (posedge ap_clk) if (!_setup) op_14_internal <= op_14;
reg op_18_internal;
always @ (posedge ap_clk) if (!_setup) op_18_internal <= op_18;
reg [3:0] op_19_internal;
always @ (posedge ap_clk) if (!_setup) op_19_internal <= op_19;
reg [3:0] op_2_internal;
always @ (posedge ap_clk) if (!_setup) op_2_internal <= op_2;
reg [1:0] op_3_internal;
always @ (posedge ap_clk) if (!_setup) op_3_internal <= op_3;
reg [15:0] op_4_internal;
always @ (posedge ap_clk) if (!_setup) op_4_internal <= op_4;
reg [1:0] op_5_internal;
always @ (posedge ap_clk) if (!_setup) op_5_internal <= op_5;
wire ap_done_A;
wire ap_done_B;
wire ap_done_eq;
assign ap_done_eq = ap_done_A == ap_done_B;
wire ap_idle_A;
wire ap_idle_B;
wire ap_idle_eq;
assign ap_idle_eq = ap_idle_A == ap_idle_B;
wire ap_ready_A;
wire ap_ready_B;
wire ap_ready_eq;
assign ap_ready_eq = ap_ready_A == ap_ready_B;
wire [31:0] op_32_A;
wire [31:0] op_32_B;
wire op_32_eq;
assign op_32_eq = op_32_A == op_32_B;
wire op_32_ap_vld_A;
wire op_32_ap_vld_B;
wire clk_enable_A;
wire clk_enable_B;
assign clk_enable_A = _setup & (~op_32_ap_vld_A | op_32_ap_vld_B);
assign clk_enable_B = _setup;
wire divergent;
assign divergent = ~(ap_done_eq & ap_idle_eq & ap_ready_eq & op_32_eq);
assign unsafe_signal = op_32_ap_vld_A & op_32_ap_vld_B & divergent;
top_A instance_A (
    .ap_clk(ap_clk),
    .clk_enable(clk_enable_A),
    .ap_start(ap_start_internal),
    .op_0(op_0_internal),
    .op_1(op_1_internal),
    .op_10(op_10_internal),
    .op_12(op_12_internal),
    .op_13(op_13_internal),
    .op_14(op_14_internal),
    .op_18(op_18_internal),
    .op_19(op_19_internal),
    .op_2(op_2_internal),
    .op_3(op_3_internal),
    .op_4(op_4_internal),
    .op_5(op_5_internal),
    .ap_done(ap_done_A),
    .ap_idle(ap_idle_A),
    .ap_ready(ap_ready_A),
    .op_32(op_32_A),
    .op_32_ap_vld(op_32_ap_vld_A)
);
top_B instance_B (
    .ap_clk(ap_clk),
    .clk_enable(clk_enable_B),
    .ap_start(ap_start_internal),
    .op_0(op_0_internal),
    .op_1(op_1_internal),
    .op_10(op_10_internal),
    .op_12(op_12_internal),
    .op_13(op_13_internal),
    .op_14(op_14_internal),
    .op_18(op_18_internal),
    .op_19(op_19_internal),
    .op_2(op_2_internal),
    .op_3(op_3_internal),
    .op_4(op_4_internal),
    .op_5(op_5_internal),
    .ap_done(ap_done_B),
    .ap_idle(ap_idle_B),
    .ap_ready(ap_ready_B),
    .op_32(op_32_B),
    .op_32_ap_vld(op_32_ap_vld_B)
);
endmodule
