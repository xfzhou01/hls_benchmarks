// Processed by function `construct_kairos` in `verilog_tricks.py`.
// Machine A:
// Processed by function `add_clk_enable_signal` in `verilog_tricks.py`.
// Processed by function `remove_reset_signal` in `verilog_tricks.py`.
module top_A (
  ap_clk,
  ap_start,
  ap_done,
  ap_idle,
  ap_ready,
  op_0,
  op_2,
  op_3,
  op_5,
  op_6,
  op_8,
  op_9,
  op_10,
  op_13,
  op_14,
  op_15,
  op_17,
  op_18,
  op_30,
  op_30_ap_vld,
clk_enable
);
input clk_enable;


input ap_clk;
wire ap_rst;
assign ap_rst = op_30_ap_vld;
input ap_start;
input [3:0] op_0;
input [7:0] op_10;
input [1:0] op_13;
input [1:0] op_14;
input [31:0] op_15;
input [1:0] op_17;
input [1:0] op_18;
input [15:0] op_2;
input [3:0] op_3;
input [3:0] op_5;
input [7:0] op_6;
input [3:0] op_8;
input [3:0] op_9;
output ap_done;
output ap_idle;
output ap_ready;
output [31:0] op_30;
output op_30_ap_vld;


reg Range1_all_ones_reg_1444;
reg Range1_all_zeros_reg_1451;
reg Range2_all_ones_reg_1439;
reg [8:0] \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.ain_s1 ;
reg [8:0] \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.bin_s1 ;
reg \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.carry_s1 ;
reg [7:0] \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.sum_s1 ;
reg [8:0] \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.ain_s1 ;
reg [8:0] \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.bin_s1 ;
reg \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.carry_s1 ;
reg [7:0] \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.sum_s1 ;
reg [8:0] \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.ain_s1 ;
reg [8:0] \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.bin_s1 ;
reg \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.carry_s1 ;
reg [7:0] \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.sum_s1 ;
reg \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.ain_s1 ;
reg \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.bin_s1 ;
reg \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.carry_s1 ;
reg \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.sum_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.ain_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.bin_s1 ;
reg \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.carry_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.sum_s1 ;
reg [15:0] \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.ain_s1 ;
reg [15:0] \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.bin_s1 ;
reg \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.carry_s1 ;
reg [15:0] \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.sum_s1 ;
reg [15:0] \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.ain_s1 ;
reg [15:0] \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.bin_s1 ;
reg \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.carry_s1 ;
reg [15:0] \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.sum_s1 ;
reg [15:0] \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.ain_s1 ;
reg [15:0] \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.bin_s1 ;
reg \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.carry_s1 ;
reg [15:0] \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.sum_s1 ;
reg [16:0] \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.ain_s1 ;
reg [16:0] \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.bin_s1 ;
reg \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.carry_s1 ;
reg [16:0] \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.sum_s1 ;
reg [1:0] \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.ain_s1 ;
reg [1:0] \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.bin_s1 ;
reg \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.carry_s1 ;
reg \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.sum_s1 ;
reg [1:0] \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.ain_s1 ;
reg [1:0] \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.bin_s1 ;
reg \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.carry_s1 ;
reg \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.sum_s1 ;
reg [1:0] \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.ain_s1 ;
reg [1:0] \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.bin_s1 ;
reg \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.carry_s1 ;
reg [1:0] \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.sum_s1 ;
reg [1:0] \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.ain_s1 ;
reg [1:0] \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.bin_s1 ;
reg \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.carry_s1 ;
reg [1:0] \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.sum_s1 ;
reg [2:0] \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.ain_s1 ;
reg [2:0] \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.bin_s1 ;
reg \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.carry_s1 ;
reg [2:0] \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.sum_s1 ;
reg [3:0] \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.ain_s1 ;
reg [3:0] \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.bin_s1 ;
reg \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.carry_s1 ;
reg [2:0] \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.sum_s1 ;
reg [3:0] \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.ain_s1 ;
reg [3:0] \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.bin_s1 ;
reg \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.carry_s1 ;
reg [2:0] \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.sum_s1 ;
reg [3:0] \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.ain_s1 ;
reg [3:0] \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.bin_s1 ;
reg \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.carry_s1 ;
reg [2:0] \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.sum_s1 ;
reg [3:0] add_ln1192_1_reg_1387;
reg [2:0] add_ln1192_2_reg_1327;
reg [31:0] add_ln691_reg_1570;
reg [6:0] add_ln69_1_reg_1342;
reg [31:0] add_ln69_3_reg_1492;
reg [31:0] add_ln69_4_reg_1528;
reg [2:0] add_ln69_5_reg_1497;
reg [3:0] add_ln69_6_reg_1533;
reg [16:0] add_ln69_reg_1337;
reg and_ln786_reg_1169;
reg and_ln788_1_reg_1482;
reg [24:0] ap_CS_fsm = 25'h0000001;
reg [15:0] \ashr_16s_16ns_16_7_1_U3.din1_cast_array[0] ;
reg [15:0] \ashr_16s_16ns_16_7_1_U3.din1_cast_array[1] ;
reg [15:0] \ashr_16s_16ns_16_7_1_U3.din1_cast_array[2] ;
reg [15:0] \ashr_16s_16ns_16_7_1_U3.din1_cast_array[3] ;
reg [15:0] \ashr_16s_16ns_16_7_1_U3.din1_cast_array[4] ;
reg [15:0] \ashr_16s_16ns_16_7_1_U3.din1_cast_array[5] ;
reg [15:0] \ashr_16s_16ns_16_7_1_U3.dout_array[0] ;
reg [15:0] \ashr_16s_16ns_16_7_1_U3.dout_array[1] ;
reg [15:0] \ashr_16s_16ns_16_7_1_U3.dout_array[2] ;
reg [15:0] \ashr_16s_16ns_16_7_1_U3.dout_array[3] ;
reg [15:0] \ashr_16s_16ns_16_7_1_U3.dout_array[4] ;
reg [15:0] \ashr_16s_16ns_16_7_1_U3.dout_array[5] ;
reg [7:0] \ashr_32s_8ns_32_7_1_U7.din1_cast_array[0] ;
reg [7:0] \ashr_32s_8ns_32_7_1_U7.din1_cast_array[1] ;
reg [7:0] \ashr_32s_8ns_32_7_1_U7.din1_cast_array[2] ;
reg [7:0] \ashr_32s_8ns_32_7_1_U7.din1_cast_array[3] ;
reg [7:0] \ashr_32s_8ns_32_7_1_U7.din1_cast_array[4] ;
reg [7:0] \ashr_32s_8ns_32_7_1_U7.din1_cast_array[5] ;
reg [31:0] \ashr_32s_8ns_32_7_1_U7.dout_array[0] ;
reg [31:0] \ashr_32s_8ns_32_7_1_U7.dout_array[1] ;
reg [31:0] \ashr_32s_8ns_32_7_1_U7.dout_array[2] ;
reg [31:0] \ashr_32s_8ns_32_7_1_U7.dout_array[3] ;
reg [31:0] \ashr_32s_8ns_32_7_1_U7.dout_array[4] ;
reg [31:0] \ashr_32s_8ns_32_7_1_U7.dout_array[5] ;
reg [15:0] ashr_ln1497_reg_1251;
reg carry_1_reg_1432;
reg icmp_ln213_reg_1266;
reg icmp_ln768_reg_1130;
reg icmp_ln786_reg_1135;
reg op_12_V_reg_1297;
reg [1:0] op_16_V_reg_1382;
reg [1:0] op_19_V_reg_1522;
reg [16:0] op_23_V_reg_1422;
reg [31:0] op_29_V_reg_1543;
reg [3:0] op_7_V_reg_1271;
reg or_ln340_reg_1190;
reg or_ln384_reg_1502;
reg or_ln785_reg_1151;
reg or_ln786_reg_1163;
reg overflow_1_reg_1476;
reg p_Result_10_reg_1098;
reg p_Result_11_reg_1110;
reg p_Result_13_reg_1141;
reg p_Result_14_reg_1392;
reg p_Result_16_reg_1404;
reg [14:0] p_Result_1_reg_1117;
reg [2:0] p_Result_2_reg_1411;
reg [3:0] p_Result_3_reg_1416;
reg [3:0] p_Val2_1_reg_1224;
reg [1:0] p_Val2_5_reg_1332;
reg [1:0] p_Val2_6_reg_1398;
reg [15:0] r_reg_1277;
reg [16:0] ret_V_11_reg_1487;
reg [33:0] ret_V_12_reg_1558;
reg [5:0] ret_V_2_reg_1261;
reg [31:0] ret_V_6_cast_reg_1563;
reg [6:0] ret_V_8_reg_1212;
reg [5:0] ret_V_9_reg_1282;
reg [5:0] ret_V_reg_1217;
reg [16:0] ret_reg_1091;
reg sel_tmp11_reg_1235;
reg [3:0] select_ln340_reg_1230;
reg [3:0] select_ln785_reg_1246;
reg [7:0] sh_V_reg_1175;
reg [15:0] \shl_16s_16ns_16_7_1_U4.din1_cast_array[0] ;
reg [15:0] \shl_16s_16ns_16_7_1_U4.din1_cast_array[1] ;
reg [15:0] \shl_16s_16ns_16_7_1_U4.din1_cast_array[2] ;
reg [15:0] \shl_16s_16ns_16_7_1_U4.din1_cast_array[3] ;
reg [15:0] \shl_16s_16ns_16_7_1_U4.din1_cast_array[4] ;
reg [15:0] \shl_16s_16ns_16_7_1_U4.din1_cast_array[5] ;
reg [15:0] \shl_16s_16ns_16_7_1_U4.dout_array[0] ;
reg [15:0] \shl_16s_16ns_16_7_1_U4.dout_array[1] ;
reg [15:0] \shl_16s_16ns_16_7_1_U4.dout_array[2] ;
reg [15:0] \shl_16s_16ns_16_7_1_U4.dout_array[3] ;
reg [15:0] \shl_16s_16ns_16_7_1_U4.dout_array[4] ;
reg [15:0] \shl_16s_16ns_16_7_1_U4.dout_array[5] ;
reg [7:0] \shl_32s_8ns_32_7_1_U8.din1_cast_array[0] ;
reg [7:0] \shl_32s_8ns_32_7_1_U8.din1_cast_array[1] ;
reg [7:0] \shl_32s_8ns_32_7_1_U8.din1_cast_array[2] ;
reg [7:0] \shl_32s_8ns_32_7_1_U8.din1_cast_array[3] ;
reg [7:0] \shl_32s_8ns_32_7_1_U8.din1_cast_array[4] ;
reg [7:0] \shl_32s_8ns_32_7_1_U8.din1_cast_array[5] ;
reg [31:0] \shl_32s_8ns_32_7_1_U8.dout_array[0] ;
reg [31:0] \shl_32s_8ns_32_7_1_U8.dout_array[1] ;
reg [31:0] \shl_32s_8ns_32_7_1_U8.dout_array[2] ;
reg [31:0] \shl_32s_8ns_32_7_1_U8.dout_array[3] ;
reg [31:0] \shl_32s_8ns_32_7_1_U8.dout_array[4] ;
reg [31:0] \shl_32s_8ns_32_7_1_U8.dout_array[5] ;
reg [15:0] shl_ln1497_reg_1256;
reg [8:0] \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.ain_s1 ;
reg [8:0] \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.bin_s1 ;
reg \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.carry_s1 ;
reg [7:0] \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.sum_s1 ;
reg [2:0] \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.ain_s1 ;
reg [2:0] \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.bin_s1 ;
reg \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.carry_s1 ;
reg [1:0] \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.sum_s1 ;
reg [3:0] \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.ain_s1 ;
reg [3:0] \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.bin_s1 ;
reg \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.carry_s1 ;
reg [3:0] \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.sum_s1 ;
reg [4:0] sub_ln1497_reg_1048;
reg tmp_4_reg_1043;
reg trunc_ln1192_1_reg_1287;
reg [2:0] trunc_ln1192_2_reg_1292;
reg trunc_ln1192_4_reg_1085;
reg [1:0] trunc_ln69_1_reg_1352;
reg [1:0] trunc_ln69_reg_1347;
reg [1:0] trunc_ln731_reg_1105;
reg xor_ln785_reg_1157;
wire _000_;
wire _001_;
wire _002_;
wire [3:0] _003_;
wire [2:0] _004_;
wire [31:0] _005_;
wire [6:0] _006_;
wire [31:0] _007_;
wire [31:0] _008_;
wire [2:0] _009_;
wire [3:0] _010_;
wire [16:0] _011_;
wire _012_;
wire _013_;
wire [24:0] _014_;
wire [15:0] _015_;
wire _016_;
wire _017_;
wire _018_;
wire _019_;
wire _020_;
wire [1:0] _021_;
wire [1:0] _022_;
wire [16:0] _023_;
wire [31:0] _024_;
wire [3:0] _025_;
wire _026_;
wire _027_;
wire _028_;
wire _029_;
wire _030_;
wire _031_;
wire _032_;
wire _033_;
wire _034_;
wire _035_;
wire [14:0] _036_;
wire [2:0] _037_;
wire [3:0] _038_;
wire [1:0] _039_;
wire [1:0] _040_;
wire [1:0] _041_;
wire [15:0] _042_;
wire [16:0] _043_;
wire [33:0] _044_;
wire [5:0] _045_;
wire [31:0] _046_;
wire [6:0] _047_;
wire [5:0] _048_;
wire [5:0] _049_;
wire [16:0] _050_;
wire _051_;
wire [3:0] _052_;
wire [3:0] _053_;
wire [7:0] _054_;
wire [15:0] _055_;
wire [4:0] _056_;
wire _057_;
wire _058_;
wire [2:0] _059_;
wire _060_;
wire [1:0] _061_;
wire [1:0] _062_;
wire [1:0] _063_;
wire _064_;
wire [1:0] _065_;
wire _066_;
wire _067_;
wire _068_;
wire _069_;
wire _070_;
wire _071_;
wire _072_;
wire _073_;
wire _074_;
wire _075_;
wire _076_;
wire _077_;
wire _078_;
wire _079_;
wire [8:0] _080_;
wire [8:0] _081_;
wire _082_;
wire [7:0] _083_;
wire [8:0] _084_;
wire [9:0] _085_;
wire [8:0] _086_;
wire [8:0] _087_;
wire _088_;
wire [7:0] _089_;
wire [8:0] _090_;
wire [9:0] _091_;
wire [8:0] _092_;
wire [8:0] _093_;
wire _094_;
wire [7:0] _095_;
wire [8:0] _096_;
wire [9:0] _097_;
wire _098_;
wire _099_;
wire _100_;
wire _101_;
wire [1:0] _102_;
wire [1:0] _103_;
wire [15:0] _104_;
wire [15:0] _105_;
wire _106_;
wire [15:0] _107_;
wire [16:0] _108_;
wire [16:0] _109_;
wire [15:0] _110_;
wire [15:0] _111_;
wire _112_;
wire [15:0] _113_;
wire [16:0] _114_;
wire [16:0] _115_;
wire [15:0] _116_;
wire [15:0] _117_;
wire _118_;
wire [15:0] _119_;
wire [16:0] _120_;
wire [16:0] _121_;
wire [15:0] _122_;
wire [15:0] _123_;
wire _124_;
wire [15:0] _125_;
wire [16:0] _126_;
wire [16:0] _127_;
wire [16:0] _128_;
wire [16:0] _129_;
wire _130_;
wire [16:0] _131_;
wire [17:0] _132_;
wire [17:0] _133_;
wire [1:0] _134_;
wire [1:0] _135_;
wire _136_;
wire _137_;
wire [1:0] _138_;
wire [2:0] _139_;
wire [1:0] _140_;
wire [1:0] _141_;
wire _142_;
wire _143_;
wire [1:0] _144_;
wire [2:0] _145_;
wire [1:0] _146_;
wire [1:0] _147_;
wire _148_;
wire [1:0] _149_;
wire [2:0] _150_;
wire [2:0] _151_;
wire [1:0] _152_;
wire [1:0] _153_;
wire _154_;
wire [1:0] _155_;
wire [2:0] _156_;
wire [2:0] _157_;
wire [2:0] _158_;
wire [2:0] _159_;
wire _160_;
wire [2:0] _161_;
wire [3:0] _162_;
wire [3:0] _163_;
wire [3:0] _164_;
wire [3:0] _165_;
wire _166_;
wire [2:0] _167_;
wire [3:0] _168_;
wire [4:0] _169_;
wire [3:0] _170_;
wire [3:0] _171_;
wire _172_;
wire [2:0] _173_;
wire [3:0] _174_;
wire [4:0] _175_;
wire [3:0] _176_;
wire [3:0] _177_;
wire _178_;
wire [2:0] _179_;
wire [3:0] _180_;
wire [4:0] _181_;
wire [15:0] _182_;
wire [15:0] _183_;
wire [15:0] _184_;
wire [15:0] _185_;
wire [15:0] _186_;
wire [15:0] _187_;
wire [15:0] _188_;
wire [15:0] _189_;
wire [15:0] _190_;
wire [15:0] _191_;
wire [15:0] _192_;
wire [15:0] _193_;
wire [15:0] _194_;
wire [15:0] _195_;
wire [15:0] _196_;
wire [15:0] _197_;
wire [15:0] _198_;
wire [15:0] _199_;
wire [15:0] _200_;
wire [15:0] _201_;
wire [15:0] _202_;
wire [15:0] _203_;
wire [15:0] _204_;
wire [15:0] _205_;
wire [15:0] _206_;
wire [15:0] _207_;
wire [15:0] _208_;
wire [15:0] _209_;
wire [15:0] _210_;
wire [7:0] _211_;
wire [7:0] _212_;
wire [7:0] _213_;
wire [7:0] _214_;
wire [7:0] _215_;
wire [7:0] _216_;
wire [31:0] _217_;
wire [31:0] _218_;
wire [31:0] _219_;
wire [31:0] _220_;
wire [31:0] _221_;
wire [31:0] _222_;
wire [7:0] _223_;
wire [31:0] _224_;
wire [7:0] _225_;
wire [31:0] _226_;
wire [7:0] _227_;
wire [31:0] _228_;
wire [7:0] _229_;
wire [31:0] _230_;
wire [7:0] _231_;
wire [31:0] _232_;
wire [7:0] _233_;
wire [31:0] _234_;
wire [31:0] _235_;
wire [31:0] _236_;
wire [31:0] _237_;
wire [15:0] _238_;
wire [15:0] _239_;
wire [15:0] _240_;
wire [15:0] _241_;
wire [15:0] _242_;
wire [15:0] _243_;
wire [15:0] _244_;
wire [15:0] _245_;
wire [15:0] _246_;
wire [15:0] _247_;
wire [15:0] _248_;
wire [15:0] _249_;
wire [15:0] _250_;
wire [15:0] _251_;
wire [15:0] _252_;
wire [15:0] _253_;
wire [15:0] _254_;
wire [15:0] _255_;
wire [15:0] _256_;
wire [15:0] _257_;
wire [15:0] _258_;
wire [15:0] _259_;
wire [15:0] _260_;
wire [15:0] _261_;
wire [15:0] _262_;
wire [15:0] _263_;
wire [15:0] _264_;
wire [15:0] _265_;
wire [15:0] _266_;
wire [7:0] _267_;
wire [7:0] _268_;
wire [7:0] _269_;
wire [7:0] _270_;
wire [7:0] _271_;
wire [7:0] _272_;
wire [31:0] _273_;
wire [31:0] _274_;
wire [31:0] _275_;
wire [31:0] _276_;
wire [31:0] _277_;
wire [31:0] _278_;
wire [7:0] _279_;
wire [31:0] _280_;
wire [7:0] _281_;
wire [31:0] _282_;
wire [7:0] _283_;
wire [31:0] _284_;
wire [7:0] _285_;
wire [31:0] _286_;
wire [7:0] _287_;
wire [31:0] _288_;
wire [7:0] _289_;
wire [31:0] _290_;
wire [31:0] _291_;
wire [31:0] _292_;
wire [31:0] _293_;
wire [8:0] _294_;
wire [8:0] _295_;
wire _296_;
wire [7:0] _297_;
wire [8:0] _298_;
wire [9:0] _299_;
wire [2:0] _300_;
wire [2:0] _301_;
wire _302_;
wire [1:0] _303_;
wire [2:0] _304_;
wire [3:0] _305_;
wire [3:0] _306_;
wire [3:0] _307_;
wire _308_;
wire [3:0] _309_;
wire [4:0] _310_;
wire [4:0] _311_;
wire _312_;
wire _313_;
wire _314_;
wire _315_;
wire _316_;
wire _317_;
wire _318_;
wire _319_;
wire _320_;
wire _321_;
wire _322_;
wire _323_;
wire _324_;
wire _325_;
wire _326_;
wire _327_;
wire _328_;
wire _329_;
wire _330_;
wire _331_;
wire _332_;
wire _333_;
wire _334_;
wire _335_;
wire _336_;
wire _337_;
wire _338_;
wire _339_;
wire Range1_all_ones_fu_800_p2;
wire Range1_all_zeros_fu_805_p2;
wire Range2_all_ones_fu_795_p2;
wire \add_17ns_17s_17_2_1_U17.ce ;
wire \add_17ns_17s_17_2_1_U17.clk ;
wire [16:0] \add_17ns_17s_17_2_1_U17.din0 ;
wire [16:0] \add_17ns_17s_17_2_1_U17.din1 ;
wire [16:0] \add_17ns_17s_17_2_1_U17.dout ;
wire \add_17ns_17s_17_2_1_U17.reset ;
wire [16:0] \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.a ;
wire [16:0] \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.ain_s0 ;
wire [16:0] \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.b ;
wire [16:0] \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.bin_s0 ;
wire \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.ce ;
wire \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.clk ;
wire \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.facout_s1 ;
wire \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.facout_s2 ;
wire [7:0] \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.fas_s1 ;
wire [8:0] \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.fas_s2 ;
wire \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.reset ;
wire [16:0] \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.s ;
wire [7:0] \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.u1.a ;
wire [7:0] \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.u1.b ;
wire \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.u1.cin ;
wire \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.u1.cout ;
wire [7:0] \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.u1.s ;
wire [8:0] \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.u2.a ;
wire [8:0] \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.u2.b ;
wire \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.u2.cin ;
wire \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.u2.cout ;
wire [8:0] \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.u2.s ;
wire \add_17s_17ns_17_2_1_U16.ce ;
wire \add_17s_17ns_17_2_1_U16.clk ;
wire [16:0] \add_17s_17ns_17_2_1_U16.din0 ;
wire [16:0] \add_17s_17ns_17_2_1_U16.din1 ;
wire [16:0] \add_17s_17ns_17_2_1_U16.dout ;
wire \add_17s_17ns_17_2_1_U16.reset ;
wire [16:0] \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.a ;
wire [16:0] \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.ain_s0 ;
wire [16:0] \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.b ;
wire [16:0] \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.bin_s0 ;
wire \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.ce ;
wire \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.clk ;
wire \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.facout_s1 ;
wire \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.facout_s2 ;
wire [7:0] \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.fas_s1 ;
wire [8:0] \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.fas_s2 ;
wire \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.reset ;
wire [16:0] \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.s ;
wire [7:0] \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.u1.a ;
wire [7:0] \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.u1.b ;
wire \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.u1.cin ;
wire \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.u1.cout ;
wire [7:0] \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.u1.s ;
wire [8:0] \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.u2.a ;
wire [8:0] \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.u2.b ;
wire \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.u2.cin ;
wire \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.u2.cout ;
wire [8:0] \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.u2.s ;
wire \add_17s_17s_17_2_1_U11.ce ;
wire \add_17s_17s_17_2_1_U11.clk ;
wire [16:0] \add_17s_17s_17_2_1_U11.din0 ;
wire [16:0] \add_17s_17s_17_2_1_U11.din1 ;
wire [16:0] \add_17s_17s_17_2_1_U11.dout ;
wire \add_17s_17s_17_2_1_U11.reset ;
wire [16:0] \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.a ;
wire [16:0] \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.ain_s0 ;
wire [16:0] \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.b ;
wire [16:0] \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.bin_s0 ;
wire \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.ce ;
wire \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.clk ;
wire \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.facout_s1 ;
wire \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.facout_s2 ;
wire [7:0] \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.fas_s1 ;
wire [8:0] \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.fas_s2 ;
wire \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.reset ;
wire [16:0] \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.s ;
wire [7:0] \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.u1.a ;
wire [7:0] \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.u1.b ;
wire \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.u1.cin ;
wire \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.u1.cout ;
wire [7:0] \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.u1.s ;
wire [8:0] \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.u2.a ;
wire [8:0] \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.u2.b ;
wire \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.u2.cin ;
wire \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.u2.cout ;
wire [8:0] \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.u2.s ;
wire \add_2ns_2ns_2_2_1_U15.ce ;
wire \add_2ns_2ns_2_2_1_U15.clk ;
wire [1:0] \add_2ns_2ns_2_2_1_U15.din0 ;
wire [1:0] \add_2ns_2ns_2_2_1_U15.din1 ;
wire [1:0] \add_2ns_2ns_2_2_1_U15.dout ;
wire \add_2ns_2ns_2_2_1_U15.reset ;
wire [1:0] \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.a ;
wire [1:0] \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.ain_s0 ;
wire [1:0] \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.b ;
wire [1:0] \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.bin_s0 ;
wire \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.ce ;
wire \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.clk ;
wire \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.facout_s1 ;
wire \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.facout_s2 ;
wire \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.fas_s1 ;
wire \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.fas_s2 ;
wire \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.reset ;
wire [1:0] \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.s ;
wire \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.u1.a ;
wire \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.u1.b ;
wire \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.u1.cin ;
wire \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.u1.cout ;
wire \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.u1.s ;
wire \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.u2.a ;
wire \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.u2.b ;
wire \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.u2.cin ;
wire \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.u2.cout ;
wire \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.u2.s ;
wire \add_32ns_32ns_32_2_1_U24.ce ;
wire \add_32ns_32ns_32_2_1_U24.clk ;
wire [31:0] \add_32ns_32ns_32_2_1_U24.din0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U24.din1 ;
wire [31:0] \add_32ns_32ns_32_2_1_U24.dout ;
wire \add_32ns_32ns_32_2_1_U24.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.a ;
wire [31:0] \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.ain_s0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.b ;
wire [31:0] \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.bin_s0 ;
wire \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.ce ;
wire \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.clk ;
wire \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.facout_s1 ;
wire \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.facout_s2 ;
wire [15:0] \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.fas_s1 ;
wire [15:0] \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.fas_s2 ;
wire \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.u1.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.u1.b ;
wire \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.u1.cin ;
wire \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.u1.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.u1.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.u2.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.u2.b ;
wire \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.u2.cin ;
wire \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.u2.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.u2.s ;
wire \add_32ns_32s_32_2_1_U20.ce ;
wire \add_32ns_32s_32_2_1_U20.clk ;
wire [31:0] \add_32ns_32s_32_2_1_U20.din0 ;
wire [31:0] \add_32ns_32s_32_2_1_U20.din1 ;
wire [31:0] \add_32ns_32s_32_2_1_U20.dout ;
wire \add_32ns_32s_32_2_1_U20.reset ;
wire [31:0] \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.a ;
wire [31:0] \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.ain_s0 ;
wire [31:0] \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.b ;
wire [31:0] \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.bin_s0 ;
wire \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.ce ;
wire \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.clk ;
wire \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.facout_s1 ;
wire \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.facout_s2 ;
wire [15:0] \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.fas_s1 ;
wire [15:0] \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.fas_s2 ;
wire \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.reset ;
wire [31:0] \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.s ;
wire [15:0] \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.u1.a ;
wire [15:0] \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.u1.b ;
wire \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.u1.cin ;
wire \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.u1.cout ;
wire [15:0] \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.u1.s ;
wire [15:0] \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.u2.a ;
wire [15:0] \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.u2.b ;
wire \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.u2.cin ;
wire \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.u2.cout ;
wire [15:0] \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.u2.s ;
wire \add_32s_32ns_32_2_1_U18.ce ;
wire \add_32s_32ns_32_2_1_U18.clk ;
wire [31:0] \add_32s_32ns_32_2_1_U18.din0 ;
wire [31:0] \add_32s_32ns_32_2_1_U18.din1 ;
wire [31:0] \add_32s_32ns_32_2_1_U18.dout ;
wire \add_32s_32ns_32_2_1_U18.reset ;
wire [31:0] \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.a ;
wire [31:0] \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.ain_s0 ;
wire [31:0] \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.b ;
wire [31:0] \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.bin_s0 ;
wire \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.ce ;
wire \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.clk ;
wire \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.facout_s1 ;
wire \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.facout_s2 ;
wire [15:0] \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.fas_s1 ;
wire [15:0] \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.fas_s2 ;
wire \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.reset ;
wire [31:0] \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.s ;
wire [15:0] \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.u1.a ;
wire [15:0] \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.u1.b ;
wire \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.u1.cin ;
wire \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.u1.cout ;
wire [15:0] \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.u1.s ;
wire [15:0] \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.u2.a ;
wire [15:0] \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.u2.b ;
wire \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.u2.cin ;
wire \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.u2.cout ;
wire [15:0] \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.u2.s ;
wire \add_32s_32ns_32_2_1_U22.ce ;
wire \add_32s_32ns_32_2_1_U22.clk ;
wire [31:0] \add_32s_32ns_32_2_1_U22.din0 ;
wire [31:0] \add_32s_32ns_32_2_1_U22.din1 ;
wire [31:0] \add_32s_32ns_32_2_1_U22.dout ;
wire \add_32s_32ns_32_2_1_U22.reset ;
wire [31:0] \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.a ;
wire [31:0] \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.ain_s0 ;
wire [31:0] \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.b ;
wire [31:0] \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.bin_s0 ;
wire \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.ce ;
wire \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.clk ;
wire \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.facout_s1 ;
wire \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.facout_s2 ;
wire [15:0] \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.fas_s1 ;
wire [15:0] \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.fas_s2 ;
wire \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.reset ;
wire [31:0] \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.s ;
wire [15:0] \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.u1.a ;
wire [15:0] \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.u1.b ;
wire \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.u1.cin ;
wire \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.u1.cout ;
wire [15:0] \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.u1.s ;
wire [15:0] \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.u2.a ;
wire [15:0] \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.u2.b ;
wire \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.u2.cin ;
wire \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.u2.cout ;
wire [15:0] \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.u2.s ;
wire \add_34s_34s_34_2_1_U23.ce ;
wire \add_34s_34s_34_2_1_U23.clk ;
wire [33:0] \add_34s_34s_34_2_1_U23.din0 ;
wire [33:0] \add_34s_34s_34_2_1_U23.din1 ;
wire [33:0] \add_34s_34s_34_2_1_U23.dout ;
wire \add_34s_34s_34_2_1_U23.reset ;
wire [33:0] \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.a ;
wire [33:0] \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.ain_s0 ;
wire [33:0] \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.b ;
wire [33:0] \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.bin_s0 ;
wire \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.ce ;
wire \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.clk ;
wire \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.facout_s1 ;
wire \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.facout_s2 ;
wire [16:0] \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.fas_s1 ;
wire [16:0] \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.fas_s2 ;
wire \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.reset ;
wire [33:0] \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.s ;
wire [16:0] \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.u1.a ;
wire [16:0] \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.u1.b ;
wire \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.u1.cin ;
wire \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.u1.cout ;
wire [16:0] \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.u1.s ;
wire [16:0] \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.u2.a ;
wire [16:0] \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.u2.b ;
wire \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.u2.cin ;
wire \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.u2.cout ;
wire [16:0] \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.u2.s ;
wire \add_3ns_3ns_3_2_1_U10.ce ;
wire \add_3ns_3ns_3_2_1_U10.clk ;
wire [2:0] \add_3ns_3ns_3_2_1_U10.din0 ;
wire [2:0] \add_3ns_3ns_3_2_1_U10.din1 ;
wire [2:0] \add_3ns_3ns_3_2_1_U10.dout ;
wire \add_3ns_3ns_3_2_1_U10.reset ;
wire [2:0] \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.a ;
wire [2:0] \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.ain_s0 ;
wire [2:0] \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.b ;
wire [2:0] \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.bin_s0 ;
wire \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.ce ;
wire \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.clk ;
wire \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.facout_s1 ;
wire \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.facout_s2 ;
wire \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.fas_s1 ;
wire [1:0] \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.fas_s2 ;
wire \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.reset ;
wire [2:0] \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.s ;
wire \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.u1.a ;
wire \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.u1.b ;
wire \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.u1.cin ;
wire \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.u1.cout ;
wire \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.u1.s ;
wire [1:0] \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.u2.a ;
wire [1:0] \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.u2.b ;
wire \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.u2.cin ;
wire \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.u2.cout ;
wire [1:0] \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.u2.s ;
wire \add_3s_3s_3_2_1_U19.ce ;
wire \add_3s_3s_3_2_1_U19.clk ;
wire [2:0] \add_3s_3s_3_2_1_U19.din0 ;
wire [2:0] \add_3s_3s_3_2_1_U19.din1 ;
wire [2:0] \add_3s_3s_3_2_1_U19.dout ;
wire \add_3s_3s_3_2_1_U19.reset ;
wire [2:0] \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.a ;
wire [2:0] \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.ain_s0 ;
wire [2:0] \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.b ;
wire [2:0] \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.bin_s0 ;
wire \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.ce ;
wire \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.clk ;
wire \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.facout_s1 ;
wire \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.facout_s2 ;
wire \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.fas_s1 ;
wire [1:0] \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.fas_s2 ;
wire \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.reset ;
wire [2:0] \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.s ;
wire \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.u1.a ;
wire \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.u1.b ;
wire \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.u1.cin ;
wire \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.u1.cout ;
wire \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.u1.s ;
wire [1:0] \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.u2.a ;
wire [1:0] \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.u2.b ;
wire \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.u2.cin ;
wire \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.u2.cout ;
wire [1:0] \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.u2.s ;
wire \add_4ns_4s_4_2_1_U14.ce ;
wire \add_4ns_4s_4_2_1_U14.clk ;
wire [3:0] \add_4ns_4s_4_2_1_U14.din0 ;
wire [3:0] \add_4ns_4s_4_2_1_U14.din1 ;
wire [3:0] \add_4ns_4s_4_2_1_U14.dout ;
wire \add_4ns_4s_4_2_1_U14.reset ;
wire [3:0] \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.a ;
wire [3:0] \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.ain_s0 ;
wire [3:0] \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.b ;
wire [3:0] \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.bin_s0 ;
wire \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.ce ;
wire \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.clk ;
wire \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.facout_s1 ;
wire \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.facout_s2 ;
wire [1:0] \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.fas_s1 ;
wire [1:0] \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.fas_s2 ;
wire \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.reset ;
wire [3:0] \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.s ;
wire [1:0] \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.u1.a ;
wire [1:0] \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.u1.b ;
wire \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.u1.cin ;
wire \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.u1.cout ;
wire [1:0] \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.u1.s ;
wire [1:0] \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.u2.a ;
wire [1:0] \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.u2.b ;
wire \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.u2.cin ;
wire \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.u2.cout ;
wire [1:0] \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.u2.s ;
wire \add_4s_4s_4_2_1_U21.ce ;
wire \add_4s_4s_4_2_1_U21.clk ;
wire [3:0] \add_4s_4s_4_2_1_U21.din0 ;
wire [3:0] \add_4s_4s_4_2_1_U21.din1 ;
wire [3:0] \add_4s_4s_4_2_1_U21.dout ;
wire \add_4s_4s_4_2_1_U21.reset ;
wire [3:0] \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.a ;
wire [3:0] \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.ain_s0 ;
wire [3:0] \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.b ;
wire [3:0] \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.bin_s0 ;
wire \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.ce ;
wire \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.clk ;
wire \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.facout_s1 ;
wire \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.facout_s2 ;
wire [1:0] \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.fas_s1 ;
wire [1:0] \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.fas_s2 ;
wire \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.reset ;
wire [3:0] \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.s ;
wire [1:0] \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.u1.a ;
wire [1:0] \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.u1.b ;
wire \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.u1.cin ;
wire \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.u1.cout ;
wire [1:0] \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.u1.s ;
wire [1:0] \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.u2.a ;
wire [1:0] \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.u2.b ;
wire \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.u2.cin ;
wire \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.u2.cout ;
wire [1:0] \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.u2.s ;
wire \add_6ns_6ns_6_2_1_U9.ce ;
wire \add_6ns_6ns_6_2_1_U9.clk ;
wire [5:0] \add_6ns_6ns_6_2_1_U9.din0 ;
wire [5:0] \add_6ns_6ns_6_2_1_U9.din1 ;
wire [5:0] \add_6ns_6ns_6_2_1_U9.dout ;
wire \add_6ns_6ns_6_2_1_U9.reset ;
wire [5:0] \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.a ;
wire [5:0] \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.ain_s0 ;
wire [5:0] \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.b ;
wire [5:0] \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.bin_s0 ;
wire \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.ce ;
wire \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.clk ;
wire \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.facout_s1 ;
wire \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.facout_s2 ;
wire [2:0] \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.fas_s1 ;
wire [2:0] \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.fas_s2 ;
wire \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.reset ;
wire [5:0] \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.s ;
wire [2:0] \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.u1.a ;
wire [2:0] \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.u1.b ;
wire \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.u1.cin ;
wire \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.u1.cout ;
wire [2:0] \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.u1.s ;
wire [2:0] \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.u2.a ;
wire [2:0] \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.u2.b ;
wire \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.u2.cin ;
wire \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.u2.cout ;
wire [2:0] \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.u2.s ;
wire \add_7ns_7s_7_2_1_U6.ce ;
wire \add_7ns_7s_7_2_1_U6.clk ;
wire [6:0] \add_7ns_7s_7_2_1_U6.din0 ;
wire [6:0] \add_7ns_7s_7_2_1_U6.din1 ;
wire [6:0] \add_7ns_7s_7_2_1_U6.dout ;
wire \add_7ns_7s_7_2_1_U6.reset ;
wire [6:0] \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.a ;
wire [6:0] \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.ain_s0 ;
wire [6:0] \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.b ;
wire [6:0] \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.bin_s0 ;
wire \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.ce ;
wire \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.clk ;
wire \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.facout_s1 ;
wire \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.facout_s2 ;
wire [2:0] \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.fas_s1 ;
wire [3:0] \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.fas_s2 ;
wire \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.reset ;
wire [6:0] \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.s ;
wire [2:0] \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.u1.a ;
wire [2:0] \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.u1.b ;
wire \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.u1.cin ;
wire \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.u1.cout ;
wire [2:0] \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.u1.s ;
wire [3:0] \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.u2.a ;
wire [3:0] \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.u2.b ;
wire \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.u2.cin ;
wire \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.u2.cout ;
wire [3:0] \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.u2.s ;
wire \add_7s_7ns_7_2_1_U12.ce ;
wire \add_7s_7ns_7_2_1_U12.clk ;
wire [6:0] \add_7s_7ns_7_2_1_U12.din0 ;
wire [6:0] \add_7s_7ns_7_2_1_U12.din1 ;
wire [6:0] \add_7s_7ns_7_2_1_U12.dout ;
wire \add_7s_7ns_7_2_1_U12.reset ;
wire [6:0] \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.a ;
wire [6:0] \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.ain_s0 ;
wire [6:0] \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.b ;
wire [6:0] \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.bin_s0 ;
wire \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.ce ;
wire \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.clk ;
wire \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.facout_s1 ;
wire \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.facout_s2 ;
wire [2:0] \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.fas_s1 ;
wire [3:0] \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.fas_s2 ;
wire \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.reset ;
wire [6:0] \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.s ;
wire [2:0] \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.u1.a ;
wire [2:0] \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.u1.b ;
wire \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.u1.cin ;
wire \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.u1.cout ;
wire [2:0] \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.u1.s ;
wire [3:0] \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.u2.a ;
wire [3:0] \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.u2.b ;
wire \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.u2.cin ;
wire \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.u2.cout ;
wire [3:0] \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.u2.s ;
wire \add_7s_7s_7_2_1_U13.ce ;
wire \add_7s_7s_7_2_1_U13.clk ;
wire [6:0] \add_7s_7s_7_2_1_U13.din0 ;
wire [6:0] \add_7s_7s_7_2_1_U13.din1 ;
wire [6:0] \add_7s_7s_7_2_1_U13.dout ;
wire \add_7s_7s_7_2_1_U13.reset ;
wire [6:0] \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.a ;
wire [6:0] \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.ain_s0 ;
wire [6:0] \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.b ;
wire [6:0] \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.bin_s0 ;
wire \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.ce ;
wire \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.clk ;
wire \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.facout_s1 ;
wire \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.facout_s2 ;
wire [2:0] \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.fas_s1 ;
wire [3:0] \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.fas_s2 ;
wire \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.reset ;
wire [6:0] \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.s ;
wire [2:0] \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.u1.a ;
wire [2:0] \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.u1.b ;
wire \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.u1.cin ;
wire \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.u1.cout ;
wire [2:0] \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.u1.s ;
wire [3:0] \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.u2.a ;
wire [3:0] \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.u2.b ;
wire \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.u2.cin ;
wire \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.u2.cout ;
wire [3:0] \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.u2.s ;
wire and_ln213_fu_624_p2;
wire and_ln340_1_fu_506_p2;
wire and_ln340_fu_493_p2;
wire and_ln780_fu_860_p2;
wire and_ln781_fu_907_p2;
wire and_ln785_1_fu_510_p2;
wire and_ln785_fu_551_p2;
wire and_ln786_fu_365_p2;
wire and_ln788_1_fu_902_p2;
wire and_ln788_fu_896_p2;
wire ap_CS_fsm_state1;
wire ap_CS_fsm_state10;
wire ap_CS_fsm_state11;
wire ap_CS_fsm_state12;
wire ap_CS_fsm_state13;
wire ap_CS_fsm_state14;
wire ap_CS_fsm_state15;
wire ap_CS_fsm_state16;
wire ap_CS_fsm_state17;
wire ap_CS_fsm_state18;
wire ap_CS_fsm_state19;
wire ap_CS_fsm_state2;
wire ap_CS_fsm_state20;
wire ap_CS_fsm_state21;
wire ap_CS_fsm_state22;
wire ap_CS_fsm_state23;
wire ap_CS_fsm_state24;
wire ap_CS_fsm_state25;
wire ap_CS_fsm_state3;
wire ap_CS_fsm_state4;
wire ap_CS_fsm_state5;
wire ap_CS_fsm_state6;
wire ap_CS_fsm_state7;
wire ap_CS_fsm_state8;
wire ap_CS_fsm_state9;
wire [24:0] ap_NS_fsm;
wire ap_clk;
wire ap_done;
wire ap_idle;
wire ap_ready;
wire ap_rst;
wire ap_start;
wire \ashr_16s_16ns_16_7_1_U3.ce ;
wire \ashr_16s_16ns_16_7_1_U3.clk ;
wire [15:0] \ashr_16s_16ns_16_7_1_U3.din0 ;
wire [15:0] \ashr_16s_16ns_16_7_1_U3.din1 ;
wire [15:0] \ashr_16s_16ns_16_7_1_U3.din1_cast ;
wire [15:0] \ashr_16s_16ns_16_7_1_U3.din1_mask ;
wire [15:0] \ashr_16s_16ns_16_7_1_U3.dout ;
wire \ashr_16s_16ns_16_7_1_U3.reset ;
wire \ashr_32s_8ns_32_7_1_U7.ce ;
wire \ashr_32s_8ns_32_7_1_U7.clk ;
wire [31:0] \ashr_32s_8ns_32_7_1_U7.din0 ;
wire [31:0] \ashr_32s_8ns_32_7_1_U7.din1 ;
wire [7:0] \ashr_32s_8ns_32_7_1_U7.din1_cast ;
wire [7:0] \ashr_32s_8ns_32_7_1_U7.din1_mask ;
wire [31:0] \ashr_32s_8ns_32_7_1_U7.dout ;
wire \ashr_32s_8ns_32_7_1_U7.reset ;
wire carry_1_fu_789_p2;
wire deleted_ones_fu_865_p3;
wire deleted_zeros_fu_842_p3;
wire [31:0] grp_fu_1004_p2;
wire [4:0] grp_fu_237_p1;
wire [4:0] grp_fu_237_p2;
wire [16:0] grp_fu_251_p0;
wire [16:0] grp_fu_251_p1;
wire [16:0] grp_fu_251_p2;
wire [15:0] grp_fu_264_p1;
wire [15:0] grp_fu_264_p2;
wire [15:0] grp_fu_277_p1;
wire [15:0] grp_fu_277_p2;
wire [7:0] grp_fu_335_p2;
wire [6:0] grp_fu_386_p0;
wire [6:0] grp_fu_386_p1;
wire [6:0] grp_fu_386_p2;
wire [31:0] grp_fu_407_p1;
wire [31:0] grp_fu_407_p2;
wire [31:0] grp_fu_416_p1;
wire [31:0] grp_fu_416_p2;
wire [5:0] grp_fu_526_p2;
wire [2:0] grp_fu_648_p0;
wire [2:0] grp_fu_648_p2;
wire [16:0] grp_fu_660_p0;
wire [16:0] grp_fu_660_p1;
wire [16:0] grp_fu_660_p2;
wire [6:0] grp_fu_666_p0;
wire [6:0] grp_fu_666_p1;
wire [6:0] grp_fu_666_p2;
wire [6:0] grp_fu_709_p0;
wire [6:0] grp_fu_709_p1;
wire [6:0] grp_fu_709_p2;
wire [3:0] grp_fu_715_p0;
wire [3:0] grp_fu_715_p2;
wire [1:0] grp_fu_723_p1;
wire [1:0] grp_fu_723_p2;
wire [16:0] grp_fu_731_p0;
wire [16:0] grp_fu_731_p2;
wire [16:0] grp_fu_814_p1;
wire [16:0] grp_fu_814_p2;
wire [31:0] grp_fu_830_p0;
wire [31:0] grp_fu_830_p2;
wire [2:0] grp_fu_836_p0;
wire [2:0] grp_fu_836_p1;
wire [2:0] grp_fu_836_p2;
wire [31:0] grp_fu_939_p1;
wire [31:0] grp_fu_939_p2;
wire [3:0] grp_fu_947_p0;
wire [3:0] grp_fu_947_p1;
wire [3:0] grp_fu_947_p2;
wire [31:0] grp_fu_969_p0;
wire [31:0] grp_fu_969_p2;
wire [33:0] grp_fu_988_p0;
wire [33:0] grp_fu_988_p1;
wire [33:0] grp_fu_988_p2;
wire icmp_ln213_fu_562_p2;
wire icmp_ln768_fu_317_p2;
wire icmp_ln786_fu_322_p2;
wire [3:0] lhs_V_1_fu_690_p1;
wire [5:0] lhs_V_1_fu_690_p3;
wire [4:0] lhs_V_fu_370_p3;
wire [3:0] op_0;
wire [7:0] op_10;
wire op_12_V_fu_629_p2;
wire [1:0] op_13;
wire [1:0] op_14;
wire [31:0] op_15;
wire [1:0] op_16_V_fu_736_p3;
wire [1:0] op_17;
wire [1:0] op_18;
wire [1:0] op_19_V_fu_960_p3;
wire [15:0] op_2;
wire [3:0] op_3;
wire [31:0] op_30;
wire op_30_ap_vld;
wire [3:0] op_5;
wire [7:0] op_6;
wire [3:0] op_7_V_fu_568_p3;
wire [3:0] op_8;
wire [3:0] op_9;
wire or_ln213_fu_619_p2;
wire or_ln340_fu_396_p2;
wire or_ln384_fu_927_p2;
wire or_ln785_1_fu_877_p2;
wire or_ln785_2_fu_546_p2;
wire or_ln785_3_fu_514_p2;
wire or_ln785_fu_341_p2;
wire or_ln786_fu_355_p2;
wire or_ln788_fu_911_p2;
wire overflow_1_fu_887_p2;
wire overflow_fu_392_p2;
wire p_Result_12_fu_439_p3;
wire [7:0] p_Result_13_fu_327_p1;
wire p_Result_15_fu_777_p3;
wire p_Result_5_fu_578_p3;
wire p_Result_9_fu_1009_p3;
wire [3:0] p_Result_s_14_fu_478_p4;
wire [1:0] p_Result_s_fu_531_p4;
wire [3:0] p_Val2_1_fu_432_p3;
wire [2:0] p_Val2_2_fu_472_p2;
wire [15:0] r_fu_573_p3;
wire [5:0] ret_V_9_fu_594_p3;
wire [32:0] rhs_3_fu_977_p3;
wire sel_tmp11_fu_520_p2;
wire [3:0] select_ln340_fu_498_p3;
wire [1:0] select_ln384_fu_953_p3;
wire [3:0] select_ln785_fu_556_p3;
wire [31:0] select_ln850_1_fu_1019_p3;
wire [5:0] select_ln850_fu_588_p3;
wire [31:0] sext_ln1497_1_fu_270_p1;
wire [3:0] sext_ln1497_fu_225_p0;
wire [3:0] sext_ln215_1_fu_247_p0;
wire [15:0] sext_ln215_fu_243_p0;
wire [3:0] sext_ln545_fu_257_p0;
wire [31:0] sext_ln545_fu_257_p1;
wire [3:0] sext_ln703_fu_382_p0;
wire [7:0] sext_ln781_fu_401_p0;
wire [31:0] sext_ln781_fu_401_p1;
wire \shl_16s_16ns_16_7_1_U4.ce ;
wire \shl_16s_16ns_16_7_1_U4.clk ;
wire [15:0] \shl_16s_16ns_16_7_1_U4.din0 ;
wire [15:0] \shl_16s_16ns_16_7_1_U4.din1 ;
wire [15:0] \shl_16s_16ns_16_7_1_U4.din1_cast ;
wire [15:0] \shl_16s_16ns_16_7_1_U4.din1_mask ;
wire [15:0] \shl_16s_16ns_16_7_1_U4.dout ;
wire \shl_16s_16ns_16_7_1_U4.reset ;
wire \shl_32s_8ns_32_7_1_U8.ce ;
wire \shl_32s_8ns_32_7_1_U8.clk ;
wire [31:0] \shl_32s_8ns_32_7_1_U8.din0 ;
wire [31:0] \shl_32s_8ns_32_7_1_U8.din1 ;
wire [7:0] \shl_32s_8ns_32_7_1_U8.din1_cast ;
wire [7:0] \shl_32s_8ns_32_7_1_U8.din1_mask ;
wire [31:0] \shl_32s_8ns_32_7_1_U8.dout ;
wire \shl_32s_8ns_32_7_1_U8.reset ;
wire [3:0] shl_ln1192_fu_704_p0;
wire \sub_17s_17s_17_2_1_U2.ce ;
wire \sub_17s_17s_17_2_1_U2.clk ;
wire [16:0] \sub_17s_17s_17_2_1_U2.din0 ;
wire [16:0] \sub_17s_17s_17_2_1_U2.din1 ;
wire [16:0] \sub_17s_17s_17_2_1_U2.dout ;
wire \sub_17s_17s_17_2_1_U2.reset ;
wire [16:0] \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.a ;
wire [16:0] \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.ain_s0 ;
wire [16:0] \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.b ;
wire [16:0] \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.bin_s0 ;
wire \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.ce ;
wire \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.clk ;
wire \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.facout_s1 ;
wire \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.facout_s2 ;
wire [7:0] \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.fas_s1 ;
wire [8:0] \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.fas_s2 ;
wire \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.reset ;
wire [16:0] \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.s ;
wire [7:0] \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.u1.a ;
wire [7:0] \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.u1.b ;
wire \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.u1.cin ;
wire \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.u1.cout ;
wire [7:0] \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.u1.s ;
wire [8:0] \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.u2.a ;
wire [8:0] \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.u2.b ;
wire \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.u2.cin ;
wire \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.u2.cout ;
wire [8:0] \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.u2.s ;
wire \sub_5ns_5s_5_2_1_U1.ce ;
wire \sub_5ns_5s_5_2_1_U1.clk ;
wire [4:0] \sub_5ns_5s_5_2_1_U1.din0 ;
wire [4:0] \sub_5ns_5s_5_2_1_U1.din1 ;
wire [4:0] \sub_5ns_5s_5_2_1_U1.dout ;
wire \sub_5ns_5s_5_2_1_U1.reset ;
wire [4:0] \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.a ;
wire [4:0] \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.ain_s0 ;
wire [4:0] \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.b ;
wire [4:0] \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.bin_s0 ;
wire \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.ce ;
wire \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.clk ;
wire \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.facout_s1 ;
wire \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.facout_s2 ;
wire [1:0] \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.fas_s1 ;
wire [2:0] \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.fas_s2 ;
wire \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.reset ;
wire [4:0] \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.s ;
wire [1:0] \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.u1.a ;
wire [1:0] \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.u1.b ;
wire \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.u1.cin ;
wire \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.u1.cout ;
wire [1:0] \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.u1.s ;
wire [2:0] \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.u2.a ;
wire [2:0] \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.u2.b ;
wire \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.u2.cin ;
wire \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.u2.cout ;
wire [2:0] \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.u2.s ;
wire \sub_8ns_8s_8_2_1_U5.ce ;
wire \sub_8ns_8s_8_2_1_U5.clk ;
wire [7:0] \sub_8ns_8s_8_2_1_U5.din0 ;
wire [7:0] \sub_8ns_8s_8_2_1_U5.din1 ;
wire [7:0] \sub_8ns_8s_8_2_1_U5.dout ;
wire \sub_8ns_8s_8_2_1_U5.reset ;
wire [7:0] \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.a ;
wire [7:0] \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.ain_s0 ;
wire [7:0] \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.b ;
wire [7:0] \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.bin_s0 ;
wire \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.ce ;
wire \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.clk ;
wire \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.facout_s1 ;
wire \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.facout_s2 ;
wire [3:0] \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.fas_s1 ;
wire [3:0] \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.fas_s2 ;
wire \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.reset ;
wire [7:0] \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.s ;
wire [3:0] \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.u1.a ;
wire [3:0] \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.u1.b ;
wire \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.u1.cin ;
wire \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.u1.cout ;
wire [3:0] \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.u1.s ;
wire [3:0] \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.u2.a ;
wire [3:0] \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.u2.b ;
wire \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.u2.cin ;
wire \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.u2.cout ;
wire [3:0] \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.u2.s ;
wire tmp_10_fu_612_p3;
wire tmp_1_fu_453_p3;
wire [3:0] tmp_4_fu_229_p1;
wire tmp_9_fu_847_p3;
wire tmp_fu_446_p3;
wire trunc_ln1192_1_fu_604_p1;
wire [2:0] trunc_ln1192_2_fu_608_p1;
wire [3:0] trunc_ln1192_4_fu_283_p0;
wire trunc_ln1192_4_fu_283_p1;
wire trunc_ln1192_fu_601_p1;
wire [1:0] trunc_ln69_1_fu_686_p1;
wire [1:0] trunc_ln69_fu_682_p1;
wire [1:0] trunc_ln731_fu_295_p1;
wire trunc_ln790_fu_893_p1;
wire trunc_ln851_1_fu_1016_p1;
wire [3:0] trunc_ln851_fu_585_p0;
wire trunc_ln851_fu_585_p1;
wire underflow_1_fu_922_p2;
wire xor_ln340_fu_488_p2;
wire xor_ln365_1_fu_466_p2;
wire xor_ln365_fu_460_p2;
wire xor_ln416_fu_784_p2;
wire xor_ln780_fu_854_p2;
wire xor_ln785_1_fu_871_p2;
wire xor_ln785_2_fu_882_p2;
wire xor_ln785_3_fu_541_p2;
wire xor_ln785_fu_345_p2;
wire xor_ln786_1_fu_360_p2;
wire xor_ln786_fu_350_p2;
wire xor_ln788_fu_916_p2;
wire [7:0] zext_ln546_1_fu_413_p0;


assign _066_ = _073_ & ap_CS_fsm[8];
assign _067_ = ap_CS_fsm[8] & _074_;
assign _068_ = tmp_4_reg_1043 & ap_CS_fsm[8];
assign _069_ = ap_CS_fsm[12] & _075_;
assign _070_ = ap_CS_fsm[12] & p_Result_13_reg_1141;
assign _071_ = _076_ & ap_CS_fsm[0];
assign _072_ = ap_start & ap_CS_fsm[0];
assign and_ln213_fu_624_p2 = trunc_ln1192_4_reg_1085 & or_ln213_fu_619_p2;
assign and_ln340_1_fu_506_p2 = or_ln786_reg_1163 & or_ln340_reg_1190;
assign and_ln340_fu_493_p2 = xor_ln340_fu_488_p2 & or_ln786_reg_1163;
assign and_ln780_fu_860_p2 = xor_ln780_fu_854_p2 & Range2_all_ones_reg_1439;
assign and_ln781_fu_907_p2 = carry_1_reg_1432 & Range1_all_ones_reg_1444;
assign and_ln785_1_fu_510_p2 = xor_ln785_reg_1157 & and_ln786_reg_1169;
assign and_ln785_fu_551_p2 = or_ln785_2_fu_546_p2 & and_ln786_reg_1169;
assign and_ln786_fu_365_p2 = xor_ln786_1_fu_360_p2 & p_Result_11_reg_1110;
assign and_ln788_1_fu_902_p2 = p_Result_16_reg_1404 & and_ln788_fu_896_p2;
assign and_ln788_fu_896_p2 = p_Val2_6_reg_1398[0] & deleted_ones_fu_865_p3;
assign carry_1_fu_789_p2 = xor_ln416_fu_784_p2 & add_ln1192_2_reg_1327[2];
assign op_12_V_fu_629_p2 = op_0[0] & and_ln213_fu_624_p2;
assign overflow_1_fu_887_p2 = xor_ln785_2_fu_882_p2 & or_ln785_1_fu_877_p2;
assign overflow_fu_392_p2 = xor_ln785_reg_1157 & or_ln785_reg_1151;
assign sel_tmp11_fu_520_p2 = xor_ln365_1_fu_466_p2 & or_ln785_3_fu_514_p2;
assign underflow_1_fu_922_p2 = xor_ln788_fu_916_p2 & p_Result_14_reg_1392;
assign xor_ln340_fu_488_p2 = ~ or_ln340_reg_1190;
assign xor_ln780_fu_854_p2 = ~ add_ln1192_1_reg_1387[3];
assign xor_ln785_3_fu_541_p2 = ~ or_ln785_reg_1151;
assign xor_ln786_1_fu_360_p2 = ~ icmp_ln786_reg_1135;
assign xor_ln416_fu_784_p2 = ~ p_Result_16_reg_1404;
assign xor_ln788_fu_916_p2 = ~ or_ln788_fu_911_p2;
assign xor_ln785_1_fu_871_p2 = ~ deleted_zeros_fu_842_p3;
assign xor_ln786_fu_350_p2 = ~ p_Result_11_reg_1110;
assign xor_ln785_2_fu_882_p2 = ~ p_Result_14_reg_1392;
assign xor_ln365_1_fu_466_p2 = ~ xor_ln365_fu_460_p2;
assign xor_ln785_fu_345_p2 = ~ p_Result_10_reg_1098;
assign p_Val2_2_fu_472_p2 = ~ { trunc_ln731_reg_1105[0], 2'h0 };
assign _073_ = ~ tmp_4_reg_1043;
assign _074_ = ~ sel_tmp11_reg_1235;
assign _075_ = ~ p_Result_13_reg_1141;
assign _076_ = ~ ap_start;
assign _077_ = p_Result_3_reg_1416 == 4'hf;
assign _078_ = ! p_Result_3_reg_1416;
assign _079_ = p_Result_2_reg_1411 == 3'h7;
always @(posedge \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.clk )
\add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.bin_s1  <= _081_;
always @(posedge \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.clk )
\add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.ain_s1  <= _080_;
always @(posedge \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.clk )
\add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.sum_s1  <= _083_;
always @(posedge \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.clk )
\add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.carry_s1  <= _082_;
assign _081_ = \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.ce  ? \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.b [16:8] : \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.bin_s1 ;
assign _080_ = \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.ce  ? \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.a [16:8] : \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.ain_s1 ;
assign _082_ = \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.ce  ? \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.facout_s1  : \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.carry_s1 ;
assign _083_ = \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.ce  ? \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.fas_s1  : \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.sum_s1 ;
assign _084_ = \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.u1.a  + \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.u1.b ;
assign { \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.u1.cout , \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.u1.s  } = _084_ + \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.u1.cin ;
assign _085_ = \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.u2.a  + \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.u2.b ;
assign { \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.u2.cout , \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.u2.s  } = _085_ + \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.u2.cin ;
always @(posedge \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.clk )
\add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.bin_s1  <= _087_;
always @(posedge \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.clk )
\add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.ain_s1  <= _086_;
always @(posedge \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.clk )
\add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.sum_s1  <= _089_;
always @(posedge \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.clk )
\add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.carry_s1  <= _088_;
assign _087_ = \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.ce  ? \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.b [16:8] : \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.bin_s1 ;
assign _086_ = \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.ce  ? \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.a [16:8] : \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.ain_s1 ;
assign _088_ = \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.ce  ? \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.facout_s1  : \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.carry_s1 ;
assign _089_ = \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.ce  ? \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.fas_s1  : \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.sum_s1 ;
assign _090_ = \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.u1.a  + \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.u1.b ;
assign { \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.u1.cout , \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.u1.s  } = _090_ + \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.u1.cin ;
assign _091_ = \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.u2.a  + \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.u2.b ;
assign { \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.u2.cout , \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.u2.s  } = _091_ + \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.u2.cin ;
always @(posedge \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.clk )
\add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.bin_s1  <= _093_;
always @(posedge \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.clk )
\add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.ain_s1  <= _092_;
always @(posedge \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.clk )
\add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.sum_s1  <= _095_;
always @(posedge \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.clk )
\add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.carry_s1  <= _094_;
assign _093_ = \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.ce  ? \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.b [16:8] : \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.bin_s1 ;
assign _092_ = \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.ce  ? \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.a [16:8] : \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.ain_s1 ;
assign _094_ = \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.ce  ? \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.facout_s1  : \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.carry_s1 ;
assign _095_ = \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.ce  ? \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.fas_s1  : \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.sum_s1 ;
assign _096_ = \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.u1.a  + \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.u1.b ;
assign { \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.u1.cout , \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.u1.s  } = _096_ + \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.u1.cin ;
assign _097_ = \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.u2.a  + \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.u2.b ;
assign { \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.u2.cout , \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.u2.s  } = _097_ + \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.u2.cin ;
always @(posedge \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.clk )
\add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.bin_s1  <= _099_;
always @(posedge \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.clk )
\add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.ain_s1  <= _098_;
always @(posedge \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.clk )
\add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.sum_s1  <= _101_;
always @(posedge \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.clk )
\add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.carry_s1  <= _100_;
assign _099_ = \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.ce  ? \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.b [1] : \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.bin_s1 ;
assign _098_ = \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.ce  ? \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.a [1] : \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.ain_s1 ;
assign _100_ = \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.ce  ? \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.facout_s1  : \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.carry_s1 ;
assign _101_ = \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.ce  ? \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.fas_s1  : \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.sum_s1 ;
assign _102_ = \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.u1.a  + \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.u1.b ;
assign { \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.u1.cout , \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.u1.s  } = _102_ + \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.u1.cin ;
assign _103_ = \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.u2.a  + \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.u2.b ;
assign { \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.u2.cout , \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.u2.s  } = _103_ + \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.u2.cin ;
always @(posedge \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.clk )
\add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.bin_s1  <= _105_;
always @(posedge \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.clk )
\add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.ain_s1  <= _104_;
always @(posedge \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.clk )
\add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.sum_s1  <= _107_;
always @(posedge \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.clk )
\add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.carry_s1  <= _106_;
assign _105_ = \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.ce  ? \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.b [31:16] : \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.bin_s1 ;
assign _104_ = \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.ce  ? \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.a [31:16] : \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.ain_s1 ;
assign _106_ = \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.ce  ? \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.facout_s1  : \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.carry_s1 ;
assign _107_ = \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.ce  ? \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.fas_s1  : \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.sum_s1 ;
assign _108_ = \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.u1.a  + \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.u1.b ;
assign { \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.u1.cout , \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.u1.s  } = _108_ + \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.u1.cin ;
assign _109_ = \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.u2.a  + \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.u2.b ;
assign { \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.u2.cout , \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.u2.s  } = _109_ + \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.u2.cin ;
always @(posedge \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.clk )
\add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.bin_s1  <= _111_;
always @(posedge \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.clk )
\add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.ain_s1  <= _110_;
always @(posedge \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.clk )
\add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.sum_s1  <= _113_;
always @(posedge \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.clk )
\add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.carry_s1  <= _112_;
assign _111_ = \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.ce  ? \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.b [31:16] : \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.bin_s1 ;
assign _110_ = \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.ce  ? \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.a [31:16] : \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.ain_s1 ;
assign _112_ = \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.ce  ? \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.facout_s1  : \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.carry_s1 ;
assign _113_ = \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.ce  ? \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.fas_s1  : \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.sum_s1 ;
assign _114_ = \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.u1.a  + \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.u1.b ;
assign { \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.u1.cout , \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.u1.s  } = _114_ + \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.u1.cin ;
assign _115_ = \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.u2.a  + \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.u2.b ;
assign { \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.u2.cout , \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.u2.s  } = _115_ + \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.u2.cin ;
always @(posedge \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.clk )
\add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.bin_s1  <= _117_;
always @(posedge \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.clk )
\add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.ain_s1  <= _116_;
always @(posedge \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.clk )
\add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.sum_s1  <= _119_;
always @(posedge \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.clk )
\add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.carry_s1  <= _118_;
assign _117_ = \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.ce  ? \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.b [31:16] : \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.bin_s1 ;
assign _116_ = \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.ce  ? \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.a [31:16] : \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.ain_s1 ;
assign _118_ = \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.ce  ? \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.facout_s1  : \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.carry_s1 ;
assign _119_ = \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.ce  ? \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.fas_s1  : \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.sum_s1 ;
assign _120_ = \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.u1.a  + \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.u1.b ;
assign { \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.u1.cout , \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.u1.s  } = _120_ + \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.u1.cin ;
assign _121_ = \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.u2.a  + \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.u2.b ;
assign { \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.u2.cout , \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.u2.s  } = _121_ + \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.u2.cin ;
always @(posedge \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.clk )
\add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.bin_s1  <= _123_;
always @(posedge \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.clk )
\add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.ain_s1  <= _122_;
always @(posedge \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.clk )
\add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.sum_s1  <= _125_;
always @(posedge \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.clk )
\add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.carry_s1  <= _124_;
assign _123_ = \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.ce  ? \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.b [31:16] : \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.bin_s1 ;
assign _122_ = \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.ce  ? \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.a [31:16] : \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.ain_s1 ;
assign _124_ = \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.ce  ? \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.facout_s1  : \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.carry_s1 ;
assign _125_ = \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.ce  ? \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.fas_s1  : \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.sum_s1 ;
assign _126_ = \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.u1.a  + \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.u1.b ;
assign { \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.u1.cout , \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.u1.s  } = _126_ + \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.u1.cin ;
assign _127_ = \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.u2.a  + \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.u2.b ;
assign { \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.u2.cout , \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.u2.s  } = _127_ + \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.u2.cin ;
always @(posedge \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.clk )
\add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.bin_s1  <= _129_;
always @(posedge \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.clk )
\add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.ain_s1  <= _128_;
always @(posedge \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.clk )
\add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.sum_s1  <= _131_;
always @(posedge \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.clk )
\add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.carry_s1  <= _130_;
assign _129_ = \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.ce  ? \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.b [33:17] : \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.bin_s1 ;
assign _128_ = \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.ce  ? \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.a [33:17] : \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.ain_s1 ;
assign _130_ = \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.ce  ? \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.facout_s1  : \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.carry_s1 ;
assign _131_ = \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.ce  ? \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.fas_s1  : \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.sum_s1 ;
assign _132_ = \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.u1.a  + \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.u1.b ;
assign { \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.u1.cout , \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.u1.s  } = _132_ + \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.u1.cin ;
assign _133_ = \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.u2.a  + \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.u2.b ;
assign { \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.u2.cout , \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.u2.s  } = _133_ + \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.u2.cin ;
always @(posedge \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.clk )
\add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.bin_s1  <= _135_;
always @(posedge \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.clk )
\add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.ain_s1  <= _134_;
always @(posedge \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.clk )
\add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.sum_s1  <= _137_;
always @(posedge \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.clk )
\add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.carry_s1  <= _136_;
assign _135_ = \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.ce  ? \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.b [2:1] : \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.bin_s1 ;
assign _134_ = \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.ce  ? \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.a [2:1] : \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.ain_s1 ;
assign _136_ = \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.ce  ? \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.facout_s1  : \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.carry_s1 ;
assign _137_ = \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.ce  ? \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.fas_s1  : \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.sum_s1 ;
assign _138_ = \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.u1.a  + \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.u1.b ;
assign { \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.u1.cout , \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.u1.s  } = _138_ + \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.u1.cin ;
assign _139_ = \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.u2.a  + \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.u2.b ;
assign { \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.u2.cout , \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.u2.s  } = _139_ + \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.u2.cin ;
always @(posedge \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.clk )
\add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.bin_s1  <= _141_;
always @(posedge \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.clk )
\add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.ain_s1  <= _140_;
always @(posedge \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.clk )
\add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.sum_s1  <= _143_;
always @(posedge \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.clk )
\add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.carry_s1  <= _142_;
assign _141_ = \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.ce  ? \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.b [2:1] : \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.bin_s1 ;
assign _140_ = \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.ce  ? \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.a [2:1] : \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.ain_s1 ;
assign _142_ = \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.ce  ? \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.facout_s1  : \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.carry_s1 ;
assign _143_ = \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.ce  ? \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.fas_s1  : \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.sum_s1 ;
assign _144_ = \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.u1.a  + \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.u1.b ;
assign { \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.u1.cout , \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.u1.s  } = _144_ + \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.u1.cin ;
assign _145_ = \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.u2.a  + \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.u2.b ;
assign { \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.u2.cout , \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.u2.s  } = _145_ + \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.u2.cin ;
always @(posedge \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.clk )
\add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.bin_s1  <= _147_;
always @(posedge \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.clk )
\add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.ain_s1  <= _146_;
always @(posedge \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.clk )
\add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.sum_s1  <= _149_;
always @(posedge \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.clk )
\add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.carry_s1  <= _148_;
assign _147_ = \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.ce  ? \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.b [3:2] : \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.bin_s1 ;
assign _146_ = \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.ce  ? \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.a [3:2] : \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.ain_s1 ;
assign _148_ = \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.ce  ? \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.facout_s1  : \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.carry_s1 ;
assign _149_ = \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.ce  ? \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.fas_s1  : \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.sum_s1 ;
assign _150_ = \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.u1.a  + \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.u1.b ;
assign { \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.u1.cout , \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.u1.s  } = _150_ + \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.u1.cin ;
assign _151_ = \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.u2.a  + \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.u2.b ;
assign { \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.u2.cout , \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.u2.s  } = _151_ + \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.u2.cin ;
always @(posedge \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.clk )
\add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.bin_s1  <= _153_;
always @(posedge \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.clk )
\add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.ain_s1  <= _152_;
always @(posedge \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.clk )
\add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.sum_s1  <= _155_;
always @(posedge \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.clk )
\add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.carry_s1  <= _154_;
assign _153_ = \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.ce  ? \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.b [3:2] : \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.bin_s1 ;
assign _152_ = \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.ce  ? \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.a [3:2] : \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.ain_s1 ;
assign _154_ = \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.ce  ? \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.facout_s1  : \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.carry_s1 ;
assign _155_ = \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.ce  ? \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.fas_s1  : \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.sum_s1 ;
assign _156_ = \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.u1.a  + \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.u1.b ;
assign { \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.u1.cout , \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.u1.s  } = _156_ + \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.u1.cin ;
assign _157_ = \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.u2.a  + \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.u2.b ;
assign { \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.u2.cout , \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.u2.s  } = _157_ + \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.u2.cin ;
always @(posedge \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.clk )
\add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.bin_s1  <= _159_;
always @(posedge \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.clk )
\add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.ain_s1  <= _158_;
always @(posedge \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.clk )
\add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.sum_s1  <= _161_;
always @(posedge \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.clk )
\add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.carry_s1  <= _160_;
assign _159_ = \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.ce  ? \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.b [5:3] : \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.bin_s1 ;
assign _158_ = \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.ce  ? \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.a [5:3] : \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.ain_s1 ;
assign _160_ = \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.ce  ? \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.facout_s1  : \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.carry_s1 ;
assign _161_ = \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.ce  ? \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.fas_s1  : \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.sum_s1 ;
assign _162_ = \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.u1.a  + \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.u1.b ;
assign { \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.u1.cout , \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.u1.s  } = _162_ + \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.u1.cin ;
assign _163_ = \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.u2.a  + \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.u2.b ;
assign { \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.u2.cout , \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.u2.s  } = _163_ + \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.u2.cin ;
always @(posedge \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.clk )
\add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.bin_s1  <= _165_;
always @(posedge \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.clk )
\add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.ain_s1  <= _164_;
always @(posedge \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.clk )
\add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.sum_s1  <= _167_;
always @(posedge \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.clk )
\add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.carry_s1  <= _166_;
assign _165_ = \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.ce  ? \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.b [6:3] : \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.bin_s1 ;
assign _164_ = \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.ce  ? \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.a [6:3] : \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.ain_s1 ;
assign _166_ = \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.ce  ? \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.facout_s1  : \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.carry_s1 ;
assign _167_ = \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.ce  ? \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.fas_s1  : \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.sum_s1 ;
assign _168_ = \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.u1.a  + \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.u1.b ;
assign { \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.u1.cout , \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.u1.s  } = _168_ + \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.u1.cin ;
assign _169_ = \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.u2.a  + \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.u2.b ;
assign { \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.u2.cout , \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.u2.s  } = _169_ + \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.u2.cin ;
always @(posedge \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.clk )
\add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.bin_s1  <= _171_;
always @(posedge \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.clk )
\add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.ain_s1  <= _170_;
always @(posedge \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.clk )
\add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.sum_s1  <= _173_;
always @(posedge \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.clk )
\add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.carry_s1  <= _172_;
assign _171_ = \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.ce  ? \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.b [6:3] : \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.bin_s1 ;
assign _170_ = \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.ce  ? \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.a [6:3] : \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.ain_s1 ;
assign _172_ = \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.ce  ? \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.facout_s1  : \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.carry_s1 ;
assign _173_ = \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.ce  ? \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.fas_s1  : \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.sum_s1 ;
assign _174_ = \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.u1.a  + \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.u1.b ;
assign { \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.u1.cout , \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.u1.s  } = _174_ + \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.u1.cin ;
assign _175_ = \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.u2.a  + \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.u2.b ;
assign { \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.u2.cout , \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.u2.s  } = _175_ + \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.u2.cin ;
always @(posedge \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.clk )
\add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.bin_s1  <= _177_;
always @(posedge \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.clk )
\add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.ain_s1  <= _176_;
always @(posedge \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.clk )
\add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.sum_s1  <= _179_;
always @(posedge \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.clk )
\add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.carry_s1  <= _178_;
assign _177_ = \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.ce  ? \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.b [6:3] : \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.bin_s1 ;
assign _176_ = \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.ce  ? \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.a [6:3] : \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.ain_s1 ;
assign _178_ = \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.ce  ? \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.facout_s1  : \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.carry_s1 ;
assign _179_ = \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.ce  ? \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.fas_s1  : \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.sum_s1 ;
assign _180_ = \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.u1.a  + \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.u1.b ;
assign { \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.u1.cout , \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.u1.s  } = _180_ + \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.u1.cin ;
assign _181_ = \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.u2.a  + \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.u2.b ;
assign { \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.u2.cout , \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.u2.s  } = _181_ + \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.u2.cin ;
always @(posedge \ashr_16s_16ns_16_7_1_U3.clk )
\ashr_16s_16ns_16_7_1_U3.dout_array[5]  <= _193_;
always @(posedge \ashr_16s_16ns_16_7_1_U3.clk )
\ashr_16s_16ns_16_7_1_U3.din1_cast_array[5]  <= _187_;
always @(posedge \ashr_16s_16ns_16_7_1_U3.clk )
\ashr_16s_16ns_16_7_1_U3.dout_array[4]  <= _192_;
always @(posedge \ashr_16s_16ns_16_7_1_U3.clk )
\ashr_16s_16ns_16_7_1_U3.din1_cast_array[4]  <= _186_;
always @(posedge \ashr_16s_16ns_16_7_1_U3.clk )
\ashr_16s_16ns_16_7_1_U3.dout_array[3]  <= _191_;
always @(posedge \ashr_16s_16ns_16_7_1_U3.clk )
\ashr_16s_16ns_16_7_1_U3.din1_cast_array[3]  <= _185_;
always @(posedge \ashr_16s_16ns_16_7_1_U3.clk )
\ashr_16s_16ns_16_7_1_U3.dout_array[2]  <= _190_;
always @(posedge \ashr_16s_16ns_16_7_1_U3.clk )
\ashr_16s_16ns_16_7_1_U3.din1_cast_array[2]  <= _184_;
always @(posedge \ashr_16s_16ns_16_7_1_U3.clk )
\ashr_16s_16ns_16_7_1_U3.dout_array[1]  <= _189_;
always @(posedge \ashr_16s_16ns_16_7_1_U3.clk )
\ashr_16s_16ns_16_7_1_U3.din1_cast_array[1]  <= _183_;
always @(posedge \ashr_16s_16ns_16_7_1_U3.clk )
\ashr_16s_16ns_16_7_1_U3.dout_array[0]  <= _188_;
always @(posedge \ashr_16s_16ns_16_7_1_U3.clk )
\ashr_16s_16ns_16_7_1_U3.din1_cast_array[0]  <= _182_;
assign _194_ = \ashr_16s_16ns_16_7_1_U3.ce  ? \ashr_16s_16ns_16_7_1_U3.din1_cast_array[4]  : \ashr_16s_16ns_16_7_1_U3.din1_cast_array[5] ;
assign _187_ = \ashr_16s_16ns_16_7_1_U3.reset  ? 16'h0000 : _194_;
assign _195_ = \ashr_16s_16ns_16_7_1_U3.ce  ? _210_ : \ashr_16s_16ns_16_7_1_U3.dout_array[5] ;
assign _193_ = \ashr_16s_16ns_16_7_1_U3.reset  ? 16'h0000 : _195_;
assign _196_ = \ashr_16s_16ns_16_7_1_U3.ce  ? \ashr_16s_16ns_16_7_1_U3.din1_cast_array[3]  : \ashr_16s_16ns_16_7_1_U3.din1_cast_array[4] ;
assign _186_ = \ashr_16s_16ns_16_7_1_U3.reset  ? 16'h0000 : _196_;
assign _197_ = \ashr_16s_16ns_16_7_1_U3.ce  ? _209_ : \ashr_16s_16ns_16_7_1_U3.dout_array[4] ;
assign _192_ = \ashr_16s_16ns_16_7_1_U3.reset  ? 16'h0000 : _197_;
assign _198_ = \ashr_16s_16ns_16_7_1_U3.ce  ? \ashr_16s_16ns_16_7_1_U3.din1_cast_array[2]  : \ashr_16s_16ns_16_7_1_U3.din1_cast_array[3] ;
assign _185_ = \ashr_16s_16ns_16_7_1_U3.reset  ? 16'h0000 : _198_;
assign _199_ = \ashr_16s_16ns_16_7_1_U3.ce  ? _208_ : \ashr_16s_16ns_16_7_1_U3.dout_array[3] ;
assign _191_ = \ashr_16s_16ns_16_7_1_U3.reset  ? 16'h0000 : _199_;
assign _200_ = \ashr_16s_16ns_16_7_1_U3.ce  ? \ashr_16s_16ns_16_7_1_U3.din1_cast_array[1]  : \ashr_16s_16ns_16_7_1_U3.din1_cast_array[2] ;
assign _184_ = \ashr_16s_16ns_16_7_1_U3.reset  ? 16'h0000 : _200_;
assign _201_ = \ashr_16s_16ns_16_7_1_U3.ce  ? _207_ : \ashr_16s_16ns_16_7_1_U3.dout_array[2] ;
assign _190_ = \ashr_16s_16ns_16_7_1_U3.reset  ? 16'h0000 : _201_;
assign _202_ = \ashr_16s_16ns_16_7_1_U3.ce  ? \ashr_16s_16ns_16_7_1_U3.din1_cast_array[0]  : \ashr_16s_16ns_16_7_1_U3.din1_cast_array[1] ;
assign _183_ = \ashr_16s_16ns_16_7_1_U3.reset  ? 16'h0000 : _202_;
assign _203_ = \ashr_16s_16ns_16_7_1_U3.ce  ? _206_ : \ashr_16s_16ns_16_7_1_U3.dout_array[1] ;
assign _189_ = \ashr_16s_16ns_16_7_1_U3.reset  ? 16'h0000 : _203_;
assign _204_ = \ashr_16s_16ns_16_7_1_U3.ce  ? \ashr_16s_16ns_16_7_1_U3.din1  : \ashr_16s_16ns_16_7_1_U3.din1_cast_array[0] ;
assign _182_ = \ashr_16s_16ns_16_7_1_U3.reset  ? 16'h0000 : _204_;
assign _205_ = \ashr_16s_16ns_16_7_1_U3.ce  ? \ashr_16s_16ns_16_7_1_U3.din0  : \ashr_16s_16ns_16_7_1_U3.dout_array[0] ;
assign _188_ = \ashr_16s_16ns_16_7_1_U3.reset  ? 16'h0000 : _205_;
assign _206_ = $signed(\ashr_16s_16ns_16_7_1_U3.dout_array[0] ) >>> { \ashr_16s_16ns_16_7_1_U3.din1_cast_array[0] [15], 15'h0000 };
assign _207_ = $signed(\ashr_16s_16ns_16_7_1_U3.dout_array[1] ) >>> { \ashr_16s_16ns_16_7_1_U3.din1_cast_array[1] [14:12], 12'h000 };
assign _208_ = $signed(\ashr_16s_16ns_16_7_1_U3.dout_array[2] ) >>> { \ashr_16s_16ns_16_7_1_U3.din1_cast_array[2] [11:9], 9'h000 };
assign _209_ = $signed(\ashr_16s_16ns_16_7_1_U3.dout_array[3] ) >>> { \ashr_16s_16ns_16_7_1_U3.din1_cast_array[3] [8:6], 6'h00 };
assign _210_ = $signed(\ashr_16s_16ns_16_7_1_U3.dout_array[4] ) >>> { \ashr_16s_16ns_16_7_1_U3.din1_cast_array[4] [5:3], 3'h0 };
assign \ashr_16s_16ns_16_7_1_U3.dout  = $signed(\ashr_16s_16ns_16_7_1_U3.dout_array[5] ) >>> \ashr_16s_16ns_16_7_1_U3.din1_cast_array[5] [2:0];
always @(posedge \ashr_32s_8ns_32_7_1_U7.clk )
\ashr_32s_8ns_32_7_1_U7.dout_array[5]  <= _222_;
always @(posedge \ashr_32s_8ns_32_7_1_U7.clk )
\ashr_32s_8ns_32_7_1_U7.din1_cast_array[5]  <= _216_;
always @(posedge \ashr_32s_8ns_32_7_1_U7.clk )
\ashr_32s_8ns_32_7_1_U7.dout_array[4]  <= _221_;
always @(posedge \ashr_32s_8ns_32_7_1_U7.clk )
\ashr_32s_8ns_32_7_1_U7.din1_cast_array[4]  <= _215_;
always @(posedge \ashr_32s_8ns_32_7_1_U7.clk )
\ashr_32s_8ns_32_7_1_U7.dout_array[3]  <= _220_;
always @(posedge \ashr_32s_8ns_32_7_1_U7.clk )
\ashr_32s_8ns_32_7_1_U7.din1_cast_array[3]  <= _214_;
always @(posedge \ashr_32s_8ns_32_7_1_U7.clk )
\ashr_32s_8ns_32_7_1_U7.dout_array[2]  <= _219_;
always @(posedge \ashr_32s_8ns_32_7_1_U7.clk )
\ashr_32s_8ns_32_7_1_U7.din1_cast_array[2]  <= _213_;
always @(posedge \ashr_32s_8ns_32_7_1_U7.clk )
\ashr_32s_8ns_32_7_1_U7.dout_array[1]  <= _218_;
always @(posedge \ashr_32s_8ns_32_7_1_U7.clk )
\ashr_32s_8ns_32_7_1_U7.din1_cast_array[1]  <= _212_;
always @(posedge \ashr_32s_8ns_32_7_1_U7.clk )
\ashr_32s_8ns_32_7_1_U7.dout_array[0]  <= _217_;
always @(posedge \ashr_32s_8ns_32_7_1_U7.clk )
\ashr_32s_8ns_32_7_1_U7.din1_cast_array[0]  <= _211_;
assign _223_ = \ashr_32s_8ns_32_7_1_U7.ce  ? \ashr_32s_8ns_32_7_1_U7.din1_cast_array[4]  : \ashr_32s_8ns_32_7_1_U7.din1_cast_array[5] ;
assign _216_ = \ashr_32s_8ns_32_7_1_U7.reset  ? 8'h00 : _223_;
assign _224_ = \ashr_32s_8ns_32_7_1_U7.ce  ? _237_ : \ashr_32s_8ns_32_7_1_U7.dout_array[5] ;
assign _222_ = \ashr_32s_8ns_32_7_1_U7.reset  ? 32'd0 : _224_;
assign _225_ = \ashr_32s_8ns_32_7_1_U7.ce  ? \ashr_32s_8ns_32_7_1_U7.din1_cast_array[3]  : \ashr_32s_8ns_32_7_1_U7.din1_cast_array[4] ;
assign _215_ = \ashr_32s_8ns_32_7_1_U7.reset  ? 8'h00 : _225_;
assign _226_ = \ashr_32s_8ns_32_7_1_U7.ce  ? _236_ : \ashr_32s_8ns_32_7_1_U7.dout_array[4] ;
assign _221_ = \ashr_32s_8ns_32_7_1_U7.reset  ? 32'd0 : _226_;
assign _227_ = \ashr_32s_8ns_32_7_1_U7.ce  ? \ashr_32s_8ns_32_7_1_U7.din1_cast_array[2]  : \ashr_32s_8ns_32_7_1_U7.din1_cast_array[3] ;
assign _214_ = \ashr_32s_8ns_32_7_1_U7.reset  ? 8'h00 : _227_;
assign _228_ = \ashr_32s_8ns_32_7_1_U7.ce  ? _235_ : \ashr_32s_8ns_32_7_1_U7.dout_array[3] ;
assign _220_ = \ashr_32s_8ns_32_7_1_U7.reset  ? 32'd0 : _228_;
assign _229_ = \ashr_32s_8ns_32_7_1_U7.ce  ? \ashr_32s_8ns_32_7_1_U7.din1_cast_array[1]  : \ashr_32s_8ns_32_7_1_U7.din1_cast_array[2] ;
assign _213_ = \ashr_32s_8ns_32_7_1_U7.reset  ? 8'h00 : _229_;
assign _230_ = \ashr_32s_8ns_32_7_1_U7.ce  ? \ashr_32s_8ns_32_7_1_U7.dout_array[1]  : \ashr_32s_8ns_32_7_1_U7.dout_array[2] ;
assign _219_ = \ashr_32s_8ns_32_7_1_U7.reset  ? 32'd0 : _230_;
assign _231_ = \ashr_32s_8ns_32_7_1_U7.ce  ? \ashr_32s_8ns_32_7_1_U7.din1_cast_array[0]  : \ashr_32s_8ns_32_7_1_U7.din1_cast_array[1] ;
assign _212_ = \ashr_32s_8ns_32_7_1_U7.reset  ? 8'h00 : _231_;
assign _232_ = \ashr_32s_8ns_32_7_1_U7.ce  ? \ashr_32s_8ns_32_7_1_U7.dout_array[0]  : \ashr_32s_8ns_32_7_1_U7.dout_array[1] ;
assign _218_ = \ashr_32s_8ns_32_7_1_U7.reset  ? 32'd0 : _232_;
assign _233_ = \ashr_32s_8ns_32_7_1_U7.ce  ? \ashr_32s_8ns_32_7_1_U7.din1 [7:0] : \ashr_32s_8ns_32_7_1_U7.din1_cast_array[0] ;
assign _211_ = \ashr_32s_8ns_32_7_1_U7.reset  ? 8'h00 : _233_;
assign _234_ = \ashr_32s_8ns_32_7_1_U7.ce  ? \ashr_32s_8ns_32_7_1_U7.din0  : \ashr_32s_8ns_32_7_1_U7.dout_array[0] ;
assign _217_ = \ashr_32s_8ns_32_7_1_U7.reset  ? 32'd0 : _234_;
assign _235_ = $signed(\ashr_32s_8ns_32_7_1_U7.dout_array[2] ) >>> { \ashr_32s_8ns_32_7_1_U7.din1_cast_array[2] [7:6], 6'h00 };
assign _236_ = $signed(\ashr_32s_8ns_32_7_1_U7.dout_array[3] ) >>> { \ashr_32s_8ns_32_7_1_U7.din1_cast_array[3] [5:4], 4'h0 };
assign _237_ = $signed(\ashr_32s_8ns_32_7_1_U7.dout_array[4] ) >>> { \ashr_32s_8ns_32_7_1_U7.din1_cast_array[4] [3:2], 2'h0 };
assign \ashr_32s_8ns_32_7_1_U7.dout  = $signed(\ashr_32s_8ns_32_7_1_U7.dout_array[5] ) >>> \ashr_32s_8ns_32_7_1_U7.din1_cast_array[5] [1:0];
always @(posedge \shl_16s_16ns_16_7_1_U4.clk )
\shl_16s_16ns_16_7_1_U4.dout_array[5]  <= _249_;
always @(posedge \shl_16s_16ns_16_7_1_U4.clk )
\shl_16s_16ns_16_7_1_U4.din1_cast_array[5]  <= _243_;
always @(posedge \shl_16s_16ns_16_7_1_U4.clk )
\shl_16s_16ns_16_7_1_U4.dout_array[4]  <= _248_;
always @(posedge \shl_16s_16ns_16_7_1_U4.clk )
\shl_16s_16ns_16_7_1_U4.din1_cast_array[4]  <= _242_;
always @(posedge \shl_16s_16ns_16_7_1_U4.clk )
\shl_16s_16ns_16_7_1_U4.dout_array[3]  <= _247_;
always @(posedge \shl_16s_16ns_16_7_1_U4.clk )
\shl_16s_16ns_16_7_1_U4.din1_cast_array[3]  <= _241_;
always @(posedge \shl_16s_16ns_16_7_1_U4.clk )
\shl_16s_16ns_16_7_1_U4.dout_array[2]  <= _246_;
always @(posedge \shl_16s_16ns_16_7_1_U4.clk )
\shl_16s_16ns_16_7_1_U4.din1_cast_array[2]  <= _240_;
always @(posedge \shl_16s_16ns_16_7_1_U4.clk )
\shl_16s_16ns_16_7_1_U4.dout_array[1]  <= _245_;
always @(posedge \shl_16s_16ns_16_7_1_U4.clk )
\shl_16s_16ns_16_7_1_U4.din1_cast_array[1]  <= _239_;
always @(posedge \shl_16s_16ns_16_7_1_U4.clk )
\shl_16s_16ns_16_7_1_U4.dout_array[0]  <= _244_;
always @(posedge \shl_16s_16ns_16_7_1_U4.clk )
\shl_16s_16ns_16_7_1_U4.din1_cast_array[0]  <= _238_;
assign _250_ = \shl_16s_16ns_16_7_1_U4.ce  ? \shl_16s_16ns_16_7_1_U4.din1_cast_array[4]  : \shl_16s_16ns_16_7_1_U4.din1_cast_array[5] ;
assign _243_ = \shl_16s_16ns_16_7_1_U4.reset  ? 16'h0000 : _250_;
assign _251_ = \shl_16s_16ns_16_7_1_U4.ce  ? _266_ : \shl_16s_16ns_16_7_1_U4.dout_array[5] ;
assign _249_ = \shl_16s_16ns_16_7_1_U4.reset  ? 16'h0000 : _251_;
assign _252_ = \shl_16s_16ns_16_7_1_U4.ce  ? \shl_16s_16ns_16_7_1_U4.din1_cast_array[3]  : \shl_16s_16ns_16_7_1_U4.din1_cast_array[4] ;
assign _242_ = \shl_16s_16ns_16_7_1_U4.reset  ? 16'h0000 : _252_;
assign _253_ = \shl_16s_16ns_16_7_1_U4.ce  ? _265_ : \shl_16s_16ns_16_7_1_U4.dout_array[4] ;
assign _248_ = \shl_16s_16ns_16_7_1_U4.reset  ? 16'h0000 : _253_;
assign _254_ = \shl_16s_16ns_16_7_1_U4.ce  ? \shl_16s_16ns_16_7_1_U4.din1_cast_array[2]  : \shl_16s_16ns_16_7_1_U4.din1_cast_array[3] ;
assign _241_ = \shl_16s_16ns_16_7_1_U4.reset  ? 16'h0000 : _254_;
assign _255_ = \shl_16s_16ns_16_7_1_U4.ce  ? _264_ : \shl_16s_16ns_16_7_1_U4.dout_array[3] ;
assign _247_ = \shl_16s_16ns_16_7_1_U4.reset  ? 16'h0000 : _255_;
assign _256_ = \shl_16s_16ns_16_7_1_U4.ce  ? \shl_16s_16ns_16_7_1_U4.din1_cast_array[1]  : \shl_16s_16ns_16_7_1_U4.din1_cast_array[2] ;
assign _240_ = \shl_16s_16ns_16_7_1_U4.reset  ? 16'h0000 : _256_;
assign _257_ = \shl_16s_16ns_16_7_1_U4.ce  ? _263_ : \shl_16s_16ns_16_7_1_U4.dout_array[2] ;
assign _246_ = \shl_16s_16ns_16_7_1_U4.reset  ? 16'h0000 : _257_;
assign _258_ = \shl_16s_16ns_16_7_1_U4.ce  ? \shl_16s_16ns_16_7_1_U4.din1_cast_array[0]  : \shl_16s_16ns_16_7_1_U4.din1_cast_array[1] ;
assign _239_ = \shl_16s_16ns_16_7_1_U4.reset  ? 16'h0000 : _258_;
assign _259_ = \shl_16s_16ns_16_7_1_U4.ce  ? _262_ : \shl_16s_16ns_16_7_1_U4.dout_array[1] ;
assign _245_ = \shl_16s_16ns_16_7_1_U4.reset  ? 16'h0000 : _259_;
assign _260_ = \shl_16s_16ns_16_7_1_U4.ce  ? \shl_16s_16ns_16_7_1_U4.din1  : \shl_16s_16ns_16_7_1_U4.din1_cast_array[0] ;
assign _238_ = \shl_16s_16ns_16_7_1_U4.reset  ? 16'h0000 : _260_;
assign _261_ = \shl_16s_16ns_16_7_1_U4.ce  ? \shl_16s_16ns_16_7_1_U4.din0  : \shl_16s_16ns_16_7_1_U4.dout_array[0] ;
assign _244_ = \shl_16s_16ns_16_7_1_U4.reset  ? 16'h0000 : _261_;
assign _262_ = \shl_16s_16ns_16_7_1_U4.dout_array[0]  << { \shl_16s_16ns_16_7_1_U4.din1_cast_array[0] [15], 15'h0000 };
assign _263_ = \shl_16s_16ns_16_7_1_U4.dout_array[1]  << { \shl_16s_16ns_16_7_1_U4.din1_cast_array[1] [14:12], 12'h000 };
assign _264_ = \shl_16s_16ns_16_7_1_U4.dout_array[2]  << { \shl_16s_16ns_16_7_1_U4.din1_cast_array[2] [11:9], 9'h000 };
assign _265_ = \shl_16s_16ns_16_7_1_U4.dout_array[3]  << { \shl_16s_16ns_16_7_1_U4.din1_cast_array[3] [8:6], 6'h00 };
assign _266_ = \shl_16s_16ns_16_7_1_U4.dout_array[4]  << { \shl_16s_16ns_16_7_1_U4.din1_cast_array[4] [5:3], 3'h0 };
assign \shl_16s_16ns_16_7_1_U4.dout  = \shl_16s_16ns_16_7_1_U4.dout_array[5]  << \shl_16s_16ns_16_7_1_U4.din1_cast_array[5] [2:0];
always @(posedge \shl_32s_8ns_32_7_1_U8.clk )
\shl_32s_8ns_32_7_1_U8.dout_array[5]  <= _278_;
always @(posedge \shl_32s_8ns_32_7_1_U8.clk )
\shl_32s_8ns_32_7_1_U8.din1_cast_array[5]  <= _272_;
always @(posedge \shl_32s_8ns_32_7_1_U8.clk )
\shl_32s_8ns_32_7_1_U8.dout_array[4]  <= _277_;
always @(posedge \shl_32s_8ns_32_7_1_U8.clk )
\shl_32s_8ns_32_7_1_U8.din1_cast_array[4]  <= _271_;
always @(posedge \shl_32s_8ns_32_7_1_U8.clk )
\shl_32s_8ns_32_7_1_U8.dout_array[3]  <= _276_;
always @(posedge \shl_32s_8ns_32_7_1_U8.clk )
\shl_32s_8ns_32_7_1_U8.din1_cast_array[3]  <= _270_;
always @(posedge \shl_32s_8ns_32_7_1_U8.clk )
\shl_32s_8ns_32_7_1_U8.dout_array[2]  <= _275_;
always @(posedge \shl_32s_8ns_32_7_1_U8.clk )
\shl_32s_8ns_32_7_1_U8.din1_cast_array[2]  <= _269_;
always @(posedge \shl_32s_8ns_32_7_1_U8.clk )
\shl_32s_8ns_32_7_1_U8.dout_array[1]  <= _274_;
always @(posedge \shl_32s_8ns_32_7_1_U8.clk )
\shl_32s_8ns_32_7_1_U8.din1_cast_array[1]  <= _268_;
always @(posedge \shl_32s_8ns_32_7_1_U8.clk )
\shl_32s_8ns_32_7_1_U8.dout_array[0]  <= _273_;
always @(posedge \shl_32s_8ns_32_7_1_U8.clk )
\shl_32s_8ns_32_7_1_U8.din1_cast_array[0]  <= _267_;
assign _279_ = \shl_32s_8ns_32_7_1_U8.ce  ? \shl_32s_8ns_32_7_1_U8.din1_cast_array[4]  : \shl_32s_8ns_32_7_1_U8.din1_cast_array[5] ;
assign _272_ = \shl_32s_8ns_32_7_1_U8.reset  ? 8'h00 : _279_;
assign _280_ = \shl_32s_8ns_32_7_1_U8.ce  ? _293_ : \shl_32s_8ns_32_7_1_U8.dout_array[5] ;
assign _278_ = \shl_32s_8ns_32_7_1_U8.reset  ? 32'd0 : _280_;
assign _281_ = \shl_32s_8ns_32_7_1_U8.ce  ? \shl_32s_8ns_32_7_1_U8.din1_cast_array[3]  : \shl_32s_8ns_32_7_1_U8.din1_cast_array[4] ;
assign _271_ = \shl_32s_8ns_32_7_1_U8.reset  ? 8'h00 : _281_;
assign _282_ = \shl_32s_8ns_32_7_1_U8.ce  ? _292_ : \shl_32s_8ns_32_7_1_U8.dout_array[4] ;
assign _277_ = \shl_32s_8ns_32_7_1_U8.reset  ? 32'd0 : _282_;
assign _283_ = \shl_32s_8ns_32_7_1_U8.ce  ? \shl_32s_8ns_32_7_1_U8.din1_cast_array[2]  : \shl_32s_8ns_32_7_1_U8.din1_cast_array[3] ;
assign _270_ = \shl_32s_8ns_32_7_1_U8.reset  ? 8'h00 : _283_;
assign _284_ = \shl_32s_8ns_32_7_1_U8.ce  ? _291_ : \shl_32s_8ns_32_7_1_U8.dout_array[3] ;
assign _276_ = \shl_32s_8ns_32_7_1_U8.reset  ? 32'd0 : _284_;
assign _285_ = \shl_32s_8ns_32_7_1_U8.ce  ? \shl_32s_8ns_32_7_1_U8.din1_cast_array[1]  : \shl_32s_8ns_32_7_1_U8.din1_cast_array[2] ;
assign _269_ = \shl_32s_8ns_32_7_1_U8.reset  ? 8'h00 : _285_;
assign _286_ = \shl_32s_8ns_32_7_1_U8.ce  ? \shl_32s_8ns_32_7_1_U8.dout_array[1]  : \shl_32s_8ns_32_7_1_U8.dout_array[2] ;
assign _275_ = \shl_32s_8ns_32_7_1_U8.reset  ? 32'd0 : _286_;
assign _287_ = \shl_32s_8ns_32_7_1_U8.ce  ? \shl_32s_8ns_32_7_1_U8.din1_cast_array[0]  : \shl_32s_8ns_32_7_1_U8.din1_cast_array[1] ;
assign _268_ = \shl_32s_8ns_32_7_1_U8.reset  ? 8'h00 : _287_;
assign _288_ = \shl_32s_8ns_32_7_1_U8.ce  ? \shl_32s_8ns_32_7_1_U8.dout_array[0]  : \shl_32s_8ns_32_7_1_U8.dout_array[1] ;
assign _274_ = \shl_32s_8ns_32_7_1_U8.reset  ? 32'd0 : _288_;
assign _289_ = \shl_32s_8ns_32_7_1_U8.ce  ? \shl_32s_8ns_32_7_1_U8.din1 [7:0] : \shl_32s_8ns_32_7_1_U8.din1_cast_array[0] ;
assign _267_ = \shl_32s_8ns_32_7_1_U8.reset  ? 8'h00 : _289_;
assign _290_ = \shl_32s_8ns_32_7_1_U8.ce  ? \shl_32s_8ns_32_7_1_U8.din0  : \shl_32s_8ns_32_7_1_U8.dout_array[0] ;
assign _273_ = \shl_32s_8ns_32_7_1_U8.reset  ? 32'd0 : _290_;
assign _291_ = \shl_32s_8ns_32_7_1_U8.dout_array[2]  << { \shl_32s_8ns_32_7_1_U8.din1_cast_array[2] [7:6], 6'h00 };
assign _292_ = \shl_32s_8ns_32_7_1_U8.dout_array[3]  << { \shl_32s_8ns_32_7_1_U8.din1_cast_array[3] [5:4], 4'h0 };
assign _293_ = \shl_32s_8ns_32_7_1_U8.dout_array[4]  << { \shl_32s_8ns_32_7_1_U8.din1_cast_array[4] [3:2], 2'h0 };
assign \shl_32s_8ns_32_7_1_U8.dout  = \shl_32s_8ns_32_7_1_U8.dout_array[5]  << \shl_32s_8ns_32_7_1_U8.din1_cast_array[5] [1:0];
assign \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.bin_s0  = ~ \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.b ;
always @(posedge \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.clk )
\sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.bin_s1  <= _295_;
always @(posedge \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.clk )
\sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.ain_s1  <= _294_;
always @(posedge \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.clk )
\sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.sum_s1  <= _297_;
always @(posedge \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.clk )
\sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.carry_s1  <= _296_;
assign _295_ = \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.ce  ? \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.bin_s0 [16:8] : \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.bin_s1 ;
assign _294_ = \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.ce  ? \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.a [16:8] : \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.ain_s1 ;
assign _296_ = \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.ce  ? \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.facout_s1  : \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.carry_s1 ;
assign _297_ = \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.ce  ? \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.fas_s1  : \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.sum_s1 ;
assign _298_ = \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.u1.a  + \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.u1.b ;
assign { \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.u1.cout , \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.u1.s  } = _298_ + \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.u1.cin ;
assign _299_ = \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.u2.a  + \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.u2.b ;
assign { \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.u2.cout , \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.u2.s  } = _299_ + \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.u2.cin ;
assign \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.bin_s0  = ~ \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.b ;
always @(posedge \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.clk )
\sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.bin_s1  <= _301_;
always @(posedge \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.clk )
\sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.ain_s1  <= _300_;
always @(posedge \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.clk )
\sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.sum_s1  <= _303_;
always @(posedge \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.clk )
\sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.carry_s1  <= _302_;
assign _301_ = \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.ce  ? \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.bin_s0 [4:2] : \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.bin_s1 ;
assign _300_ = \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.ce  ? \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.a [4:2] : \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.ain_s1 ;
assign _302_ = \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.ce  ? \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.facout_s1  : \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.carry_s1 ;
assign _303_ = \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.ce  ? \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.fas_s1  : \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.sum_s1 ;
assign _304_ = \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.u1.a  + \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.u1.b ;
assign { \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.u1.cout , \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.u1.s  } = _304_ + \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.u1.cin ;
assign _305_ = \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.u2.a  + \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.u2.b ;
assign { \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.u2.cout , \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.u2.s  } = _305_ + \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.u2.cin ;
assign \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.bin_s0  = ~ \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.b ;
always @(posedge \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.clk )
\sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.bin_s1  <= _307_;
always @(posedge \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.clk )
\sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.ain_s1  <= _306_;
always @(posedge \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.clk )
\sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.sum_s1  <= _309_;
always @(posedge \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.clk )
\sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.carry_s1  <= _308_;
assign _307_ = \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.ce  ? \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.bin_s0 [7:4] : \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.bin_s1 ;
assign _306_ = \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.ce  ? \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.a [7:4] : \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.ain_s1 ;
assign _308_ = \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.ce  ? \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.facout_s1  : \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.carry_s1 ;
assign _309_ = \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.ce  ? \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.fas_s1  : \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.sum_s1 ;
assign _310_ = \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.u1.a  + \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.u1.b ;
assign { \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.u1.cout , \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.u1.s  } = _310_ + \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.u1.cin ;
assign _311_ = \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.u2.a  + \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.u2.b ;
assign { \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.u2.cout , \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.u2.s  } = _311_ + \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.u2.cin ;
assign _312_ = | op_0[3:2];
assign _313_ = | p_Result_1_reg_1117;
assign _314_ = p_Result_1_reg_1117 != 15'h7fff;
assign or_ln213_fu_619_p2 = op_0[1] | icmp_ln213_reg_1266;
assign or_ln340_fu_396_p2 = p_Result_10_reg_1098 | overflow_fu_392_p2;
assign or_ln384_fu_927_p2 = underflow_1_fu_922_p2 | overflow_1_reg_1476;
assign or_ln785_1_fu_877_p2 = xor_ln785_1_fu_871_p2 | p_Result_16_reg_1404;
assign or_ln785_2_fu_546_p2 = xor_ln785_3_fu_541_p2 | p_Result_10_reg_1098;
assign or_ln785_3_fu_514_p2 = and_ln785_1_fu_510_p2 | and_ln340_1_fu_506_p2;
assign or_ln785_fu_341_p2 = p_Result_11_reg_1110 | icmp_ln768_reg_1130;
assign or_ln786_fu_355_p2 = xor_ln786_fu_350_p2 | icmp_ln786_reg_1135;
assign or_ln788_fu_911_p2 = and_ln788_1_reg_1482 | and_ln781_fu_907_p2;
always @(posedge ap_clk)
trunc_ln1192_4_reg_1085 <= _060_;
always @(posedge ap_clk)
tmp_4_reg_1043 <= _057_;
always @(posedge ap_clk)
sub_ln1497_reg_1048 <= _056_;
always @(posedge ap_clk)
shl_ln1497_reg_1256 <= _055_;
always @(posedge ap_clk)
select_ln785_reg_1246 <= _053_;
always @(posedge ap_clk)
ret_V_12_reg_1558 <= _044_;
always @(posedge ap_clk)
ret_V_6_cast_reg_1563 <= _046_;
always @(posedge ap_clk)
p_Val2_1_reg_1224[3:2] <= _039_;
always @(posedge ap_clk)
select_ln340_reg_1230 <= _052_;
always @(posedge ap_clk)
sel_tmp11_reg_1235 <= _051_;
always @(posedge ap_clk)
ret_reg_1091 <= _050_;
always @(posedge ap_clk)
p_Result_10_reg_1098 <= _031_;
always @(posedge ap_clk)
trunc_ln731_reg_1105 <= _063_;
always @(posedge ap_clk)
p_Result_11_reg_1110 <= _032_;
always @(posedge ap_clk)
p_Result_1_reg_1117 <= _036_;
always @(posedge ap_clk)
or_ln384_reg_1502 <= _027_;
always @(posedge ap_clk)
or_ln340_reg_1190 <= _026_;
always @(posedge ap_clk)
ret_V_8_reg_1212 <= _047_;
always @(posedge ap_clk)
ret_V_reg_1217 <= _049_;
always @(posedge ap_clk)
op_29_V_reg_1543 <= _024_;
always @(posedge ap_clk)
op_7_V_reg_1271 <= _025_;
always @(posedge ap_clk)
r_reg_1277 <= _042_;
always @(posedge ap_clk)
ret_V_9_reg_1282 <= _048_;
always @(posedge ap_clk)
trunc_ln1192_1_reg_1287 <= _058_;
always @(posedge ap_clk)
trunc_ln1192_2_reg_1292 <= _059_;
always @(posedge ap_clk)
op_12_V_reg_1297 <= _020_;
always @(posedge ap_clk)
icmp_ln768_reg_1130 <= _018_;
always @(posedge ap_clk)
icmp_ln786_reg_1135 <= _019_;
always @(posedge ap_clk)
p_Result_13_reg_1141 <= _033_;
always @(posedge ap_clk)
ret_V_2_reg_1261 <= _045_;
always @(posedge ap_clk)
icmp_ln213_reg_1266 <= _017_;
always @(posedge ap_clk)
ashr_ln1497_reg_1251 <= _015_;
always @(posedge ap_clk)
or_ln785_reg_1151 <= _028_;
always @(posedge ap_clk)
xor_ln785_reg_1157 <= _064_;
always @(posedge ap_clk)
or_ln786_reg_1163 <= _029_;
always @(posedge ap_clk)
and_ln786_reg_1169 <= _012_;
always @(posedge ap_clk)
sh_V_reg_1175 <= _054_;
always @(posedge ap_clk)
op_19_V_reg_1522 <= _022_;
always @(posedge ap_clk)
add_ln69_4_reg_1528 <= _008_;
always @(posedge ap_clk)
add_ln69_6_reg_1533 <= _010_;
always @(posedge ap_clk)
overflow_1_reg_1476 <= _030_;
always @(posedge ap_clk)
and_ln788_1_reg_1482 <= _013_;
always @(posedge ap_clk)
ret_V_11_reg_1487 <= _043_;
always @(posedge ap_clk)
add_ln69_3_reg_1492 <= _007_;
always @(posedge ap_clk)
add_ln69_5_reg_1497 <= _009_;
always @(posedge ap_clk)
add_ln691_reg_1570 <= _005_;
always @(posedge ap_clk)
add_ln1192_2_reg_1327 <= _004_;
always @(posedge ap_clk)
p_Val2_5_reg_1332 <= _040_;
always @(posedge ap_clk)
add_ln69_reg_1337 <= _011_;
always @(posedge ap_clk)
add_ln69_1_reg_1342 <= _006_;
always @(posedge ap_clk)
op_16_V_reg_1382 <= _021_;
always @(posedge ap_clk)
add_ln1192_1_reg_1387 <= _003_;
always @(posedge ap_clk)
p_Result_14_reg_1392 <= _034_;
always @(posedge ap_clk)
p_Val2_6_reg_1398 <= _041_;
always @(posedge ap_clk)
p_Result_16_reg_1404 <= _035_;
always @(posedge ap_clk)
p_Result_2_reg_1411 <= _037_;
always @(posedge ap_clk)
p_Result_3_reg_1416 <= _038_;
always @(posedge ap_clk)
op_23_V_reg_1422 <= _023_;
always @(posedge ap_clk)
carry_1_reg_1432 <= _016_;
always @(posedge ap_clk)
Range2_all_ones_reg_1439 <= _002_;
always @(posedge ap_clk)
Range1_all_ones_reg_1444 <= _000_;
always @(posedge ap_clk)
Range1_all_zeros_reg_1451 <= _001_;
always @(posedge ap_clk)
ap_CS_fsm <= _014_;
always @(posedge ap_clk)
p_Val2_1_reg_1224[1:0] <= 2'h0;
always @(posedge ap_clk)
trunc_ln69_reg_1347 <= _062_;
always @(posedge ap_clk)
trunc_ln69_1_reg_1352 <= _061_;
assign _065_ = _072_ ? 2'h2 : 2'h1;
assign _315_ = ap_CS_fsm == 1'h1;
function [24:0] _869_;
input [24:0] a;
input [624:0] b;
input [24:0] s;
case (s)
25'b0000000000000000000000001:
_869_ = b[24:0];
25'b0000000000000000000000010:
_869_ = b[49:25];
25'b0000000000000000000000100:
_869_ = b[74:50];
25'b0000000000000000000001000:
_869_ = b[99:75];
25'b0000000000000000000010000:
_869_ = b[124:100];
25'b0000000000000000000100000:
_869_ = b[149:125];
25'b0000000000000000001000000:
_869_ = b[174:150];
25'b0000000000000000010000000:
_869_ = b[199:175];
25'b0000000000000000100000000:
_869_ = b[224:200];
25'b0000000000000001000000000:
_869_ = b[249:225];
25'b0000000000000010000000000:
_869_ = b[274:250];
25'b0000000000000100000000000:
_869_ = b[299:275];
25'b0000000000001000000000000:
_869_ = b[324:300];
25'b0000000000010000000000000:
_869_ = b[349:325];
25'b0000000000100000000000000:
_869_ = b[374:350];
25'b0000000001000000000000000:
_869_ = b[399:375];
25'b0000000010000000000000000:
_869_ = b[424:400];
25'b0000000100000000000000000:
_869_ = b[449:425];
25'b0000001000000000000000000:
_869_ = b[474:450];
25'b0000010000000000000000000:
_869_ = b[499:475];
25'b0000100000000000000000000:
_869_ = b[524:500];
25'b0001000000000000000000000:
_869_ = b[549:525];
25'b0010000000000000000000000:
_869_ = b[574:550];
25'b0100000000000000000000000:
_869_ = b[599:575];
25'b1000000000000000000000000:
_869_ = b[624:600];
25'b0000000000000000000000000:
_869_ = a;
default:
_869_ = 25'bx;
endcase
endfunction
assign ap_NS_fsm = _869_(25'hxxxxxxx, { 23'h000000, _065_, 600'h000002000002000002000002000002000002000002000002000002000002000002000002000002000002000002000002000002000002000002000002000002000002000002000000000001 }, { _315_, _339_, _338_, _337_, _336_, _335_, _334_, _333_, _332_, _331_, _330_, _329_, _328_, _327_, _326_, _325_, _324_, _323_, _322_, _321_, _320_, _319_, _318_, _317_, _316_ });
assign _316_ = ap_CS_fsm == 25'h1000000;
assign _317_ = ap_CS_fsm == 24'h800000;
assign _318_ = ap_CS_fsm == 23'h400000;
assign _319_ = ap_CS_fsm == 22'h200000;
assign _320_ = ap_CS_fsm == 21'h100000;
assign _321_ = ap_CS_fsm == 20'h80000;
assign _322_ = ap_CS_fsm == 19'h40000;
assign _323_ = ap_CS_fsm == 18'h20000;
assign _324_ = ap_CS_fsm == 17'h10000;
assign _325_ = ap_CS_fsm == 16'h8000;
assign _326_ = ap_CS_fsm == 15'h4000;
assign _327_ = ap_CS_fsm == 14'h2000;
assign _328_ = ap_CS_fsm == 13'h1000;
assign _329_ = ap_CS_fsm == 12'h800;
assign _330_ = ap_CS_fsm == 11'h400;
assign _331_ = ap_CS_fsm == 10'h200;
assign _332_ = ap_CS_fsm == 9'h100;
assign _333_ = ap_CS_fsm == 8'h80;
assign _334_ = ap_CS_fsm == 7'h40;
assign _335_ = ap_CS_fsm == 6'h20;
assign _336_ = ap_CS_fsm == 5'h10;
assign _337_ = ap_CS_fsm == 4'h8;
assign _338_ = ap_CS_fsm == 3'h4;
assign _339_ = ap_CS_fsm == 2'h2;
assign op_30_ap_vld = ap_CS_fsm[24] ? 1'h1 : 1'h0;
assign ap_idle = _071_ ? 1'h1 : 1'h0;
assign _062_ = _070_ ? grp_fu_407_p2[1:0] : trunc_ln69_reg_1347;
assign _061_ = _069_ ? grp_fu_416_p2[1:0] : trunc_ln69_1_reg_1352;
assign _060_ = ap_CS_fsm[2] ? op_5[0] : trunc_ln1192_4_reg_1085;
assign _057_ = ap_CS_fsm[0] ? op_8[3] : tmp_4_reg_1043;
assign _056_ = ap_CS_fsm[1] ? grp_fu_237_p2 : sub_ln1497_reg_1048;
assign _055_ = _068_ ? grp_fu_277_p2 : shl_ln1497_reg_1256;
assign _053_ = _067_ ? select_ln785_fu_556_p3 : select_ln785_reg_1246;
assign _046_ = ap_CS_fsm[21] ? grp_fu_988_p2[32:1] : ret_V_6_cast_reg_1563;
assign _044_ = ap_CS_fsm[21] ? grp_fu_988_p2 : ret_V_12_reg_1558;
assign _051_ = ap_CS_fsm[7] ? sel_tmp11_fu_520_p2 : sel_tmp11_reg_1235;
assign _052_ = ap_CS_fsm[7] ? select_ln340_fu_498_p3 : select_ln340_reg_1230;
assign _039_ = ap_CS_fsm[7] ? trunc_ln731_reg_1105 : p_Val2_1_reg_1224[3:2];
assign _036_ = ap_CS_fsm[3] ? grp_fu_251_p2[16:2] : p_Result_1_reg_1117;
assign _032_ = ap_CS_fsm[3] ? grp_fu_251_p2[1] : p_Result_11_reg_1110;
assign _063_ = ap_CS_fsm[3] ? grp_fu_251_p2[1:0] : trunc_ln731_reg_1105;
assign _031_ = ap_CS_fsm[3] ? grp_fu_251_p2[16] : p_Result_10_reg_1098;
assign _050_ = ap_CS_fsm[3] ? grp_fu_251_p2 : ret_reg_1091;
assign _027_ = ap_CS_fsm[16] ? or_ln384_fu_927_p2 : or_ln384_reg_1502;
assign _049_ = ap_CS_fsm[6] ? grp_fu_386_p2[6:1] : ret_V_reg_1217;
assign _047_ = ap_CS_fsm[6] ? grp_fu_386_p2 : ret_V_8_reg_1212;
assign _026_ = ap_CS_fsm[6] ? or_ln340_fu_396_p2 : or_ln340_reg_1190;
assign _024_ = ap_CS_fsm[19] ? grp_fu_969_p2 : op_29_V_reg_1543;
assign _020_ = ap_CS_fsm[9] ? op_12_V_fu_629_p2 : op_12_V_reg_1297;
assign _059_ = ap_CS_fsm[9] ? op_7_V_fu_568_p3[2:0] : trunc_ln1192_2_reg_1292;
assign _058_ = ap_CS_fsm[9] ? op_7_V_fu_568_p3[0] : trunc_ln1192_1_reg_1287;
assign _048_ = ap_CS_fsm[9] ? ret_V_9_fu_594_p3 : ret_V_9_reg_1282;
assign _042_ = ap_CS_fsm[9] ? r_fu_573_p3 : r_reg_1277;
assign _025_ = ap_CS_fsm[9] ? op_7_V_fu_568_p3 : op_7_V_reg_1271;
assign _033_ = ap_CS_fsm[4] ? op_6[7] : p_Result_13_reg_1141;
assign _019_ = ap_CS_fsm[4] ? icmp_ln786_fu_322_p2 : icmp_ln786_reg_1135;
assign _018_ = ap_CS_fsm[4] ? icmp_ln768_fu_317_p2 : icmp_ln768_reg_1130;
assign _017_ = ap_CS_fsm[8] ? icmp_ln213_fu_562_p2 : icmp_ln213_reg_1266;
assign _045_ = ap_CS_fsm[8] ? grp_fu_526_p2 : ret_V_2_reg_1261;
assign _015_ = _066_ ? grp_fu_264_p2 : ashr_ln1497_reg_1251;
assign _054_ = ap_CS_fsm[5] ? grp_fu_335_p2 : sh_V_reg_1175;
assign _012_ = ap_CS_fsm[5] ? and_ln786_fu_365_p2 : and_ln786_reg_1169;
assign _029_ = ap_CS_fsm[5] ? or_ln786_fu_355_p2 : or_ln786_reg_1163;
assign _064_ = ap_CS_fsm[5] ? xor_ln785_fu_345_p2 : xor_ln785_reg_1157;
assign _028_ = ap_CS_fsm[5] ? or_ln785_fu_341_p2 : or_ln785_reg_1151;
assign _010_ = ap_CS_fsm[17] ? grp_fu_947_p2 : add_ln69_6_reg_1533;
assign _008_ = ap_CS_fsm[17] ? grp_fu_939_p2 : add_ln69_4_reg_1528;
assign _022_ = ap_CS_fsm[17] ? op_19_V_fu_960_p3 : op_19_V_reg_1522;
assign _009_ = ap_CS_fsm[15] ? grp_fu_836_p2 : add_ln69_5_reg_1497;
assign _007_ = ap_CS_fsm[15] ? grp_fu_830_p2 : add_ln69_3_reg_1492;
assign _043_ = ap_CS_fsm[15] ? grp_fu_814_p2 : ret_V_11_reg_1487;
assign _013_ = ap_CS_fsm[15] ? and_ln788_1_fu_902_p2 : and_ln788_1_reg_1482;
assign _030_ = ap_CS_fsm[15] ? overflow_1_fu_887_p2 : overflow_1_reg_1476;
assign _005_ = ap_CS_fsm[23] ? grp_fu_1004_p2 : add_ln691_reg_1570;
assign _006_ = ap_CS_fsm[11] ? grp_fu_666_p2 : add_ln69_1_reg_1342;
assign _011_ = ap_CS_fsm[11] ? grp_fu_660_p2 : add_ln69_reg_1337;
assign _040_ = ap_CS_fsm[11] ? grp_fu_648_p2[2:1] : p_Val2_5_reg_1332;
assign _004_ = ap_CS_fsm[11] ? grp_fu_648_p2 : add_ln1192_2_reg_1327;
assign _023_ = ap_CS_fsm[13] ? grp_fu_731_p2 : op_23_V_reg_1422;
assign _038_ = ap_CS_fsm[13] ? grp_fu_709_p2[6:3] : p_Result_3_reg_1416;
assign _037_ = ap_CS_fsm[13] ? grp_fu_709_p2[6:4] : p_Result_2_reg_1411;
assign _035_ = ap_CS_fsm[13] ? grp_fu_723_p2[1] : p_Result_16_reg_1404;
assign _041_ = ap_CS_fsm[13] ? grp_fu_723_p2 : p_Val2_6_reg_1398;
assign _034_ = ap_CS_fsm[13] ? grp_fu_709_p2[6] : p_Result_14_reg_1392;
assign _003_ = ap_CS_fsm[13] ? grp_fu_715_p2 : add_ln1192_1_reg_1387;
assign _021_ = ap_CS_fsm[13] ? op_16_V_fu_736_p3 : op_16_V_reg_1382;
assign _001_ = ap_CS_fsm[14] ? Range1_all_zeros_fu_805_p2 : Range1_all_zeros_reg_1451;
assign _000_ = ap_CS_fsm[14] ? Range1_all_ones_fu_800_p2 : Range1_all_ones_reg_1444;
assign _002_ = ap_CS_fsm[14] ? Range2_all_ones_fu_795_p2 : Range2_all_ones_reg_1439;
assign _016_ = ap_CS_fsm[14] ? carry_1_fu_789_p2 : carry_1_reg_1432;
assign _014_ = ap_rst ? 25'h0000001 : ap_NS_fsm;
assign Range1_all_ones_fu_800_p2 = _077_ ? 1'h1 : 1'h0;
assign Range1_all_zeros_fu_805_p2 = _078_ ? 1'h1 : 1'h0;
assign Range2_all_ones_fu_795_p2 = _079_ ? 1'h1 : 1'h0;
assign deleted_ones_fu_865_p3 = carry_1_reg_1432 ? and_ln780_fu_860_p2 : Range1_all_ones_reg_1444;
assign deleted_zeros_fu_842_p3 = carry_1_reg_1432 ? Range1_all_ones_reg_1444 : Range1_all_zeros_reg_1451;
assign icmp_ln213_fu_562_p2 = _312_ ? 1'h1 : 1'h0;
assign icmp_ln768_fu_317_p2 = _313_ ? 1'h1 : 1'h0;
assign icmp_ln786_fu_322_p2 = _314_ ? 1'h1 : 1'h0;
assign op_16_V_fu_736_p3 = p_Result_13_reg_1141 ? trunc_ln69_reg_1347 : trunc_ln69_1_reg_1352;
assign op_19_V_fu_960_p3 = or_ln384_reg_1502 ? select_ln384_fu_953_p3 : p_Val2_6_reg_1398;
assign op_30 = ret_V_12_reg_1558[33] ? select_ln850_1_fu_1019_p3 : ret_V_6_cast_reg_1563;
assign op_7_V_fu_568_p3 = sel_tmp11_reg_1235 ? p_Val2_1_reg_1224 : select_ln785_reg_1246;
assign r_fu_573_p3 = tmp_4_reg_1043 ? shl_ln1497_reg_1256 : ashr_ln1497_reg_1251;
assign ret_V_9_fu_594_p3 = ret_V_8_reg_1212[6] ? select_ln850_fu_588_p3 : ret_V_reg_1217;
assign select_ln340_fu_498_p3 = and_ln340_fu_493_p2 ? { trunc_ln731_reg_1105, 2'h0 } : { ret_reg_1091[2], p_Val2_2_fu_472_p2 };
assign select_ln384_fu_953_p3 = overflow_1_reg_1476 ? 2'h1 : 2'h3;
assign select_ln785_fu_556_p3 = and_ln785_fu_551_p2 ? p_Val2_1_reg_1224 : select_ln340_reg_1230;
assign select_ln850_1_fu_1019_p3 = op_19_V_reg_1522[0] ? add_ln691_reg_1570 : ret_V_6_cast_reg_1563;
assign select_ln850_fu_588_p3 = op_9[0] ? ret_V_2_reg_1261 : ret_V_reg_1217;
assign xor_ln365_fu_460_p2 = ret_reg_1091[2] ^ ret_reg_1091[1];
assign ap_CS_fsm_state1 = ap_CS_fsm[0];
assign ap_CS_fsm_state10 = ap_CS_fsm[9];
assign ap_CS_fsm_state11 = ap_CS_fsm[10];
assign ap_CS_fsm_state12 = ap_CS_fsm[11];
assign ap_CS_fsm_state13 = ap_CS_fsm[12];
assign ap_CS_fsm_state14 = ap_CS_fsm[13];
assign ap_CS_fsm_state15 = ap_CS_fsm[14];
assign ap_CS_fsm_state16 = ap_CS_fsm[15];
assign ap_CS_fsm_state17 = ap_CS_fsm[16];
assign ap_CS_fsm_state18 = ap_CS_fsm[17];
assign ap_CS_fsm_state19 = ap_CS_fsm[18];
assign ap_CS_fsm_state2 = ap_CS_fsm[1];
assign ap_CS_fsm_state20 = ap_CS_fsm[19];
assign ap_CS_fsm_state21 = ap_CS_fsm[20];
assign ap_CS_fsm_state22 = ap_CS_fsm[21];
assign ap_CS_fsm_state23 = ap_CS_fsm[22];
assign ap_CS_fsm_state24 = ap_CS_fsm[23];
assign ap_CS_fsm_state25 = ap_CS_fsm[24];
assign ap_CS_fsm_state3 = ap_CS_fsm[2];
assign ap_CS_fsm_state4 = ap_CS_fsm[3];
assign ap_CS_fsm_state5 = ap_CS_fsm[4];
assign ap_CS_fsm_state6 = ap_CS_fsm[5];
assign ap_CS_fsm_state7 = ap_CS_fsm[6];
assign ap_CS_fsm_state8 = ap_CS_fsm[7];
assign ap_CS_fsm_state9 = ap_CS_fsm[8];
assign ap_done = op_30_ap_vld;
assign ap_ready = op_30_ap_vld;
assign grp_fu_237_p1 = { op_8[3], op_8 };
assign grp_fu_251_p0 = { op_2[15], op_2 };
assign grp_fu_251_p1 = { op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5 };
assign grp_fu_264_p1 = { op_8[3], op_8[3], op_8[3], op_8[3], op_8[3], op_8[3], op_8[3], op_8[3], op_8[3], op_8[3], op_8[3], op_8[3], op_8 };
assign grp_fu_277_p1 = { sub_ln1497_reg_1048[4], sub_ln1497_reg_1048[4], sub_ln1497_reg_1048[4], sub_ln1497_reg_1048[4], sub_ln1497_reg_1048[4], sub_ln1497_reg_1048[4], sub_ln1497_reg_1048[4], sub_ln1497_reg_1048[4], sub_ln1497_reg_1048[4], sub_ln1497_reg_1048[4], sub_ln1497_reg_1048[4], sub_ln1497_reg_1048 };
assign grp_fu_386_p0 = { 2'h0, op_3, 1'h0 };
assign grp_fu_386_p1 = { op_9[3], op_9[3], op_9[3], op_9 };
assign grp_fu_407_p1 = { 24'h000000, sh_V_reg_1175 };
assign grp_fu_416_p1 = { 24'h000000, op_6 };
assign grp_fu_648_p0 = { trunc_ln1192_4_reg_1085, 2'h0 };
assign grp_fu_660_p0 = { r_reg_1277[15], r_reg_1277 };
assign grp_fu_660_p1 = { op_10[7], op_10[7], op_10[7], op_10[7], op_10[7], op_10[7], op_10[7], op_10[7], op_10[7], op_10 };
assign grp_fu_666_p0 = { ret_V_9_reg_1282[5], ret_V_9_reg_1282 };
assign grp_fu_666_p1 = { 6'h00, op_12_V_reg_1297 };
assign grp_fu_709_p0 = { op_5[3], op_5, 2'h0 };
assign grp_fu_709_p1 = { op_7_V_reg_1271[3], op_7_V_reg_1271[3], op_7_V_reg_1271[3], op_7_V_reg_1271 };
assign grp_fu_715_p0 = { op_5[1:0], 2'h0 };
assign grp_fu_723_p1 = { 1'h0, trunc_ln1192_1_reg_1287 };
assign grp_fu_731_p0 = { add_ln69_1_reg_1342[6], add_ln69_1_reg_1342[6], add_ln69_1_reg_1342[6], add_ln69_1_reg_1342[6], add_ln69_1_reg_1342[6], add_ln69_1_reg_1342[6], add_ln69_1_reg_1342[6], add_ln69_1_reg_1342[6], add_ln69_1_reg_1342[6], add_ln69_1_reg_1342[6], add_ln69_1_reg_1342 };
assign grp_fu_814_p1 = { op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13 };
assign grp_fu_830_p0 = { op_14[1], op_14[1], op_14[1], op_14[1], op_14[1], op_14[1], op_14[1], op_14[1], op_14[1], op_14[1], op_14[1], op_14[1], op_14[1], op_14[1], op_14[1], op_14[1], op_14[1], op_14[1], op_14[1], op_14[1], op_14[1], op_14[1], op_14[1], op_14[1], op_14[1], op_14[1], op_14[1], op_14[1], op_14[1], op_14[1], op_14 };
assign grp_fu_836_p0 = { op_18[1], op_18 };
assign grp_fu_836_p1 = { op_16_V_reg_1382[1], op_16_V_reg_1382 };
assign grp_fu_939_p1 = { ret_V_11_reg_1487[16], ret_V_11_reg_1487[16], ret_V_11_reg_1487[16], ret_V_11_reg_1487[16], ret_V_11_reg_1487[16], ret_V_11_reg_1487[16], ret_V_11_reg_1487[16], ret_V_11_reg_1487[16], ret_V_11_reg_1487[16], ret_V_11_reg_1487[16], ret_V_11_reg_1487[16], ret_V_11_reg_1487[16], ret_V_11_reg_1487[16], ret_V_11_reg_1487[16], ret_V_11_reg_1487[16], ret_V_11_reg_1487 };
assign grp_fu_947_p0 = { add_ln69_5_reg_1497[2], add_ln69_5_reg_1497 };
assign grp_fu_947_p1 = { op_17[1], op_17[1], op_17 };
assign grp_fu_969_p0 = { add_ln69_6_reg_1533[3], add_ln69_6_reg_1533[3], add_ln69_6_reg_1533[3], add_ln69_6_reg_1533[3], add_ln69_6_reg_1533[3], add_ln69_6_reg_1533[3], add_ln69_6_reg_1533[3], add_ln69_6_reg_1533[3], add_ln69_6_reg_1533[3], add_ln69_6_reg_1533[3], add_ln69_6_reg_1533[3], add_ln69_6_reg_1533[3], add_ln69_6_reg_1533[3], add_ln69_6_reg_1533[3], add_ln69_6_reg_1533[3], add_ln69_6_reg_1533[3], add_ln69_6_reg_1533[3], add_ln69_6_reg_1533[3], add_ln69_6_reg_1533[3], add_ln69_6_reg_1533[3], add_ln69_6_reg_1533[3], add_ln69_6_reg_1533[3], add_ln69_6_reg_1533[3], add_ln69_6_reg_1533[3], add_ln69_6_reg_1533[3], add_ln69_6_reg_1533[3], add_ln69_6_reg_1533[3], add_ln69_6_reg_1533[3], add_ln69_6_reg_1533 };
assign grp_fu_988_p0 = { op_29_V_reg_1543[31], op_29_V_reg_1543, 1'h0 };
assign grp_fu_988_p1 = { op_19_V_reg_1522[1], op_19_V_reg_1522[1], op_19_V_reg_1522[1], op_19_V_reg_1522[1], op_19_V_reg_1522[1], op_19_V_reg_1522[1], op_19_V_reg_1522[1], op_19_V_reg_1522[1], op_19_V_reg_1522[1], op_19_V_reg_1522[1], op_19_V_reg_1522[1], op_19_V_reg_1522[1], op_19_V_reg_1522[1], op_19_V_reg_1522[1], op_19_V_reg_1522[1], op_19_V_reg_1522[1], op_19_V_reg_1522[1], op_19_V_reg_1522[1], op_19_V_reg_1522[1], op_19_V_reg_1522[1], op_19_V_reg_1522[1], op_19_V_reg_1522[1], op_19_V_reg_1522[1], op_19_V_reg_1522[1], op_19_V_reg_1522[1], op_19_V_reg_1522[1], op_19_V_reg_1522[1], op_19_V_reg_1522[1], op_19_V_reg_1522[1], op_19_V_reg_1522[1], op_19_V_reg_1522[1], op_19_V_reg_1522[1], op_19_V_reg_1522 };
assign lhs_V_1_fu_690_p1 = op_5;
assign lhs_V_1_fu_690_p3 = { op_5, 2'h0 };
assign lhs_V_fu_370_p3 = { op_3, 1'h0 };
assign p_Result_12_fu_439_p3 = ret_reg_1091[2];
assign p_Result_13_fu_327_p1 = op_6;
assign p_Result_15_fu_777_p3 = add_ln1192_2_reg_1327[2];
assign p_Result_5_fu_578_p3 = ret_V_8_reg_1212[6];
assign p_Result_9_fu_1009_p3 = ret_V_12_reg_1558[33];
assign p_Result_s_14_fu_478_p4 = { ret_reg_1091[2], p_Val2_2_fu_472_p2 };
assign p_Result_s_fu_531_p4 = op_0[3:2];
assign p_Val2_1_fu_432_p3 = { trunc_ln731_reg_1105, 2'h0 };
assign rhs_3_fu_977_p3 = { op_29_V_reg_1543, 1'h0 };
assign sext_ln1497_1_fu_270_p1 = { sub_ln1497_reg_1048[4], sub_ln1497_reg_1048[4], sub_ln1497_reg_1048[4], sub_ln1497_reg_1048[4], sub_ln1497_reg_1048[4], sub_ln1497_reg_1048[4], sub_ln1497_reg_1048[4], sub_ln1497_reg_1048[4], sub_ln1497_reg_1048[4], sub_ln1497_reg_1048[4], sub_ln1497_reg_1048[4], sub_ln1497_reg_1048[4], sub_ln1497_reg_1048[4], sub_ln1497_reg_1048[4], sub_ln1497_reg_1048[4], sub_ln1497_reg_1048[4], sub_ln1497_reg_1048[4], sub_ln1497_reg_1048[4], sub_ln1497_reg_1048[4], sub_ln1497_reg_1048[4], sub_ln1497_reg_1048[4], sub_ln1497_reg_1048[4], sub_ln1497_reg_1048[4], sub_ln1497_reg_1048[4], sub_ln1497_reg_1048[4], sub_ln1497_reg_1048[4], sub_ln1497_reg_1048[4], sub_ln1497_reg_1048 };
assign sext_ln1497_fu_225_p0 = op_8;
assign sext_ln215_1_fu_247_p0 = op_5;
assign sext_ln215_fu_243_p0 = op_2;
assign sext_ln545_fu_257_p0 = op_8;
assign sext_ln545_fu_257_p1 = { op_8[3], op_8[3], op_8[3], op_8[3], op_8[3], op_8[3], op_8[3], op_8[3], op_8[3], op_8[3], op_8[3], op_8[3], op_8[3], op_8[3], op_8[3], op_8[3], op_8[3], op_8[3], op_8[3], op_8[3], op_8[3], op_8[3], op_8[3], op_8[3], op_8[3], op_8[3], op_8[3], op_8[3], op_8 };
assign sext_ln703_fu_382_p0 = op_9;
assign sext_ln781_fu_401_p0 = op_6;
assign sext_ln781_fu_401_p1 = { op_6[7], op_6[7], op_6[7], op_6[7], op_6[7], op_6[7], op_6[7], op_6[7], op_6[7], op_6[7], op_6[7], op_6[7], op_6[7], op_6[7], op_6[7], op_6[7], op_6[7], op_6[7], op_6[7], op_6[7], op_6[7], op_6[7], op_6[7], op_6[7], op_6 };
assign shl_ln1192_fu_704_p0 = op_5;
assign tmp_10_fu_612_p3 = op_0[1];
assign tmp_1_fu_453_p3 = ret_reg_1091[1];
assign tmp_4_fu_229_p1 = op_8;
assign tmp_9_fu_847_p3 = add_ln1192_1_reg_1387[3];
assign tmp_fu_446_p3 = ret_reg_1091[2];
assign trunc_ln1192_1_fu_604_p1 = op_7_V_fu_568_p3[0];
assign trunc_ln1192_2_fu_608_p1 = op_7_V_fu_568_p3[2:0];
assign trunc_ln1192_4_fu_283_p0 = op_5;
assign trunc_ln1192_4_fu_283_p1 = op_5[0];
assign trunc_ln1192_fu_601_p1 = op_0[0];
assign trunc_ln69_1_fu_686_p1 = grp_fu_416_p2[1:0];
assign trunc_ln69_fu_682_p1 = grp_fu_407_p2[1:0];
assign trunc_ln731_fu_295_p1 = grp_fu_251_p2[1:0];
assign trunc_ln790_fu_893_p1 = p_Val2_6_reg_1398[0];
assign trunc_ln851_1_fu_1016_p1 = op_19_V_reg_1522[0];
assign trunc_ln851_fu_585_p0 = op_9;
assign trunc_ln851_fu_585_p1 = op_9[0];
assign zext_ln546_1_fu_413_p0 = op_6;
assign \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.ain_s0  = \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.a ;
assign \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.s  = { \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.fas_s2 , \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.sum_s1  };
assign \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.u2.a  = \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.ain_s1 ;
assign \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.u2.b  = \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.bin_s1 ;
assign \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.u2.cin  = \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.carry_s1 ;
assign \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.facout_s2  = \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.u2.cout ;
assign \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.fas_s2  = \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.u2.s ;
assign \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.u1.a  = \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.a [3:0];
assign \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.u1.b  = \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.bin_s0 [3:0];
assign \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.u1.cin  = 1'h1;
assign \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.facout_s1  = \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.u1.cout ;
assign \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.fas_s1  = \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.u1.s ;
assign \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.a  = \sub_8ns_8s_8_2_1_U5.din0 ;
assign \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.b  = \sub_8ns_8s_8_2_1_U5.din1 ;
assign \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.ce  = \sub_8ns_8s_8_2_1_U5.ce ;
assign \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.clk  = \sub_8ns_8s_8_2_1_U5.clk ;
assign \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.reset  = \sub_8ns_8s_8_2_1_U5.reset ;
assign \sub_8ns_8s_8_2_1_U5.dout  = \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.s ;
assign \sub_8ns_8s_8_2_1_U5.ce  = 1'h1;
assign \sub_8ns_8s_8_2_1_U5.clk  = ap_clk;
assign \sub_8ns_8s_8_2_1_U5.din0  = 8'h00;
assign \sub_8ns_8s_8_2_1_U5.din1  = op_6;
assign grp_fu_335_p2 = \sub_8ns_8s_8_2_1_U5.dout ;
assign \sub_8ns_8s_8_2_1_U5.reset  = ap_rst;
assign \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.ain_s0  = \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.a ;
assign \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.s  = { \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.fas_s2 , \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.sum_s1  };
assign \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.u2.a  = \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.ain_s1 ;
assign \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.u2.b  = \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.bin_s1 ;
assign \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.u2.cin  = \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.carry_s1 ;
assign \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.facout_s2  = \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.u2.cout ;
assign \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.fas_s2  = \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.u2.s ;
assign \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.u1.a  = \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.a [1:0];
assign \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.u1.b  = \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.bin_s0 [1:0];
assign \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.u1.cin  = 1'h1;
assign \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.facout_s1  = \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.u1.cout ;
assign \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.fas_s1  = \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.u1.s ;
assign \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.a  = \sub_5ns_5s_5_2_1_U1.din0 ;
assign \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.b  = \sub_5ns_5s_5_2_1_U1.din1 ;
assign \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.ce  = \sub_5ns_5s_5_2_1_U1.ce ;
assign \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.clk  = \sub_5ns_5s_5_2_1_U1.clk ;
assign \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.reset  = \sub_5ns_5s_5_2_1_U1.reset ;
assign \sub_5ns_5s_5_2_1_U1.dout  = \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.s ;
assign \sub_5ns_5s_5_2_1_U1.ce  = 1'h1;
assign \sub_5ns_5s_5_2_1_U1.clk  = ap_clk;
assign \sub_5ns_5s_5_2_1_U1.din0  = 5'h00;
assign \sub_5ns_5s_5_2_1_U1.din1  = { op_8[3], op_8 };
assign grp_fu_237_p2 = \sub_5ns_5s_5_2_1_U1.dout ;
assign \sub_5ns_5s_5_2_1_U1.reset  = ap_rst;
assign \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.ain_s0  = \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.a ;
assign \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.s  = { \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.fas_s2 , \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.sum_s1  };
assign \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.u2.a  = \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.ain_s1 ;
assign \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.u2.b  = \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.bin_s1 ;
assign \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.u2.cin  = \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.carry_s1 ;
assign \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.facout_s2  = \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.u2.cout ;
assign \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.fas_s2  = \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.u2.s ;
assign \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.u1.a  = \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.a [7:0];
assign \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.u1.b  = \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.bin_s0 [7:0];
assign \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.u1.cin  = 1'h1;
assign \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.facout_s1  = \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.u1.cout ;
assign \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.fas_s1  = \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.u1.s ;
assign \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.a  = \sub_17s_17s_17_2_1_U2.din0 ;
assign \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.b  = \sub_17s_17s_17_2_1_U2.din1 ;
assign \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.ce  = \sub_17s_17s_17_2_1_U2.ce ;
assign \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.clk  = \sub_17s_17s_17_2_1_U2.clk ;
assign \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.reset  = \sub_17s_17s_17_2_1_U2.reset ;
assign \sub_17s_17s_17_2_1_U2.dout  = \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.s ;
assign \sub_17s_17s_17_2_1_U2.ce  = 1'h1;
assign \sub_17s_17s_17_2_1_U2.clk  = ap_clk;
assign \sub_17s_17s_17_2_1_U2.din0  = { op_2[15], op_2 };
assign \sub_17s_17s_17_2_1_U2.din1  = { op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5 };
assign grp_fu_251_p2 = \sub_17s_17s_17_2_1_U2.dout ;
assign \sub_17s_17s_17_2_1_U2.reset  = ap_rst;
assign \shl_32s_8ns_32_7_1_U8.din1_cast  = \shl_32s_8ns_32_7_1_U8.din1 [7:0];
assign \shl_32s_8ns_32_7_1_U8.din1_mask  = 8'h03;
assign \shl_32s_8ns_32_7_1_U8.ce  = 1'h1;
assign \shl_32s_8ns_32_7_1_U8.clk  = ap_clk;
assign \shl_32s_8ns_32_7_1_U8.din0  = { op_6[7], op_6[7], op_6[7], op_6[7], op_6[7], op_6[7], op_6[7], op_6[7], op_6[7], op_6[7], op_6[7], op_6[7], op_6[7], op_6[7], op_6[7], op_6[7], op_6[7], op_6[7], op_6[7], op_6[7], op_6[7], op_6[7], op_6[7], op_6[7], op_6 };
assign \shl_32s_8ns_32_7_1_U8.din1  = { 24'h000000, op_6 };
assign grp_fu_416_p2 = \shl_32s_8ns_32_7_1_U8.dout ;
assign \shl_32s_8ns_32_7_1_U8.reset  = ap_rst;
assign \shl_16s_16ns_16_7_1_U4.din1_cast  = \shl_16s_16ns_16_7_1_U4.din1 ;
assign \shl_16s_16ns_16_7_1_U4.din1_mask  = 16'h0007;
assign \shl_16s_16ns_16_7_1_U4.ce  = 1'h1;
assign \shl_16s_16ns_16_7_1_U4.clk  = ap_clk;
assign \shl_16s_16ns_16_7_1_U4.din0  = op_2;
assign \shl_16s_16ns_16_7_1_U4.din1  = { sub_ln1497_reg_1048[4], sub_ln1497_reg_1048[4], sub_ln1497_reg_1048[4], sub_ln1497_reg_1048[4], sub_ln1497_reg_1048[4], sub_ln1497_reg_1048[4], sub_ln1497_reg_1048[4], sub_ln1497_reg_1048[4], sub_ln1497_reg_1048[4], sub_ln1497_reg_1048[4], sub_ln1497_reg_1048[4], sub_ln1497_reg_1048 };
assign grp_fu_277_p2 = \shl_16s_16ns_16_7_1_U4.dout ;
assign \shl_16s_16ns_16_7_1_U4.reset  = ap_rst;
assign \ashr_32s_8ns_32_7_1_U7.din1_cast  = \ashr_32s_8ns_32_7_1_U7.din1 [7:0];
assign \ashr_32s_8ns_32_7_1_U7.din1_mask  = 8'h03;
assign \ashr_32s_8ns_32_7_1_U7.ce  = 1'h1;
assign \ashr_32s_8ns_32_7_1_U7.clk  = ap_clk;
assign \ashr_32s_8ns_32_7_1_U7.din0  = { op_6[7], op_6[7], op_6[7], op_6[7], op_6[7], op_6[7], op_6[7], op_6[7], op_6[7], op_6[7], op_6[7], op_6[7], op_6[7], op_6[7], op_6[7], op_6[7], op_6[7], op_6[7], op_6[7], op_6[7], op_6[7], op_6[7], op_6[7], op_6[7], op_6 };
assign \ashr_32s_8ns_32_7_1_U7.din1  = { 24'h000000, sh_V_reg_1175 };
assign grp_fu_407_p2 = \ashr_32s_8ns_32_7_1_U7.dout ;
assign \ashr_32s_8ns_32_7_1_U7.reset  = ap_rst;
assign \ashr_16s_16ns_16_7_1_U3.din1_cast  = \ashr_16s_16ns_16_7_1_U3.din1 ;
assign \ashr_16s_16ns_16_7_1_U3.din1_mask  = 16'h0007;
assign \ashr_16s_16ns_16_7_1_U3.ce  = 1'h1;
assign \ashr_16s_16ns_16_7_1_U3.clk  = ap_clk;
assign \ashr_16s_16ns_16_7_1_U3.din0  = op_2;
assign \ashr_16s_16ns_16_7_1_U3.din1  = { op_8[3], op_8[3], op_8[3], op_8[3], op_8[3], op_8[3], op_8[3], op_8[3], op_8[3], op_8[3], op_8[3], op_8[3], op_8 };
assign grp_fu_264_p2 = \ashr_16s_16ns_16_7_1_U3.dout ;
assign \ashr_16s_16ns_16_7_1_U3.reset  = ap_rst;
assign \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.ain_s0  = \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.a ;
assign \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.bin_s0  = \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.b ;
assign \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.s  = { \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.fas_s2 , \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.sum_s1  };
assign \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.u2.a  = \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.ain_s1 ;
assign \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.u2.b  = \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.bin_s1 ;
assign \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.u2.cin  = \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.carry_s1 ;
assign \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.facout_s2  = \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.u2.cout ;
assign \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.fas_s2  = \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.u2.s ;
assign \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.u1.a  = \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.a [2:0];
assign \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.u1.b  = \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.b [2:0];
assign \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.u1.cin  = 1'h0;
assign \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.facout_s1  = \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.u1.cout ;
assign \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.fas_s1  = \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.u1.s ;
assign \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.a  = \add_7s_7s_7_2_1_U13.din0 ;
assign \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.b  = \add_7s_7s_7_2_1_U13.din1 ;
assign \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.ce  = \add_7s_7s_7_2_1_U13.ce ;
assign \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.clk  = \add_7s_7s_7_2_1_U13.clk ;
assign \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.reset  = \add_7s_7s_7_2_1_U13.reset ;
assign \add_7s_7s_7_2_1_U13.dout  = \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.s ;
assign \add_7s_7s_7_2_1_U13.ce  = 1'h1;
assign \add_7s_7s_7_2_1_U13.clk  = ap_clk;
assign \add_7s_7s_7_2_1_U13.din0  = { op_5[3], op_5, 2'h0 };
assign \add_7s_7s_7_2_1_U13.din1  = { op_7_V_reg_1271[3], op_7_V_reg_1271[3], op_7_V_reg_1271[3], op_7_V_reg_1271 };
assign grp_fu_709_p2 = \add_7s_7s_7_2_1_U13.dout ;
assign \add_7s_7s_7_2_1_U13.reset  = ap_rst;
assign \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.ain_s0  = \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.a ;
assign \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.bin_s0  = \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.b ;
assign \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.s  = { \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.fas_s2 , \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.sum_s1  };
assign \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.u2.a  = \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.ain_s1 ;
assign \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.u2.b  = \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.bin_s1 ;
assign \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.u2.cin  = \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.carry_s1 ;
assign \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.facout_s2  = \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.u2.cout ;
assign \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.fas_s2  = \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.u2.s ;
assign \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.u1.a  = \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.a [2:0];
assign \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.u1.b  = \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.b [2:0];
assign \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.u1.cin  = 1'h0;
assign \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.facout_s1  = \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.u1.cout ;
assign \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.fas_s1  = \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.u1.s ;
assign \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.a  = \add_7s_7ns_7_2_1_U12.din0 ;
assign \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.b  = \add_7s_7ns_7_2_1_U12.din1 ;
assign \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.ce  = \add_7s_7ns_7_2_1_U12.ce ;
assign \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.clk  = \add_7s_7ns_7_2_1_U12.clk ;
assign \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.reset  = \add_7s_7ns_7_2_1_U12.reset ;
assign \add_7s_7ns_7_2_1_U12.dout  = \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.s ;
assign \add_7s_7ns_7_2_1_U12.ce  = 1'h1;
assign \add_7s_7ns_7_2_1_U12.clk  = ap_clk;
assign \add_7s_7ns_7_2_1_U12.din0  = { ret_V_9_reg_1282[5], ret_V_9_reg_1282 };
assign \add_7s_7ns_7_2_1_U12.din1  = { 6'h00, op_12_V_reg_1297 };
assign grp_fu_666_p2 = \add_7s_7ns_7_2_1_U12.dout ;
assign \add_7s_7ns_7_2_1_U12.reset  = ap_rst;
assign \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.ain_s0  = \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.a ;
assign \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.bin_s0  = \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.b ;
assign \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.s  = { \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.fas_s2 , \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.sum_s1  };
assign \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.u2.a  = \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.ain_s1 ;
assign \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.u2.b  = \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.bin_s1 ;
assign \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.u2.cin  = \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.carry_s1 ;
assign \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.facout_s2  = \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.u2.cout ;
assign \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.fas_s2  = \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.u2.s ;
assign \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.u1.a  = \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.a [2:0];
assign \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.u1.b  = \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.b [2:0];
assign \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.u1.cin  = 1'h0;
assign \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.facout_s1  = \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.u1.cout ;
assign \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.fas_s1  = \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.u1.s ;
assign \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.a  = \add_7ns_7s_7_2_1_U6.din0 ;
assign \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.b  = \add_7ns_7s_7_2_1_U6.din1 ;
assign \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.ce  = \add_7ns_7s_7_2_1_U6.ce ;
assign \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.clk  = \add_7ns_7s_7_2_1_U6.clk ;
assign \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.reset  = \add_7ns_7s_7_2_1_U6.reset ;
assign \add_7ns_7s_7_2_1_U6.dout  = \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.s ;
assign \add_7ns_7s_7_2_1_U6.ce  = 1'h1;
assign \add_7ns_7s_7_2_1_U6.clk  = ap_clk;
assign \add_7ns_7s_7_2_1_U6.din0  = { 2'h0, op_3, 1'h0 };
assign \add_7ns_7s_7_2_1_U6.din1  = { op_9[3], op_9[3], op_9[3], op_9 };
assign grp_fu_386_p2 = \add_7ns_7s_7_2_1_U6.dout ;
assign \add_7ns_7s_7_2_1_U6.reset  = ap_rst;
assign \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.ain_s0  = \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.a ;
assign \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.bin_s0  = \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.b ;
assign \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.s  = { \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.fas_s2 , \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.sum_s1  };
assign \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.u2.a  = \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.ain_s1 ;
assign \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.u2.b  = \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.bin_s1 ;
assign \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.u2.cin  = \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.carry_s1 ;
assign \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.facout_s2  = \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.u2.cout ;
assign \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.fas_s2  = \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.u2.s ;
assign \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.u1.a  = \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.a [2:0];
assign \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.u1.b  = \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.b [2:0];
assign \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.u1.cin  = 1'h0;
assign \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.facout_s1  = \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.u1.cout ;
assign \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.fas_s1  = \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.u1.s ;
assign \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.a  = \add_6ns_6ns_6_2_1_U9.din0 ;
assign \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.b  = \add_6ns_6ns_6_2_1_U9.din1 ;
assign \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.ce  = \add_6ns_6ns_6_2_1_U9.ce ;
assign \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.clk  = \add_6ns_6ns_6_2_1_U9.clk ;
assign \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.reset  = \add_6ns_6ns_6_2_1_U9.reset ;
assign \add_6ns_6ns_6_2_1_U9.dout  = \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.s ;
assign \add_6ns_6ns_6_2_1_U9.ce  = 1'h1;
assign \add_6ns_6ns_6_2_1_U9.clk  = ap_clk;
assign \add_6ns_6ns_6_2_1_U9.din0  = ret_V_reg_1217;
assign \add_6ns_6ns_6_2_1_U9.din1  = 6'h01;
assign grp_fu_526_p2 = \add_6ns_6ns_6_2_1_U9.dout ;
assign \add_6ns_6ns_6_2_1_U9.reset  = ap_rst;
assign \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.ain_s0  = \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.a ;
assign \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.bin_s0  = \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.b ;
assign \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.s  = { \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.fas_s2 , \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.sum_s1  };
assign \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.u2.a  = \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.ain_s1 ;
assign \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.u2.b  = \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.bin_s1 ;
assign \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.u2.cin  = \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.carry_s1 ;
assign \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.facout_s2  = \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.u2.cout ;
assign \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.fas_s2  = \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.u2.s ;
assign \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.u1.a  = \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.a [1:0];
assign \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.u1.b  = \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.b [1:0];
assign \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.u1.cin  = 1'h0;
assign \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.facout_s1  = \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.u1.cout ;
assign \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.fas_s1  = \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.u1.s ;
assign \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.a  = \add_4s_4s_4_2_1_U21.din0 ;
assign \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.b  = \add_4s_4s_4_2_1_U21.din1 ;
assign \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.ce  = \add_4s_4s_4_2_1_U21.ce ;
assign \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.clk  = \add_4s_4s_4_2_1_U21.clk ;
assign \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.reset  = \add_4s_4s_4_2_1_U21.reset ;
assign \add_4s_4s_4_2_1_U21.dout  = \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.s ;
assign \add_4s_4s_4_2_1_U21.ce  = 1'h1;
assign \add_4s_4s_4_2_1_U21.clk  = ap_clk;
assign \add_4s_4s_4_2_1_U21.din0  = { add_ln69_5_reg_1497[2], add_ln69_5_reg_1497 };
assign \add_4s_4s_4_2_1_U21.din1  = { op_17[1], op_17[1], op_17 };
assign grp_fu_947_p2 = \add_4s_4s_4_2_1_U21.dout ;
assign \add_4s_4s_4_2_1_U21.reset  = ap_rst;
assign \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.ain_s0  = \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.a ;
assign \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.bin_s0  = \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.b ;
assign \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.s  = { \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.fas_s2 , \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.sum_s1  };
assign \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.u2.a  = \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.ain_s1 ;
assign \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.u2.b  = \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.bin_s1 ;
assign \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.u2.cin  = \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.carry_s1 ;
assign \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.facout_s2  = \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.u2.cout ;
assign \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.fas_s2  = \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.u2.s ;
assign \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.u1.a  = \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.a [1:0];
assign \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.u1.b  = \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.b [1:0];
assign \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.u1.cin  = 1'h0;
assign \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.facout_s1  = \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.u1.cout ;
assign \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.fas_s1  = \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.u1.s ;
assign \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.a  = \add_4ns_4s_4_2_1_U14.din0 ;
assign \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.b  = \add_4ns_4s_4_2_1_U14.din1 ;
assign \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.ce  = \add_4ns_4s_4_2_1_U14.ce ;
assign \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.clk  = \add_4ns_4s_4_2_1_U14.clk ;
assign \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.reset  = \add_4ns_4s_4_2_1_U14.reset ;
assign \add_4ns_4s_4_2_1_U14.dout  = \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.s ;
assign \add_4ns_4s_4_2_1_U14.ce  = 1'h1;
assign \add_4ns_4s_4_2_1_U14.clk  = ap_clk;
assign \add_4ns_4s_4_2_1_U14.din0  = { op_5[1:0], 2'h0 };
assign \add_4ns_4s_4_2_1_U14.din1  = op_7_V_reg_1271;
assign grp_fu_715_p2 = \add_4ns_4s_4_2_1_U14.dout ;
assign \add_4ns_4s_4_2_1_U14.reset  = ap_rst;
assign \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.ain_s0  = \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.a ;
assign \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.bin_s0  = \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.b ;
assign \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.s  = { \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.fas_s2 , \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.sum_s1  };
assign \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.u2.a  = \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.ain_s1 ;
assign \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.u2.b  = \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.bin_s1 ;
assign \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.u2.cin  = \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.carry_s1 ;
assign \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.facout_s2  = \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.u2.cout ;
assign \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.fas_s2  = \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.u2.s ;
assign \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.u1.a  = \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.a [0];
assign \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.u1.b  = \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.b [0];
assign \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.u1.cin  = 1'h0;
assign \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.facout_s1  = \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.u1.cout ;
assign \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.fas_s1  = \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.u1.s ;
assign \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.a  = \add_3s_3s_3_2_1_U19.din0 ;
assign \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.b  = \add_3s_3s_3_2_1_U19.din1 ;
assign \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.ce  = \add_3s_3s_3_2_1_U19.ce ;
assign \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.clk  = \add_3s_3s_3_2_1_U19.clk ;
assign \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.reset  = \add_3s_3s_3_2_1_U19.reset ;
assign \add_3s_3s_3_2_1_U19.dout  = \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.s ;
assign \add_3s_3s_3_2_1_U19.ce  = 1'h1;
assign \add_3s_3s_3_2_1_U19.clk  = ap_clk;
assign \add_3s_3s_3_2_1_U19.din0  = { op_18[1], op_18 };
assign \add_3s_3s_3_2_1_U19.din1  = { op_16_V_reg_1382[1], op_16_V_reg_1382 };
assign grp_fu_836_p2 = \add_3s_3s_3_2_1_U19.dout ;
assign \add_3s_3s_3_2_1_U19.reset  = ap_rst;
assign \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.ain_s0  = \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.a ;
assign \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.bin_s0  = \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.b ;
assign \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.s  = { \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.fas_s2 , \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.sum_s1  };
assign \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.u2.a  = \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.ain_s1 ;
assign \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.u2.b  = \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.bin_s1 ;
assign \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.u2.cin  = \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.carry_s1 ;
assign \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.facout_s2  = \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.u2.cout ;
assign \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.fas_s2  = \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.u2.s ;
assign \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.u1.a  = \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.a [0];
assign \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.u1.b  = \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.b [0];
assign \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.u1.cin  = 1'h0;
assign \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.facout_s1  = \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.u1.cout ;
assign \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.fas_s1  = \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.u1.s ;
assign \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.a  = \add_3ns_3ns_3_2_1_U10.din0 ;
assign \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.b  = \add_3ns_3ns_3_2_1_U10.din1 ;
assign \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.ce  = \add_3ns_3ns_3_2_1_U10.ce ;
assign \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.clk  = \add_3ns_3ns_3_2_1_U10.clk ;
assign \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.reset  = \add_3ns_3ns_3_2_1_U10.reset ;
assign \add_3ns_3ns_3_2_1_U10.dout  = \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.s ;
assign \add_3ns_3ns_3_2_1_U10.ce  = 1'h1;
assign \add_3ns_3ns_3_2_1_U10.clk  = ap_clk;
assign \add_3ns_3ns_3_2_1_U10.din0  = { trunc_ln1192_4_reg_1085, 2'h0 };
assign \add_3ns_3ns_3_2_1_U10.din1  = trunc_ln1192_2_reg_1292;
assign grp_fu_648_p2 = \add_3ns_3ns_3_2_1_U10.dout ;
assign \add_3ns_3ns_3_2_1_U10.reset  = ap_rst;
assign \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.ain_s0  = \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.a ;
assign \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.bin_s0  = \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.b ;
assign \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.s  = { \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.fas_s2 , \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.sum_s1  };
assign \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.u2.a  = \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.ain_s1 ;
assign \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.u2.b  = \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.bin_s1 ;
assign \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.u2.cin  = \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.carry_s1 ;
assign \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.facout_s2  = \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.u2.cout ;
assign \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.fas_s2  = \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.u2.s ;
assign \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.u1.a  = \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.a [16:0];
assign \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.u1.b  = \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.b [16:0];
assign \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.u1.cin  = 1'h0;
assign \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.facout_s1  = \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.u1.cout ;
assign \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.fas_s1  = \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.u1.s ;
assign \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.a  = \add_34s_34s_34_2_1_U23.din0 ;
assign \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.b  = \add_34s_34s_34_2_1_U23.din1 ;
assign \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.ce  = \add_34s_34s_34_2_1_U23.ce ;
assign \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.clk  = \add_34s_34s_34_2_1_U23.clk ;
assign \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.reset  = \add_34s_34s_34_2_1_U23.reset ;
assign \add_34s_34s_34_2_1_U23.dout  = \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.s ;
assign \add_34s_34s_34_2_1_U23.ce  = 1'h1;
assign \add_34s_34s_34_2_1_U23.clk  = ap_clk;
assign \add_34s_34s_34_2_1_U23.din0  = { op_29_V_reg_1543[31], op_29_V_reg_1543, 1'h0 };
assign \add_34s_34s_34_2_1_U23.din1  = { op_19_V_reg_1522[1], op_19_V_reg_1522[1], op_19_V_reg_1522[1], op_19_V_reg_1522[1], op_19_V_reg_1522[1], op_19_V_reg_1522[1], op_19_V_reg_1522[1], op_19_V_reg_1522[1], op_19_V_reg_1522[1], op_19_V_reg_1522[1], op_19_V_reg_1522[1], op_19_V_reg_1522[1], op_19_V_reg_1522[1], op_19_V_reg_1522[1], op_19_V_reg_1522[1], op_19_V_reg_1522[1], op_19_V_reg_1522[1], op_19_V_reg_1522[1], op_19_V_reg_1522[1], op_19_V_reg_1522[1], op_19_V_reg_1522[1], op_19_V_reg_1522[1], op_19_V_reg_1522[1], op_19_V_reg_1522[1], op_19_V_reg_1522[1], op_19_V_reg_1522[1], op_19_V_reg_1522[1], op_19_V_reg_1522[1], op_19_V_reg_1522[1], op_19_V_reg_1522[1], op_19_V_reg_1522[1], op_19_V_reg_1522[1], op_19_V_reg_1522 };
assign grp_fu_988_p2 = \add_34s_34s_34_2_1_U23.dout ;
assign \add_34s_34s_34_2_1_U23.reset  = ap_rst;
assign \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.ain_s0  = \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.a ;
assign \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.bin_s0  = \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.b ;
assign \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.s  = { \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.fas_s2 , \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.sum_s1  };
assign \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.u2.a  = \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.ain_s1 ;
assign \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.u2.b  = \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.bin_s1 ;
assign \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.u2.cin  = \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.carry_s1 ;
assign \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.facout_s2  = \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.u2.cout ;
assign \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.fas_s2  = \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.u2.s ;
assign \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.u1.a  = \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.a [15:0];
assign \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.u1.b  = \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.b [15:0];
assign \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.u1.cin  = 1'h0;
assign \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.facout_s1  = \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.u1.cout ;
assign \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.fas_s1  = \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.u1.s ;
assign \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.a  = \add_32s_32ns_32_2_1_U22.din0 ;
assign \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.b  = \add_32s_32ns_32_2_1_U22.din1 ;
assign \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.ce  = \add_32s_32ns_32_2_1_U22.ce ;
assign \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.clk  = \add_32s_32ns_32_2_1_U22.clk ;
assign \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.reset  = \add_32s_32ns_32_2_1_U22.reset ;
assign \add_32s_32ns_32_2_1_U22.dout  = \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.s ;
assign \add_32s_32ns_32_2_1_U22.ce  = 1'h1;
assign \add_32s_32ns_32_2_1_U22.clk  = ap_clk;
assign \add_32s_32ns_32_2_1_U22.din0  = { add_ln69_6_reg_1533[3], add_ln69_6_reg_1533[3], add_ln69_6_reg_1533[3], add_ln69_6_reg_1533[3], add_ln69_6_reg_1533[3], add_ln69_6_reg_1533[3], add_ln69_6_reg_1533[3], add_ln69_6_reg_1533[3], add_ln69_6_reg_1533[3], add_ln69_6_reg_1533[3], add_ln69_6_reg_1533[3], add_ln69_6_reg_1533[3], add_ln69_6_reg_1533[3], add_ln69_6_reg_1533[3], add_ln69_6_reg_1533[3], add_ln69_6_reg_1533[3], add_ln69_6_reg_1533[3], add_ln69_6_reg_1533[3], add_ln69_6_reg_1533[3], add_ln69_6_reg_1533[3], add_ln69_6_reg_1533[3], add_ln69_6_reg_1533[3], add_ln69_6_reg_1533[3], add_ln69_6_reg_1533[3], add_ln69_6_reg_1533[3], add_ln69_6_reg_1533[3], add_ln69_6_reg_1533[3], add_ln69_6_reg_1533[3], add_ln69_6_reg_1533 };
assign \add_32s_32ns_32_2_1_U22.din1  = add_ln69_4_reg_1528;
assign grp_fu_969_p2 = \add_32s_32ns_32_2_1_U22.dout ;
assign \add_32s_32ns_32_2_1_U22.reset  = ap_rst;
assign \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.ain_s0  = \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.a ;
assign \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.bin_s0  = \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.b ;
assign \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.s  = { \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.fas_s2 , \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.sum_s1  };
assign \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.u2.a  = \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.ain_s1 ;
assign \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.u2.b  = \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.bin_s1 ;
assign \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.u2.cin  = \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.carry_s1 ;
assign \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.facout_s2  = \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.u2.cout ;
assign \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.fas_s2  = \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.u2.s ;
assign \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.u1.a  = \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.a [15:0];
assign \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.u1.b  = \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.b [15:0];
assign \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.u1.cin  = 1'h0;
assign \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.facout_s1  = \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.u1.cout ;
assign \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.fas_s1  = \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.u1.s ;
assign \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.a  = \add_32s_32ns_32_2_1_U18.din0 ;
assign \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.b  = \add_32s_32ns_32_2_1_U18.din1 ;
assign \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.ce  = \add_32s_32ns_32_2_1_U18.ce ;
assign \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.clk  = \add_32s_32ns_32_2_1_U18.clk ;
assign \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.reset  = \add_32s_32ns_32_2_1_U18.reset ;
assign \add_32s_32ns_32_2_1_U18.dout  = \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.s ;
assign \add_32s_32ns_32_2_1_U18.ce  = 1'h1;
assign \add_32s_32ns_32_2_1_U18.clk  = ap_clk;
assign \add_32s_32ns_32_2_1_U18.din0  = { op_14[1], op_14[1], op_14[1], op_14[1], op_14[1], op_14[1], op_14[1], op_14[1], op_14[1], op_14[1], op_14[1], op_14[1], op_14[1], op_14[1], op_14[1], op_14[1], op_14[1], op_14[1], op_14[1], op_14[1], op_14[1], op_14[1], op_14[1], op_14[1], op_14[1], op_14[1], op_14[1], op_14[1], op_14[1], op_14[1], op_14 };
assign \add_32s_32ns_32_2_1_U18.din1  = op_15;
assign grp_fu_830_p2 = \add_32s_32ns_32_2_1_U18.dout ;
assign \add_32s_32ns_32_2_1_U18.reset  = ap_rst;
assign \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.ain_s0  = \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.a ;
assign \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.bin_s0  = \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.b ;
assign \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.s  = { \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.fas_s2 , \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.sum_s1  };
assign \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.u2.a  = \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.ain_s1 ;
assign \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.u2.b  = \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.bin_s1 ;
assign \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.u2.cin  = \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.carry_s1 ;
assign \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.facout_s2  = \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.u2.cout ;
assign \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.fas_s2  = \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.u2.s ;
assign \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.u1.a  = \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.a [15:0];
assign \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.u1.b  = \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.b [15:0];
assign \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.u1.cin  = 1'h0;
assign \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.facout_s1  = \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.u1.cout ;
assign \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.fas_s1  = \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.u1.s ;
assign \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.a  = \add_32ns_32s_32_2_1_U20.din0 ;
assign \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.b  = \add_32ns_32s_32_2_1_U20.din1 ;
assign \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.ce  = \add_32ns_32s_32_2_1_U20.ce ;
assign \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.clk  = \add_32ns_32s_32_2_1_U20.clk ;
assign \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.reset  = \add_32ns_32s_32_2_1_U20.reset ;
assign \add_32ns_32s_32_2_1_U20.dout  = \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.s ;
assign \add_32ns_32s_32_2_1_U20.ce  = 1'h1;
assign \add_32ns_32s_32_2_1_U20.clk  = ap_clk;
assign \add_32ns_32s_32_2_1_U20.din0  = add_ln69_3_reg_1492;
assign \add_32ns_32s_32_2_1_U20.din1  = { ret_V_11_reg_1487[16], ret_V_11_reg_1487[16], ret_V_11_reg_1487[16], ret_V_11_reg_1487[16], ret_V_11_reg_1487[16], ret_V_11_reg_1487[16], ret_V_11_reg_1487[16], ret_V_11_reg_1487[16], ret_V_11_reg_1487[16], ret_V_11_reg_1487[16], ret_V_11_reg_1487[16], ret_V_11_reg_1487[16], ret_V_11_reg_1487[16], ret_V_11_reg_1487[16], ret_V_11_reg_1487[16], ret_V_11_reg_1487 };
assign grp_fu_939_p2 = \add_32ns_32s_32_2_1_U20.dout ;
assign \add_32ns_32s_32_2_1_U20.reset  = ap_rst;
assign \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.ain_s0  = \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.a ;
assign \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.bin_s0  = \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.b ;
assign \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.s  = { \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.fas_s2 , \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.sum_s1  };
assign \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.u2.a  = \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.ain_s1 ;
assign \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.u2.b  = \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.bin_s1 ;
assign \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.u2.cin  = \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.carry_s1 ;
assign \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.facout_s2  = \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.u2.cout ;
assign \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.fas_s2  = \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.u2.s ;
assign \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.u1.a  = \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.a [15:0];
assign \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.u1.b  = \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.b [15:0];
assign \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.u1.cin  = 1'h0;
assign \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.facout_s1  = \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.u1.cout ;
assign \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.fas_s1  = \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.u1.s ;
assign \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.a  = \add_32ns_32ns_32_2_1_U24.din0 ;
assign \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.b  = \add_32ns_32ns_32_2_1_U24.din1 ;
assign \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.ce  = \add_32ns_32ns_32_2_1_U24.ce ;
assign \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.clk  = \add_32ns_32ns_32_2_1_U24.clk ;
assign \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.reset  = \add_32ns_32ns_32_2_1_U24.reset ;
assign \add_32ns_32ns_32_2_1_U24.dout  = \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.s ;
assign \add_32ns_32ns_32_2_1_U24.ce  = 1'h1;
assign \add_32ns_32ns_32_2_1_U24.clk  = ap_clk;
assign \add_32ns_32ns_32_2_1_U24.din0  = ret_V_6_cast_reg_1563;
assign \add_32ns_32ns_32_2_1_U24.din1  = 32'd1;
assign grp_fu_1004_p2 = \add_32ns_32ns_32_2_1_U24.dout ;
assign \add_32ns_32ns_32_2_1_U24.reset  = ap_rst;
assign \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.ain_s0  = \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.a ;
assign \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.bin_s0  = \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.b ;
assign \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.s  = { \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.fas_s2 , \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.sum_s1  };
assign \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.u2.a  = \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.ain_s1 ;
assign \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.u2.b  = \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.bin_s1 ;
assign \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.u2.cin  = \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.carry_s1 ;
assign \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.facout_s2  = \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.u2.cout ;
assign \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.fas_s2  = \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.u2.s ;
assign \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.u1.a  = \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.a [0];
assign \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.u1.b  = \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.b [0];
assign \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.u1.cin  = 1'h0;
assign \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.facout_s1  = \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.u1.cout ;
assign \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.fas_s1  = \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.u1.s ;
assign \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.a  = \add_2ns_2ns_2_2_1_U15.din0 ;
assign \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.b  = \add_2ns_2ns_2_2_1_U15.din1 ;
assign \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.ce  = \add_2ns_2ns_2_2_1_U15.ce ;
assign \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.clk  = \add_2ns_2ns_2_2_1_U15.clk ;
assign \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.reset  = \add_2ns_2ns_2_2_1_U15.reset ;
assign \add_2ns_2ns_2_2_1_U15.dout  = \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.s ;
assign \add_2ns_2ns_2_2_1_U15.ce  = 1'h1;
assign \add_2ns_2ns_2_2_1_U15.clk  = ap_clk;
assign \add_2ns_2ns_2_2_1_U15.din0  = p_Val2_5_reg_1332;
assign \add_2ns_2ns_2_2_1_U15.din1  = { 1'h0, trunc_ln1192_1_reg_1287 };
assign grp_fu_723_p2 = \add_2ns_2ns_2_2_1_U15.dout ;
assign \add_2ns_2ns_2_2_1_U15.reset  = ap_rst;
assign \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.ain_s0  = \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.a ;
assign \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.bin_s0  = \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.b ;
assign \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.s  = { \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.fas_s2 , \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.sum_s1  };
assign \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.u2.a  = \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.ain_s1 ;
assign \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.u2.b  = \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.bin_s1 ;
assign \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.u2.cin  = \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.carry_s1 ;
assign \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.facout_s2  = \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.u2.cout ;
assign \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.fas_s2  = \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.u2.s ;
assign \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.u1.a  = \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.a [7:0];
assign \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.u1.b  = \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.b [7:0];
assign \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.u1.cin  = 1'h0;
assign \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.facout_s1  = \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.u1.cout ;
assign \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.fas_s1  = \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.u1.s ;
assign \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.a  = \add_17s_17s_17_2_1_U11.din0 ;
assign \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.b  = \add_17s_17s_17_2_1_U11.din1 ;
assign \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.ce  = \add_17s_17s_17_2_1_U11.ce ;
assign \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.clk  = \add_17s_17s_17_2_1_U11.clk ;
assign \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.reset  = \add_17s_17s_17_2_1_U11.reset ;
assign \add_17s_17s_17_2_1_U11.dout  = \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.s ;
assign \add_17s_17s_17_2_1_U11.ce  = 1'h1;
assign \add_17s_17s_17_2_1_U11.clk  = ap_clk;
assign \add_17s_17s_17_2_1_U11.din0  = { r_reg_1277[15], r_reg_1277 };
assign \add_17s_17s_17_2_1_U11.din1  = { op_10[7], op_10[7], op_10[7], op_10[7], op_10[7], op_10[7], op_10[7], op_10[7], op_10[7], op_10 };
assign grp_fu_660_p2 = \add_17s_17s_17_2_1_U11.dout ;
assign \add_17s_17s_17_2_1_U11.reset  = ap_rst;
assign \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.ain_s0  = \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.a ;
assign \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.bin_s0  = \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.b ;
assign \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.s  = { \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.fas_s2 , \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.sum_s1  };
assign \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.u2.a  = \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.ain_s1 ;
assign \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.u2.b  = \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.bin_s1 ;
assign \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.u2.cin  = \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.carry_s1 ;
assign \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.facout_s2  = \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.u2.cout ;
assign \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.fas_s2  = \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.u2.s ;
assign \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.u1.a  = \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.a [7:0];
assign \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.u1.b  = \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.b [7:0];
assign \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.u1.cin  = 1'h0;
assign \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.facout_s1  = \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.u1.cout ;
assign \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.fas_s1  = \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.u1.s ;
assign \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.a  = \add_17s_17ns_17_2_1_U16.din0 ;
assign \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.b  = \add_17s_17ns_17_2_1_U16.din1 ;
assign \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.ce  = \add_17s_17ns_17_2_1_U16.ce ;
assign \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.clk  = \add_17s_17ns_17_2_1_U16.clk ;
assign \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.reset  = \add_17s_17ns_17_2_1_U16.reset ;
assign \add_17s_17ns_17_2_1_U16.dout  = \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.s ;
assign \add_17s_17ns_17_2_1_U16.ce  = 1'h1;
assign \add_17s_17ns_17_2_1_U16.clk  = ap_clk;
assign \add_17s_17ns_17_2_1_U16.din0  = { add_ln69_1_reg_1342[6], add_ln69_1_reg_1342[6], add_ln69_1_reg_1342[6], add_ln69_1_reg_1342[6], add_ln69_1_reg_1342[6], add_ln69_1_reg_1342[6], add_ln69_1_reg_1342[6], add_ln69_1_reg_1342[6], add_ln69_1_reg_1342[6], add_ln69_1_reg_1342[6], add_ln69_1_reg_1342 };
assign \add_17s_17ns_17_2_1_U16.din1  = add_ln69_reg_1337;
assign grp_fu_731_p2 = \add_17s_17ns_17_2_1_U16.dout ;
assign \add_17s_17ns_17_2_1_U16.reset  = ap_rst;
assign \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.ain_s0  = \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.a ;
assign \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.bin_s0  = \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.b ;
assign \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.s  = { \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.fas_s2 , \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.sum_s1  };
assign \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.u2.a  = \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.ain_s1 ;
assign \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.u2.b  = \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.bin_s1 ;
assign \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.u2.cin  = \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.carry_s1 ;
assign \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.facout_s2  = \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.u2.cout ;
assign \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.fas_s2  = \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.u2.s ;
assign \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.u1.a  = \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.a [7:0];
assign \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.u1.b  = \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.b [7:0];
assign \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.u1.cin  = 1'h0;
assign \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.facout_s1  = \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.u1.cout ;
assign \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.fas_s1  = \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.u1.s ;
assign \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.a  = \add_17ns_17s_17_2_1_U17.din0 ;
assign \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.b  = \add_17ns_17s_17_2_1_U17.din1 ;
assign \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.ce  = \add_17ns_17s_17_2_1_U17.ce ;
assign \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.clk  = \add_17ns_17s_17_2_1_U17.clk ;
assign \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.reset  = \add_17ns_17s_17_2_1_U17.reset ;
assign \add_17ns_17s_17_2_1_U17.dout  = \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.s ;
assign \add_17ns_17s_17_2_1_U17.ce  = 1'h1;
assign \add_17ns_17s_17_2_1_U17.clk  = ap_clk;
assign \add_17ns_17s_17_2_1_U17.din0  = op_23_V_reg_1422;
assign \add_17ns_17s_17_2_1_U17.din1  = { op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13 };
assign grp_fu_814_p2 = \add_17ns_17s_17_2_1_U17.dout ;
assign \add_17ns_17s_17_2_1_U17.reset  = ap_rst;
endmodule


// Machine B:
// Processed by function `add_clk_enable_signal` in `verilog_tricks.py`.
// Processed by function `remove_reset_signal` in `verilog_tricks.py`.
module top_B (
  ap_clk,
  ap_start,
  ap_done,
  ap_idle,
  ap_ready,
  op_0,
  op_2,
  op_3,
  op_5,
  op_6,
  op_8,
  op_9,
  op_10,
  op_13,
  op_14,
  op_15,
  op_17,
  op_18,
  op_30,
  op_30_ap_vld,
clk_enable
);
input clk_enable;


input ap_clk;
wire ap_rst;
assign ap_rst = op_30_ap_vld;
input ap_start;
input [3:0] op_0;
input [7:0] op_10;
input [1:0] op_13;
input [1:0] op_14;
input [31:0] op_15;
input [1:0] op_17;
input [1:0] op_18;
input [15:0] op_2;
input [3:0] op_3;
input [3:0] op_5;
input [7:0] op_6;
input [3:0] op_8;
input [3:0] op_9;
output ap_done;
output ap_idle;
output ap_ready;
output [31:0] op_30;
output op_30_ap_vld;


reg Range1_all_ones_reg_1444;
reg Range1_all_zeros_reg_1451;
reg Range2_all_ones_reg_1439;
reg [8:0] \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.ain_s1 ;
reg [8:0] \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.bin_s1 ;
reg \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.carry_s1 ;
reg [7:0] \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.sum_s1 ;
reg [8:0] \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.ain_s1 ;
reg [8:0] \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.bin_s1 ;
reg \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.carry_s1 ;
reg [7:0] \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.sum_s1 ;
reg [8:0] \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.ain_s1 ;
reg [8:0] \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.bin_s1 ;
reg \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.carry_s1 ;
reg [7:0] \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.sum_s1 ;
reg \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.ain_s1 ;
reg \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.bin_s1 ;
reg \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.carry_s1 ;
reg \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.sum_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.ain_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.bin_s1 ;
reg \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.carry_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.sum_s1 ;
reg [15:0] \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.ain_s1 ;
reg [15:0] \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.bin_s1 ;
reg \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.carry_s1 ;
reg [15:0] \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.sum_s1 ;
reg [15:0] \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.ain_s1 ;
reg [15:0] \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.bin_s1 ;
reg \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.carry_s1 ;
reg [15:0] \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.sum_s1 ;
reg [15:0] \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.ain_s1 ;
reg [15:0] \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.bin_s1 ;
reg \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.carry_s1 ;
reg [15:0] \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.sum_s1 ;
reg [16:0] \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.ain_s1 ;
reg [16:0] \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.bin_s1 ;
reg \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.carry_s1 ;
reg [16:0] \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.sum_s1 ;
reg [1:0] \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.ain_s1 ;
reg [1:0] \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.bin_s1 ;
reg \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.carry_s1 ;
reg \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.sum_s1 ;
reg [1:0] \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.ain_s1 ;
reg [1:0] \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.bin_s1 ;
reg \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.carry_s1 ;
reg \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.sum_s1 ;
reg [1:0] \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.ain_s1 ;
reg [1:0] \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.bin_s1 ;
reg \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.carry_s1 ;
reg [1:0] \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.sum_s1 ;
reg [1:0] \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.ain_s1 ;
reg [1:0] \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.bin_s1 ;
reg \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.carry_s1 ;
reg [1:0] \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.sum_s1 ;
reg [2:0] \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.ain_s1 ;
reg [2:0] \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.bin_s1 ;
reg \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.carry_s1 ;
reg [2:0] \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.sum_s1 ;
reg [3:0] \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.ain_s1 ;
reg [3:0] \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.bin_s1 ;
reg \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.carry_s1 ;
reg [2:0] \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.sum_s1 ;
reg [3:0] \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.ain_s1 ;
reg [3:0] \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.bin_s1 ;
reg \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.carry_s1 ;
reg [2:0] \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.sum_s1 ;
reg [3:0] \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.ain_s1 ;
reg [3:0] \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.bin_s1 ;
reg \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.carry_s1 ;
reg [2:0] \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.sum_s1 ;
reg [3:0] add_ln1192_1_reg_1387;
reg [2:0] add_ln1192_2_reg_1327;
reg [31:0] add_ln691_reg_1570;
reg [6:0] add_ln69_1_reg_1342;
reg [31:0] add_ln69_3_reg_1492;
reg [31:0] add_ln69_4_reg_1528;
reg [2:0] add_ln69_5_reg_1497;
reg [3:0] add_ln69_6_reg_1533;
reg [16:0] add_ln69_reg_1337;
reg and_ln786_reg_1169;
reg and_ln788_1_reg_1482;
reg [24:0] ap_CS_fsm = 25'h0000001;
reg [15:0] \ashr_16s_16ns_16_7_1_U3.din1_cast_array[0] ;
reg [15:0] \ashr_16s_16ns_16_7_1_U3.din1_cast_array[1] ;
reg [15:0] \ashr_16s_16ns_16_7_1_U3.din1_cast_array[2] ;
reg [15:0] \ashr_16s_16ns_16_7_1_U3.din1_cast_array[3] ;
reg [15:0] \ashr_16s_16ns_16_7_1_U3.din1_cast_array[4] ;
reg [15:0] \ashr_16s_16ns_16_7_1_U3.din1_cast_array[5] ;
reg [15:0] \ashr_16s_16ns_16_7_1_U3.dout_array[0] ;
reg [15:0] \ashr_16s_16ns_16_7_1_U3.dout_array[1] ;
reg [15:0] \ashr_16s_16ns_16_7_1_U3.dout_array[2] ;
reg [15:0] \ashr_16s_16ns_16_7_1_U3.dout_array[3] ;
reg [15:0] \ashr_16s_16ns_16_7_1_U3.dout_array[4] ;
reg [15:0] \ashr_16s_16ns_16_7_1_U3.dout_array[5] ;
reg [7:0] \ashr_32s_8ns_32_7_1_U7.din1_cast_array[0] ;
reg [7:0] \ashr_32s_8ns_32_7_1_U7.din1_cast_array[1] ;
reg [7:0] \ashr_32s_8ns_32_7_1_U7.din1_cast_array[2] ;
reg [7:0] \ashr_32s_8ns_32_7_1_U7.din1_cast_array[3] ;
reg [7:0] \ashr_32s_8ns_32_7_1_U7.din1_cast_array[4] ;
reg [7:0] \ashr_32s_8ns_32_7_1_U7.din1_cast_array[5] ;
reg [31:0] \ashr_32s_8ns_32_7_1_U7.dout_array[0] ;
reg [31:0] \ashr_32s_8ns_32_7_1_U7.dout_array[1] ;
reg [31:0] \ashr_32s_8ns_32_7_1_U7.dout_array[2] ;
reg [31:0] \ashr_32s_8ns_32_7_1_U7.dout_array[3] ;
reg [31:0] \ashr_32s_8ns_32_7_1_U7.dout_array[4] ;
reg [31:0] \ashr_32s_8ns_32_7_1_U7.dout_array[5] ;
reg [15:0] ashr_ln1497_reg_1251;
reg carry_1_reg_1432;
reg icmp_ln213_reg_1266;
reg icmp_ln768_reg_1130;
reg icmp_ln786_reg_1135;
reg op_12_V_reg_1297;
reg [1:0] op_16_V_reg_1382;
reg [1:0] op_19_V_reg_1522;
reg [16:0] op_23_V_reg_1422;
reg [31:0] op_29_V_reg_1543;
reg [3:0] op_7_V_reg_1271;
reg or_ln340_reg_1190;
reg or_ln384_reg_1502;
reg or_ln785_reg_1151;
reg or_ln786_reg_1163;
reg overflow_1_reg_1476;
reg p_Result_10_reg_1098;
reg p_Result_11_reg_1110;
reg p_Result_13_reg_1141;
reg p_Result_14_reg_1392;
reg p_Result_16_reg_1404;
reg [14:0] p_Result_1_reg_1117;
reg [2:0] p_Result_2_reg_1411;
reg [3:0] p_Result_3_reg_1416;
reg [3:0] p_Val2_1_reg_1224;
reg [1:0] p_Val2_5_reg_1332;
reg [1:0] p_Val2_6_reg_1398;
reg [15:0] r_reg_1277;
reg [16:0] ret_V_11_reg_1487;
reg [33:0] ret_V_12_reg_1558;
reg [5:0] ret_V_2_reg_1261;
reg [31:0] ret_V_6_cast_reg_1563;
reg [6:0] ret_V_8_reg_1212;
reg [5:0] ret_V_9_reg_1282;
reg [5:0] ret_V_reg_1217;
reg [16:0] ret_reg_1091;
reg sel_tmp11_reg_1235;
reg [3:0] select_ln340_reg_1230;
reg [3:0] select_ln785_reg_1246;
reg [7:0] sh_V_reg_1175;
reg [15:0] \shl_16s_16ns_16_7_1_U4.din1_cast_array[0] ;
reg [15:0] \shl_16s_16ns_16_7_1_U4.din1_cast_array[1] ;
reg [15:0] \shl_16s_16ns_16_7_1_U4.din1_cast_array[2] ;
reg [15:0] \shl_16s_16ns_16_7_1_U4.din1_cast_array[3] ;
reg [15:0] \shl_16s_16ns_16_7_1_U4.din1_cast_array[4] ;
reg [15:0] \shl_16s_16ns_16_7_1_U4.din1_cast_array[5] ;
reg [15:0] \shl_16s_16ns_16_7_1_U4.dout_array[0] ;
reg [15:0] \shl_16s_16ns_16_7_1_U4.dout_array[1] ;
reg [15:0] \shl_16s_16ns_16_7_1_U4.dout_array[2] ;
reg [15:0] \shl_16s_16ns_16_7_1_U4.dout_array[3] ;
reg [15:0] \shl_16s_16ns_16_7_1_U4.dout_array[4] ;
reg [15:0] \shl_16s_16ns_16_7_1_U4.dout_array[5] ;
reg [7:0] \shl_32s_8ns_32_7_1_U8.din1_cast_array[0] ;
reg [7:0] \shl_32s_8ns_32_7_1_U8.din1_cast_array[1] ;
reg [7:0] \shl_32s_8ns_32_7_1_U8.din1_cast_array[2] ;
reg [7:0] \shl_32s_8ns_32_7_1_U8.din1_cast_array[3] ;
reg [7:0] \shl_32s_8ns_32_7_1_U8.din1_cast_array[4] ;
reg [7:0] \shl_32s_8ns_32_7_1_U8.din1_cast_array[5] ;
reg [31:0] \shl_32s_8ns_32_7_1_U8.dout_array[0] ;
reg [31:0] \shl_32s_8ns_32_7_1_U8.dout_array[1] ;
reg [31:0] \shl_32s_8ns_32_7_1_U8.dout_array[2] ;
reg [31:0] \shl_32s_8ns_32_7_1_U8.dout_array[3] ;
reg [31:0] \shl_32s_8ns_32_7_1_U8.dout_array[4] ;
reg [31:0] \shl_32s_8ns_32_7_1_U8.dout_array[5] ;
reg [15:0] shl_ln1497_reg_1256;
reg [8:0] \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.ain_s1 ;
reg [8:0] \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.bin_s1 ;
reg \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.carry_s1 ;
reg [7:0] \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.sum_s1 ;
reg [2:0] \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.ain_s1 ;
reg [2:0] \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.bin_s1 ;
reg \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.carry_s1 ;
reg [1:0] \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.sum_s1 ;
reg [3:0] \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.ain_s1 ;
reg [3:0] \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.bin_s1 ;
reg \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.carry_s1 ;
reg [3:0] \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.sum_s1 ;
reg [4:0] sub_ln1497_reg_1048;
reg tmp_4_reg_1043;
reg trunc_ln1192_1_reg_1287;
reg [2:0] trunc_ln1192_2_reg_1292;
reg trunc_ln1192_4_reg_1085;
reg [1:0] trunc_ln69_1_reg_1352;
reg [1:0] trunc_ln69_reg_1347;
reg [1:0] trunc_ln731_reg_1105;
reg xor_ln785_reg_1157;
wire _000_;
wire _001_;
wire _002_;
wire [3:0] _003_;
wire [2:0] _004_;
wire [31:0] _005_;
wire [6:0] _006_;
wire [31:0] _007_;
wire [31:0] _008_;
wire [2:0] _009_;
wire [3:0] _010_;
wire [16:0] _011_;
wire _012_;
wire _013_;
wire [24:0] _014_;
wire [15:0] _015_;
wire _016_;
wire _017_;
wire _018_;
wire _019_;
wire _020_;
wire [1:0] _021_;
wire [1:0] _022_;
wire [16:0] _023_;
wire [31:0] _024_;
wire [3:0] _025_;
wire _026_;
wire _027_;
wire _028_;
wire _029_;
wire _030_;
wire _031_;
wire _032_;
wire _033_;
wire _034_;
wire _035_;
wire [14:0] _036_;
wire [2:0] _037_;
wire [3:0] _038_;
wire [1:0] _039_;
wire [1:0] _040_;
wire [1:0] _041_;
wire [15:0] _042_;
wire [16:0] _043_;
wire [33:0] _044_;
wire [5:0] _045_;
wire [31:0] _046_;
wire [6:0] _047_;
wire [5:0] _048_;
wire [5:0] _049_;
wire [16:0] _050_;
wire _051_;
wire [3:0] _052_;
wire [3:0] _053_;
wire [7:0] _054_;
wire [15:0] _055_;
wire [4:0] _056_;
wire _057_;
wire _058_;
wire [2:0] _059_;
wire _060_;
wire [1:0] _061_;
wire [1:0] _062_;
wire [1:0] _063_;
wire _064_;
wire [1:0] _065_;
wire _066_;
wire _067_;
wire _068_;
wire _069_;
wire _070_;
wire _071_;
wire _072_;
wire _073_;
wire _074_;
wire _075_;
wire _076_;
wire _077_;
wire _078_;
wire _079_;
wire [8:0] _080_;
wire [8:0] _081_;
wire _082_;
wire [7:0] _083_;
wire [8:0] _084_;
wire [9:0] _085_;
wire [8:0] _086_;
wire [8:0] _087_;
wire _088_;
wire [7:0] _089_;
wire [8:0] _090_;
wire [9:0] _091_;
wire [8:0] _092_;
wire [8:0] _093_;
wire _094_;
wire [7:0] _095_;
wire [8:0] _096_;
wire [9:0] _097_;
wire _098_;
wire _099_;
wire _100_;
wire _101_;
wire [1:0] _102_;
wire [1:0] _103_;
wire [15:0] _104_;
wire [15:0] _105_;
wire _106_;
wire [15:0] _107_;
wire [16:0] _108_;
wire [16:0] _109_;
wire [15:0] _110_;
wire [15:0] _111_;
wire _112_;
wire [15:0] _113_;
wire [16:0] _114_;
wire [16:0] _115_;
wire [15:0] _116_;
wire [15:0] _117_;
wire _118_;
wire [15:0] _119_;
wire [16:0] _120_;
wire [16:0] _121_;
wire [15:0] _122_;
wire [15:0] _123_;
wire _124_;
wire [15:0] _125_;
wire [16:0] _126_;
wire [16:0] _127_;
wire [16:0] _128_;
wire [16:0] _129_;
wire _130_;
wire [16:0] _131_;
wire [17:0] _132_;
wire [17:0] _133_;
wire [1:0] _134_;
wire [1:0] _135_;
wire _136_;
wire _137_;
wire [1:0] _138_;
wire [2:0] _139_;
wire [1:0] _140_;
wire [1:0] _141_;
wire _142_;
wire _143_;
wire [1:0] _144_;
wire [2:0] _145_;
wire [1:0] _146_;
wire [1:0] _147_;
wire _148_;
wire [1:0] _149_;
wire [2:0] _150_;
wire [2:0] _151_;
wire [1:0] _152_;
wire [1:0] _153_;
wire _154_;
wire [1:0] _155_;
wire [2:0] _156_;
wire [2:0] _157_;
wire [2:0] _158_;
wire [2:0] _159_;
wire _160_;
wire [2:0] _161_;
wire [3:0] _162_;
wire [3:0] _163_;
wire [3:0] _164_;
wire [3:0] _165_;
wire _166_;
wire [2:0] _167_;
wire [3:0] _168_;
wire [4:0] _169_;
wire [3:0] _170_;
wire [3:0] _171_;
wire _172_;
wire [2:0] _173_;
wire [3:0] _174_;
wire [4:0] _175_;
wire [3:0] _176_;
wire [3:0] _177_;
wire _178_;
wire [2:0] _179_;
wire [3:0] _180_;
wire [4:0] _181_;
wire [15:0] _182_;
wire [15:0] _183_;
wire [15:0] _184_;
wire [15:0] _185_;
wire [15:0] _186_;
wire [15:0] _187_;
wire [15:0] _188_;
wire [15:0] _189_;
wire [15:0] _190_;
wire [15:0] _191_;
wire [15:0] _192_;
wire [15:0] _193_;
wire [15:0] _194_;
wire [15:0] _195_;
wire [15:0] _196_;
wire [15:0] _197_;
wire [15:0] _198_;
wire [15:0] _199_;
wire [15:0] _200_;
wire [15:0] _201_;
wire [15:0] _202_;
wire [15:0] _203_;
wire [15:0] _204_;
wire [15:0] _205_;
wire [15:0] _206_;
wire [15:0] _207_;
wire [15:0] _208_;
wire [15:0] _209_;
wire [15:0] _210_;
wire [7:0] _211_;
wire [7:0] _212_;
wire [7:0] _213_;
wire [7:0] _214_;
wire [7:0] _215_;
wire [7:0] _216_;
wire [31:0] _217_;
wire [31:0] _218_;
wire [31:0] _219_;
wire [31:0] _220_;
wire [31:0] _221_;
wire [31:0] _222_;
wire [7:0] _223_;
wire [31:0] _224_;
wire [7:0] _225_;
wire [31:0] _226_;
wire [7:0] _227_;
wire [31:0] _228_;
wire [7:0] _229_;
wire [31:0] _230_;
wire [7:0] _231_;
wire [31:0] _232_;
wire [7:0] _233_;
wire [31:0] _234_;
wire [31:0] _235_;
wire [31:0] _236_;
wire [31:0] _237_;
wire [15:0] _238_;
wire [15:0] _239_;
wire [15:0] _240_;
wire [15:0] _241_;
wire [15:0] _242_;
wire [15:0] _243_;
wire [15:0] _244_;
wire [15:0] _245_;
wire [15:0] _246_;
wire [15:0] _247_;
wire [15:0] _248_;
wire [15:0] _249_;
wire [15:0] _250_;
wire [15:0] _251_;
wire [15:0] _252_;
wire [15:0] _253_;
wire [15:0] _254_;
wire [15:0] _255_;
wire [15:0] _256_;
wire [15:0] _257_;
wire [15:0] _258_;
wire [15:0] _259_;
wire [15:0] _260_;
wire [15:0] _261_;
wire [15:0] _262_;
wire [15:0] _263_;
wire [15:0] _264_;
wire [15:0] _265_;
wire [15:0] _266_;
wire [7:0] _267_;
wire [7:0] _268_;
wire [7:0] _269_;
wire [7:0] _270_;
wire [7:0] _271_;
wire [7:0] _272_;
wire [31:0] _273_;
wire [31:0] _274_;
wire [31:0] _275_;
wire [31:0] _276_;
wire [31:0] _277_;
wire [31:0] _278_;
wire [7:0] _279_;
wire [31:0] _280_;
wire [7:0] _281_;
wire [31:0] _282_;
wire [7:0] _283_;
wire [31:0] _284_;
wire [7:0] _285_;
wire [31:0] _286_;
wire [7:0] _287_;
wire [31:0] _288_;
wire [7:0] _289_;
wire [31:0] _290_;
wire [31:0] _291_;
wire [31:0] _292_;
wire [31:0] _293_;
wire [8:0] _294_;
wire [8:0] _295_;
wire _296_;
wire [7:0] _297_;
wire [8:0] _298_;
wire [9:0] _299_;
wire [2:0] _300_;
wire [2:0] _301_;
wire _302_;
wire [1:0] _303_;
wire [2:0] _304_;
wire [3:0] _305_;
wire [3:0] _306_;
wire [3:0] _307_;
wire _308_;
wire [3:0] _309_;
wire [4:0] _310_;
wire [4:0] _311_;
wire _312_;
wire _313_;
wire _314_;
wire _315_;
wire _316_;
wire _317_;
wire _318_;
wire _319_;
wire _320_;
wire _321_;
wire _322_;
wire _323_;
wire _324_;
wire _325_;
wire _326_;
wire _327_;
wire _328_;
wire _329_;
wire _330_;
wire _331_;
wire _332_;
wire _333_;
wire _334_;
wire _335_;
wire _336_;
wire _337_;
wire _338_;
wire _339_;
wire Range1_all_ones_fu_800_p2;
wire Range1_all_zeros_fu_805_p2;
wire Range2_all_ones_fu_795_p2;
wire \add_17ns_17s_17_2_1_U17.ce ;
wire \add_17ns_17s_17_2_1_U17.clk ;
wire [16:0] \add_17ns_17s_17_2_1_U17.din0 ;
wire [16:0] \add_17ns_17s_17_2_1_U17.din1 ;
wire [16:0] \add_17ns_17s_17_2_1_U17.dout ;
wire \add_17ns_17s_17_2_1_U17.reset ;
wire [16:0] \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.a ;
wire [16:0] \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.ain_s0 ;
wire [16:0] \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.b ;
wire [16:0] \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.bin_s0 ;
wire \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.ce ;
wire \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.clk ;
wire \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.facout_s1 ;
wire \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.facout_s2 ;
wire [7:0] \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.fas_s1 ;
wire [8:0] \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.fas_s2 ;
wire \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.reset ;
wire [16:0] \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.s ;
wire [7:0] \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.u1.a ;
wire [7:0] \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.u1.b ;
wire \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.u1.cin ;
wire \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.u1.cout ;
wire [7:0] \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.u1.s ;
wire [8:0] \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.u2.a ;
wire [8:0] \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.u2.b ;
wire \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.u2.cin ;
wire \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.u2.cout ;
wire [8:0] \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.u2.s ;
wire \add_17s_17ns_17_2_1_U16.ce ;
wire \add_17s_17ns_17_2_1_U16.clk ;
wire [16:0] \add_17s_17ns_17_2_1_U16.din0 ;
wire [16:0] \add_17s_17ns_17_2_1_U16.din1 ;
wire [16:0] \add_17s_17ns_17_2_1_U16.dout ;
wire \add_17s_17ns_17_2_1_U16.reset ;
wire [16:0] \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.a ;
wire [16:0] \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.ain_s0 ;
wire [16:0] \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.b ;
wire [16:0] \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.bin_s0 ;
wire \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.ce ;
wire \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.clk ;
wire \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.facout_s1 ;
wire \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.facout_s2 ;
wire [7:0] \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.fas_s1 ;
wire [8:0] \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.fas_s2 ;
wire \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.reset ;
wire [16:0] \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.s ;
wire [7:0] \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.u1.a ;
wire [7:0] \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.u1.b ;
wire \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.u1.cin ;
wire \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.u1.cout ;
wire [7:0] \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.u1.s ;
wire [8:0] \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.u2.a ;
wire [8:0] \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.u2.b ;
wire \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.u2.cin ;
wire \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.u2.cout ;
wire [8:0] \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.u2.s ;
wire \add_17s_17s_17_2_1_U11.ce ;
wire \add_17s_17s_17_2_1_U11.clk ;
wire [16:0] \add_17s_17s_17_2_1_U11.din0 ;
wire [16:0] \add_17s_17s_17_2_1_U11.din1 ;
wire [16:0] \add_17s_17s_17_2_1_U11.dout ;
wire \add_17s_17s_17_2_1_U11.reset ;
wire [16:0] \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.a ;
wire [16:0] \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.ain_s0 ;
wire [16:0] \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.b ;
wire [16:0] \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.bin_s0 ;
wire \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.ce ;
wire \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.clk ;
wire \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.facout_s1 ;
wire \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.facout_s2 ;
wire [7:0] \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.fas_s1 ;
wire [8:0] \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.fas_s2 ;
wire \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.reset ;
wire [16:0] \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.s ;
wire [7:0] \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.u1.a ;
wire [7:0] \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.u1.b ;
wire \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.u1.cin ;
wire \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.u1.cout ;
wire [7:0] \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.u1.s ;
wire [8:0] \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.u2.a ;
wire [8:0] \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.u2.b ;
wire \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.u2.cin ;
wire \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.u2.cout ;
wire [8:0] \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.u2.s ;
wire \add_2ns_2ns_2_2_1_U15.ce ;
wire \add_2ns_2ns_2_2_1_U15.clk ;
wire [1:0] \add_2ns_2ns_2_2_1_U15.din0 ;
wire [1:0] \add_2ns_2ns_2_2_1_U15.din1 ;
wire [1:0] \add_2ns_2ns_2_2_1_U15.dout ;
wire \add_2ns_2ns_2_2_1_U15.reset ;
wire [1:0] \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.a ;
wire [1:0] \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.ain_s0 ;
wire [1:0] \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.b ;
wire [1:0] \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.bin_s0 ;
wire \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.ce ;
wire \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.clk ;
wire \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.facout_s1 ;
wire \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.facout_s2 ;
wire \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.fas_s1 ;
wire \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.fas_s2 ;
wire \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.reset ;
wire [1:0] \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.s ;
wire \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.u1.a ;
wire \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.u1.b ;
wire \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.u1.cin ;
wire \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.u1.cout ;
wire \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.u1.s ;
wire \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.u2.a ;
wire \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.u2.b ;
wire \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.u2.cin ;
wire \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.u2.cout ;
wire \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.u2.s ;
wire \add_32ns_32ns_32_2_1_U24.ce ;
wire \add_32ns_32ns_32_2_1_U24.clk ;
wire [31:0] \add_32ns_32ns_32_2_1_U24.din0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U24.din1 ;
wire [31:0] \add_32ns_32ns_32_2_1_U24.dout ;
wire \add_32ns_32ns_32_2_1_U24.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.a ;
wire [31:0] \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.ain_s0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.b ;
wire [31:0] \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.bin_s0 ;
wire \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.ce ;
wire \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.clk ;
wire \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.facout_s1 ;
wire \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.facout_s2 ;
wire [15:0] \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.fas_s1 ;
wire [15:0] \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.fas_s2 ;
wire \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.u1.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.u1.b ;
wire \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.u1.cin ;
wire \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.u1.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.u1.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.u2.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.u2.b ;
wire \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.u2.cin ;
wire \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.u2.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.u2.s ;
wire \add_32ns_32s_32_2_1_U20.ce ;
wire \add_32ns_32s_32_2_1_U20.clk ;
wire [31:0] \add_32ns_32s_32_2_1_U20.din0 ;
wire [31:0] \add_32ns_32s_32_2_1_U20.din1 ;
wire [31:0] \add_32ns_32s_32_2_1_U20.dout ;
wire \add_32ns_32s_32_2_1_U20.reset ;
wire [31:0] \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.a ;
wire [31:0] \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.ain_s0 ;
wire [31:0] \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.b ;
wire [31:0] \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.bin_s0 ;
wire \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.ce ;
wire \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.clk ;
wire \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.facout_s1 ;
wire \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.facout_s2 ;
wire [15:0] \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.fas_s1 ;
wire [15:0] \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.fas_s2 ;
wire \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.reset ;
wire [31:0] \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.s ;
wire [15:0] \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.u1.a ;
wire [15:0] \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.u1.b ;
wire \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.u1.cin ;
wire \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.u1.cout ;
wire [15:0] \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.u1.s ;
wire [15:0] \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.u2.a ;
wire [15:0] \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.u2.b ;
wire \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.u2.cin ;
wire \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.u2.cout ;
wire [15:0] \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.u2.s ;
wire \add_32s_32ns_32_2_1_U18.ce ;
wire \add_32s_32ns_32_2_1_U18.clk ;
wire [31:0] \add_32s_32ns_32_2_1_U18.din0 ;
wire [31:0] \add_32s_32ns_32_2_1_U18.din1 ;
wire [31:0] \add_32s_32ns_32_2_1_U18.dout ;
wire \add_32s_32ns_32_2_1_U18.reset ;
wire [31:0] \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.a ;
wire [31:0] \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.ain_s0 ;
wire [31:0] \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.b ;
wire [31:0] \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.bin_s0 ;
wire \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.ce ;
wire \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.clk ;
wire \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.facout_s1 ;
wire \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.facout_s2 ;
wire [15:0] \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.fas_s1 ;
wire [15:0] \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.fas_s2 ;
wire \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.reset ;
wire [31:0] \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.s ;
wire [15:0] \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.u1.a ;
wire [15:0] \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.u1.b ;
wire \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.u1.cin ;
wire \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.u1.cout ;
wire [15:0] \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.u1.s ;
wire [15:0] \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.u2.a ;
wire [15:0] \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.u2.b ;
wire \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.u2.cin ;
wire \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.u2.cout ;
wire [15:0] \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.u2.s ;
wire \add_32s_32ns_32_2_1_U22.ce ;
wire \add_32s_32ns_32_2_1_U22.clk ;
wire [31:0] \add_32s_32ns_32_2_1_U22.din0 ;
wire [31:0] \add_32s_32ns_32_2_1_U22.din1 ;
wire [31:0] \add_32s_32ns_32_2_1_U22.dout ;
wire \add_32s_32ns_32_2_1_U22.reset ;
wire [31:0] \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.a ;
wire [31:0] \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.ain_s0 ;
wire [31:0] \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.b ;
wire [31:0] \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.bin_s0 ;
wire \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.ce ;
wire \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.clk ;
wire \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.facout_s1 ;
wire \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.facout_s2 ;
wire [15:0] \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.fas_s1 ;
wire [15:0] \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.fas_s2 ;
wire \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.reset ;
wire [31:0] \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.s ;
wire [15:0] \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.u1.a ;
wire [15:0] \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.u1.b ;
wire \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.u1.cin ;
wire \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.u1.cout ;
wire [15:0] \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.u1.s ;
wire [15:0] \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.u2.a ;
wire [15:0] \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.u2.b ;
wire \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.u2.cin ;
wire \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.u2.cout ;
wire [15:0] \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.u2.s ;
wire \add_34s_34s_34_2_1_U23.ce ;
wire \add_34s_34s_34_2_1_U23.clk ;
wire [33:0] \add_34s_34s_34_2_1_U23.din0 ;
wire [33:0] \add_34s_34s_34_2_1_U23.din1 ;
wire [33:0] \add_34s_34s_34_2_1_U23.dout ;
wire \add_34s_34s_34_2_1_U23.reset ;
wire [33:0] \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.a ;
wire [33:0] \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.ain_s0 ;
wire [33:0] \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.b ;
wire [33:0] \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.bin_s0 ;
wire \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.ce ;
wire \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.clk ;
wire \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.facout_s1 ;
wire \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.facout_s2 ;
wire [16:0] \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.fas_s1 ;
wire [16:0] \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.fas_s2 ;
wire \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.reset ;
wire [33:0] \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.s ;
wire [16:0] \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.u1.a ;
wire [16:0] \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.u1.b ;
wire \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.u1.cin ;
wire \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.u1.cout ;
wire [16:0] \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.u1.s ;
wire [16:0] \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.u2.a ;
wire [16:0] \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.u2.b ;
wire \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.u2.cin ;
wire \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.u2.cout ;
wire [16:0] \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.u2.s ;
wire \add_3ns_3ns_3_2_1_U10.ce ;
wire \add_3ns_3ns_3_2_1_U10.clk ;
wire [2:0] \add_3ns_3ns_3_2_1_U10.din0 ;
wire [2:0] \add_3ns_3ns_3_2_1_U10.din1 ;
wire [2:0] \add_3ns_3ns_3_2_1_U10.dout ;
wire \add_3ns_3ns_3_2_1_U10.reset ;
wire [2:0] \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.a ;
wire [2:0] \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.ain_s0 ;
wire [2:0] \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.b ;
wire [2:0] \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.bin_s0 ;
wire \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.ce ;
wire \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.clk ;
wire \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.facout_s1 ;
wire \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.facout_s2 ;
wire \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.fas_s1 ;
wire [1:0] \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.fas_s2 ;
wire \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.reset ;
wire [2:0] \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.s ;
wire \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.u1.a ;
wire \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.u1.b ;
wire \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.u1.cin ;
wire \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.u1.cout ;
wire \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.u1.s ;
wire [1:0] \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.u2.a ;
wire [1:0] \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.u2.b ;
wire \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.u2.cin ;
wire \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.u2.cout ;
wire [1:0] \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.u2.s ;
wire \add_3s_3s_3_2_1_U19.ce ;
wire \add_3s_3s_3_2_1_U19.clk ;
wire [2:0] \add_3s_3s_3_2_1_U19.din0 ;
wire [2:0] \add_3s_3s_3_2_1_U19.din1 ;
wire [2:0] \add_3s_3s_3_2_1_U19.dout ;
wire \add_3s_3s_3_2_1_U19.reset ;
wire [2:0] \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.a ;
wire [2:0] \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.ain_s0 ;
wire [2:0] \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.b ;
wire [2:0] \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.bin_s0 ;
wire \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.ce ;
wire \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.clk ;
wire \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.facout_s1 ;
wire \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.facout_s2 ;
wire \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.fas_s1 ;
wire [1:0] \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.fas_s2 ;
wire \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.reset ;
wire [2:0] \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.s ;
wire \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.u1.a ;
wire \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.u1.b ;
wire \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.u1.cin ;
wire \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.u1.cout ;
wire \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.u1.s ;
wire [1:0] \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.u2.a ;
wire [1:0] \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.u2.b ;
wire \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.u2.cin ;
wire \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.u2.cout ;
wire [1:0] \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.u2.s ;
wire \add_4ns_4s_4_2_1_U14.ce ;
wire \add_4ns_4s_4_2_1_U14.clk ;
wire [3:0] \add_4ns_4s_4_2_1_U14.din0 ;
wire [3:0] \add_4ns_4s_4_2_1_U14.din1 ;
wire [3:0] \add_4ns_4s_4_2_1_U14.dout ;
wire \add_4ns_4s_4_2_1_U14.reset ;
wire [3:0] \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.a ;
wire [3:0] \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.ain_s0 ;
wire [3:0] \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.b ;
wire [3:0] \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.bin_s0 ;
wire \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.ce ;
wire \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.clk ;
wire \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.facout_s1 ;
wire \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.facout_s2 ;
wire [1:0] \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.fas_s1 ;
wire [1:0] \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.fas_s2 ;
wire \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.reset ;
wire [3:0] \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.s ;
wire [1:0] \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.u1.a ;
wire [1:0] \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.u1.b ;
wire \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.u1.cin ;
wire \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.u1.cout ;
wire [1:0] \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.u1.s ;
wire [1:0] \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.u2.a ;
wire [1:0] \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.u2.b ;
wire \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.u2.cin ;
wire \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.u2.cout ;
wire [1:0] \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.u2.s ;
wire \add_4s_4s_4_2_1_U21.ce ;
wire \add_4s_4s_4_2_1_U21.clk ;
wire [3:0] \add_4s_4s_4_2_1_U21.din0 ;
wire [3:0] \add_4s_4s_4_2_1_U21.din1 ;
wire [3:0] \add_4s_4s_4_2_1_U21.dout ;
wire \add_4s_4s_4_2_1_U21.reset ;
wire [3:0] \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.a ;
wire [3:0] \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.ain_s0 ;
wire [3:0] \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.b ;
wire [3:0] \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.bin_s0 ;
wire \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.ce ;
wire \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.clk ;
wire \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.facout_s1 ;
wire \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.facout_s2 ;
wire [1:0] \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.fas_s1 ;
wire [1:0] \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.fas_s2 ;
wire \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.reset ;
wire [3:0] \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.s ;
wire [1:0] \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.u1.a ;
wire [1:0] \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.u1.b ;
wire \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.u1.cin ;
wire \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.u1.cout ;
wire [1:0] \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.u1.s ;
wire [1:0] \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.u2.a ;
wire [1:0] \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.u2.b ;
wire \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.u2.cin ;
wire \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.u2.cout ;
wire [1:0] \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.u2.s ;
wire \add_6ns_6ns_6_2_1_U9.ce ;
wire \add_6ns_6ns_6_2_1_U9.clk ;
wire [5:0] \add_6ns_6ns_6_2_1_U9.din0 ;
wire [5:0] \add_6ns_6ns_6_2_1_U9.din1 ;
wire [5:0] \add_6ns_6ns_6_2_1_U9.dout ;
wire \add_6ns_6ns_6_2_1_U9.reset ;
wire [5:0] \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.a ;
wire [5:0] \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.ain_s0 ;
wire [5:0] \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.b ;
wire [5:0] \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.bin_s0 ;
wire \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.ce ;
wire \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.clk ;
wire \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.facout_s1 ;
wire \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.facout_s2 ;
wire [2:0] \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.fas_s1 ;
wire [2:0] \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.fas_s2 ;
wire \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.reset ;
wire [5:0] \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.s ;
wire [2:0] \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.u1.a ;
wire [2:0] \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.u1.b ;
wire \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.u1.cin ;
wire \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.u1.cout ;
wire [2:0] \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.u1.s ;
wire [2:0] \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.u2.a ;
wire [2:0] \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.u2.b ;
wire \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.u2.cin ;
wire \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.u2.cout ;
wire [2:0] \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.u2.s ;
wire \add_7ns_7s_7_2_1_U6.ce ;
wire \add_7ns_7s_7_2_1_U6.clk ;
wire [6:0] \add_7ns_7s_7_2_1_U6.din0 ;
wire [6:0] \add_7ns_7s_7_2_1_U6.din1 ;
wire [6:0] \add_7ns_7s_7_2_1_U6.dout ;
wire \add_7ns_7s_7_2_1_U6.reset ;
wire [6:0] \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.a ;
wire [6:0] \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.ain_s0 ;
wire [6:0] \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.b ;
wire [6:0] \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.bin_s0 ;
wire \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.ce ;
wire \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.clk ;
wire \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.facout_s1 ;
wire \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.facout_s2 ;
wire [2:0] \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.fas_s1 ;
wire [3:0] \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.fas_s2 ;
wire \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.reset ;
wire [6:0] \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.s ;
wire [2:0] \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.u1.a ;
wire [2:0] \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.u1.b ;
wire \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.u1.cin ;
wire \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.u1.cout ;
wire [2:0] \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.u1.s ;
wire [3:0] \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.u2.a ;
wire [3:0] \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.u2.b ;
wire \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.u2.cin ;
wire \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.u2.cout ;
wire [3:0] \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.u2.s ;
wire \add_7s_7ns_7_2_1_U12.ce ;
wire \add_7s_7ns_7_2_1_U12.clk ;
wire [6:0] \add_7s_7ns_7_2_1_U12.din0 ;
wire [6:0] \add_7s_7ns_7_2_1_U12.din1 ;
wire [6:0] \add_7s_7ns_7_2_1_U12.dout ;
wire \add_7s_7ns_7_2_1_U12.reset ;
wire [6:0] \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.a ;
wire [6:0] \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.ain_s0 ;
wire [6:0] \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.b ;
wire [6:0] \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.bin_s0 ;
wire \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.ce ;
wire \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.clk ;
wire \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.facout_s1 ;
wire \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.facout_s2 ;
wire [2:0] \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.fas_s1 ;
wire [3:0] \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.fas_s2 ;
wire \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.reset ;
wire [6:0] \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.s ;
wire [2:0] \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.u1.a ;
wire [2:0] \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.u1.b ;
wire \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.u1.cin ;
wire \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.u1.cout ;
wire [2:0] \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.u1.s ;
wire [3:0] \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.u2.a ;
wire [3:0] \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.u2.b ;
wire \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.u2.cin ;
wire \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.u2.cout ;
wire [3:0] \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.u2.s ;
wire \add_7s_7s_7_2_1_U13.ce ;
wire \add_7s_7s_7_2_1_U13.clk ;
wire [6:0] \add_7s_7s_7_2_1_U13.din0 ;
wire [6:0] \add_7s_7s_7_2_1_U13.din1 ;
wire [6:0] \add_7s_7s_7_2_1_U13.dout ;
wire \add_7s_7s_7_2_1_U13.reset ;
wire [6:0] \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.a ;
wire [6:0] \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.ain_s0 ;
wire [6:0] \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.b ;
wire [6:0] \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.bin_s0 ;
wire \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.ce ;
wire \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.clk ;
wire \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.facout_s1 ;
wire \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.facout_s2 ;
wire [2:0] \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.fas_s1 ;
wire [3:0] \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.fas_s2 ;
wire \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.reset ;
wire [6:0] \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.s ;
wire [2:0] \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.u1.a ;
wire [2:0] \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.u1.b ;
wire \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.u1.cin ;
wire \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.u1.cout ;
wire [2:0] \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.u1.s ;
wire [3:0] \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.u2.a ;
wire [3:0] \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.u2.b ;
wire \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.u2.cin ;
wire \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.u2.cout ;
wire [3:0] \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.u2.s ;
wire and_ln213_fu_624_p2;
wire and_ln340_1_fu_506_p2;
wire and_ln340_fu_493_p2;
wire and_ln780_fu_860_p2;
wire and_ln781_fu_907_p2;
wire and_ln785_1_fu_510_p2;
wire and_ln785_fu_551_p2;
wire and_ln786_fu_365_p2;
wire and_ln788_1_fu_902_p2;
wire and_ln788_fu_896_p2;
wire ap_CS_fsm_state1;
wire ap_CS_fsm_state10;
wire ap_CS_fsm_state11;
wire ap_CS_fsm_state12;
wire ap_CS_fsm_state13;
wire ap_CS_fsm_state14;
wire ap_CS_fsm_state15;
wire ap_CS_fsm_state16;
wire ap_CS_fsm_state17;
wire ap_CS_fsm_state18;
wire ap_CS_fsm_state19;
wire ap_CS_fsm_state2;
wire ap_CS_fsm_state20;
wire ap_CS_fsm_state21;
wire ap_CS_fsm_state22;
wire ap_CS_fsm_state23;
wire ap_CS_fsm_state24;
wire ap_CS_fsm_state25;
wire ap_CS_fsm_state3;
wire ap_CS_fsm_state4;
wire ap_CS_fsm_state5;
wire ap_CS_fsm_state6;
wire ap_CS_fsm_state7;
wire ap_CS_fsm_state8;
wire ap_CS_fsm_state9;
wire [24:0] ap_NS_fsm;
wire ap_clk;
wire ap_done;
wire ap_idle;
wire ap_ready;
wire ap_rst;
wire ap_start;
wire \ashr_16s_16ns_16_7_1_U3.ce ;
wire \ashr_16s_16ns_16_7_1_U3.clk ;
wire [15:0] \ashr_16s_16ns_16_7_1_U3.din0 ;
wire [15:0] \ashr_16s_16ns_16_7_1_U3.din1 ;
wire [15:0] \ashr_16s_16ns_16_7_1_U3.din1_cast ;
wire [15:0] \ashr_16s_16ns_16_7_1_U3.din1_mask ;
wire [15:0] \ashr_16s_16ns_16_7_1_U3.dout ;
wire \ashr_16s_16ns_16_7_1_U3.reset ;
wire \ashr_32s_8ns_32_7_1_U7.ce ;
wire \ashr_32s_8ns_32_7_1_U7.clk ;
wire [31:0] \ashr_32s_8ns_32_7_1_U7.din0 ;
wire [31:0] \ashr_32s_8ns_32_7_1_U7.din1 ;
wire [7:0] \ashr_32s_8ns_32_7_1_U7.din1_cast ;
wire [7:0] \ashr_32s_8ns_32_7_1_U7.din1_mask ;
wire [31:0] \ashr_32s_8ns_32_7_1_U7.dout ;
wire \ashr_32s_8ns_32_7_1_U7.reset ;
wire carry_1_fu_789_p2;
wire deleted_ones_fu_865_p3;
wire deleted_zeros_fu_842_p3;
wire [31:0] grp_fu_1004_p2;
wire [4:0] grp_fu_237_p1;
wire [4:0] grp_fu_237_p2;
wire [16:0] grp_fu_251_p0;
wire [16:0] grp_fu_251_p1;
wire [16:0] grp_fu_251_p2;
wire [15:0] grp_fu_264_p1;
wire [15:0] grp_fu_264_p2;
wire [15:0] grp_fu_277_p1;
wire [15:0] grp_fu_277_p2;
wire [7:0] grp_fu_335_p2;
wire [6:0] grp_fu_386_p0;
wire [6:0] grp_fu_386_p1;
wire [6:0] grp_fu_386_p2;
wire [31:0] grp_fu_407_p1;
wire [31:0] grp_fu_407_p2;
wire [31:0] grp_fu_416_p1;
wire [31:0] grp_fu_416_p2;
wire [5:0] grp_fu_526_p2;
wire [2:0] grp_fu_648_p0;
wire [2:0] grp_fu_648_p2;
wire [16:0] grp_fu_660_p0;
wire [16:0] grp_fu_660_p1;
wire [16:0] grp_fu_660_p2;
wire [6:0] grp_fu_666_p0;
wire [6:0] grp_fu_666_p1;
wire [6:0] grp_fu_666_p2;
wire [6:0] grp_fu_709_p0;
wire [6:0] grp_fu_709_p1;
wire [6:0] grp_fu_709_p2;
wire [3:0] grp_fu_715_p0;
wire [3:0] grp_fu_715_p2;
wire [1:0] grp_fu_723_p1;
wire [1:0] grp_fu_723_p2;
wire [16:0] grp_fu_731_p0;
wire [16:0] grp_fu_731_p2;
wire [16:0] grp_fu_814_p1;
wire [16:0] grp_fu_814_p2;
wire [31:0] grp_fu_830_p0;
wire [31:0] grp_fu_830_p2;
wire [2:0] grp_fu_836_p0;
wire [2:0] grp_fu_836_p1;
wire [2:0] grp_fu_836_p2;
wire [31:0] grp_fu_939_p1;
wire [31:0] grp_fu_939_p2;
wire [3:0] grp_fu_947_p0;
wire [3:0] grp_fu_947_p1;
wire [3:0] grp_fu_947_p2;
wire [31:0] grp_fu_969_p0;
wire [31:0] grp_fu_969_p2;
wire [33:0] grp_fu_988_p0;
wire [33:0] grp_fu_988_p1;
wire [33:0] grp_fu_988_p2;
wire icmp_ln213_fu_562_p2;
wire icmp_ln768_fu_317_p2;
wire icmp_ln786_fu_322_p2;
wire [3:0] lhs_V_1_fu_690_p1;
wire [5:0] lhs_V_1_fu_690_p3;
wire [4:0] lhs_V_fu_370_p3;
wire [3:0] op_0;
wire [7:0] op_10;
wire op_12_V_fu_629_p2;
wire [1:0] op_13;
wire [1:0] op_14;
wire [31:0] op_15;
wire [1:0] op_16_V_fu_736_p3;
wire [1:0] op_17;
wire [1:0] op_18;
wire [1:0] op_19_V_fu_960_p3;
wire [15:0] op_2;
wire [3:0] op_3;
wire [31:0] op_30;
wire op_30_ap_vld;
wire [3:0] op_5;
wire [7:0] op_6;
wire [3:0] op_7_V_fu_568_p3;
wire [3:0] op_8;
wire [3:0] op_9;
wire or_ln213_fu_619_p2;
wire or_ln340_fu_396_p2;
wire or_ln384_fu_927_p2;
wire or_ln785_1_fu_877_p2;
wire or_ln785_2_fu_546_p2;
wire or_ln785_3_fu_514_p2;
wire or_ln785_fu_341_p2;
wire or_ln786_fu_355_p2;
wire or_ln788_fu_911_p2;
wire overflow_1_fu_887_p2;
wire overflow_fu_392_p2;
wire p_Result_12_fu_439_p3;
wire [7:0] p_Result_13_fu_327_p1;
wire p_Result_15_fu_777_p3;
wire p_Result_5_fu_578_p3;
wire p_Result_9_fu_1009_p3;
wire [3:0] p_Result_s_14_fu_478_p4;
wire [1:0] p_Result_s_fu_531_p4;
wire [3:0] p_Val2_1_fu_432_p3;
wire [2:0] p_Val2_2_fu_472_p2;
wire [15:0] r_fu_573_p3;
wire [5:0] ret_V_9_fu_594_p3;
wire [32:0] rhs_3_fu_977_p3;
wire sel_tmp11_fu_520_p2;
wire [3:0] select_ln340_fu_498_p3;
wire [1:0] select_ln384_fu_953_p3;
wire [3:0] select_ln785_fu_556_p3;
wire [31:0] select_ln850_1_fu_1019_p3;
wire [5:0] select_ln850_fu_588_p3;
wire [31:0] sext_ln1497_1_fu_270_p1;
wire [3:0] sext_ln1497_fu_225_p0;
wire [3:0] sext_ln215_1_fu_247_p0;
wire [15:0] sext_ln215_fu_243_p0;
wire [3:0] sext_ln545_fu_257_p0;
wire [31:0] sext_ln545_fu_257_p1;
wire [3:0] sext_ln703_fu_382_p0;
wire [7:0] sext_ln781_fu_401_p0;
wire [31:0] sext_ln781_fu_401_p1;
wire \shl_16s_16ns_16_7_1_U4.ce ;
wire \shl_16s_16ns_16_7_1_U4.clk ;
wire [15:0] \shl_16s_16ns_16_7_1_U4.din0 ;
wire [15:0] \shl_16s_16ns_16_7_1_U4.din1 ;
wire [15:0] \shl_16s_16ns_16_7_1_U4.din1_cast ;
wire [15:0] \shl_16s_16ns_16_7_1_U4.din1_mask ;
wire [15:0] \shl_16s_16ns_16_7_1_U4.dout ;
wire \shl_16s_16ns_16_7_1_U4.reset ;
wire \shl_32s_8ns_32_7_1_U8.ce ;
wire \shl_32s_8ns_32_7_1_U8.clk ;
wire [31:0] \shl_32s_8ns_32_7_1_U8.din0 ;
wire [31:0] \shl_32s_8ns_32_7_1_U8.din1 ;
wire [7:0] \shl_32s_8ns_32_7_1_U8.din1_cast ;
wire [7:0] \shl_32s_8ns_32_7_1_U8.din1_mask ;
wire [31:0] \shl_32s_8ns_32_7_1_U8.dout ;
wire \shl_32s_8ns_32_7_1_U8.reset ;
wire [3:0] shl_ln1192_fu_704_p0;
wire \sub_17s_17s_17_2_1_U2.ce ;
wire \sub_17s_17s_17_2_1_U2.clk ;
wire [16:0] \sub_17s_17s_17_2_1_U2.din0 ;
wire [16:0] \sub_17s_17s_17_2_1_U2.din1 ;
wire [16:0] \sub_17s_17s_17_2_1_U2.dout ;
wire \sub_17s_17s_17_2_1_U2.reset ;
wire [16:0] \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.a ;
wire [16:0] \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.ain_s0 ;
wire [16:0] \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.b ;
wire [16:0] \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.bin_s0 ;
wire \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.ce ;
wire \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.clk ;
wire \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.facout_s1 ;
wire \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.facout_s2 ;
wire [7:0] \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.fas_s1 ;
wire [8:0] \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.fas_s2 ;
wire \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.reset ;
wire [16:0] \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.s ;
wire [7:0] \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.u1.a ;
wire [7:0] \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.u1.b ;
wire \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.u1.cin ;
wire \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.u1.cout ;
wire [7:0] \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.u1.s ;
wire [8:0] \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.u2.a ;
wire [8:0] \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.u2.b ;
wire \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.u2.cin ;
wire \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.u2.cout ;
wire [8:0] \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.u2.s ;
wire \sub_5ns_5s_5_2_1_U1.ce ;
wire \sub_5ns_5s_5_2_1_U1.clk ;
wire [4:0] \sub_5ns_5s_5_2_1_U1.din0 ;
wire [4:0] \sub_5ns_5s_5_2_1_U1.din1 ;
wire [4:0] \sub_5ns_5s_5_2_1_U1.dout ;
wire \sub_5ns_5s_5_2_1_U1.reset ;
wire [4:0] \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.a ;
wire [4:0] \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.ain_s0 ;
wire [4:0] \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.b ;
wire [4:0] \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.bin_s0 ;
wire \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.ce ;
wire \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.clk ;
wire \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.facout_s1 ;
wire \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.facout_s2 ;
wire [1:0] \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.fas_s1 ;
wire [2:0] \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.fas_s2 ;
wire \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.reset ;
wire [4:0] \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.s ;
wire [1:0] \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.u1.a ;
wire [1:0] \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.u1.b ;
wire \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.u1.cin ;
wire \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.u1.cout ;
wire [1:0] \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.u1.s ;
wire [2:0] \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.u2.a ;
wire [2:0] \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.u2.b ;
wire \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.u2.cin ;
wire \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.u2.cout ;
wire [2:0] \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.u2.s ;
wire \sub_8ns_8s_8_2_1_U5.ce ;
wire \sub_8ns_8s_8_2_1_U5.clk ;
wire [7:0] \sub_8ns_8s_8_2_1_U5.din0 ;
wire [7:0] \sub_8ns_8s_8_2_1_U5.din1 ;
wire [7:0] \sub_8ns_8s_8_2_1_U5.dout ;
wire \sub_8ns_8s_8_2_1_U5.reset ;
wire [7:0] \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.a ;
wire [7:0] \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.ain_s0 ;
wire [7:0] \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.b ;
wire [7:0] \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.bin_s0 ;
wire \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.ce ;
wire \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.clk ;
wire \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.facout_s1 ;
wire \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.facout_s2 ;
wire [3:0] \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.fas_s1 ;
wire [3:0] \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.fas_s2 ;
wire \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.reset ;
wire [7:0] \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.s ;
wire [3:0] \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.u1.a ;
wire [3:0] \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.u1.b ;
wire \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.u1.cin ;
wire \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.u1.cout ;
wire [3:0] \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.u1.s ;
wire [3:0] \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.u2.a ;
wire [3:0] \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.u2.b ;
wire \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.u2.cin ;
wire \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.u2.cout ;
wire [3:0] \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.u2.s ;
wire tmp_10_fu_612_p3;
wire tmp_1_fu_453_p3;
wire [3:0] tmp_4_fu_229_p1;
wire tmp_9_fu_847_p3;
wire tmp_fu_446_p3;
wire trunc_ln1192_1_fu_604_p1;
wire [2:0] trunc_ln1192_2_fu_608_p1;
wire [3:0] trunc_ln1192_4_fu_283_p0;
wire trunc_ln1192_4_fu_283_p1;
wire trunc_ln1192_fu_601_p1;
wire [1:0] trunc_ln69_1_fu_686_p1;
wire [1:0] trunc_ln69_fu_682_p1;
wire [1:0] trunc_ln731_fu_295_p1;
wire trunc_ln790_fu_893_p1;
wire trunc_ln851_1_fu_1016_p1;
wire [3:0] trunc_ln851_fu_585_p0;
wire trunc_ln851_fu_585_p1;
wire underflow_1_fu_922_p2;
wire xor_ln340_fu_488_p2;
wire xor_ln365_1_fu_466_p2;
wire xor_ln365_fu_460_p2;
wire xor_ln416_fu_784_p2;
wire xor_ln780_fu_854_p2;
wire xor_ln785_1_fu_871_p2;
wire xor_ln785_2_fu_882_p2;
wire xor_ln785_3_fu_541_p2;
wire xor_ln785_fu_345_p2;
wire xor_ln786_1_fu_360_p2;
wire xor_ln786_fu_350_p2;
wire xor_ln788_fu_916_p2;
wire [7:0] zext_ln546_1_fu_413_p0;


assign _066_ = _073_ & ap_CS_fsm[8];
assign _067_ = ap_CS_fsm[8] & _074_;
assign _068_ = tmp_4_reg_1043 & ap_CS_fsm[8];
assign _069_ = ap_CS_fsm[12] & _075_;
assign _070_ = ap_CS_fsm[12] & p_Result_13_reg_1141;
assign _071_ = _076_ & ap_CS_fsm[0];
assign _072_ = ap_start & ap_CS_fsm[0];
assign and_ln213_fu_624_p2 = trunc_ln1192_4_reg_1085 & or_ln213_fu_619_p2;
assign and_ln340_1_fu_506_p2 = or_ln786_reg_1163 & or_ln340_reg_1190;
assign and_ln340_fu_493_p2 = xor_ln340_fu_488_p2 & or_ln786_reg_1163;
assign and_ln780_fu_860_p2 = xor_ln780_fu_854_p2 & Range2_all_ones_reg_1439;
assign and_ln781_fu_907_p2 = carry_1_reg_1432 & Range1_all_ones_reg_1444;
assign and_ln785_1_fu_510_p2 = xor_ln785_reg_1157 & and_ln786_reg_1169;
assign and_ln785_fu_551_p2 = or_ln785_2_fu_546_p2 & and_ln786_reg_1169;
assign and_ln786_fu_365_p2 = xor_ln786_1_fu_360_p2 & p_Result_11_reg_1110;
assign and_ln788_1_fu_902_p2 = p_Result_16_reg_1404 & and_ln788_fu_896_p2;
assign and_ln788_fu_896_p2 = p_Val2_6_reg_1398[0] & deleted_ones_fu_865_p3;
assign carry_1_fu_789_p2 = xor_ln416_fu_784_p2 & add_ln1192_2_reg_1327[2];
assign op_12_V_fu_629_p2 = op_0[0] & and_ln213_fu_624_p2;
assign overflow_1_fu_887_p2 = xor_ln785_2_fu_882_p2 & or_ln785_1_fu_877_p2;
assign overflow_fu_392_p2 = xor_ln785_reg_1157 & or_ln785_reg_1151;
assign sel_tmp11_fu_520_p2 = xor_ln365_1_fu_466_p2 & or_ln785_3_fu_514_p2;
assign underflow_1_fu_922_p2 = xor_ln788_fu_916_p2 & p_Result_14_reg_1392;
assign xor_ln340_fu_488_p2 = ~ or_ln340_reg_1190;
assign xor_ln780_fu_854_p2 = ~ add_ln1192_1_reg_1387[3];
assign xor_ln785_3_fu_541_p2 = ~ or_ln785_reg_1151;
assign xor_ln786_1_fu_360_p2 = ~ icmp_ln786_reg_1135;
assign xor_ln416_fu_784_p2 = ~ p_Result_16_reg_1404;
assign xor_ln788_fu_916_p2 = ~ or_ln788_fu_911_p2;
assign xor_ln785_1_fu_871_p2 = ~ deleted_zeros_fu_842_p3;
assign xor_ln786_fu_350_p2 = ~ p_Result_11_reg_1110;
assign xor_ln785_2_fu_882_p2 = ~ p_Result_14_reg_1392;
assign xor_ln365_1_fu_466_p2 = ~ xor_ln365_fu_460_p2;
assign xor_ln785_fu_345_p2 = ~ p_Result_10_reg_1098;
assign p_Val2_2_fu_472_p2 = ~ { trunc_ln731_reg_1105[0], 2'h0 };
assign _073_ = ~ tmp_4_reg_1043;
assign _074_ = ~ sel_tmp11_reg_1235;
assign _075_ = ~ p_Result_13_reg_1141;
assign _076_ = ~ ap_start;
assign _077_ = p_Result_3_reg_1416 == 4'hf;
assign _078_ = ! p_Result_3_reg_1416;
assign _079_ = p_Result_2_reg_1411 == 3'h7;
always @(posedge \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.clk )
\add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.bin_s1  <= _081_;
always @(posedge \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.clk )
\add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.ain_s1  <= _080_;
always @(posedge \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.clk )
\add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.sum_s1  <= _083_;
always @(posedge \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.clk )
\add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.carry_s1  <= _082_;
assign _081_ = \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.ce  ? \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.b [16:8] : \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.bin_s1 ;
assign _080_ = \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.ce  ? \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.a [16:8] : \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.ain_s1 ;
assign _082_ = \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.ce  ? \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.facout_s1  : \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.carry_s1 ;
assign _083_ = \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.ce  ? \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.fas_s1  : \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.sum_s1 ;
assign _084_ = \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.u1.a  + \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.u1.b ;
assign { \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.u1.cout , \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.u1.s  } = _084_ + \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.u1.cin ;
assign _085_ = \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.u2.a  + \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.u2.b ;
assign { \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.u2.cout , \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.u2.s  } = _085_ + \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.u2.cin ;
always @(posedge \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.clk )
\add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.bin_s1  <= _087_;
always @(posedge \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.clk )
\add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.ain_s1  <= _086_;
always @(posedge \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.clk )
\add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.sum_s1  <= _089_;
always @(posedge \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.clk )
\add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.carry_s1  <= _088_;
assign _087_ = \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.ce  ? \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.b [16:8] : \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.bin_s1 ;
assign _086_ = \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.ce  ? \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.a [16:8] : \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.ain_s1 ;
assign _088_ = \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.ce  ? \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.facout_s1  : \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.carry_s1 ;
assign _089_ = \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.ce  ? \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.fas_s1  : \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.sum_s1 ;
assign _090_ = \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.u1.a  + \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.u1.b ;
assign { \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.u1.cout , \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.u1.s  } = _090_ + \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.u1.cin ;
assign _091_ = \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.u2.a  + \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.u2.b ;
assign { \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.u2.cout , \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.u2.s  } = _091_ + \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.u2.cin ;
always @(posedge \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.clk )
\add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.bin_s1  <= _093_;
always @(posedge \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.clk )
\add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.ain_s1  <= _092_;
always @(posedge \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.clk )
\add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.sum_s1  <= _095_;
always @(posedge \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.clk )
\add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.carry_s1  <= _094_;
assign _093_ = \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.ce  ? \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.b [16:8] : \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.bin_s1 ;
assign _092_ = \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.ce  ? \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.a [16:8] : \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.ain_s1 ;
assign _094_ = \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.ce  ? \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.facout_s1  : \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.carry_s1 ;
assign _095_ = \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.ce  ? \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.fas_s1  : \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.sum_s1 ;
assign _096_ = \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.u1.a  + \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.u1.b ;
assign { \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.u1.cout , \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.u1.s  } = _096_ + \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.u1.cin ;
assign _097_ = \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.u2.a  + \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.u2.b ;
assign { \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.u2.cout , \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.u2.s  } = _097_ + \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.u2.cin ;
always @(posedge \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.clk )
\add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.bin_s1  <= _099_;
always @(posedge \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.clk )
\add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.ain_s1  <= _098_;
always @(posedge \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.clk )
\add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.sum_s1  <= _101_;
always @(posedge \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.clk )
\add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.carry_s1  <= _100_;
assign _099_ = \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.ce  ? \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.b [1] : \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.bin_s1 ;
assign _098_ = \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.ce  ? \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.a [1] : \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.ain_s1 ;
assign _100_ = \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.ce  ? \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.facout_s1  : \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.carry_s1 ;
assign _101_ = \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.ce  ? \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.fas_s1  : \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.sum_s1 ;
assign _102_ = \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.u1.a  + \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.u1.b ;
assign { \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.u1.cout , \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.u1.s  } = _102_ + \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.u1.cin ;
assign _103_ = \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.u2.a  + \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.u2.b ;
assign { \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.u2.cout , \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.u2.s  } = _103_ + \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.u2.cin ;
always @(posedge \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.clk )
\add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.bin_s1  <= _105_;
always @(posedge \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.clk )
\add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.ain_s1  <= _104_;
always @(posedge \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.clk )
\add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.sum_s1  <= _107_;
always @(posedge \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.clk )
\add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.carry_s1  <= _106_;
assign _105_ = \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.ce  ? \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.b [31:16] : \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.bin_s1 ;
assign _104_ = \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.ce  ? \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.a [31:16] : \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.ain_s1 ;
assign _106_ = \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.ce  ? \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.facout_s1  : \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.carry_s1 ;
assign _107_ = \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.ce  ? \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.fas_s1  : \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.sum_s1 ;
assign _108_ = \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.u1.a  + \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.u1.b ;
assign { \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.u1.cout , \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.u1.s  } = _108_ + \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.u1.cin ;
assign _109_ = \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.u2.a  + \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.u2.b ;
assign { \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.u2.cout , \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.u2.s  } = _109_ + \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.u2.cin ;
always @(posedge \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.clk )
\add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.bin_s1  <= _111_;
always @(posedge \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.clk )
\add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.ain_s1  <= _110_;
always @(posedge \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.clk )
\add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.sum_s1  <= _113_;
always @(posedge \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.clk )
\add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.carry_s1  <= _112_;
assign _111_ = \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.ce  ? \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.b [31:16] : \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.bin_s1 ;
assign _110_ = \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.ce  ? \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.a [31:16] : \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.ain_s1 ;
assign _112_ = \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.ce  ? \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.facout_s1  : \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.carry_s1 ;
assign _113_ = \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.ce  ? \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.fas_s1  : \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.sum_s1 ;
assign _114_ = \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.u1.a  + \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.u1.b ;
assign { \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.u1.cout , \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.u1.s  } = _114_ + \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.u1.cin ;
assign _115_ = \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.u2.a  + \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.u2.b ;
assign { \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.u2.cout , \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.u2.s  } = _115_ + \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.u2.cin ;
always @(posedge \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.clk )
\add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.bin_s1  <= _117_;
always @(posedge \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.clk )
\add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.ain_s1  <= _116_;
always @(posedge \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.clk )
\add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.sum_s1  <= _119_;
always @(posedge \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.clk )
\add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.carry_s1  <= _118_;
assign _117_ = \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.ce  ? \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.b [31:16] : \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.bin_s1 ;
assign _116_ = \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.ce  ? \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.a [31:16] : \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.ain_s1 ;
assign _118_ = \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.ce  ? \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.facout_s1  : \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.carry_s1 ;
assign _119_ = \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.ce  ? \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.fas_s1  : \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.sum_s1 ;
assign _120_ = \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.u1.a  + \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.u1.b ;
assign { \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.u1.cout , \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.u1.s  } = _120_ + \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.u1.cin ;
assign _121_ = \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.u2.a  + \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.u2.b ;
assign { \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.u2.cout , \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.u2.s  } = _121_ + \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.u2.cin ;
always @(posedge \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.clk )
\add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.bin_s1  <= _123_;
always @(posedge \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.clk )
\add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.ain_s1  <= _122_;
always @(posedge \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.clk )
\add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.sum_s1  <= _125_;
always @(posedge \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.clk )
\add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.carry_s1  <= _124_;
assign _123_ = \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.ce  ? \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.b [31:16] : \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.bin_s1 ;
assign _122_ = \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.ce  ? \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.a [31:16] : \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.ain_s1 ;
assign _124_ = \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.ce  ? \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.facout_s1  : \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.carry_s1 ;
assign _125_ = \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.ce  ? \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.fas_s1  : \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.sum_s1 ;
assign _126_ = \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.u1.a  + \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.u1.b ;
assign { \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.u1.cout , \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.u1.s  } = _126_ + \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.u1.cin ;
assign _127_ = \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.u2.a  + \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.u2.b ;
assign { \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.u2.cout , \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.u2.s  } = _127_ + \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.u2.cin ;
always @(posedge \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.clk )
\add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.bin_s1  <= _129_;
always @(posedge \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.clk )
\add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.ain_s1  <= _128_;
always @(posedge \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.clk )
\add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.sum_s1  <= _131_;
always @(posedge \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.clk )
\add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.carry_s1  <= _130_;
assign _129_ = \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.ce  ? \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.b [33:17] : \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.bin_s1 ;
assign _128_ = \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.ce  ? \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.a [33:17] : \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.ain_s1 ;
assign _130_ = \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.ce  ? \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.facout_s1  : \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.carry_s1 ;
assign _131_ = \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.ce  ? \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.fas_s1  : \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.sum_s1 ;
assign _132_ = \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.u1.a  + \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.u1.b ;
assign { \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.u1.cout , \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.u1.s  } = _132_ + \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.u1.cin ;
assign _133_ = \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.u2.a  + \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.u2.b ;
assign { \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.u2.cout , \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.u2.s  } = _133_ + \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.u2.cin ;
always @(posedge \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.clk )
\add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.bin_s1  <= _135_;
always @(posedge \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.clk )
\add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.ain_s1  <= _134_;
always @(posedge \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.clk )
\add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.sum_s1  <= _137_;
always @(posedge \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.clk )
\add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.carry_s1  <= _136_;
assign _135_ = \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.ce  ? \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.b [2:1] : \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.bin_s1 ;
assign _134_ = \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.ce  ? \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.a [2:1] : \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.ain_s1 ;
assign _136_ = \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.ce  ? \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.facout_s1  : \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.carry_s1 ;
assign _137_ = \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.ce  ? \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.fas_s1  : \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.sum_s1 ;
assign _138_ = \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.u1.a  + \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.u1.b ;
assign { \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.u1.cout , \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.u1.s  } = _138_ + \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.u1.cin ;
assign _139_ = \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.u2.a  + \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.u2.b ;
assign { \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.u2.cout , \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.u2.s  } = _139_ + \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.u2.cin ;
always @(posedge \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.clk )
\add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.bin_s1  <= _141_;
always @(posedge \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.clk )
\add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.ain_s1  <= _140_;
always @(posedge \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.clk )
\add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.sum_s1  <= _143_;
always @(posedge \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.clk )
\add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.carry_s1  <= _142_;
assign _141_ = \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.ce  ? \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.b [2:1] : \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.bin_s1 ;
assign _140_ = \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.ce  ? \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.a [2:1] : \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.ain_s1 ;
assign _142_ = \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.ce  ? \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.facout_s1  : \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.carry_s1 ;
assign _143_ = \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.ce  ? \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.fas_s1  : \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.sum_s1 ;
assign _144_ = \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.u1.a  + \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.u1.b ;
assign { \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.u1.cout , \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.u1.s  } = _144_ + \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.u1.cin ;
assign _145_ = \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.u2.a  + \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.u2.b ;
assign { \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.u2.cout , \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.u2.s  } = _145_ + \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.u2.cin ;
always @(posedge \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.clk )
\add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.bin_s1  <= _147_;
always @(posedge \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.clk )
\add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.ain_s1  <= _146_;
always @(posedge \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.clk )
\add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.sum_s1  <= _149_;
always @(posedge \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.clk )
\add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.carry_s1  <= _148_;
assign _147_ = \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.ce  ? \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.b [3:2] : \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.bin_s1 ;
assign _146_ = \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.ce  ? \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.a [3:2] : \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.ain_s1 ;
assign _148_ = \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.ce  ? \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.facout_s1  : \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.carry_s1 ;
assign _149_ = \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.ce  ? \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.fas_s1  : \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.sum_s1 ;
assign _150_ = \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.u1.a  + \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.u1.b ;
assign { \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.u1.cout , \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.u1.s  } = _150_ + \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.u1.cin ;
assign _151_ = \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.u2.a  + \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.u2.b ;
assign { \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.u2.cout , \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.u2.s  } = _151_ + \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.u2.cin ;
always @(posedge \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.clk )
\add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.bin_s1  <= _153_;
always @(posedge \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.clk )
\add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.ain_s1  <= _152_;
always @(posedge \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.clk )
\add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.sum_s1  <= _155_;
always @(posedge \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.clk )
\add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.carry_s1  <= _154_;
assign _153_ = \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.ce  ? \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.b [3:2] : \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.bin_s1 ;
assign _152_ = \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.ce  ? \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.a [3:2] : \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.ain_s1 ;
assign _154_ = \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.ce  ? \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.facout_s1  : \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.carry_s1 ;
assign _155_ = \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.ce  ? \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.fas_s1  : \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.sum_s1 ;
assign _156_ = \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.u1.a  + \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.u1.b ;
assign { \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.u1.cout , \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.u1.s  } = _156_ + \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.u1.cin ;
assign _157_ = \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.u2.a  + \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.u2.b ;
assign { \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.u2.cout , \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.u2.s  } = _157_ + \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.u2.cin ;
always @(posedge \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.clk )
\add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.bin_s1  <= _159_;
always @(posedge \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.clk )
\add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.ain_s1  <= _158_;
always @(posedge \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.clk )
\add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.sum_s1  <= _161_;
always @(posedge \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.clk )
\add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.carry_s1  <= _160_;
assign _159_ = \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.ce  ? \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.b [5:3] : \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.bin_s1 ;
assign _158_ = \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.ce  ? \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.a [5:3] : \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.ain_s1 ;
assign _160_ = \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.ce  ? \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.facout_s1  : \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.carry_s1 ;
assign _161_ = \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.ce  ? \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.fas_s1  : \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.sum_s1 ;
assign _162_ = \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.u1.a  + \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.u1.b ;
assign { \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.u1.cout , \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.u1.s  } = _162_ + \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.u1.cin ;
assign _163_ = \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.u2.a  + \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.u2.b ;
assign { \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.u2.cout , \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.u2.s  } = _163_ + \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.u2.cin ;
always @(posedge \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.clk )
\add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.bin_s1  <= _165_;
always @(posedge \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.clk )
\add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.ain_s1  <= _164_;
always @(posedge \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.clk )
\add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.sum_s1  <= _167_;
always @(posedge \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.clk )
\add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.carry_s1  <= _166_;
assign _165_ = \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.ce  ? \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.b [6:3] : \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.bin_s1 ;
assign _164_ = \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.ce  ? \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.a [6:3] : \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.ain_s1 ;
assign _166_ = \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.ce  ? \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.facout_s1  : \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.carry_s1 ;
assign _167_ = \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.ce  ? \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.fas_s1  : \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.sum_s1 ;
assign _168_ = \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.u1.a  + \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.u1.b ;
assign { \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.u1.cout , \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.u1.s  } = _168_ + \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.u1.cin ;
assign _169_ = \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.u2.a  + \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.u2.b ;
assign { \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.u2.cout , \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.u2.s  } = _169_ + \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.u2.cin ;
always @(posedge \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.clk )
\add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.bin_s1  <= _171_;
always @(posedge \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.clk )
\add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.ain_s1  <= _170_;
always @(posedge \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.clk )
\add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.sum_s1  <= _173_;
always @(posedge \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.clk )
\add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.carry_s1  <= _172_;
assign _171_ = \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.ce  ? \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.b [6:3] : \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.bin_s1 ;
assign _170_ = \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.ce  ? \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.a [6:3] : \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.ain_s1 ;
assign _172_ = \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.ce  ? \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.facout_s1  : \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.carry_s1 ;
assign _173_ = \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.ce  ? \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.fas_s1  : \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.sum_s1 ;
assign _174_ = \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.u1.a  + \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.u1.b ;
assign { \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.u1.cout , \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.u1.s  } = _174_ + \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.u1.cin ;
assign _175_ = \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.u2.a  + \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.u2.b ;
assign { \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.u2.cout , \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.u2.s  } = _175_ + \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.u2.cin ;
always @(posedge \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.clk )
\add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.bin_s1  <= _177_;
always @(posedge \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.clk )
\add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.ain_s1  <= _176_;
always @(posedge \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.clk )
\add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.sum_s1  <= _179_;
always @(posedge \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.clk )
\add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.carry_s1  <= _178_;
assign _177_ = \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.ce  ? \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.b [6:3] : \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.bin_s1 ;
assign _176_ = \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.ce  ? \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.a [6:3] : \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.ain_s1 ;
assign _178_ = \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.ce  ? \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.facout_s1  : \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.carry_s1 ;
assign _179_ = \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.ce  ? \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.fas_s1  : \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.sum_s1 ;
assign _180_ = \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.u1.a  + \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.u1.b ;
assign { \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.u1.cout , \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.u1.s  } = _180_ + \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.u1.cin ;
assign _181_ = \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.u2.a  + \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.u2.b ;
assign { \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.u2.cout , \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.u2.s  } = _181_ + \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.u2.cin ;
always @(posedge \ashr_16s_16ns_16_7_1_U3.clk )
\ashr_16s_16ns_16_7_1_U3.dout_array[5]  <= _193_;
always @(posedge \ashr_16s_16ns_16_7_1_U3.clk )
\ashr_16s_16ns_16_7_1_U3.din1_cast_array[5]  <= _187_;
always @(posedge \ashr_16s_16ns_16_7_1_U3.clk )
\ashr_16s_16ns_16_7_1_U3.dout_array[4]  <= _192_;
always @(posedge \ashr_16s_16ns_16_7_1_U3.clk )
\ashr_16s_16ns_16_7_1_U3.din1_cast_array[4]  <= _186_;
always @(posedge \ashr_16s_16ns_16_7_1_U3.clk )
\ashr_16s_16ns_16_7_1_U3.dout_array[3]  <= _191_;
always @(posedge \ashr_16s_16ns_16_7_1_U3.clk )
\ashr_16s_16ns_16_7_1_U3.din1_cast_array[3]  <= _185_;
always @(posedge \ashr_16s_16ns_16_7_1_U3.clk )
\ashr_16s_16ns_16_7_1_U3.dout_array[2]  <= _190_;
always @(posedge \ashr_16s_16ns_16_7_1_U3.clk )
\ashr_16s_16ns_16_7_1_U3.din1_cast_array[2]  <= _184_;
always @(posedge \ashr_16s_16ns_16_7_1_U3.clk )
\ashr_16s_16ns_16_7_1_U3.dout_array[1]  <= _189_;
always @(posedge \ashr_16s_16ns_16_7_1_U3.clk )
\ashr_16s_16ns_16_7_1_U3.din1_cast_array[1]  <= _183_;
always @(posedge \ashr_16s_16ns_16_7_1_U3.clk )
\ashr_16s_16ns_16_7_1_U3.dout_array[0]  <= _188_;
always @(posedge \ashr_16s_16ns_16_7_1_U3.clk )
\ashr_16s_16ns_16_7_1_U3.din1_cast_array[0]  <= _182_;
assign _194_ = \ashr_16s_16ns_16_7_1_U3.ce  ? \ashr_16s_16ns_16_7_1_U3.din1_cast_array[4]  : \ashr_16s_16ns_16_7_1_U3.din1_cast_array[5] ;
assign _187_ = \ashr_16s_16ns_16_7_1_U3.reset  ? 16'h0000 : _194_;
assign _195_ = \ashr_16s_16ns_16_7_1_U3.ce  ? _210_ : \ashr_16s_16ns_16_7_1_U3.dout_array[5] ;
assign _193_ = \ashr_16s_16ns_16_7_1_U3.reset  ? 16'h0000 : _195_;
assign _196_ = \ashr_16s_16ns_16_7_1_U3.ce  ? \ashr_16s_16ns_16_7_1_U3.din1_cast_array[3]  : \ashr_16s_16ns_16_7_1_U3.din1_cast_array[4] ;
assign _186_ = \ashr_16s_16ns_16_7_1_U3.reset  ? 16'h0000 : _196_;
assign _197_ = \ashr_16s_16ns_16_7_1_U3.ce  ? _209_ : \ashr_16s_16ns_16_7_1_U3.dout_array[4] ;
assign _192_ = \ashr_16s_16ns_16_7_1_U3.reset  ? 16'h0000 : _197_;
assign _198_ = \ashr_16s_16ns_16_7_1_U3.ce  ? \ashr_16s_16ns_16_7_1_U3.din1_cast_array[2]  : \ashr_16s_16ns_16_7_1_U3.din1_cast_array[3] ;
assign _185_ = \ashr_16s_16ns_16_7_1_U3.reset  ? 16'h0000 : _198_;
assign _199_ = \ashr_16s_16ns_16_7_1_U3.ce  ? _208_ : \ashr_16s_16ns_16_7_1_U3.dout_array[3] ;
assign _191_ = \ashr_16s_16ns_16_7_1_U3.reset  ? 16'h0000 : _199_;
assign _200_ = \ashr_16s_16ns_16_7_1_U3.ce  ? \ashr_16s_16ns_16_7_1_U3.din1_cast_array[1]  : \ashr_16s_16ns_16_7_1_U3.din1_cast_array[2] ;
assign _184_ = \ashr_16s_16ns_16_7_1_U3.reset  ? 16'h0000 : _200_;
assign _201_ = \ashr_16s_16ns_16_7_1_U3.ce  ? _207_ : \ashr_16s_16ns_16_7_1_U3.dout_array[2] ;
assign _190_ = \ashr_16s_16ns_16_7_1_U3.reset  ? 16'h0000 : _201_;
assign _202_ = \ashr_16s_16ns_16_7_1_U3.ce  ? \ashr_16s_16ns_16_7_1_U3.din1_cast_array[0]  : \ashr_16s_16ns_16_7_1_U3.din1_cast_array[1] ;
assign _183_ = \ashr_16s_16ns_16_7_1_U3.reset  ? 16'h0000 : _202_;
assign _203_ = \ashr_16s_16ns_16_7_1_U3.ce  ? _206_ : \ashr_16s_16ns_16_7_1_U3.dout_array[1] ;
assign _189_ = \ashr_16s_16ns_16_7_1_U3.reset  ? 16'h0000 : _203_;
assign _204_ = \ashr_16s_16ns_16_7_1_U3.ce  ? \ashr_16s_16ns_16_7_1_U3.din1  : \ashr_16s_16ns_16_7_1_U3.din1_cast_array[0] ;
assign _182_ = \ashr_16s_16ns_16_7_1_U3.reset  ? 16'h0000 : _204_;
assign _205_ = \ashr_16s_16ns_16_7_1_U3.ce  ? \ashr_16s_16ns_16_7_1_U3.din0  : \ashr_16s_16ns_16_7_1_U3.dout_array[0] ;
assign _188_ = \ashr_16s_16ns_16_7_1_U3.reset  ? 16'h0000 : _205_;
assign _206_ = $signed(\ashr_16s_16ns_16_7_1_U3.dout_array[0] ) >>> { \ashr_16s_16ns_16_7_1_U3.din1_cast_array[0] [15], 15'h0000 };
assign _207_ = $signed(\ashr_16s_16ns_16_7_1_U3.dout_array[1] ) >>> { \ashr_16s_16ns_16_7_1_U3.din1_cast_array[1] [14:12], 12'h000 };
assign _208_ = $signed(\ashr_16s_16ns_16_7_1_U3.dout_array[2] ) >>> { \ashr_16s_16ns_16_7_1_U3.din1_cast_array[2] [11:9], 9'h000 };
assign _209_ = $signed(\ashr_16s_16ns_16_7_1_U3.dout_array[3] ) >>> { \ashr_16s_16ns_16_7_1_U3.din1_cast_array[3] [8:6], 6'h00 };
assign _210_ = $signed(\ashr_16s_16ns_16_7_1_U3.dout_array[4] ) >>> { \ashr_16s_16ns_16_7_1_U3.din1_cast_array[4] [5:3], 3'h0 };
assign \ashr_16s_16ns_16_7_1_U3.dout  = $signed(\ashr_16s_16ns_16_7_1_U3.dout_array[5] ) >>> \ashr_16s_16ns_16_7_1_U3.din1_cast_array[5] [2:0];
always @(posedge \ashr_32s_8ns_32_7_1_U7.clk )
\ashr_32s_8ns_32_7_1_U7.dout_array[5]  <= _222_;
always @(posedge \ashr_32s_8ns_32_7_1_U7.clk )
\ashr_32s_8ns_32_7_1_U7.din1_cast_array[5]  <= _216_;
always @(posedge \ashr_32s_8ns_32_7_1_U7.clk )
\ashr_32s_8ns_32_7_1_U7.dout_array[4]  <= _221_;
always @(posedge \ashr_32s_8ns_32_7_1_U7.clk )
\ashr_32s_8ns_32_7_1_U7.din1_cast_array[4]  <= _215_;
always @(posedge \ashr_32s_8ns_32_7_1_U7.clk )
\ashr_32s_8ns_32_7_1_U7.dout_array[3]  <= _220_;
always @(posedge \ashr_32s_8ns_32_7_1_U7.clk )
\ashr_32s_8ns_32_7_1_U7.din1_cast_array[3]  <= _214_;
always @(posedge \ashr_32s_8ns_32_7_1_U7.clk )
\ashr_32s_8ns_32_7_1_U7.dout_array[2]  <= _219_;
always @(posedge \ashr_32s_8ns_32_7_1_U7.clk )
\ashr_32s_8ns_32_7_1_U7.din1_cast_array[2]  <= _213_;
always @(posedge \ashr_32s_8ns_32_7_1_U7.clk )
\ashr_32s_8ns_32_7_1_U7.dout_array[1]  <= _218_;
always @(posedge \ashr_32s_8ns_32_7_1_U7.clk )
\ashr_32s_8ns_32_7_1_U7.din1_cast_array[1]  <= _212_;
always @(posedge \ashr_32s_8ns_32_7_1_U7.clk )
\ashr_32s_8ns_32_7_1_U7.dout_array[0]  <= _217_;
always @(posedge \ashr_32s_8ns_32_7_1_U7.clk )
\ashr_32s_8ns_32_7_1_U7.din1_cast_array[0]  <= _211_;
assign _223_ = \ashr_32s_8ns_32_7_1_U7.ce  ? \ashr_32s_8ns_32_7_1_U7.din1_cast_array[4]  : \ashr_32s_8ns_32_7_1_U7.din1_cast_array[5] ;
assign _216_ = \ashr_32s_8ns_32_7_1_U7.reset  ? 8'h00 : _223_;
assign _224_ = \ashr_32s_8ns_32_7_1_U7.ce  ? _237_ : \ashr_32s_8ns_32_7_1_U7.dout_array[5] ;
assign _222_ = \ashr_32s_8ns_32_7_1_U7.reset  ? 32'd0 : _224_;
assign _225_ = \ashr_32s_8ns_32_7_1_U7.ce  ? \ashr_32s_8ns_32_7_1_U7.din1_cast_array[3]  : \ashr_32s_8ns_32_7_1_U7.din1_cast_array[4] ;
assign _215_ = \ashr_32s_8ns_32_7_1_U7.reset  ? 8'h00 : _225_;
assign _226_ = \ashr_32s_8ns_32_7_1_U7.ce  ? _236_ : \ashr_32s_8ns_32_7_1_U7.dout_array[4] ;
assign _221_ = \ashr_32s_8ns_32_7_1_U7.reset  ? 32'd0 : _226_;
assign _227_ = \ashr_32s_8ns_32_7_1_U7.ce  ? \ashr_32s_8ns_32_7_1_U7.din1_cast_array[2]  : \ashr_32s_8ns_32_7_1_U7.din1_cast_array[3] ;
assign _214_ = \ashr_32s_8ns_32_7_1_U7.reset  ? 8'h00 : _227_;
assign _228_ = \ashr_32s_8ns_32_7_1_U7.ce  ? _235_ : \ashr_32s_8ns_32_7_1_U7.dout_array[3] ;
assign _220_ = \ashr_32s_8ns_32_7_1_U7.reset  ? 32'd0 : _228_;
assign _229_ = \ashr_32s_8ns_32_7_1_U7.ce  ? \ashr_32s_8ns_32_7_1_U7.din1_cast_array[1]  : \ashr_32s_8ns_32_7_1_U7.din1_cast_array[2] ;
assign _213_ = \ashr_32s_8ns_32_7_1_U7.reset  ? 8'h00 : _229_;
assign _230_ = \ashr_32s_8ns_32_7_1_U7.ce  ? \ashr_32s_8ns_32_7_1_U7.dout_array[1]  : \ashr_32s_8ns_32_7_1_U7.dout_array[2] ;
assign _219_ = \ashr_32s_8ns_32_7_1_U7.reset  ? 32'd0 : _230_;
assign _231_ = \ashr_32s_8ns_32_7_1_U7.ce  ? \ashr_32s_8ns_32_7_1_U7.din1_cast_array[0]  : \ashr_32s_8ns_32_7_1_U7.din1_cast_array[1] ;
assign _212_ = \ashr_32s_8ns_32_7_1_U7.reset  ? 8'h00 : _231_;
assign _232_ = \ashr_32s_8ns_32_7_1_U7.ce  ? \ashr_32s_8ns_32_7_1_U7.dout_array[0]  : \ashr_32s_8ns_32_7_1_U7.dout_array[1] ;
assign _218_ = \ashr_32s_8ns_32_7_1_U7.reset  ? 32'd0 : _232_;
assign _233_ = \ashr_32s_8ns_32_7_1_U7.ce  ? \ashr_32s_8ns_32_7_1_U7.din1 [7:0] : \ashr_32s_8ns_32_7_1_U7.din1_cast_array[0] ;
assign _211_ = \ashr_32s_8ns_32_7_1_U7.reset  ? 8'h00 : _233_;
assign _234_ = \ashr_32s_8ns_32_7_1_U7.ce  ? \ashr_32s_8ns_32_7_1_U7.din0  : \ashr_32s_8ns_32_7_1_U7.dout_array[0] ;
assign _217_ = \ashr_32s_8ns_32_7_1_U7.reset  ? 32'd0 : _234_;
assign _235_ = $signed(\ashr_32s_8ns_32_7_1_U7.dout_array[2] ) >>> { \ashr_32s_8ns_32_7_1_U7.din1_cast_array[2] [7:6], 6'h00 };
assign _236_ = $signed(\ashr_32s_8ns_32_7_1_U7.dout_array[3] ) >>> { \ashr_32s_8ns_32_7_1_U7.din1_cast_array[3] [5:4], 4'h0 };
assign _237_ = $signed(\ashr_32s_8ns_32_7_1_U7.dout_array[4] ) >>> { \ashr_32s_8ns_32_7_1_U7.din1_cast_array[4] [3:2], 2'h0 };
assign \ashr_32s_8ns_32_7_1_U7.dout  = $signed(\ashr_32s_8ns_32_7_1_U7.dout_array[5] ) >>> \ashr_32s_8ns_32_7_1_U7.din1_cast_array[5] [1:0];
always @(posedge \shl_16s_16ns_16_7_1_U4.clk )
\shl_16s_16ns_16_7_1_U4.dout_array[5]  <= _249_;
always @(posedge \shl_16s_16ns_16_7_1_U4.clk )
\shl_16s_16ns_16_7_1_U4.din1_cast_array[5]  <= _243_;
always @(posedge \shl_16s_16ns_16_7_1_U4.clk )
\shl_16s_16ns_16_7_1_U4.dout_array[4]  <= _248_;
always @(posedge \shl_16s_16ns_16_7_1_U4.clk )
\shl_16s_16ns_16_7_1_U4.din1_cast_array[4]  <= _242_;
always @(posedge \shl_16s_16ns_16_7_1_U4.clk )
\shl_16s_16ns_16_7_1_U4.dout_array[3]  <= _247_;
always @(posedge \shl_16s_16ns_16_7_1_U4.clk )
\shl_16s_16ns_16_7_1_U4.din1_cast_array[3]  <= _241_;
always @(posedge \shl_16s_16ns_16_7_1_U4.clk )
\shl_16s_16ns_16_7_1_U4.dout_array[2]  <= _246_;
always @(posedge \shl_16s_16ns_16_7_1_U4.clk )
\shl_16s_16ns_16_7_1_U4.din1_cast_array[2]  <= _240_;
always @(posedge \shl_16s_16ns_16_7_1_U4.clk )
\shl_16s_16ns_16_7_1_U4.dout_array[1]  <= _245_;
always @(posedge \shl_16s_16ns_16_7_1_U4.clk )
\shl_16s_16ns_16_7_1_U4.din1_cast_array[1]  <= _239_;
always @(posedge \shl_16s_16ns_16_7_1_U4.clk )
\shl_16s_16ns_16_7_1_U4.dout_array[0]  <= _244_;
always @(posedge \shl_16s_16ns_16_7_1_U4.clk )
\shl_16s_16ns_16_7_1_U4.din1_cast_array[0]  <= _238_;
assign _250_ = \shl_16s_16ns_16_7_1_U4.ce  ? \shl_16s_16ns_16_7_1_U4.din1_cast_array[4]  : \shl_16s_16ns_16_7_1_U4.din1_cast_array[5] ;
assign _243_ = \shl_16s_16ns_16_7_1_U4.reset  ? 16'h0000 : _250_;
assign _251_ = \shl_16s_16ns_16_7_1_U4.ce  ? _266_ : \shl_16s_16ns_16_7_1_U4.dout_array[5] ;
assign _249_ = \shl_16s_16ns_16_7_1_U4.reset  ? 16'h0000 : _251_;
assign _252_ = \shl_16s_16ns_16_7_1_U4.ce  ? \shl_16s_16ns_16_7_1_U4.din1_cast_array[3]  : \shl_16s_16ns_16_7_1_U4.din1_cast_array[4] ;
assign _242_ = \shl_16s_16ns_16_7_1_U4.reset  ? 16'h0000 : _252_;
assign _253_ = \shl_16s_16ns_16_7_1_U4.ce  ? _265_ : \shl_16s_16ns_16_7_1_U4.dout_array[4] ;
assign _248_ = \shl_16s_16ns_16_7_1_U4.reset  ? 16'h0000 : _253_;
assign _254_ = \shl_16s_16ns_16_7_1_U4.ce  ? \shl_16s_16ns_16_7_1_U4.din1_cast_array[2]  : \shl_16s_16ns_16_7_1_U4.din1_cast_array[3] ;
assign _241_ = \shl_16s_16ns_16_7_1_U4.reset  ? 16'h0000 : _254_;
assign _255_ = \shl_16s_16ns_16_7_1_U4.ce  ? _264_ : \shl_16s_16ns_16_7_1_U4.dout_array[3] ;
assign _247_ = \shl_16s_16ns_16_7_1_U4.reset  ? 16'h0000 : _255_;
assign _256_ = \shl_16s_16ns_16_7_1_U4.ce  ? \shl_16s_16ns_16_7_1_U4.din1_cast_array[1]  : \shl_16s_16ns_16_7_1_U4.din1_cast_array[2] ;
assign _240_ = \shl_16s_16ns_16_7_1_U4.reset  ? 16'h0000 : _256_;
assign _257_ = \shl_16s_16ns_16_7_1_U4.ce  ? _263_ : \shl_16s_16ns_16_7_1_U4.dout_array[2] ;
assign _246_ = \shl_16s_16ns_16_7_1_U4.reset  ? 16'h0000 : _257_;
assign _258_ = \shl_16s_16ns_16_7_1_U4.ce  ? \shl_16s_16ns_16_7_1_U4.din1_cast_array[0]  : \shl_16s_16ns_16_7_1_U4.din1_cast_array[1] ;
assign _239_ = \shl_16s_16ns_16_7_1_U4.reset  ? 16'h0000 : _258_;
assign _259_ = \shl_16s_16ns_16_7_1_U4.ce  ? _262_ : \shl_16s_16ns_16_7_1_U4.dout_array[1] ;
assign _245_ = \shl_16s_16ns_16_7_1_U4.reset  ? 16'h0000 : _259_;
assign _260_ = \shl_16s_16ns_16_7_1_U4.ce  ? \shl_16s_16ns_16_7_1_U4.din1  : \shl_16s_16ns_16_7_1_U4.din1_cast_array[0] ;
assign _238_ = \shl_16s_16ns_16_7_1_U4.reset  ? 16'h0000 : _260_;
assign _261_ = \shl_16s_16ns_16_7_1_U4.ce  ? \shl_16s_16ns_16_7_1_U4.din0  : \shl_16s_16ns_16_7_1_U4.dout_array[0] ;
assign _244_ = \shl_16s_16ns_16_7_1_U4.reset  ? 16'h0000 : _261_;
assign _262_ = \shl_16s_16ns_16_7_1_U4.dout_array[0]  << { \shl_16s_16ns_16_7_1_U4.din1_cast_array[0] [15], 15'h0000 };
assign _263_ = \shl_16s_16ns_16_7_1_U4.dout_array[1]  << { \shl_16s_16ns_16_7_1_U4.din1_cast_array[1] [14:12], 12'h000 };
assign _264_ = \shl_16s_16ns_16_7_1_U4.dout_array[2]  << { \shl_16s_16ns_16_7_1_U4.din1_cast_array[2] [11:9], 9'h000 };
assign _265_ = \shl_16s_16ns_16_7_1_U4.dout_array[3]  << { \shl_16s_16ns_16_7_1_U4.din1_cast_array[3] [8:6], 6'h00 };
assign _266_ = \shl_16s_16ns_16_7_1_U4.dout_array[4]  << { \shl_16s_16ns_16_7_1_U4.din1_cast_array[4] [5:3], 3'h0 };
assign \shl_16s_16ns_16_7_1_U4.dout  = \shl_16s_16ns_16_7_1_U4.dout_array[5]  << \shl_16s_16ns_16_7_1_U4.din1_cast_array[5] [2:0];
always @(posedge \shl_32s_8ns_32_7_1_U8.clk )
\shl_32s_8ns_32_7_1_U8.dout_array[5]  <= _278_;
always @(posedge \shl_32s_8ns_32_7_1_U8.clk )
\shl_32s_8ns_32_7_1_U8.din1_cast_array[5]  <= _272_;
always @(posedge \shl_32s_8ns_32_7_1_U8.clk )
\shl_32s_8ns_32_7_1_U8.dout_array[4]  <= _277_;
always @(posedge \shl_32s_8ns_32_7_1_U8.clk )
\shl_32s_8ns_32_7_1_U8.din1_cast_array[4]  <= _271_;
always @(posedge \shl_32s_8ns_32_7_1_U8.clk )
\shl_32s_8ns_32_7_1_U8.dout_array[3]  <= _276_;
always @(posedge \shl_32s_8ns_32_7_1_U8.clk )
\shl_32s_8ns_32_7_1_U8.din1_cast_array[3]  <= _270_;
always @(posedge \shl_32s_8ns_32_7_1_U8.clk )
\shl_32s_8ns_32_7_1_U8.dout_array[2]  <= _275_;
always @(posedge \shl_32s_8ns_32_7_1_U8.clk )
\shl_32s_8ns_32_7_1_U8.din1_cast_array[2]  <= _269_;
always @(posedge \shl_32s_8ns_32_7_1_U8.clk )
\shl_32s_8ns_32_7_1_U8.dout_array[1]  <= _274_;
always @(posedge \shl_32s_8ns_32_7_1_U8.clk )
\shl_32s_8ns_32_7_1_U8.din1_cast_array[1]  <= _268_;
always @(posedge \shl_32s_8ns_32_7_1_U8.clk )
\shl_32s_8ns_32_7_1_U8.dout_array[0]  <= _273_;
always @(posedge \shl_32s_8ns_32_7_1_U8.clk )
\shl_32s_8ns_32_7_1_U8.din1_cast_array[0]  <= _267_;
assign _279_ = \shl_32s_8ns_32_7_1_U8.ce  ? \shl_32s_8ns_32_7_1_U8.din1_cast_array[4]  : \shl_32s_8ns_32_7_1_U8.din1_cast_array[5] ;
assign _272_ = \shl_32s_8ns_32_7_1_U8.reset  ? 8'h00 : _279_;
assign _280_ = \shl_32s_8ns_32_7_1_U8.ce  ? _293_ : \shl_32s_8ns_32_7_1_U8.dout_array[5] ;
assign _278_ = \shl_32s_8ns_32_7_1_U8.reset  ? 32'd0 : _280_;
assign _281_ = \shl_32s_8ns_32_7_1_U8.ce  ? \shl_32s_8ns_32_7_1_U8.din1_cast_array[3]  : \shl_32s_8ns_32_7_1_U8.din1_cast_array[4] ;
assign _271_ = \shl_32s_8ns_32_7_1_U8.reset  ? 8'h00 : _281_;
assign _282_ = \shl_32s_8ns_32_7_1_U8.ce  ? _292_ : \shl_32s_8ns_32_7_1_U8.dout_array[4] ;
assign _277_ = \shl_32s_8ns_32_7_1_U8.reset  ? 32'd0 : _282_;
assign _283_ = \shl_32s_8ns_32_7_1_U8.ce  ? \shl_32s_8ns_32_7_1_U8.din1_cast_array[2]  : \shl_32s_8ns_32_7_1_U8.din1_cast_array[3] ;
assign _270_ = \shl_32s_8ns_32_7_1_U8.reset  ? 8'h00 : _283_;
assign _284_ = \shl_32s_8ns_32_7_1_U8.ce  ? _291_ : \shl_32s_8ns_32_7_1_U8.dout_array[3] ;
assign _276_ = \shl_32s_8ns_32_7_1_U8.reset  ? 32'd0 : _284_;
assign _285_ = \shl_32s_8ns_32_7_1_U8.ce  ? \shl_32s_8ns_32_7_1_U8.din1_cast_array[1]  : \shl_32s_8ns_32_7_1_U8.din1_cast_array[2] ;
assign _269_ = \shl_32s_8ns_32_7_1_U8.reset  ? 8'h00 : _285_;
assign _286_ = \shl_32s_8ns_32_7_1_U8.ce  ? \shl_32s_8ns_32_7_1_U8.dout_array[1]  : \shl_32s_8ns_32_7_1_U8.dout_array[2] ;
assign _275_ = \shl_32s_8ns_32_7_1_U8.reset  ? 32'd0 : _286_;
assign _287_ = \shl_32s_8ns_32_7_1_U8.ce  ? \shl_32s_8ns_32_7_1_U8.din1_cast_array[0]  : \shl_32s_8ns_32_7_1_U8.din1_cast_array[1] ;
assign _268_ = \shl_32s_8ns_32_7_1_U8.reset  ? 8'h00 : _287_;
assign _288_ = \shl_32s_8ns_32_7_1_U8.ce  ? \shl_32s_8ns_32_7_1_U8.dout_array[0]  : \shl_32s_8ns_32_7_1_U8.dout_array[1] ;
assign _274_ = \shl_32s_8ns_32_7_1_U8.reset  ? 32'd0 : _288_;
assign _289_ = \shl_32s_8ns_32_7_1_U8.ce  ? \shl_32s_8ns_32_7_1_U8.din1 [7:0] : \shl_32s_8ns_32_7_1_U8.din1_cast_array[0] ;
assign _267_ = \shl_32s_8ns_32_7_1_U8.reset  ? 8'h00 : _289_;
assign _290_ = \shl_32s_8ns_32_7_1_U8.ce  ? \shl_32s_8ns_32_7_1_U8.din0  : \shl_32s_8ns_32_7_1_U8.dout_array[0] ;
assign _273_ = \shl_32s_8ns_32_7_1_U8.reset  ? 32'd0 : _290_;
assign _291_ = \shl_32s_8ns_32_7_1_U8.dout_array[2]  << { \shl_32s_8ns_32_7_1_U8.din1_cast_array[2] [7:6], 6'h00 };
assign _292_ = \shl_32s_8ns_32_7_1_U8.dout_array[3]  << { \shl_32s_8ns_32_7_1_U8.din1_cast_array[3] [5:4], 4'h0 };
assign _293_ = \shl_32s_8ns_32_7_1_U8.dout_array[4]  << { \shl_32s_8ns_32_7_1_U8.din1_cast_array[4] [3:2], 2'h0 };
assign \shl_32s_8ns_32_7_1_U8.dout  = \shl_32s_8ns_32_7_1_U8.dout_array[5]  << \shl_32s_8ns_32_7_1_U8.din1_cast_array[5] [1:0];
assign \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.bin_s0  = ~ \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.b ;
always @(posedge \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.clk )
\sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.bin_s1  <= _295_;
always @(posedge \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.clk )
\sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.ain_s1  <= _294_;
always @(posedge \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.clk )
\sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.sum_s1  <= _297_;
always @(posedge \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.clk )
\sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.carry_s1  <= _296_;
assign _295_ = \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.ce  ? \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.bin_s0 [16:8] : \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.bin_s1 ;
assign _294_ = \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.ce  ? \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.a [16:8] : \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.ain_s1 ;
assign _296_ = \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.ce  ? \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.facout_s1  : \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.carry_s1 ;
assign _297_ = \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.ce  ? \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.fas_s1  : \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.sum_s1 ;
assign _298_ = \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.u1.a  + \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.u1.b ;
assign { \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.u1.cout , \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.u1.s  } = _298_ + \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.u1.cin ;
assign _299_ = \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.u2.a  + \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.u2.b ;
assign { \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.u2.cout , \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.u2.s  } = _299_ + \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.u2.cin ;
assign \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.bin_s0  = ~ \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.b ;
always @(posedge \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.clk )
\sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.bin_s1  <= _301_;
always @(posedge \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.clk )
\sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.ain_s1  <= _300_;
always @(posedge \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.clk )
\sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.sum_s1  <= _303_;
always @(posedge \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.clk )
\sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.carry_s1  <= _302_;
assign _301_ = \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.ce  ? \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.bin_s0 [4:2] : \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.bin_s1 ;
assign _300_ = \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.ce  ? \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.a [4:2] : \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.ain_s1 ;
assign _302_ = \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.ce  ? \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.facout_s1  : \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.carry_s1 ;
assign _303_ = \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.ce  ? \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.fas_s1  : \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.sum_s1 ;
assign _304_ = \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.u1.a  + \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.u1.b ;
assign { \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.u1.cout , \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.u1.s  } = _304_ + \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.u1.cin ;
assign _305_ = \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.u2.a  + \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.u2.b ;
assign { \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.u2.cout , \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.u2.s  } = _305_ + \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.u2.cin ;
assign \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.bin_s0  = ~ \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.b ;
always @(posedge \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.clk )
\sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.bin_s1  <= _307_;
always @(posedge \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.clk )
\sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.ain_s1  <= _306_;
always @(posedge \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.clk )
\sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.sum_s1  <= _309_;
always @(posedge \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.clk )
\sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.carry_s1  <= _308_;
assign _307_ = \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.ce  ? \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.bin_s0 [7:4] : \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.bin_s1 ;
assign _306_ = \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.ce  ? \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.a [7:4] : \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.ain_s1 ;
assign _308_ = \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.ce  ? \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.facout_s1  : \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.carry_s1 ;
assign _309_ = \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.ce  ? \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.fas_s1  : \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.sum_s1 ;
assign _310_ = \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.u1.a  + \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.u1.b ;
assign { \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.u1.cout , \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.u1.s  } = _310_ + \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.u1.cin ;
assign _311_ = \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.u2.a  + \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.u2.b ;
assign { \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.u2.cout , \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.u2.s  } = _311_ + \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.u2.cin ;
assign _312_ = | op_0[3:2];
assign _313_ = | p_Result_1_reg_1117;
assign _314_ = p_Result_1_reg_1117 != 15'h7fff;
assign or_ln213_fu_619_p2 = op_0[1] | icmp_ln213_reg_1266;
assign or_ln340_fu_396_p2 = p_Result_10_reg_1098 | overflow_fu_392_p2;
assign or_ln384_fu_927_p2 = underflow_1_fu_922_p2 | overflow_1_reg_1476;
assign or_ln785_1_fu_877_p2 = xor_ln785_1_fu_871_p2 | p_Result_16_reg_1404;
assign or_ln785_2_fu_546_p2 = xor_ln785_3_fu_541_p2 | p_Result_10_reg_1098;
assign or_ln785_3_fu_514_p2 = and_ln785_1_fu_510_p2 | and_ln340_1_fu_506_p2;
assign or_ln785_fu_341_p2 = p_Result_11_reg_1110 | icmp_ln768_reg_1130;
assign or_ln786_fu_355_p2 = xor_ln786_fu_350_p2 | icmp_ln786_reg_1135;
assign or_ln788_fu_911_p2 = and_ln788_1_reg_1482 | and_ln781_fu_907_p2;
always @(posedge ap_clk)
trunc_ln1192_4_reg_1085 <= _060_;
always @(posedge ap_clk)
tmp_4_reg_1043 <= _057_;
always @(posedge ap_clk)
sub_ln1497_reg_1048 <= _056_;
always @(posedge ap_clk)
shl_ln1497_reg_1256 <= _055_;
always @(posedge ap_clk)
select_ln785_reg_1246 <= _053_;
always @(posedge ap_clk)
ret_V_12_reg_1558 <= _044_;
always @(posedge ap_clk)
ret_V_6_cast_reg_1563 <= _046_;
always @(posedge ap_clk)
p_Val2_1_reg_1224[3:2] <= _039_;
always @(posedge ap_clk)
select_ln340_reg_1230 <= _052_;
always @(posedge ap_clk)
sel_tmp11_reg_1235 <= _051_;
always @(posedge ap_clk)
ret_reg_1091 <= _050_;
always @(posedge ap_clk)
p_Result_10_reg_1098 <= _031_;
always @(posedge ap_clk)
trunc_ln731_reg_1105 <= _063_;
always @(posedge ap_clk)
p_Result_11_reg_1110 <= _032_;
always @(posedge ap_clk)
p_Result_1_reg_1117 <= _036_;
always @(posedge ap_clk)
or_ln384_reg_1502 <= _027_;
always @(posedge ap_clk)
or_ln340_reg_1190 <= _026_;
always @(posedge ap_clk)
ret_V_8_reg_1212 <= _047_;
always @(posedge ap_clk)
ret_V_reg_1217 <= _049_;
always @(posedge ap_clk)
op_29_V_reg_1543 <= _024_;
always @(posedge ap_clk)
op_7_V_reg_1271 <= _025_;
always @(posedge ap_clk)
r_reg_1277 <= _042_;
always @(posedge ap_clk)
ret_V_9_reg_1282 <= _048_;
always @(posedge ap_clk)
trunc_ln1192_1_reg_1287 <= _058_;
always @(posedge ap_clk)
trunc_ln1192_2_reg_1292 <= _059_;
always @(posedge ap_clk)
op_12_V_reg_1297 <= _020_;
always @(posedge ap_clk)
icmp_ln768_reg_1130 <= _018_;
always @(posedge ap_clk)
icmp_ln786_reg_1135 <= _019_;
always @(posedge ap_clk)
p_Result_13_reg_1141 <= _033_;
always @(posedge ap_clk)
ret_V_2_reg_1261 <= _045_;
always @(posedge ap_clk)
icmp_ln213_reg_1266 <= _017_;
always @(posedge ap_clk)
ashr_ln1497_reg_1251 <= _015_;
always @(posedge ap_clk)
or_ln785_reg_1151 <= _028_;
always @(posedge ap_clk)
xor_ln785_reg_1157 <= _064_;
always @(posedge ap_clk)
or_ln786_reg_1163 <= _029_;
always @(posedge ap_clk)
and_ln786_reg_1169 <= _012_;
always @(posedge ap_clk)
sh_V_reg_1175 <= _054_;
always @(posedge ap_clk)
op_19_V_reg_1522 <= _022_;
always @(posedge ap_clk)
add_ln69_4_reg_1528 <= _008_;
always @(posedge ap_clk)
add_ln69_6_reg_1533 <= _010_;
always @(posedge ap_clk)
overflow_1_reg_1476 <= _030_;
always @(posedge ap_clk)
and_ln788_1_reg_1482 <= _013_;
always @(posedge ap_clk)
ret_V_11_reg_1487 <= _043_;
always @(posedge ap_clk)
add_ln69_3_reg_1492 <= _007_;
always @(posedge ap_clk)
add_ln69_5_reg_1497 <= _009_;
always @(posedge ap_clk)
add_ln691_reg_1570 <= _005_;
always @(posedge ap_clk)
add_ln1192_2_reg_1327 <= _004_;
always @(posedge ap_clk)
p_Val2_5_reg_1332 <= _040_;
always @(posedge ap_clk)
add_ln69_reg_1337 <= _011_;
always @(posedge ap_clk)
add_ln69_1_reg_1342 <= _006_;
always @(posedge ap_clk)
op_16_V_reg_1382 <= _021_;
always @(posedge ap_clk)
add_ln1192_1_reg_1387 <= _003_;
always @(posedge ap_clk)
p_Result_14_reg_1392 <= _034_;
always @(posedge ap_clk)
p_Val2_6_reg_1398 <= _041_;
always @(posedge ap_clk)
p_Result_16_reg_1404 <= _035_;
always @(posedge ap_clk)
p_Result_2_reg_1411 <= _037_;
always @(posedge ap_clk)
p_Result_3_reg_1416 <= _038_;
always @(posedge ap_clk)
op_23_V_reg_1422 <= _023_;
always @(posedge ap_clk)
carry_1_reg_1432 <= _016_;
always @(posedge ap_clk)
Range2_all_ones_reg_1439 <= _002_;
always @(posedge ap_clk)
Range1_all_ones_reg_1444 <= _000_;
always @(posedge ap_clk)
Range1_all_zeros_reg_1451 <= _001_;
always @(posedge ap_clk)
ap_CS_fsm <= _014_;
always @(posedge ap_clk)
p_Val2_1_reg_1224[1:0] <= 2'h0;
always @(posedge ap_clk)
trunc_ln69_reg_1347 <= _062_;
always @(posedge ap_clk)
trunc_ln69_1_reg_1352 <= _061_;
assign _065_ = _072_ ? 2'h2 : 2'h1;
assign _315_ = ap_CS_fsm == 1'h1;
function [24:0] _869_;
input [24:0] a;
input [624:0] b;
input [24:0] s;
case (s)
25'b0000000000000000000000001:
_869_ = b[24:0];
25'b0000000000000000000000010:
_869_ = b[49:25];
25'b0000000000000000000000100:
_869_ = b[74:50];
25'b0000000000000000000001000:
_869_ = b[99:75];
25'b0000000000000000000010000:
_869_ = b[124:100];
25'b0000000000000000000100000:
_869_ = b[149:125];
25'b0000000000000000001000000:
_869_ = b[174:150];
25'b0000000000000000010000000:
_869_ = b[199:175];
25'b0000000000000000100000000:
_869_ = b[224:200];
25'b0000000000000001000000000:
_869_ = b[249:225];
25'b0000000000000010000000000:
_869_ = b[274:250];
25'b0000000000000100000000000:
_869_ = b[299:275];
25'b0000000000001000000000000:
_869_ = b[324:300];
25'b0000000000010000000000000:
_869_ = b[349:325];
25'b0000000000100000000000000:
_869_ = b[374:350];
25'b0000000001000000000000000:
_869_ = b[399:375];
25'b0000000010000000000000000:
_869_ = b[424:400];
25'b0000000100000000000000000:
_869_ = b[449:425];
25'b0000001000000000000000000:
_869_ = b[474:450];
25'b0000010000000000000000000:
_869_ = b[499:475];
25'b0000100000000000000000000:
_869_ = b[524:500];
25'b0001000000000000000000000:
_869_ = b[549:525];
25'b0010000000000000000000000:
_869_ = b[574:550];
25'b0100000000000000000000000:
_869_ = b[599:575];
25'b1000000000000000000000000:
_869_ = b[624:600];
25'b0000000000000000000000000:
_869_ = a;
default:
_869_ = 25'bx;
endcase
endfunction
assign ap_NS_fsm = _869_(25'hxxxxxxx, { 23'h000000, _065_, 600'h000002000002000002000002000002000002000002000002000002000002000002000002000002000002000002000002000002000002000002000002000002000002000002000000000001 }, { _315_, _339_, _338_, _337_, _336_, _335_, _334_, _333_, _332_, _331_, _330_, _329_, _328_, _327_, _326_, _325_, _324_, _323_, _322_, _321_, _320_, _319_, _318_, _317_, _316_ });
assign _316_ = ap_CS_fsm == 25'h1000000;
assign _317_ = ap_CS_fsm == 24'h800000;
assign _318_ = ap_CS_fsm == 23'h400000;
assign _319_ = ap_CS_fsm == 22'h200000;
assign _320_ = ap_CS_fsm == 21'h100000;
assign _321_ = ap_CS_fsm == 20'h80000;
assign _322_ = ap_CS_fsm == 19'h40000;
assign _323_ = ap_CS_fsm == 18'h20000;
assign _324_ = ap_CS_fsm == 17'h10000;
assign _325_ = ap_CS_fsm == 16'h8000;
assign _326_ = ap_CS_fsm == 15'h4000;
assign _327_ = ap_CS_fsm == 14'h2000;
assign _328_ = ap_CS_fsm == 13'h1000;
assign _329_ = ap_CS_fsm == 12'h800;
assign _330_ = ap_CS_fsm == 11'h400;
assign _331_ = ap_CS_fsm == 10'h200;
assign _332_ = ap_CS_fsm == 9'h100;
assign _333_ = ap_CS_fsm == 8'h80;
assign _334_ = ap_CS_fsm == 7'h40;
assign _335_ = ap_CS_fsm == 6'h20;
assign _336_ = ap_CS_fsm == 5'h10;
assign _337_ = ap_CS_fsm == 4'h8;
assign _338_ = ap_CS_fsm == 3'h4;
assign _339_ = ap_CS_fsm == 2'h2;
assign op_30_ap_vld = ap_CS_fsm[24] ? 1'h1 : 1'h0;
assign ap_idle = _071_ ? 1'h1 : 1'h0;
assign _062_ = _070_ ? grp_fu_407_p2[1:0] : trunc_ln69_reg_1347;
assign _061_ = _069_ ? grp_fu_416_p2[1:0] : trunc_ln69_1_reg_1352;
assign _060_ = ap_CS_fsm[2] ? op_5[0] : trunc_ln1192_4_reg_1085;
assign _057_ = ap_CS_fsm[0] ? op_8[3] : tmp_4_reg_1043;
assign _056_ = ap_CS_fsm[1] ? grp_fu_237_p2 : sub_ln1497_reg_1048;
assign _055_ = _068_ ? grp_fu_277_p2 : shl_ln1497_reg_1256;
assign _053_ = _067_ ? select_ln785_fu_556_p3 : select_ln785_reg_1246;
assign _046_ = ap_CS_fsm[21] ? grp_fu_988_p2[32:1] : ret_V_6_cast_reg_1563;
assign _044_ = ap_CS_fsm[21] ? grp_fu_988_p2 : ret_V_12_reg_1558;
assign _051_ = ap_CS_fsm[7] ? sel_tmp11_fu_520_p2 : sel_tmp11_reg_1235;
assign _052_ = ap_CS_fsm[7] ? select_ln340_fu_498_p3 : select_ln340_reg_1230;
assign _039_ = ap_CS_fsm[7] ? trunc_ln731_reg_1105 : p_Val2_1_reg_1224[3:2];
assign _036_ = ap_CS_fsm[3] ? grp_fu_251_p2[16:2] : p_Result_1_reg_1117;
assign _032_ = ap_CS_fsm[3] ? grp_fu_251_p2[1] : p_Result_11_reg_1110;
assign _063_ = ap_CS_fsm[3] ? grp_fu_251_p2[1:0] : trunc_ln731_reg_1105;
assign _031_ = ap_CS_fsm[3] ? grp_fu_251_p2[16] : p_Result_10_reg_1098;
assign _050_ = ap_CS_fsm[3] ? grp_fu_251_p2 : ret_reg_1091;
assign _027_ = ap_CS_fsm[16] ? or_ln384_fu_927_p2 : or_ln384_reg_1502;
assign _049_ = ap_CS_fsm[6] ? grp_fu_386_p2[6:1] : ret_V_reg_1217;
assign _047_ = ap_CS_fsm[6] ? grp_fu_386_p2 : ret_V_8_reg_1212;
assign _026_ = ap_CS_fsm[6] ? or_ln340_fu_396_p2 : or_ln340_reg_1190;
assign _024_ = ap_CS_fsm[19] ? grp_fu_969_p2 : op_29_V_reg_1543;
assign _020_ = ap_CS_fsm[9] ? op_12_V_fu_629_p2 : op_12_V_reg_1297;
assign _059_ = ap_CS_fsm[9] ? op_7_V_fu_568_p3[2:0] : trunc_ln1192_2_reg_1292;
assign _058_ = ap_CS_fsm[9] ? op_7_V_fu_568_p3[0] : trunc_ln1192_1_reg_1287;
assign _048_ = ap_CS_fsm[9] ? ret_V_9_fu_594_p3 : ret_V_9_reg_1282;
assign _042_ = ap_CS_fsm[9] ? r_fu_573_p3 : r_reg_1277;
assign _025_ = ap_CS_fsm[9] ? op_7_V_fu_568_p3 : op_7_V_reg_1271;
assign _033_ = ap_CS_fsm[4] ? op_6[7] : p_Result_13_reg_1141;
assign _019_ = ap_CS_fsm[4] ? icmp_ln786_fu_322_p2 : icmp_ln786_reg_1135;
assign _018_ = ap_CS_fsm[4] ? icmp_ln768_fu_317_p2 : icmp_ln768_reg_1130;
assign _017_ = ap_CS_fsm[8] ? icmp_ln213_fu_562_p2 : icmp_ln213_reg_1266;
assign _045_ = ap_CS_fsm[8] ? grp_fu_526_p2 : ret_V_2_reg_1261;
assign _015_ = _066_ ? grp_fu_264_p2 : ashr_ln1497_reg_1251;
assign _054_ = ap_CS_fsm[5] ? grp_fu_335_p2 : sh_V_reg_1175;
assign _012_ = ap_CS_fsm[5] ? and_ln786_fu_365_p2 : and_ln786_reg_1169;
assign _029_ = ap_CS_fsm[5] ? or_ln786_fu_355_p2 : or_ln786_reg_1163;
assign _064_ = ap_CS_fsm[5] ? xor_ln785_fu_345_p2 : xor_ln785_reg_1157;
assign _028_ = ap_CS_fsm[5] ? or_ln785_fu_341_p2 : or_ln785_reg_1151;
assign _010_ = ap_CS_fsm[17] ? grp_fu_947_p2 : add_ln69_6_reg_1533;
assign _008_ = ap_CS_fsm[17] ? grp_fu_939_p2 : add_ln69_4_reg_1528;
assign _022_ = ap_CS_fsm[17] ? op_19_V_fu_960_p3 : op_19_V_reg_1522;
assign _009_ = ap_CS_fsm[15] ? grp_fu_836_p2 : add_ln69_5_reg_1497;
assign _007_ = ap_CS_fsm[15] ? grp_fu_830_p2 : add_ln69_3_reg_1492;
assign _043_ = ap_CS_fsm[15] ? grp_fu_814_p2 : ret_V_11_reg_1487;
assign _013_ = ap_CS_fsm[15] ? and_ln788_1_fu_902_p2 : and_ln788_1_reg_1482;
assign _030_ = ap_CS_fsm[15] ? overflow_1_fu_887_p2 : overflow_1_reg_1476;
assign _005_ = ap_CS_fsm[23] ? grp_fu_1004_p2 : add_ln691_reg_1570;
assign _006_ = ap_CS_fsm[11] ? grp_fu_666_p2 : add_ln69_1_reg_1342;
assign _011_ = ap_CS_fsm[11] ? grp_fu_660_p2 : add_ln69_reg_1337;
assign _040_ = ap_CS_fsm[11] ? grp_fu_648_p2[2:1] : p_Val2_5_reg_1332;
assign _004_ = ap_CS_fsm[11] ? grp_fu_648_p2 : add_ln1192_2_reg_1327;
assign _023_ = ap_CS_fsm[13] ? grp_fu_731_p2 : op_23_V_reg_1422;
assign _038_ = ap_CS_fsm[13] ? grp_fu_709_p2[6:3] : p_Result_3_reg_1416;
assign _037_ = ap_CS_fsm[13] ? grp_fu_709_p2[6:4] : p_Result_2_reg_1411;
assign _035_ = ap_CS_fsm[13] ? grp_fu_723_p2[1] : p_Result_16_reg_1404;
assign _041_ = ap_CS_fsm[13] ? grp_fu_723_p2 : p_Val2_6_reg_1398;
assign _034_ = ap_CS_fsm[13] ? grp_fu_709_p2[6] : p_Result_14_reg_1392;
assign _003_ = ap_CS_fsm[13] ? grp_fu_715_p2 : add_ln1192_1_reg_1387;
assign _021_ = ap_CS_fsm[13] ? op_16_V_fu_736_p3 : op_16_V_reg_1382;
assign _001_ = ap_CS_fsm[14] ? Range1_all_zeros_fu_805_p2 : Range1_all_zeros_reg_1451;
assign _000_ = ap_CS_fsm[14] ? Range1_all_ones_fu_800_p2 : Range1_all_ones_reg_1444;
assign _002_ = ap_CS_fsm[14] ? Range2_all_ones_fu_795_p2 : Range2_all_ones_reg_1439;
assign _016_ = ap_CS_fsm[14] ? carry_1_fu_789_p2 : carry_1_reg_1432;
assign _014_ = ap_rst ? 25'h0000001 : ap_NS_fsm;
assign Range1_all_ones_fu_800_p2 = _077_ ? 1'h1 : 1'h0;
assign Range1_all_zeros_fu_805_p2 = _078_ ? 1'h1 : 1'h0;
assign Range2_all_ones_fu_795_p2 = _079_ ? 1'h1 : 1'h0;
assign deleted_ones_fu_865_p3 = carry_1_reg_1432 ? and_ln780_fu_860_p2 : Range1_all_ones_reg_1444;
assign deleted_zeros_fu_842_p3 = carry_1_reg_1432 ? Range1_all_ones_reg_1444 : Range1_all_zeros_reg_1451;
assign icmp_ln213_fu_562_p2 = _312_ ? 1'h1 : 1'h0;
assign icmp_ln768_fu_317_p2 = _313_ ? 1'h1 : 1'h0;
assign icmp_ln786_fu_322_p2 = _314_ ? 1'h1 : 1'h0;
assign op_16_V_fu_736_p3 = p_Result_13_reg_1141 ? trunc_ln69_reg_1347 : trunc_ln69_1_reg_1352;
assign op_19_V_fu_960_p3 = or_ln384_reg_1502 ? select_ln384_fu_953_p3 : p_Val2_6_reg_1398;
assign op_30 = ret_V_12_reg_1558[33] ? select_ln850_1_fu_1019_p3 : ret_V_6_cast_reg_1563;
assign op_7_V_fu_568_p3 = sel_tmp11_reg_1235 ? p_Val2_1_reg_1224 : select_ln785_reg_1246;
assign r_fu_573_p3 = tmp_4_reg_1043 ? shl_ln1497_reg_1256 : ashr_ln1497_reg_1251;
assign ret_V_9_fu_594_p3 = ret_V_8_reg_1212[6] ? select_ln850_fu_588_p3 : ret_V_reg_1217;
assign select_ln340_fu_498_p3 = and_ln340_fu_493_p2 ? { trunc_ln731_reg_1105, 2'h0 } : { ret_reg_1091[2], p_Val2_2_fu_472_p2 };
assign select_ln384_fu_953_p3 = overflow_1_reg_1476 ? 2'h1 : 2'h3;
assign select_ln785_fu_556_p3 = and_ln785_fu_551_p2 ? p_Val2_1_reg_1224 : select_ln340_reg_1230;
assign select_ln850_1_fu_1019_p3 = op_19_V_reg_1522[0] ? add_ln691_reg_1570 : ret_V_6_cast_reg_1563;
assign select_ln850_fu_588_p3 = op_9[0] ? ret_V_2_reg_1261 : ret_V_reg_1217;
assign xor_ln365_fu_460_p2 = ret_reg_1091[2] ^ ret_reg_1091[1];
assign ap_CS_fsm_state1 = ap_CS_fsm[0];
assign ap_CS_fsm_state10 = ap_CS_fsm[9];
assign ap_CS_fsm_state11 = ap_CS_fsm[10];
assign ap_CS_fsm_state12 = ap_CS_fsm[11];
assign ap_CS_fsm_state13 = ap_CS_fsm[12];
assign ap_CS_fsm_state14 = ap_CS_fsm[13];
assign ap_CS_fsm_state15 = ap_CS_fsm[14];
assign ap_CS_fsm_state16 = ap_CS_fsm[15];
assign ap_CS_fsm_state17 = ap_CS_fsm[16];
assign ap_CS_fsm_state18 = ap_CS_fsm[17];
assign ap_CS_fsm_state19 = ap_CS_fsm[18];
assign ap_CS_fsm_state2 = ap_CS_fsm[1];
assign ap_CS_fsm_state20 = ap_CS_fsm[19];
assign ap_CS_fsm_state21 = ap_CS_fsm[20];
assign ap_CS_fsm_state22 = ap_CS_fsm[21];
assign ap_CS_fsm_state23 = ap_CS_fsm[22];
assign ap_CS_fsm_state24 = ap_CS_fsm[23];
assign ap_CS_fsm_state25 = ap_CS_fsm[24];
assign ap_CS_fsm_state3 = ap_CS_fsm[2];
assign ap_CS_fsm_state4 = ap_CS_fsm[3];
assign ap_CS_fsm_state5 = ap_CS_fsm[4];
assign ap_CS_fsm_state6 = ap_CS_fsm[5];
assign ap_CS_fsm_state7 = ap_CS_fsm[6];
assign ap_CS_fsm_state8 = ap_CS_fsm[7];
assign ap_CS_fsm_state9 = ap_CS_fsm[8];
assign ap_done = op_30_ap_vld;
assign ap_ready = op_30_ap_vld;
assign grp_fu_237_p1 = { op_8[3], op_8 };
assign grp_fu_251_p0 = { op_2[15], op_2 };
assign grp_fu_251_p1 = { op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5 };
assign grp_fu_264_p1 = { op_8[3], op_8[3], op_8[3], op_8[3], op_8[3], op_8[3], op_8[3], op_8[3], op_8[3], op_8[3], op_8[3], op_8[3], op_8 };
assign grp_fu_277_p1 = { sub_ln1497_reg_1048[4], sub_ln1497_reg_1048[4], sub_ln1497_reg_1048[4], sub_ln1497_reg_1048[4], sub_ln1497_reg_1048[4], sub_ln1497_reg_1048[4], sub_ln1497_reg_1048[4], sub_ln1497_reg_1048[4], sub_ln1497_reg_1048[4], sub_ln1497_reg_1048[4], sub_ln1497_reg_1048[4], sub_ln1497_reg_1048 };
assign grp_fu_386_p0 = { 2'h0, op_3, 1'h0 };
assign grp_fu_386_p1 = { op_9[3], op_9[3], op_9[3], op_9 };
assign grp_fu_407_p1 = { 24'h000000, sh_V_reg_1175 };
assign grp_fu_416_p1 = { 24'h000000, op_6 };
assign grp_fu_648_p0 = { trunc_ln1192_4_reg_1085, 2'h0 };
assign grp_fu_660_p0 = { r_reg_1277[15], r_reg_1277 };
assign grp_fu_660_p1 = { op_10[7], op_10[7], op_10[7], op_10[7], op_10[7], op_10[7], op_10[7], op_10[7], op_10[7], op_10 };
assign grp_fu_666_p0 = { ret_V_9_reg_1282[5], ret_V_9_reg_1282 };
assign grp_fu_666_p1 = { 6'h00, op_12_V_reg_1297 };
assign grp_fu_709_p0 = { op_5[3], op_5, 2'h0 };
assign grp_fu_709_p1 = { op_7_V_reg_1271[3], op_7_V_reg_1271[3], op_7_V_reg_1271[3], op_7_V_reg_1271 };
assign grp_fu_715_p0 = { op_5[1:0], 2'h0 };
assign grp_fu_723_p1 = { 1'h0, trunc_ln1192_1_reg_1287 };
assign grp_fu_731_p0 = { add_ln69_1_reg_1342[6], add_ln69_1_reg_1342[6], add_ln69_1_reg_1342[6], add_ln69_1_reg_1342[6], add_ln69_1_reg_1342[6], add_ln69_1_reg_1342[6], add_ln69_1_reg_1342[6], add_ln69_1_reg_1342[6], add_ln69_1_reg_1342[6], add_ln69_1_reg_1342[6], add_ln69_1_reg_1342 };
assign grp_fu_814_p1 = { op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13 };
assign grp_fu_830_p0 = { op_14[1], op_14[1], op_14[1], op_14[1], op_14[1], op_14[1], op_14[1], op_14[1], op_14[1], op_14[1], op_14[1], op_14[1], op_14[1], op_14[1], op_14[1], op_14[1], op_14[1], op_14[1], op_14[1], op_14[1], op_14[1], op_14[1], op_14[1], op_14[1], op_14[1], op_14[1], op_14[1], op_14[1], op_14[1], op_14[1], op_14 };
assign grp_fu_836_p0 = { op_18[1], op_18 };
assign grp_fu_836_p1 = { op_16_V_reg_1382[1], op_16_V_reg_1382 };
assign grp_fu_939_p1 = { ret_V_11_reg_1487[16], ret_V_11_reg_1487[16], ret_V_11_reg_1487[16], ret_V_11_reg_1487[16], ret_V_11_reg_1487[16], ret_V_11_reg_1487[16], ret_V_11_reg_1487[16], ret_V_11_reg_1487[16], ret_V_11_reg_1487[16], ret_V_11_reg_1487[16], ret_V_11_reg_1487[16], ret_V_11_reg_1487[16], ret_V_11_reg_1487[16], ret_V_11_reg_1487[16], ret_V_11_reg_1487[16], ret_V_11_reg_1487 };
assign grp_fu_947_p0 = { add_ln69_5_reg_1497[2], add_ln69_5_reg_1497 };
assign grp_fu_947_p1 = { op_17[1], op_17[1], op_17 };
assign grp_fu_969_p0 = { add_ln69_6_reg_1533[3], add_ln69_6_reg_1533[3], add_ln69_6_reg_1533[3], add_ln69_6_reg_1533[3], add_ln69_6_reg_1533[3], add_ln69_6_reg_1533[3], add_ln69_6_reg_1533[3], add_ln69_6_reg_1533[3], add_ln69_6_reg_1533[3], add_ln69_6_reg_1533[3], add_ln69_6_reg_1533[3], add_ln69_6_reg_1533[3], add_ln69_6_reg_1533[3], add_ln69_6_reg_1533[3], add_ln69_6_reg_1533[3], add_ln69_6_reg_1533[3], add_ln69_6_reg_1533[3], add_ln69_6_reg_1533[3], add_ln69_6_reg_1533[3], add_ln69_6_reg_1533[3], add_ln69_6_reg_1533[3], add_ln69_6_reg_1533[3], add_ln69_6_reg_1533[3], add_ln69_6_reg_1533[3], add_ln69_6_reg_1533[3], add_ln69_6_reg_1533[3], add_ln69_6_reg_1533[3], add_ln69_6_reg_1533[3], add_ln69_6_reg_1533 };
assign grp_fu_988_p0 = { op_29_V_reg_1543[31], op_29_V_reg_1543, 1'h0 };
assign grp_fu_988_p1 = { op_19_V_reg_1522[1], op_19_V_reg_1522[1], op_19_V_reg_1522[1], op_19_V_reg_1522[1], op_19_V_reg_1522[1], op_19_V_reg_1522[1], op_19_V_reg_1522[1], op_19_V_reg_1522[1], op_19_V_reg_1522[1], op_19_V_reg_1522[1], op_19_V_reg_1522[1], op_19_V_reg_1522[1], op_19_V_reg_1522[1], op_19_V_reg_1522[1], op_19_V_reg_1522[1], op_19_V_reg_1522[1], op_19_V_reg_1522[1], op_19_V_reg_1522[1], op_19_V_reg_1522[1], op_19_V_reg_1522[1], op_19_V_reg_1522[1], op_19_V_reg_1522[1], op_19_V_reg_1522[1], op_19_V_reg_1522[1], op_19_V_reg_1522[1], op_19_V_reg_1522[1], op_19_V_reg_1522[1], op_19_V_reg_1522[1], op_19_V_reg_1522[1], op_19_V_reg_1522[1], op_19_V_reg_1522[1], op_19_V_reg_1522[1], op_19_V_reg_1522 };
assign lhs_V_1_fu_690_p1 = op_5;
assign lhs_V_1_fu_690_p3 = { op_5, 2'h0 };
assign lhs_V_fu_370_p3 = { op_3, 1'h0 };
assign p_Result_12_fu_439_p3 = ret_reg_1091[2];
assign p_Result_13_fu_327_p1 = op_6;
assign p_Result_15_fu_777_p3 = add_ln1192_2_reg_1327[2];
assign p_Result_5_fu_578_p3 = ret_V_8_reg_1212[6];
assign p_Result_9_fu_1009_p3 = ret_V_12_reg_1558[33];
assign p_Result_s_14_fu_478_p4 = { ret_reg_1091[2], p_Val2_2_fu_472_p2 };
assign p_Result_s_fu_531_p4 = op_0[3:2];
assign p_Val2_1_fu_432_p3 = { trunc_ln731_reg_1105, 2'h0 };
assign rhs_3_fu_977_p3 = { op_29_V_reg_1543, 1'h0 };
assign sext_ln1497_1_fu_270_p1 = { sub_ln1497_reg_1048[4], sub_ln1497_reg_1048[4], sub_ln1497_reg_1048[4], sub_ln1497_reg_1048[4], sub_ln1497_reg_1048[4], sub_ln1497_reg_1048[4], sub_ln1497_reg_1048[4], sub_ln1497_reg_1048[4], sub_ln1497_reg_1048[4], sub_ln1497_reg_1048[4], sub_ln1497_reg_1048[4], sub_ln1497_reg_1048[4], sub_ln1497_reg_1048[4], sub_ln1497_reg_1048[4], sub_ln1497_reg_1048[4], sub_ln1497_reg_1048[4], sub_ln1497_reg_1048[4], sub_ln1497_reg_1048[4], sub_ln1497_reg_1048[4], sub_ln1497_reg_1048[4], sub_ln1497_reg_1048[4], sub_ln1497_reg_1048[4], sub_ln1497_reg_1048[4], sub_ln1497_reg_1048[4], sub_ln1497_reg_1048[4], sub_ln1497_reg_1048[4], sub_ln1497_reg_1048[4], sub_ln1497_reg_1048 };
assign sext_ln1497_fu_225_p0 = op_8;
assign sext_ln215_1_fu_247_p0 = op_5;
assign sext_ln215_fu_243_p0 = op_2;
assign sext_ln545_fu_257_p0 = op_8;
assign sext_ln545_fu_257_p1 = { op_8[3], op_8[3], op_8[3], op_8[3], op_8[3], op_8[3], op_8[3], op_8[3], op_8[3], op_8[3], op_8[3], op_8[3], op_8[3], op_8[3], op_8[3], op_8[3], op_8[3], op_8[3], op_8[3], op_8[3], op_8[3], op_8[3], op_8[3], op_8[3], op_8[3], op_8[3], op_8[3], op_8[3], op_8 };
assign sext_ln703_fu_382_p0 = op_9;
assign sext_ln781_fu_401_p0 = op_6;
assign sext_ln781_fu_401_p1 = { op_6[7], op_6[7], op_6[7], op_6[7], op_6[7], op_6[7], op_6[7], op_6[7], op_6[7], op_6[7], op_6[7], op_6[7], op_6[7], op_6[7], op_6[7], op_6[7], op_6[7], op_6[7], op_6[7], op_6[7], op_6[7], op_6[7], op_6[7], op_6[7], op_6 };
assign shl_ln1192_fu_704_p0 = op_5;
assign tmp_10_fu_612_p3 = op_0[1];
assign tmp_1_fu_453_p3 = ret_reg_1091[1];
assign tmp_4_fu_229_p1 = op_8;
assign tmp_9_fu_847_p3 = add_ln1192_1_reg_1387[3];
assign tmp_fu_446_p3 = ret_reg_1091[2];
assign trunc_ln1192_1_fu_604_p1 = op_7_V_fu_568_p3[0];
assign trunc_ln1192_2_fu_608_p1 = op_7_V_fu_568_p3[2:0];
assign trunc_ln1192_4_fu_283_p0 = op_5;
assign trunc_ln1192_4_fu_283_p1 = op_5[0];
assign trunc_ln1192_fu_601_p1 = op_0[0];
assign trunc_ln69_1_fu_686_p1 = grp_fu_416_p2[1:0];
assign trunc_ln69_fu_682_p1 = grp_fu_407_p2[1:0];
assign trunc_ln731_fu_295_p1 = grp_fu_251_p2[1:0];
assign trunc_ln790_fu_893_p1 = p_Val2_6_reg_1398[0];
assign trunc_ln851_1_fu_1016_p1 = op_19_V_reg_1522[0];
assign trunc_ln851_fu_585_p0 = op_9;
assign trunc_ln851_fu_585_p1 = op_9[0];
assign zext_ln546_1_fu_413_p0 = op_6;
assign \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.ain_s0  = \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.a ;
assign \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.s  = { \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.fas_s2 , \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.sum_s1  };
assign \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.u2.a  = \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.ain_s1 ;
assign \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.u2.b  = \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.bin_s1 ;
assign \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.u2.cin  = \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.carry_s1 ;
assign \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.facout_s2  = \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.u2.cout ;
assign \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.fas_s2  = \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.u2.s ;
assign \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.u1.a  = \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.a [3:0];
assign \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.u1.b  = \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.bin_s0 [3:0];
assign \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.u1.cin  = 1'h1;
assign \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.facout_s1  = \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.u1.cout ;
assign \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.fas_s1  = \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.u1.s ;
assign \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.a  = \sub_8ns_8s_8_2_1_U5.din0 ;
assign \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.b  = \sub_8ns_8s_8_2_1_U5.din1 ;
assign \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.ce  = \sub_8ns_8s_8_2_1_U5.ce ;
assign \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.clk  = \sub_8ns_8s_8_2_1_U5.clk ;
assign \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.reset  = \sub_8ns_8s_8_2_1_U5.reset ;
assign \sub_8ns_8s_8_2_1_U5.dout  = \sub_8ns_8s_8_2_1_U5.top_sub_8ns_8s_8_2_1_Adder_2_U.s ;
assign \sub_8ns_8s_8_2_1_U5.ce  = 1'h1;
assign \sub_8ns_8s_8_2_1_U5.clk  = ap_clk;
assign \sub_8ns_8s_8_2_1_U5.din0  = 8'h00;
assign \sub_8ns_8s_8_2_1_U5.din1  = op_6;
assign grp_fu_335_p2 = \sub_8ns_8s_8_2_1_U5.dout ;
assign \sub_8ns_8s_8_2_1_U5.reset  = ap_rst;
assign \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.ain_s0  = \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.a ;
assign \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.s  = { \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.fas_s2 , \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.sum_s1  };
assign \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.u2.a  = \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.ain_s1 ;
assign \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.u2.b  = \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.bin_s1 ;
assign \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.u2.cin  = \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.carry_s1 ;
assign \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.facout_s2  = \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.u2.cout ;
assign \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.fas_s2  = \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.u2.s ;
assign \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.u1.a  = \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.a [1:0];
assign \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.u1.b  = \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.bin_s0 [1:0];
assign \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.u1.cin  = 1'h1;
assign \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.facout_s1  = \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.u1.cout ;
assign \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.fas_s1  = \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.u1.s ;
assign \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.a  = \sub_5ns_5s_5_2_1_U1.din0 ;
assign \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.b  = \sub_5ns_5s_5_2_1_U1.din1 ;
assign \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.ce  = \sub_5ns_5s_5_2_1_U1.ce ;
assign \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.clk  = \sub_5ns_5s_5_2_1_U1.clk ;
assign \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.reset  = \sub_5ns_5s_5_2_1_U1.reset ;
assign \sub_5ns_5s_5_2_1_U1.dout  = \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.s ;
assign \sub_5ns_5s_5_2_1_U1.ce  = 1'h1;
assign \sub_5ns_5s_5_2_1_U1.clk  = ap_clk;
assign \sub_5ns_5s_5_2_1_U1.din0  = 5'h00;
assign \sub_5ns_5s_5_2_1_U1.din1  = { op_8[3], op_8 };
assign grp_fu_237_p2 = \sub_5ns_5s_5_2_1_U1.dout ;
assign \sub_5ns_5s_5_2_1_U1.reset  = ap_rst;
assign \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.ain_s0  = \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.a ;
assign \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.s  = { \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.fas_s2 , \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.sum_s1  };
assign \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.u2.a  = \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.ain_s1 ;
assign \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.u2.b  = \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.bin_s1 ;
assign \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.u2.cin  = \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.carry_s1 ;
assign \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.facout_s2  = \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.u2.cout ;
assign \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.fas_s2  = \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.u2.s ;
assign \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.u1.a  = \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.a [7:0];
assign \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.u1.b  = \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.bin_s0 [7:0];
assign \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.u1.cin  = 1'h1;
assign \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.facout_s1  = \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.u1.cout ;
assign \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.fas_s1  = \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.u1.s ;
assign \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.a  = \sub_17s_17s_17_2_1_U2.din0 ;
assign \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.b  = \sub_17s_17s_17_2_1_U2.din1 ;
assign \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.ce  = \sub_17s_17s_17_2_1_U2.ce ;
assign \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.clk  = \sub_17s_17s_17_2_1_U2.clk ;
assign \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.reset  = \sub_17s_17s_17_2_1_U2.reset ;
assign \sub_17s_17s_17_2_1_U2.dout  = \sub_17s_17s_17_2_1_U2.top_sub_17s_17s_17_2_1_Adder_1_U.s ;
assign \sub_17s_17s_17_2_1_U2.ce  = 1'h1;
assign \sub_17s_17s_17_2_1_U2.clk  = ap_clk;
assign \sub_17s_17s_17_2_1_U2.din0  = { op_2[15], op_2 };
assign \sub_17s_17s_17_2_1_U2.din1  = { op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5 };
assign grp_fu_251_p2 = \sub_17s_17s_17_2_1_U2.dout ;
assign \sub_17s_17s_17_2_1_U2.reset  = ap_rst;
assign \shl_32s_8ns_32_7_1_U8.din1_cast  = \shl_32s_8ns_32_7_1_U8.din1 [7:0];
assign \shl_32s_8ns_32_7_1_U8.din1_mask  = 8'h03;
assign \shl_32s_8ns_32_7_1_U8.ce  = 1'h1;
assign \shl_32s_8ns_32_7_1_U8.clk  = ap_clk;
assign \shl_32s_8ns_32_7_1_U8.din0  = { op_6[7], op_6[7], op_6[7], op_6[7], op_6[7], op_6[7], op_6[7], op_6[7], op_6[7], op_6[7], op_6[7], op_6[7], op_6[7], op_6[7], op_6[7], op_6[7], op_6[7], op_6[7], op_6[7], op_6[7], op_6[7], op_6[7], op_6[7], op_6[7], op_6 };
assign \shl_32s_8ns_32_7_1_U8.din1  = { 24'h000000, op_6 };
assign grp_fu_416_p2 = \shl_32s_8ns_32_7_1_U8.dout ;
assign \shl_32s_8ns_32_7_1_U8.reset  = ap_rst;
assign \shl_16s_16ns_16_7_1_U4.din1_cast  = \shl_16s_16ns_16_7_1_U4.din1 ;
assign \shl_16s_16ns_16_7_1_U4.din1_mask  = 16'h0007;
assign \shl_16s_16ns_16_7_1_U4.ce  = 1'h1;
assign \shl_16s_16ns_16_7_1_U4.clk  = ap_clk;
assign \shl_16s_16ns_16_7_1_U4.din0  = op_2;
assign \shl_16s_16ns_16_7_1_U4.din1  = { sub_ln1497_reg_1048[4], sub_ln1497_reg_1048[4], sub_ln1497_reg_1048[4], sub_ln1497_reg_1048[4], sub_ln1497_reg_1048[4], sub_ln1497_reg_1048[4], sub_ln1497_reg_1048[4], sub_ln1497_reg_1048[4], sub_ln1497_reg_1048[4], sub_ln1497_reg_1048[4], sub_ln1497_reg_1048[4], sub_ln1497_reg_1048 };
assign grp_fu_277_p2 = \shl_16s_16ns_16_7_1_U4.dout ;
assign \shl_16s_16ns_16_7_1_U4.reset  = ap_rst;
assign \ashr_32s_8ns_32_7_1_U7.din1_cast  = \ashr_32s_8ns_32_7_1_U7.din1 [7:0];
assign \ashr_32s_8ns_32_7_1_U7.din1_mask  = 8'h03;
assign \ashr_32s_8ns_32_7_1_U7.ce  = 1'h1;
assign \ashr_32s_8ns_32_7_1_U7.clk  = ap_clk;
assign \ashr_32s_8ns_32_7_1_U7.din0  = { op_6[7], op_6[7], op_6[7], op_6[7], op_6[7], op_6[7], op_6[7], op_6[7], op_6[7], op_6[7], op_6[7], op_6[7], op_6[7], op_6[7], op_6[7], op_6[7], op_6[7], op_6[7], op_6[7], op_6[7], op_6[7], op_6[7], op_6[7], op_6[7], op_6 };
assign \ashr_32s_8ns_32_7_1_U7.din1  = { 24'h000000, sh_V_reg_1175 };
assign grp_fu_407_p2 = \ashr_32s_8ns_32_7_1_U7.dout ;
assign \ashr_32s_8ns_32_7_1_U7.reset  = ap_rst;
assign \ashr_16s_16ns_16_7_1_U3.din1_cast  = \ashr_16s_16ns_16_7_1_U3.din1 ;
assign \ashr_16s_16ns_16_7_1_U3.din1_mask  = 16'h0007;
assign \ashr_16s_16ns_16_7_1_U3.ce  = 1'h1;
assign \ashr_16s_16ns_16_7_1_U3.clk  = ap_clk;
assign \ashr_16s_16ns_16_7_1_U3.din0  = op_2;
assign \ashr_16s_16ns_16_7_1_U3.din1  = { op_8[3], op_8[3], op_8[3], op_8[3], op_8[3], op_8[3], op_8[3], op_8[3], op_8[3], op_8[3], op_8[3], op_8[3], op_8 };
assign grp_fu_264_p2 = \ashr_16s_16ns_16_7_1_U3.dout ;
assign \ashr_16s_16ns_16_7_1_U3.reset  = ap_rst;
assign \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.ain_s0  = \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.a ;
assign \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.bin_s0  = \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.b ;
assign \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.s  = { \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.fas_s2 , \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.sum_s1  };
assign \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.u2.a  = \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.ain_s1 ;
assign \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.u2.b  = \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.bin_s1 ;
assign \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.u2.cin  = \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.carry_s1 ;
assign \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.facout_s2  = \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.u2.cout ;
assign \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.fas_s2  = \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.u2.s ;
assign \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.u1.a  = \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.a [2:0];
assign \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.u1.b  = \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.b [2:0];
assign \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.u1.cin  = 1'h0;
assign \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.facout_s1  = \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.u1.cout ;
assign \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.fas_s1  = \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.u1.s ;
assign \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.a  = \add_7s_7s_7_2_1_U13.din0 ;
assign \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.b  = \add_7s_7s_7_2_1_U13.din1 ;
assign \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.ce  = \add_7s_7s_7_2_1_U13.ce ;
assign \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.clk  = \add_7s_7s_7_2_1_U13.clk ;
assign \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.reset  = \add_7s_7s_7_2_1_U13.reset ;
assign \add_7s_7s_7_2_1_U13.dout  = \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_8_U.s ;
assign \add_7s_7s_7_2_1_U13.ce  = 1'h1;
assign \add_7s_7s_7_2_1_U13.clk  = ap_clk;
assign \add_7s_7s_7_2_1_U13.din0  = { op_5[3], op_5, 2'h0 };
assign \add_7s_7s_7_2_1_U13.din1  = { op_7_V_reg_1271[3], op_7_V_reg_1271[3], op_7_V_reg_1271[3], op_7_V_reg_1271 };
assign grp_fu_709_p2 = \add_7s_7s_7_2_1_U13.dout ;
assign \add_7s_7s_7_2_1_U13.reset  = ap_rst;
assign \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.ain_s0  = \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.a ;
assign \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.bin_s0  = \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.b ;
assign \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.s  = { \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.fas_s2 , \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.sum_s1  };
assign \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.u2.a  = \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.ain_s1 ;
assign \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.u2.b  = \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.bin_s1 ;
assign \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.u2.cin  = \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.carry_s1 ;
assign \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.facout_s2  = \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.u2.cout ;
assign \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.fas_s2  = \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.u2.s ;
assign \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.u1.a  = \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.a [2:0];
assign \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.u1.b  = \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.b [2:0];
assign \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.u1.cin  = 1'h0;
assign \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.facout_s1  = \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.u1.cout ;
assign \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.fas_s1  = \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.u1.s ;
assign \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.a  = \add_7s_7ns_7_2_1_U12.din0 ;
assign \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.b  = \add_7s_7ns_7_2_1_U12.din1 ;
assign \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.ce  = \add_7s_7ns_7_2_1_U12.ce ;
assign \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.clk  = \add_7s_7ns_7_2_1_U12.clk ;
assign \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.reset  = \add_7s_7ns_7_2_1_U12.reset ;
assign \add_7s_7ns_7_2_1_U12.dout  = \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_7_U.s ;
assign \add_7s_7ns_7_2_1_U12.ce  = 1'h1;
assign \add_7s_7ns_7_2_1_U12.clk  = ap_clk;
assign \add_7s_7ns_7_2_1_U12.din0  = { ret_V_9_reg_1282[5], ret_V_9_reg_1282 };
assign \add_7s_7ns_7_2_1_U12.din1  = { 6'h00, op_12_V_reg_1297 };
assign grp_fu_666_p2 = \add_7s_7ns_7_2_1_U12.dout ;
assign \add_7s_7ns_7_2_1_U12.reset  = ap_rst;
assign \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.ain_s0  = \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.a ;
assign \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.bin_s0  = \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.b ;
assign \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.s  = { \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.fas_s2 , \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.sum_s1  };
assign \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.u2.a  = \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.ain_s1 ;
assign \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.u2.b  = \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.bin_s1 ;
assign \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.u2.cin  = \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.carry_s1 ;
assign \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.facout_s2  = \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.u2.cout ;
assign \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.fas_s2  = \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.u2.s ;
assign \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.u1.a  = \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.a [2:0];
assign \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.u1.b  = \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.b [2:0];
assign \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.u1.cin  = 1'h0;
assign \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.facout_s1  = \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.u1.cout ;
assign \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.fas_s1  = \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.u1.s ;
assign \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.a  = \add_7ns_7s_7_2_1_U6.din0 ;
assign \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.b  = \add_7ns_7s_7_2_1_U6.din1 ;
assign \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.ce  = \add_7ns_7s_7_2_1_U6.ce ;
assign \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.clk  = \add_7ns_7s_7_2_1_U6.clk ;
assign \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.reset  = \add_7ns_7s_7_2_1_U6.reset ;
assign \add_7ns_7s_7_2_1_U6.dout  = \add_7ns_7s_7_2_1_U6.top_add_7ns_7s_7_2_1_Adder_3_U.s ;
assign \add_7ns_7s_7_2_1_U6.ce  = 1'h1;
assign \add_7ns_7s_7_2_1_U6.clk  = ap_clk;
assign \add_7ns_7s_7_2_1_U6.din0  = { 2'h0, op_3, 1'h0 };
assign \add_7ns_7s_7_2_1_U6.din1  = { op_9[3], op_9[3], op_9[3], op_9 };
assign grp_fu_386_p2 = \add_7ns_7s_7_2_1_U6.dout ;
assign \add_7ns_7s_7_2_1_U6.reset  = ap_rst;
assign \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.ain_s0  = \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.a ;
assign \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.bin_s0  = \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.b ;
assign \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.s  = { \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.fas_s2 , \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.sum_s1  };
assign \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.u2.a  = \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.ain_s1 ;
assign \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.u2.b  = \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.bin_s1 ;
assign \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.u2.cin  = \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.carry_s1 ;
assign \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.facout_s2  = \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.u2.cout ;
assign \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.fas_s2  = \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.u2.s ;
assign \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.u1.a  = \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.a [2:0];
assign \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.u1.b  = \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.b [2:0];
assign \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.u1.cin  = 1'h0;
assign \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.facout_s1  = \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.u1.cout ;
assign \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.fas_s1  = \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.u1.s ;
assign \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.a  = \add_6ns_6ns_6_2_1_U9.din0 ;
assign \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.b  = \add_6ns_6ns_6_2_1_U9.din1 ;
assign \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.ce  = \add_6ns_6ns_6_2_1_U9.ce ;
assign \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.clk  = \add_6ns_6ns_6_2_1_U9.clk ;
assign \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.reset  = \add_6ns_6ns_6_2_1_U9.reset ;
assign \add_6ns_6ns_6_2_1_U9.dout  = \add_6ns_6ns_6_2_1_U9.top_add_6ns_6ns_6_2_1_Adder_4_U.s ;
assign \add_6ns_6ns_6_2_1_U9.ce  = 1'h1;
assign \add_6ns_6ns_6_2_1_U9.clk  = ap_clk;
assign \add_6ns_6ns_6_2_1_U9.din0  = ret_V_reg_1217;
assign \add_6ns_6ns_6_2_1_U9.din1  = 6'h01;
assign grp_fu_526_p2 = \add_6ns_6ns_6_2_1_U9.dout ;
assign \add_6ns_6ns_6_2_1_U9.reset  = ap_rst;
assign \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.ain_s0  = \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.a ;
assign \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.bin_s0  = \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.b ;
assign \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.s  = { \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.fas_s2 , \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.sum_s1  };
assign \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.u2.a  = \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.ain_s1 ;
assign \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.u2.b  = \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.bin_s1 ;
assign \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.u2.cin  = \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.carry_s1 ;
assign \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.facout_s2  = \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.u2.cout ;
assign \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.fas_s2  = \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.u2.s ;
assign \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.u1.a  = \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.a [1:0];
assign \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.u1.b  = \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.b [1:0];
assign \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.u1.cin  = 1'h0;
assign \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.facout_s1  = \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.u1.cout ;
assign \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.fas_s1  = \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.u1.s ;
assign \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.a  = \add_4s_4s_4_2_1_U21.din0 ;
assign \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.b  = \add_4s_4s_4_2_1_U21.din1 ;
assign \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.ce  = \add_4s_4s_4_2_1_U21.ce ;
assign \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.clk  = \add_4s_4s_4_2_1_U21.clk ;
assign \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.reset  = \add_4s_4s_4_2_1_U21.reset ;
assign \add_4s_4s_4_2_1_U21.dout  = \add_4s_4s_4_2_1_U21.top_add_4s_4s_4_2_1_Adder_16_U.s ;
assign \add_4s_4s_4_2_1_U21.ce  = 1'h1;
assign \add_4s_4s_4_2_1_U21.clk  = ap_clk;
assign \add_4s_4s_4_2_1_U21.din0  = { add_ln69_5_reg_1497[2], add_ln69_5_reg_1497 };
assign \add_4s_4s_4_2_1_U21.din1  = { op_17[1], op_17[1], op_17 };
assign grp_fu_947_p2 = \add_4s_4s_4_2_1_U21.dout ;
assign \add_4s_4s_4_2_1_U21.reset  = ap_rst;
assign \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.ain_s0  = \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.a ;
assign \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.bin_s0  = \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.b ;
assign \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.s  = { \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.fas_s2 , \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.sum_s1  };
assign \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.u2.a  = \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.ain_s1 ;
assign \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.u2.b  = \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.bin_s1 ;
assign \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.u2.cin  = \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.carry_s1 ;
assign \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.facout_s2  = \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.u2.cout ;
assign \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.fas_s2  = \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.u2.s ;
assign \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.u1.a  = \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.a [1:0];
assign \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.u1.b  = \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.b [1:0];
assign \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.u1.cin  = 1'h0;
assign \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.facout_s1  = \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.u1.cout ;
assign \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.fas_s1  = \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.u1.s ;
assign \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.a  = \add_4ns_4s_4_2_1_U14.din0 ;
assign \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.b  = \add_4ns_4s_4_2_1_U14.din1 ;
assign \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.ce  = \add_4ns_4s_4_2_1_U14.ce ;
assign \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.clk  = \add_4ns_4s_4_2_1_U14.clk ;
assign \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.reset  = \add_4ns_4s_4_2_1_U14.reset ;
assign \add_4ns_4s_4_2_1_U14.dout  = \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_9_U.s ;
assign \add_4ns_4s_4_2_1_U14.ce  = 1'h1;
assign \add_4ns_4s_4_2_1_U14.clk  = ap_clk;
assign \add_4ns_4s_4_2_1_U14.din0  = { op_5[1:0], 2'h0 };
assign \add_4ns_4s_4_2_1_U14.din1  = op_7_V_reg_1271;
assign grp_fu_715_p2 = \add_4ns_4s_4_2_1_U14.dout ;
assign \add_4ns_4s_4_2_1_U14.reset  = ap_rst;
assign \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.ain_s0  = \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.a ;
assign \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.bin_s0  = \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.b ;
assign \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.s  = { \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.fas_s2 , \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.sum_s1  };
assign \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.u2.a  = \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.ain_s1 ;
assign \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.u2.b  = \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.bin_s1 ;
assign \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.u2.cin  = \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.carry_s1 ;
assign \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.facout_s2  = \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.u2.cout ;
assign \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.fas_s2  = \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.u2.s ;
assign \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.u1.a  = \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.a [0];
assign \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.u1.b  = \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.b [0];
assign \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.u1.cin  = 1'h0;
assign \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.facout_s1  = \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.u1.cout ;
assign \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.fas_s1  = \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.u1.s ;
assign \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.a  = \add_3s_3s_3_2_1_U19.din0 ;
assign \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.b  = \add_3s_3s_3_2_1_U19.din1 ;
assign \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.ce  = \add_3s_3s_3_2_1_U19.ce ;
assign \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.clk  = \add_3s_3s_3_2_1_U19.clk ;
assign \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.reset  = \add_3s_3s_3_2_1_U19.reset ;
assign \add_3s_3s_3_2_1_U19.dout  = \add_3s_3s_3_2_1_U19.top_add_3s_3s_3_2_1_Adder_14_U.s ;
assign \add_3s_3s_3_2_1_U19.ce  = 1'h1;
assign \add_3s_3s_3_2_1_U19.clk  = ap_clk;
assign \add_3s_3s_3_2_1_U19.din0  = { op_18[1], op_18 };
assign \add_3s_3s_3_2_1_U19.din1  = { op_16_V_reg_1382[1], op_16_V_reg_1382 };
assign grp_fu_836_p2 = \add_3s_3s_3_2_1_U19.dout ;
assign \add_3s_3s_3_2_1_U19.reset  = ap_rst;
assign \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.ain_s0  = \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.a ;
assign \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.bin_s0  = \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.b ;
assign \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.s  = { \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.fas_s2 , \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.sum_s1  };
assign \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.u2.a  = \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.ain_s1 ;
assign \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.u2.b  = \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.bin_s1 ;
assign \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.u2.cin  = \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.carry_s1 ;
assign \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.facout_s2  = \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.u2.cout ;
assign \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.fas_s2  = \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.u2.s ;
assign \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.u1.a  = \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.a [0];
assign \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.u1.b  = \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.b [0];
assign \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.u1.cin  = 1'h0;
assign \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.facout_s1  = \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.u1.cout ;
assign \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.fas_s1  = \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.u1.s ;
assign \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.a  = \add_3ns_3ns_3_2_1_U10.din0 ;
assign \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.b  = \add_3ns_3ns_3_2_1_U10.din1 ;
assign \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.ce  = \add_3ns_3ns_3_2_1_U10.ce ;
assign \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.clk  = \add_3ns_3ns_3_2_1_U10.clk ;
assign \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.reset  = \add_3ns_3ns_3_2_1_U10.reset ;
assign \add_3ns_3ns_3_2_1_U10.dout  = \add_3ns_3ns_3_2_1_U10.top_add_3ns_3ns_3_2_1_Adder_5_U.s ;
assign \add_3ns_3ns_3_2_1_U10.ce  = 1'h1;
assign \add_3ns_3ns_3_2_1_U10.clk  = ap_clk;
assign \add_3ns_3ns_3_2_1_U10.din0  = { trunc_ln1192_4_reg_1085, 2'h0 };
assign \add_3ns_3ns_3_2_1_U10.din1  = trunc_ln1192_2_reg_1292;
assign grp_fu_648_p2 = \add_3ns_3ns_3_2_1_U10.dout ;
assign \add_3ns_3ns_3_2_1_U10.reset  = ap_rst;
assign \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.ain_s0  = \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.a ;
assign \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.bin_s0  = \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.b ;
assign \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.s  = { \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.fas_s2 , \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.sum_s1  };
assign \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.u2.a  = \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.ain_s1 ;
assign \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.u2.b  = \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.bin_s1 ;
assign \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.u2.cin  = \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.carry_s1 ;
assign \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.facout_s2  = \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.u2.cout ;
assign \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.fas_s2  = \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.u2.s ;
assign \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.u1.a  = \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.a [16:0];
assign \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.u1.b  = \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.b [16:0];
assign \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.u1.cin  = 1'h0;
assign \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.facout_s1  = \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.u1.cout ;
assign \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.fas_s1  = \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.u1.s ;
assign \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.a  = \add_34s_34s_34_2_1_U23.din0 ;
assign \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.b  = \add_34s_34s_34_2_1_U23.din1 ;
assign \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.ce  = \add_34s_34s_34_2_1_U23.ce ;
assign \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.clk  = \add_34s_34s_34_2_1_U23.clk ;
assign \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.reset  = \add_34s_34s_34_2_1_U23.reset ;
assign \add_34s_34s_34_2_1_U23.dout  = \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_17_U.s ;
assign \add_34s_34s_34_2_1_U23.ce  = 1'h1;
assign \add_34s_34s_34_2_1_U23.clk  = ap_clk;
assign \add_34s_34s_34_2_1_U23.din0  = { op_29_V_reg_1543[31], op_29_V_reg_1543, 1'h0 };
assign \add_34s_34s_34_2_1_U23.din1  = { op_19_V_reg_1522[1], op_19_V_reg_1522[1], op_19_V_reg_1522[1], op_19_V_reg_1522[1], op_19_V_reg_1522[1], op_19_V_reg_1522[1], op_19_V_reg_1522[1], op_19_V_reg_1522[1], op_19_V_reg_1522[1], op_19_V_reg_1522[1], op_19_V_reg_1522[1], op_19_V_reg_1522[1], op_19_V_reg_1522[1], op_19_V_reg_1522[1], op_19_V_reg_1522[1], op_19_V_reg_1522[1], op_19_V_reg_1522[1], op_19_V_reg_1522[1], op_19_V_reg_1522[1], op_19_V_reg_1522[1], op_19_V_reg_1522[1], op_19_V_reg_1522[1], op_19_V_reg_1522[1], op_19_V_reg_1522[1], op_19_V_reg_1522[1], op_19_V_reg_1522[1], op_19_V_reg_1522[1], op_19_V_reg_1522[1], op_19_V_reg_1522[1], op_19_V_reg_1522[1], op_19_V_reg_1522[1], op_19_V_reg_1522[1], op_19_V_reg_1522 };
assign grp_fu_988_p2 = \add_34s_34s_34_2_1_U23.dout ;
assign \add_34s_34s_34_2_1_U23.reset  = ap_rst;
assign \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.ain_s0  = \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.a ;
assign \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.bin_s0  = \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.b ;
assign \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.s  = { \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.fas_s2 , \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.sum_s1  };
assign \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.u2.a  = \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.ain_s1 ;
assign \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.u2.b  = \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.bin_s1 ;
assign \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.u2.cin  = \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.carry_s1 ;
assign \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.facout_s2  = \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.u2.cout ;
assign \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.fas_s2  = \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.u2.s ;
assign \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.u1.a  = \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.a [15:0];
assign \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.u1.b  = \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.b [15:0];
assign \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.u1.cin  = 1'h0;
assign \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.facout_s1  = \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.u1.cout ;
assign \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.fas_s1  = \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.u1.s ;
assign \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.a  = \add_32s_32ns_32_2_1_U22.din0 ;
assign \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.b  = \add_32s_32ns_32_2_1_U22.din1 ;
assign \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.ce  = \add_32s_32ns_32_2_1_U22.ce ;
assign \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.clk  = \add_32s_32ns_32_2_1_U22.clk ;
assign \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.reset  = \add_32s_32ns_32_2_1_U22.reset ;
assign \add_32s_32ns_32_2_1_U22.dout  = \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_13_U.s ;
assign \add_32s_32ns_32_2_1_U22.ce  = 1'h1;
assign \add_32s_32ns_32_2_1_U22.clk  = ap_clk;
assign \add_32s_32ns_32_2_1_U22.din0  = { add_ln69_6_reg_1533[3], add_ln69_6_reg_1533[3], add_ln69_6_reg_1533[3], add_ln69_6_reg_1533[3], add_ln69_6_reg_1533[3], add_ln69_6_reg_1533[3], add_ln69_6_reg_1533[3], add_ln69_6_reg_1533[3], add_ln69_6_reg_1533[3], add_ln69_6_reg_1533[3], add_ln69_6_reg_1533[3], add_ln69_6_reg_1533[3], add_ln69_6_reg_1533[3], add_ln69_6_reg_1533[3], add_ln69_6_reg_1533[3], add_ln69_6_reg_1533[3], add_ln69_6_reg_1533[3], add_ln69_6_reg_1533[3], add_ln69_6_reg_1533[3], add_ln69_6_reg_1533[3], add_ln69_6_reg_1533[3], add_ln69_6_reg_1533[3], add_ln69_6_reg_1533[3], add_ln69_6_reg_1533[3], add_ln69_6_reg_1533[3], add_ln69_6_reg_1533[3], add_ln69_6_reg_1533[3], add_ln69_6_reg_1533[3], add_ln69_6_reg_1533 };
assign \add_32s_32ns_32_2_1_U22.din1  = add_ln69_4_reg_1528;
assign grp_fu_969_p2 = \add_32s_32ns_32_2_1_U22.dout ;
assign \add_32s_32ns_32_2_1_U22.reset  = ap_rst;
assign \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.ain_s0  = \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.a ;
assign \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.bin_s0  = \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.b ;
assign \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.s  = { \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.fas_s2 , \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.sum_s1  };
assign \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.u2.a  = \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.ain_s1 ;
assign \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.u2.b  = \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.bin_s1 ;
assign \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.u2.cin  = \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.carry_s1 ;
assign \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.facout_s2  = \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.u2.cout ;
assign \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.fas_s2  = \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.u2.s ;
assign \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.u1.a  = \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.a [15:0];
assign \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.u1.b  = \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.b [15:0];
assign \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.u1.cin  = 1'h0;
assign \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.facout_s1  = \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.u1.cout ;
assign \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.fas_s1  = \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.u1.s ;
assign \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.a  = \add_32s_32ns_32_2_1_U18.din0 ;
assign \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.b  = \add_32s_32ns_32_2_1_U18.din1 ;
assign \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.ce  = \add_32s_32ns_32_2_1_U18.ce ;
assign \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.clk  = \add_32s_32ns_32_2_1_U18.clk ;
assign \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.reset  = \add_32s_32ns_32_2_1_U18.reset ;
assign \add_32s_32ns_32_2_1_U18.dout  = \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_13_U.s ;
assign \add_32s_32ns_32_2_1_U18.ce  = 1'h1;
assign \add_32s_32ns_32_2_1_U18.clk  = ap_clk;
assign \add_32s_32ns_32_2_1_U18.din0  = { op_14[1], op_14[1], op_14[1], op_14[1], op_14[1], op_14[1], op_14[1], op_14[1], op_14[1], op_14[1], op_14[1], op_14[1], op_14[1], op_14[1], op_14[1], op_14[1], op_14[1], op_14[1], op_14[1], op_14[1], op_14[1], op_14[1], op_14[1], op_14[1], op_14[1], op_14[1], op_14[1], op_14[1], op_14[1], op_14[1], op_14 };
assign \add_32s_32ns_32_2_1_U18.din1  = op_15;
assign grp_fu_830_p2 = \add_32s_32ns_32_2_1_U18.dout ;
assign \add_32s_32ns_32_2_1_U18.reset  = ap_rst;
assign \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.ain_s0  = \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.a ;
assign \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.bin_s0  = \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.b ;
assign \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.s  = { \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.fas_s2 , \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.sum_s1  };
assign \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.u2.a  = \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.ain_s1 ;
assign \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.u2.b  = \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.bin_s1 ;
assign \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.u2.cin  = \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.carry_s1 ;
assign \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.facout_s2  = \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.u2.cout ;
assign \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.fas_s2  = \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.u2.s ;
assign \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.u1.a  = \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.a [15:0];
assign \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.u1.b  = \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.b [15:0];
assign \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.u1.cin  = 1'h0;
assign \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.facout_s1  = \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.u1.cout ;
assign \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.fas_s1  = \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.u1.s ;
assign \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.a  = \add_32ns_32s_32_2_1_U20.din0 ;
assign \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.b  = \add_32ns_32s_32_2_1_U20.din1 ;
assign \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.ce  = \add_32ns_32s_32_2_1_U20.ce ;
assign \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.clk  = \add_32ns_32s_32_2_1_U20.clk ;
assign \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.reset  = \add_32ns_32s_32_2_1_U20.reset ;
assign \add_32ns_32s_32_2_1_U20.dout  = \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_15_U.s ;
assign \add_32ns_32s_32_2_1_U20.ce  = 1'h1;
assign \add_32ns_32s_32_2_1_U20.clk  = ap_clk;
assign \add_32ns_32s_32_2_1_U20.din0  = add_ln69_3_reg_1492;
assign \add_32ns_32s_32_2_1_U20.din1  = { ret_V_11_reg_1487[16], ret_V_11_reg_1487[16], ret_V_11_reg_1487[16], ret_V_11_reg_1487[16], ret_V_11_reg_1487[16], ret_V_11_reg_1487[16], ret_V_11_reg_1487[16], ret_V_11_reg_1487[16], ret_V_11_reg_1487[16], ret_V_11_reg_1487[16], ret_V_11_reg_1487[16], ret_V_11_reg_1487[16], ret_V_11_reg_1487[16], ret_V_11_reg_1487[16], ret_V_11_reg_1487[16], ret_V_11_reg_1487 };
assign grp_fu_939_p2 = \add_32ns_32s_32_2_1_U20.dout ;
assign \add_32ns_32s_32_2_1_U20.reset  = ap_rst;
assign \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.ain_s0  = \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.a ;
assign \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.bin_s0  = \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.b ;
assign \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.s  = { \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.fas_s2 , \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.sum_s1  };
assign \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.u2.a  = \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.ain_s1 ;
assign \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.u2.b  = \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.bin_s1 ;
assign \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.u2.cin  = \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.carry_s1 ;
assign \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.facout_s2  = \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.u2.cout ;
assign \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.fas_s2  = \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.u2.s ;
assign \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.u1.a  = \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.a [15:0];
assign \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.u1.b  = \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.b [15:0];
assign \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.u1.cin  = 1'h0;
assign \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.facout_s1  = \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.u1.cout ;
assign \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.fas_s1  = \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.u1.s ;
assign \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.a  = \add_32ns_32ns_32_2_1_U24.din0 ;
assign \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.b  = \add_32ns_32ns_32_2_1_U24.din1 ;
assign \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.ce  = \add_32ns_32ns_32_2_1_U24.ce ;
assign \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.clk  = \add_32ns_32ns_32_2_1_U24.clk ;
assign \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.reset  = \add_32ns_32ns_32_2_1_U24.reset ;
assign \add_32ns_32ns_32_2_1_U24.dout  = \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_18_U.s ;
assign \add_32ns_32ns_32_2_1_U24.ce  = 1'h1;
assign \add_32ns_32ns_32_2_1_U24.clk  = ap_clk;
assign \add_32ns_32ns_32_2_1_U24.din0  = ret_V_6_cast_reg_1563;
assign \add_32ns_32ns_32_2_1_U24.din1  = 32'd1;
assign grp_fu_1004_p2 = \add_32ns_32ns_32_2_1_U24.dout ;
assign \add_32ns_32ns_32_2_1_U24.reset  = ap_rst;
assign \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.ain_s0  = \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.a ;
assign \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.bin_s0  = \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.b ;
assign \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.s  = { \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.fas_s2 , \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.sum_s1  };
assign \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.u2.a  = \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.ain_s1 ;
assign \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.u2.b  = \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.bin_s1 ;
assign \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.u2.cin  = \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.carry_s1 ;
assign \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.facout_s2  = \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.u2.cout ;
assign \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.fas_s2  = \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.u2.s ;
assign \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.u1.a  = \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.a [0];
assign \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.u1.b  = \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.b [0];
assign \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.u1.cin  = 1'h0;
assign \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.facout_s1  = \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.u1.cout ;
assign \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.fas_s1  = \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.u1.s ;
assign \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.a  = \add_2ns_2ns_2_2_1_U15.din0 ;
assign \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.b  = \add_2ns_2ns_2_2_1_U15.din1 ;
assign \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.ce  = \add_2ns_2ns_2_2_1_U15.ce ;
assign \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.clk  = \add_2ns_2ns_2_2_1_U15.clk ;
assign \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.reset  = \add_2ns_2ns_2_2_1_U15.reset ;
assign \add_2ns_2ns_2_2_1_U15.dout  = \add_2ns_2ns_2_2_1_U15.top_add_2ns_2ns_2_2_1_Adder_10_U.s ;
assign \add_2ns_2ns_2_2_1_U15.ce  = 1'h1;
assign \add_2ns_2ns_2_2_1_U15.clk  = ap_clk;
assign \add_2ns_2ns_2_2_1_U15.din0  = p_Val2_5_reg_1332;
assign \add_2ns_2ns_2_2_1_U15.din1  = { 1'h0, trunc_ln1192_1_reg_1287 };
assign grp_fu_723_p2 = \add_2ns_2ns_2_2_1_U15.dout ;
assign \add_2ns_2ns_2_2_1_U15.reset  = ap_rst;
assign \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.ain_s0  = \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.a ;
assign \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.bin_s0  = \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.b ;
assign \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.s  = { \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.fas_s2 , \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.sum_s1  };
assign \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.u2.a  = \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.ain_s1 ;
assign \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.u2.b  = \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.bin_s1 ;
assign \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.u2.cin  = \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.carry_s1 ;
assign \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.facout_s2  = \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.u2.cout ;
assign \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.fas_s2  = \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.u2.s ;
assign \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.u1.a  = \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.a [7:0];
assign \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.u1.b  = \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.b [7:0];
assign \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.u1.cin  = 1'h0;
assign \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.facout_s1  = \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.u1.cout ;
assign \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.fas_s1  = \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.u1.s ;
assign \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.a  = \add_17s_17s_17_2_1_U11.din0 ;
assign \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.b  = \add_17s_17s_17_2_1_U11.din1 ;
assign \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.ce  = \add_17s_17s_17_2_1_U11.ce ;
assign \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.clk  = \add_17s_17s_17_2_1_U11.clk ;
assign \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.reset  = \add_17s_17s_17_2_1_U11.reset ;
assign \add_17s_17s_17_2_1_U11.dout  = \add_17s_17s_17_2_1_U11.top_add_17s_17s_17_2_1_Adder_6_U.s ;
assign \add_17s_17s_17_2_1_U11.ce  = 1'h1;
assign \add_17s_17s_17_2_1_U11.clk  = ap_clk;
assign \add_17s_17s_17_2_1_U11.din0  = { r_reg_1277[15], r_reg_1277 };
assign \add_17s_17s_17_2_1_U11.din1  = { op_10[7], op_10[7], op_10[7], op_10[7], op_10[7], op_10[7], op_10[7], op_10[7], op_10[7], op_10 };
assign grp_fu_660_p2 = \add_17s_17s_17_2_1_U11.dout ;
assign \add_17s_17s_17_2_1_U11.reset  = ap_rst;
assign \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.ain_s0  = \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.a ;
assign \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.bin_s0  = \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.b ;
assign \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.s  = { \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.fas_s2 , \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.sum_s1  };
assign \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.u2.a  = \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.ain_s1 ;
assign \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.u2.b  = \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.bin_s1 ;
assign \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.u2.cin  = \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.carry_s1 ;
assign \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.facout_s2  = \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.u2.cout ;
assign \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.fas_s2  = \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.u2.s ;
assign \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.u1.a  = \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.a [7:0];
assign \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.u1.b  = \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.b [7:0];
assign \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.u1.cin  = 1'h0;
assign \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.facout_s1  = \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.u1.cout ;
assign \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.fas_s1  = \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.u1.s ;
assign \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.a  = \add_17s_17ns_17_2_1_U16.din0 ;
assign \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.b  = \add_17s_17ns_17_2_1_U16.din1 ;
assign \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.ce  = \add_17s_17ns_17_2_1_U16.ce ;
assign \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.clk  = \add_17s_17ns_17_2_1_U16.clk ;
assign \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.reset  = \add_17s_17ns_17_2_1_U16.reset ;
assign \add_17s_17ns_17_2_1_U16.dout  = \add_17s_17ns_17_2_1_U16.top_add_17s_17ns_17_2_1_Adder_11_U.s ;
assign \add_17s_17ns_17_2_1_U16.ce  = 1'h1;
assign \add_17s_17ns_17_2_1_U16.clk  = ap_clk;
assign \add_17s_17ns_17_2_1_U16.din0  = { add_ln69_1_reg_1342[6], add_ln69_1_reg_1342[6], add_ln69_1_reg_1342[6], add_ln69_1_reg_1342[6], add_ln69_1_reg_1342[6], add_ln69_1_reg_1342[6], add_ln69_1_reg_1342[6], add_ln69_1_reg_1342[6], add_ln69_1_reg_1342[6], add_ln69_1_reg_1342[6], add_ln69_1_reg_1342 };
assign \add_17s_17ns_17_2_1_U16.din1  = add_ln69_reg_1337;
assign grp_fu_731_p2 = \add_17s_17ns_17_2_1_U16.dout ;
assign \add_17s_17ns_17_2_1_U16.reset  = ap_rst;
assign \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.ain_s0  = \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.a ;
assign \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.bin_s0  = \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.b ;
assign \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.s  = { \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.fas_s2 , \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.sum_s1  };
assign \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.u2.a  = \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.ain_s1 ;
assign \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.u2.b  = \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.bin_s1 ;
assign \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.u2.cin  = \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.carry_s1 ;
assign \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.facout_s2  = \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.u2.cout ;
assign \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.fas_s2  = \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.u2.s ;
assign \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.u1.a  = \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.a [7:0];
assign \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.u1.b  = \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.b [7:0];
assign \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.u1.cin  = 1'h0;
assign \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.facout_s1  = \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.u1.cout ;
assign \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.fas_s1  = \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.u1.s ;
assign \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.a  = \add_17ns_17s_17_2_1_U17.din0 ;
assign \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.b  = \add_17ns_17s_17_2_1_U17.din1 ;
assign \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.ce  = \add_17ns_17s_17_2_1_U17.ce ;
assign \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.clk  = \add_17ns_17s_17_2_1_U17.clk ;
assign \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.reset  = \add_17ns_17s_17_2_1_U17.reset ;
assign \add_17ns_17s_17_2_1_U17.dout  = \add_17ns_17s_17_2_1_U17.top_add_17ns_17s_17_2_1_Adder_12_U.s ;
assign \add_17ns_17s_17_2_1_U17.ce  = 1'h1;
assign \add_17ns_17s_17_2_1_U17.clk  = ap_clk;
assign \add_17ns_17s_17_2_1_U17.din0  = op_23_V_reg_1422;
assign \add_17ns_17s_17_2_1_U17.din1  = { op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13 };
assign grp_fu_814_p2 = \add_17ns_17s_17_2_1_U17.dout ;
assign \add_17ns_17s_17_2_1_U17.reset  = ap_rst;
endmodule


// Product machine:
module top_A_times_top_B (ap_start, op_0, op_10, op_13, op_14, op_15, op_17, op_18, op_2, op_3, op_5, op_6, op_8, op_9, ap_clk, unsafe_signal);
input ap_start;
input [3:0] op_0;
input [7:0] op_10;
input [1:0] op_13;
input [1:0] op_14;
input [31:0] op_15;
input [1:0] op_17;
input [1:0] op_18;
input [15:0] op_2;
input [3:0] op_3;
input [3:0] op_5;
input [7:0] op_6;
input [3:0] op_8;
input [3:0] op_9;
input ap_clk;
output unsafe_signal;
reg _setup;
initial _setup = 1'b0;
always @ (posedge ap_clk) _setup <= 1'b1;
reg ap_start_internal;
always @ (posedge ap_clk) if (!_setup) ap_start_internal <= ap_start;
reg [3:0] op_0_internal;
always @ (posedge ap_clk) if (!_setup) op_0_internal <= op_0;
reg [7:0] op_10_internal;
always @ (posedge ap_clk) if (!_setup) op_10_internal <= op_10;
reg [1:0] op_13_internal;
always @ (posedge ap_clk) if (!_setup) op_13_internal <= op_13;
reg [1:0] op_14_internal;
always @ (posedge ap_clk) if (!_setup) op_14_internal <= op_14;
reg [31:0] op_15_internal;
always @ (posedge ap_clk) if (!_setup) op_15_internal <= op_15;
reg [1:0] op_17_internal;
always @ (posedge ap_clk) if (!_setup) op_17_internal <= op_17;
reg [1:0] op_18_internal;
always @ (posedge ap_clk) if (!_setup) op_18_internal <= op_18;
reg [15:0] op_2_internal;
always @ (posedge ap_clk) if (!_setup) op_2_internal <= op_2;
reg [3:0] op_3_internal;
always @ (posedge ap_clk) if (!_setup) op_3_internal <= op_3;
reg [3:0] op_5_internal;
always @ (posedge ap_clk) if (!_setup) op_5_internal <= op_5;
reg [7:0] op_6_internal;
always @ (posedge ap_clk) if (!_setup) op_6_internal <= op_6;
reg [3:0] op_8_internal;
always @ (posedge ap_clk) if (!_setup) op_8_internal <= op_8;
reg [3:0] op_9_internal;
always @ (posedge ap_clk) if (!_setup) op_9_internal <= op_9;
wire ap_done_A;
wire ap_done_B;
wire ap_done_eq;
assign ap_done_eq = ap_done_A == ap_done_B;
wire ap_idle_A;
wire ap_idle_B;
wire ap_idle_eq;
assign ap_idle_eq = ap_idle_A == ap_idle_B;
wire ap_ready_A;
wire ap_ready_B;
wire ap_ready_eq;
assign ap_ready_eq = ap_ready_A == ap_ready_B;
wire [31:0] op_30_A;
wire [31:0] op_30_B;
wire op_30_eq;
assign op_30_eq = op_30_A == op_30_B;
wire op_30_ap_vld_A;
wire op_30_ap_vld_B;
wire clk_enable_A;
wire clk_enable_B;
assign clk_enable_A = _setup & (~op_30_ap_vld_A | op_30_ap_vld_B);
assign clk_enable_B = _setup;
wire divergent;
assign divergent = ~(ap_done_eq & ap_idle_eq & ap_ready_eq & op_30_eq);
assign unsafe_signal = op_30_ap_vld_A & op_30_ap_vld_B & divergent;
top_A instance_A (
    .ap_clk(ap_clk),
    .clk_enable(clk_enable_A),
    .ap_start(ap_start_internal),
    .op_0(op_0_internal),
    .op_10(op_10_internal),
    .op_13(op_13_internal),
    .op_14(op_14_internal),
    .op_15(op_15_internal),
    .op_17(op_17_internal),
    .op_18(op_18_internal),
    .op_2(op_2_internal),
    .op_3(op_3_internal),
    .op_5(op_5_internal),
    .op_6(op_6_internal),
    .op_8(op_8_internal),
    .op_9(op_9_internal),
    .ap_done(ap_done_A),
    .ap_idle(ap_idle_A),
    .ap_ready(ap_ready_A),
    .op_30(op_30_A),
    .op_30_ap_vld(op_30_ap_vld_A)
);
top_B instance_B (
    .ap_clk(ap_clk),
    .clk_enable(clk_enable_B),
    .ap_start(ap_start_internal),
    .op_0(op_0_internal),
    .op_10(op_10_internal),
    .op_13(op_13_internal),
    .op_14(op_14_internal),
    .op_15(op_15_internal),
    .op_17(op_17_internal),
    .op_18(op_18_internal),
    .op_2(op_2_internal),
    .op_3(op_3_internal),
    .op_5(op_5_internal),
    .op_6(op_6_internal),
    .op_8(op_8_internal),
    .op_9(op_9_internal),
    .ap_done(ap_done_B),
    .ap_idle(ap_idle_B),
    .ap_ready(ap_ready_B),
    .op_30(op_30_B),
    .op_30_ap_vld(op_30_ap_vld_B)
);
endmodule
