// Processed by function `construct_kairos` in `verilog_tricks.py`.
// Machine A:
// Processed by function `add_clk_enable_signal` in `verilog_tricks.py`.
// Processed by function `remove_reset_signal` in `verilog_tricks.py`.
module top_A (
  ap_clk,
  ap_start,
  ap_done,
  ap_idle,
  ap_ready,
  op_0,
  op_1,
  op_2,
  op_3,
  op_9,
  op_12,
  op_13,
  op_14,
  op_16,
  op_17,
  op_30,
  op_30_ap_vld,
clk_enable
);
input clk_enable;


input ap_clk;
wire ap_rst;
assign ap_rst = op_30_ap_vld;
input ap_start;
input [15:0] op_0;
input op_1;
input [3:0] op_12;
input op_13;
input [1:0] op_14;
input [1:0] op_16;
input [3:0] op_17;
input [7:0] op_2;
input op_3;
input [3:0] op_9;
output ap_done;
output ap_idle;
output ap_ready;
output [31:0] op_30;
output op_30_ap_vld;


reg Range2_all_ones_reg_800;
reg [6:0] \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.ain_s1 ;
reg [6:0] \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.bin_s1 ;
reg \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.carry_s1 ;
reg [5:0] \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.sum_s1 ;
reg [6:0] \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.ain_s1 ;
reg [6:0] \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.bin_s1 ;
reg \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.carry_s1 ;
reg [6:0] \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.sum_s1 ;
reg [6:0] \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.ain_s1 ;
reg [6:0] \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.bin_s1 ;
reg \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.carry_s1 ;
reg [6:0] \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.sum_s1 ;
reg [6:0] \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.ain_s1 ;
reg [6:0] \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.bin_s1 ;
reg \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.carry_s1 ;
reg [6:0] \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.sum_s1 ;
reg [7:0] \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.ain_s1 ;
reg [7:0] \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.bin_s1 ;
reg \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.carry_s1 ;
reg [6:0] \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.sum_s1 ;
reg [7:0] \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.ain_s1 ;
reg [7:0] \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.bin_s1 ;
reg \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.carry_s1 ;
reg [6:0] \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.sum_s1 ;
reg [8:0] \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.ain_s1 ;
reg [8:0] \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.bin_s1 ;
reg \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.carry_s1 ;
reg [7:0] \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.sum_s1 ;
reg [8:0] \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.ain_s1 ;
reg [8:0] \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.bin_s1 ;
reg \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.carry_s1 ;
reg [8:0] \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.sum_s1 ;
reg [8:0] \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.ain_s1 ;
reg [8:0] \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.bin_s1 ;
reg \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.carry_s1 ;
reg [8:0] \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.sum_s1 ;
reg \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.ain_s1 ;
reg \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.bin_s1 ;
reg \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.carry_s1 ;
reg \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.sum_s1 ;
reg \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.ain_s1 ;
reg \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.bin_s1 ;
reg \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.carry_s1 ;
reg \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.sum_s1 ;
reg [1:0] \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.ain_s1 ;
reg [1:0] \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.bin_s1 ;
reg \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.carry_s1 ;
reg \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.sum_s1 ;
reg [1:0] \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.ain_s1 ;
reg [1:0] \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.bin_s1 ;
reg \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.carry_s1 ;
reg [1:0] \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.sum_s1 ;
reg [1:0] \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.ain_s1 ;
reg [1:0] \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.bin_s1 ;
reg \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.carry_s1 ;
reg [1:0] \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.sum_s1 ;
reg [2:0] \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.ain_s1 ;
reg [2:0] \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.bin_s1 ;
reg \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.carry_s1 ;
reg [1:0] \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.sum_s1 ;
reg [4:0] \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.ain_s1 ;
reg [4:0] \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.bin_s1 ;
reg \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.carry_s1 ;
reg [3:0] \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.sum_s1 ;
reg [13:0] add_ln69_1_reg_1045;
reg [2:0] add_ln69_2_reg_1030;
reg [3:0] add_ln69_3_reg_1050;
reg [17:0] add_ln69_5_reg_1115;
reg [4:0] add_ln69_7_reg_1120;
reg [13:0] add_ln69_reg_1025;
reg and_ln786_reg_867;
reg [22:0] ap_CS_fsm = 23'h000001;
reg deleted_zeros_reg_856;
reg icmp_ln851_1_reg_938;
reg icmp_ln851_2_reg_809;
reg icmp_ln851_3_reg_985;
reg icmp_ln851_reg_779;
reg neg_src_reg_862;
reg [13:0] op_25_V_reg_1060;
reg [13:0] op_26_V_reg_1075;
reg [3:0] op_6_V_reg_917;
reg or_ln778_reg_845;
reg p_Result_3_reg_771;
reg p_Result_4_reg_789;
reg p_Result_5_reg_820;
reg [3:0] p_Val2_3_reg_814;
reg [1:0] ret_V_11_reg_968;
reg [1:0] ret_V_12_reg_995;
reg [8:0] ret_V_17_reg_873;
reg [1:0] ret_V_18_reg_953;
reg [16:0] ret_V_19_reg_900;
reg [12:0] ret_V_20_reg_980;
reg [4:0] ret_V_21_reg_963;
reg [1:0] ret_V_22_reg_1015;
reg [14:0] ret_V_24_reg_1090;
reg [1:0] ret_V_2_reg_933;
reg [12:0] ret_V_4_reg_905;
reg [12:0] ret_V_6_reg_958;
reg [1:0] ret_V_reg_878;
reg [8:0] select_ln1192_reg_834;
reg [3:0] select_ln340_reg_895;
reg [13:0] select_ln69_reg_1020;
reg [4:0] select_ln703_reg_928;
reg [1:0] select_ln831_reg_922;
reg [2:0] \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.ain_s1 ;
reg [2:0] \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.bin_s1 ;
reg \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.carry_s1 ;
reg [1:0] \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.sum_s1 ;
reg [1:0] tmp_reg_948;
reg [2:0] trunc_ln851_2_reg_975;
reg [3:0] trunc_ln851_reg_912;
reg xor_ln416_reg_839;
wire _000_;
wire [13:0] _001_;
wire [2:0] _002_;
wire [3:0] _003_;
wire [17:0] _004_;
wire [4:0] _005_;
wire [13:0] _006_;
wire _007_;
wire [22:0] _008_;
wire _009_;
wire _010_;
wire _011_;
wire _012_;
wire _013_;
wire _014_;
wire [13:0] _015_;
wire [13:0] _016_;
wire [3:0] _017_;
wire _018_;
wire _019_;
wire _020_;
wire _021_;
wire [3:0] _022_;
wire [1:0] _023_;
wire [1:0] _024_;
wire [8:0] _025_;
wire [1:0] _026_;
wire [16:0] _027_;
wire [12:0] _028_;
wire [4:0] _029_;
wire [1:0] _030_;
wire [14:0] _031_;
wire [1:0] _032_;
wire [12:0] _033_;
wire [12:0] _034_;
wire [1:0] _035_;
wire [1:0] _036_;
wire [3:0] _037_;
wire [7:0] _038_;
wire [1:0] _039_;
wire [1:0] _040_;
wire [1:0] _041_;
wire [2:0] _042_;
wire [3:0] _043_;
wire _044_;
wire [1:0] _045_;
wire _046_;
wire _047_;
wire _048_;
wire _049_;
wire _050_;
wire _051_;
wire _052_;
wire _053_;
wire [6:0] _054_;
wire [6:0] _055_;
wire _056_;
wire [5:0] _057_;
wire [6:0] _058_;
wire [7:0] _059_;
wire [6:0] _060_;
wire [6:0] _061_;
wire _062_;
wire [6:0] _063_;
wire [7:0] _064_;
wire [7:0] _065_;
wire [6:0] _066_;
wire [6:0] _067_;
wire _068_;
wire [6:0] _069_;
wire [7:0] _070_;
wire [7:0] _071_;
wire [6:0] _072_;
wire [6:0] _073_;
wire _074_;
wire [6:0] _075_;
wire [7:0] _076_;
wire [7:0] _077_;
wire [7:0] _078_;
wire [7:0] _079_;
wire _080_;
wire [6:0] _081_;
wire [7:0] _082_;
wire [8:0] _083_;
wire [7:0] _084_;
wire [7:0] _085_;
wire _086_;
wire [6:0] _087_;
wire [7:0] _088_;
wire [8:0] _089_;
wire [8:0] _090_;
wire [8:0] _091_;
wire _092_;
wire [7:0] _093_;
wire [8:0] _094_;
wire [9:0] _095_;
wire [8:0] _096_;
wire [8:0] _097_;
wire _098_;
wire [8:0] _099_;
wire [9:0] _100_;
wire [9:0] _101_;
wire [8:0] _102_;
wire [8:0] _103_;
wire _104_;
wire [8:0] _105_;
wire [9:0] _106_;
wire [9:0] _107_;
wire _108_;
wire _109_;
wire _110_;
wire _111_;
wire [1:0] _112_;
wire [1:0] _113_;
wire _114_;
wire _115_;
wire _116_;
wire _117_;
wire [1:0] _118_;
wire [1:0] _119_;
wire [1:0] _120_;
wire [1:0] _121_;
wire _122_;
wire _123_;
wire [1:0] _124_;
wire [2:0] _125_;
wire [1:0] _126_;
wire [1:0] _127_;
wire _128_;
wire [1:0] _129_;
wire [2:0] _130_;
wire [2:0] _131_;
wire [1:0] _132_;
wire [1:0] _133_;
wire _134_;
wire [1:0] _135_;
wire [2:0] _136_;
wire [2:0] _137_;
wire [2:0] _138_;
wire [2:0] _139_;
wire _140_;
wire [1:0] _141_;
wire [2:0] _142_;
wire [3:0] _143_;
wire [4:0] _144_;
wire [4:0] _145_;
wire _146_;
wire [3:0] _147_;
wire [4:0] _148_;
wire [5:0] _149_;
wire [2:0] _150_;
wire [2:0] _151_;
wire _152_;
wire [1:0] _153_;
wire [2:0] _154_;
wire [3:0] _155_;
wire _156_;
wire _157_;
wire _158_;
wire _159_;
wire _160_;
wire _161_;
wire _162_;
wire _163_;
wire _164_;
wire _165_;
wire _166_;
wire _167_;
wire _168_;
wire _169_;
wire _170_;
wire _171_;
wire _172_;
wire _173_;
wire _174_;
wire _175_;
wire _176_;
wire _177_;
wire _178_;
wire [7:0] Range2_all_ones_fu_241_p1;
wire \add_13ns_13ns_13_2_1_U5.ce ;
wire \add_13ns_13ns_13_2_1_U5.clk ;
wire [12:0] \add_13ns_13ns_13_2_1_U5.din0 ;
wire [12:0] \add_13ns_13ns_13_2_1_U5.din1 ;
wire [12:0] \add_13ns_13ns_13_2_1_U5.dout ;
wire \add_13ns_13ns_13_2_1_U5.reset ;
wire [12:0] \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.a ;
wire [12:0] \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.ain_s0 ;
wire [12:0] \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.b ;
wire [12:0] \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.bin_s0 ;
wire \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.ce ;
wire \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.clk ;
wire \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.facout_s1 ;
wire \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.facout_s2 ;
wire [5:0] \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.fas_s1 ;
wire [6:0] \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.fas_s2 ;
wire \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.reset ;
wire [12:0] \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.s ;
wire [5:0] \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.u1.a ;
wire [5:0] \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.u1.b ;
wire \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.u1.cin ;
wire \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.u1.cout ;
wire [5:0] \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.u1.s ;
wire [6:0] \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.u2.a ;
wire [6:0] \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.u2.b ;
wire \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.u2.cin ;
wire \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.u2.cout ;
wire [6:0] \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.u2.s ;
wire \add_14ns_14ns_14_2_1_U10.ce ;
wire \add_14ns_14ns_14_2_1_U10.clk ;
wire [13:0] \add_14ns_14ns_14_2_1_U10.din0 ;
wire [13:0] \add_14ns_14ns_14_2_1_U10.din1 ;
wire [13:0] \add_14ns_14ns_14_2_1_U10.dout ;
wire \add_14ns_14ns_14_2_1_U10.reset ;
wire [13:0] \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.a ;
wire [13:0] \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.ain_s0 ;
wire [13:0] \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.b ;
wire [13:0] \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.bin_s0 ;
wire \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.ce ;
wire \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.clk ;
wire \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.facout_s1 ;
wire \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.facout_s2 ;
wire [6:0] \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.fas_s1 ;
wire [6:0] \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.fas_s2 ;
wire \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.reset ;
wire [13:0] \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.s ;
wire [6:0] \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.u1.a ;
wire [6:0] \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.u1.b ;
wire \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.u1.cin ;
wire \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.u1.cout ;
wire [6:0] \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.u1.s ;
wire [6:0] \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.u2.a ;
wire [6:0] \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.u2.b ;
wire \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.u2.cin ;
wire \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.u2.cout ;
wire [6:0] \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.u2.s ;
wire \add_14s_14ns_14_2_1_U12.ce ;
wire \add_14s_14ns_14_2_1_U12.clk ;
wire [13:0] \add_14s_14ns_14_2_1_U12.din0 ;
wire [13:0] \add_14s_14ns_14_2_1_U12.din1 ;
wire [13:0] \add_14s_14ns_14_2_1_U12.dout ;
wire \add_14s_14ns_14_2_1_U12.reset ;
wire [13:0] \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.a ;
wire [13:0] \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.ain_s0 ;
wire [13:0] \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.b ;
wire [13:0] \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.bin_s0 ;
wire \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.ce ;
wire \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.clk ;
wire \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.facout_s1 ;
wire \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.facout_s2 ;
wire [6:0] \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.fas_s1 ;
wire [6:0] \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.fas_s2 ;
wire \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.reset ;
wire [13:0] \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.s ;
wire [6:0] \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.u1.a ;
wire [6:0] \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.u1.b ;
wire \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.u1.cin ;
wire \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.u1.cout ;
wire [6:0] \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.u1.s ;
wire [6:0] \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.u2.a ;
wire [6:0] \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.u2.b ;
wire \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.u2.cin ;
wire \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.u2.cout ;
wire [6:0] \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.u2.s ;
wire \add_14s_14ns_14_2_1_U8.ce ;
wire \add_14s_14ns_14_2_1_U8.clk ;
wire [13:0] \add_14s_14ns_14_2_1_U8.din0 ;
wire [13:0] \add_14s_14ns_14_2_1_U8.din1 ;
wire [13:0] \add_14s_14ns_14_2_1_U8.dout ;
wire \add_14s_14ns_14_2_1_U8.reset ;
wire [13:0] \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.a ;
wire [13:0] \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.ain_s0 ;
wire [13:0] \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.b ;
wire [13:0] \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.bin_s0 ;
wire \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.ce ;
wire \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.clk ;
wire \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.facout_s1 ;
wire \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.facout_s2 ;
wire [6:0] \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.fas_s1 ;
wire [6:0] \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.fas_s2 ;
wire \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.reset ;
wire [13:0] \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.s ;
wire [6:0] \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.u1.a ;
wire [6:0] \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.u1.b ;
wire \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.u1.cin ;
wire \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.u1.cout ;
wire [6:0] \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.u1.s ;
wire [6:0] \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.u2.a ;
wire [6:0] \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.u2.b ;
wire \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.u2.cin ;
wire \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.u2.cout ;
wire [6:0] \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.u2.s ;
wire \add_15ns_15s_15_2_1_U13.ce ;
wire \add_15ns_15s_15_2_1_U13.clk ;
wire [14:0] \add_15ns_15s_15_2_1_U13.din0 ;
wire [14:0] \add_15ns_15s_15_2_1_U13.din1 ;
wire [14:0] \add_15ns_15s_15_2_1_U13.dout ;
wire \add_15ns_15s_15_2_1_U13.reset ;
wire [14:0] \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.a ;
wire [14:0] \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.ain_s0 ;
wire [14:0] \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.b ;
wire [14:0] \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.bin_s0 ;
wire \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.ce ;
wire \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.clk ;
wire \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.facout_s1 ;
wire \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.facout_s2 ;
wire [6:0] \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.fas_s1 ;
wire [7:0] \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.fas_s2 ;
wire \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.reset ;
wire [14:0] \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.s ;
wire [6:0] \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.u1.a ;
wire [6:0] \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.u1.b ;
wire \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.u1.cin ;
wire \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.u1.cout ;
wire [6:0] \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.u1.s ;
wire [7:0] \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.u2.a ;
wire [7:0] \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.u2.b ;
wire \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.u2.cin ;
wire \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.u2.cout ;
wire [7:0] \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.u2.s ;
wire \add_15s_15s_15_2_1_U14.ce ;
wire \add_15s_15s_15_2_1_U14.clk ;
wire [14:0] \add_15s_15s_15_2_1_U14.din0 ;
wire [14:0] \add_15s_15s_15_2_1_U14.din1 ;
wire [14:0] \add_15s_15s_15_2_1_U14.dout ;
wire \add_15s_15s_15_2_1_U14.reset ;
wire [14:0] \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.a ;
wire [14:0] \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.ain_s0 ;
wire [14:0] \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.b ;
wire [14:0] \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.bin_s0 ;
wire \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.ce ;
wire \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.clk ;
wire \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.facout_s1 ;
wire \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.facout_s2 ;
wire [6:0] \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.fas_s1 ;
wire [7:0] \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.fas_s2 ;
wire \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.reset ;
wire [14:0] \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.s ;
wire [6:0] \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.u1.a ;
wire [6:0] \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.u1.b ;
wire \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.u1.cin ;
wire \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.u1.cout ;
wire [6:0] \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.u1.s ;
wire [7:0] \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.u2.a ;
wire [7:0] \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.u2.b ;
wire \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.u2.cin ;
wire \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.u2.cout ;
wire [7:0] \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.u2.s ;
wire \add_17s_17s_17_2_1_U3.ce ;
wire \add_17s_17s_17_2_1_U3.clk ;
wire [16:0] \add_17s_17s_17_2_1_U3.din0 ;
wire [16:0] \add_17s_17s_17_2_1_U3.din1 ;
wire [16:0] \add_17s_17s_17_2_1_U3.dout ;
wire \add_17s_17s_17_2_1_U3.reset ;
wire [16:0] \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.a ;
wire [16:0] \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.ain_s0 ;
wire [16:0] \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.b ;
wire [16:0] \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.bin_s0 ;
wire \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.ce ;
wire \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.clk ;
wire \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.facout_s1 ;
wire \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.facout_s2 ;
wire [7:0] \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.fas_s1 ;
wire [8:0] \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.fas_s2 ;
wire \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.reset ;
wire [16:0] \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.s ;
wire [7:0] \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.u1.a ;
wire [7:0] \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.u1.b ;
wire \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.u1.cin ;
wire \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.u1.cout ;
wire [7:0] \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.u1.s ;
wire [8:0] \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.u2.a ;
wire [8:0] \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.u2.b ;
wire \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.u2.cin ;
wire \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.u2.cout ;
wire [8:0] \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.u2.s ;
wire \add_18s_18ns_18_2_1_U15.ce ;
wire \add_18s_18ns_18_2_1_U15.clk ;
wire [17:0] \add_18s_18ns_18_2_1_U15.din0 ;
wire [17:0] \add_18s_18ns_18_2_1_U15.din1 ;
wire [17:0] \add_18s_18ns_18_2_1_U15.dout ;
wire \add_18s_18ns_18_2_1_U15.reset ;
wire [17:0] \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.a ;
wire [17:0] \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.ain_s0 ;
wire [17:0] \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.b ;
wire [17:0] \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.bin_s0 ;
wire \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.ce ;
wire \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.clk ;
wire \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.facout_s1 ;
wire \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.facout_s2 ;
wire [8:0] \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.fas_s1 ;
wire [8:0] \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.fas_s2 ;
wire \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.reset ;
wire [17:0] \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.s ;
wire [8:0] \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.u1.a ;
wire [8:0] \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.u1.b ;
wire \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.u1.cin ;
wire \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.u1.cout ;
wire [8:0] \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.u1.s ;
wire [8:0] \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.u2.a ;
wire [8:0] \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.u2.b ;
wire \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.u2.cin ;
wire \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.u2.cout ;
wire [8:0] \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.u2.s ;
wire \add_18s_18ns_18_2_1_U17.ce ;
wire \add_18s_18ns_18_2_1_U17.clk ;
wire [17:0] \add_18s_18ns_18_2_1_U17.din0 ;
wire [17:0] \add_18s_18ns_18_2_1_U17.din1 ;
wire [17:0] \add_18s_18ns_18_2_1_U17.dout ;
wire \add_18s_18ns_18_2_1_U17.reset ;
wire [17:0] \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.a ;
wire [17:0] \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.ain_s0 ;
wire [17:0] \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.b ;
wire [17:0] \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.bin_s0 ;
wire \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.ce ;
wire \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.clk ;
wire \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.facout_s1 ;
wire \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.facout_s2 ;
wire [8:0] \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.fas_s1 ;
wire [8:0] \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.fas_s2 ;
wire \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.reset ;
wire [17:0] \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.s ;
wire [8:0] \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.u1.a ;
wire [8:0] \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.u1.b ;
wire \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.u1.cin ;
wire \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.u1.cout ;
wire [8:0] \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.u1.s ;
wire [8:0] \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.u2.a ;
wire [8:0] \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.u2.b ;
wire \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.u2.cin ;
wire \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.u2.cout ;
wire [8:0] \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.u2.s ;
wire \add_2ns_2ns_2_2_1_U4.ce ;
wire \add_2ns_2ns_2_2_1_U4.clk ;
wire [1:0] \add_2ns_2ns_2_2_1_U4.din0 ;
wire [1:0] \add_2ns_2ns_2_2_1_U4.din1 ;
wire [1:0] \add_2ns_2ns_2_2_1_U4.dout ;
wire \add_2ns_2ns_2_2_1_U4.reset ;
wire [1:0] \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.a ;
wire [1:0] \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.ain_s0 ;
wire [1:0] \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.b ;
wire [1:0] \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.bin_s0 ;
wire \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.ce ;
wire \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.clk ;
wire \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.facout_s1 ;
wire \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.facout_s2 ;
wire \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.fas_s1 ;
wire \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.fas_s2 ;
wire \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.reset ;
wire [1:0] \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.s ;
wire \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.u1.a ;
wire \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.u1.b ;
wire \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.u1.cin ;
wire \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.u1.cout ;
wire \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.u1.s ;
wire \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.u2.a ;
wire \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.u2.b ;
wire \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.u2.cin ;
wire \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.u2.cout ;
wire \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.u2.s ;
wire \add_2ns_2ns_2_2_1_U7.ce ;
wire \add_2ns_2ns_2_2_1_U7.clk ;
wire [1:0] \add_2ns_2ns_2_2_1_U7.din0 ;
wire [1:0] \add_2ns_2ns_2_2_1_U7.din1 ;
wire [1:0] \add_2ns_2ns_2_2_1_U7.dout ;
wire \add_2ns_2ns_2_2_1_U7.reset ;
wire [1:0] \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.a ;
wire [1:0] \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.ain_s0 ;
wire [1:0] \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.b ;
wire [1:0] \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.bin_s0 ;
wire \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.ce ;
wire \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.clk ;
wire \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.facout_s1 ;
wire \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.facout_s2 ;
wire \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.fas_s1 ;
wire \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.fas_s2 ;
wire \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.reset ;
wire [1:0] \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.s ;
wire \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.u1.a ;
wire \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.u1.b ;
wire \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.u1.cin ;
wire \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.u1.cout ;
wire \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.u1.s ;
wire \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.u2.a ;
wire \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.u2.b ;
wire \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.u2.cin ;
wire \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.u2.cout ;
wire \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.u2.s ;
wire \add_3ns_3ns_3_2_1_U9.ce ;
wire \add_3ns_3ns_3_2_1_U9.clk ;
wire [2:0] \add_3ns_3ns_3_2_1_U9.din0 ;
wire [2:0] \add_3ns_3ns_3_2_1_U9.din1 ;
wire [2:0] \add_3ns_3ns_3_2_1_U9.dout ;
wire \add_3ns_3ns_3_2_1_U9.reset ;
wire [2:0] \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.a ;
wire [2:0] \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.ain_s0 ;
wire [2:0] \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.b ;
wire [2:0] \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.bin_s0 ;
wire \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.ce ;
wire \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.clk ;
wire \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.facout_s1 ;
wire \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.facout_s2 ;
wire \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.fas_s1 ;
wire [1:0] \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.fas_s2 ;
wire \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.reset ;
wire [2:0] \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.s ;
wire \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.u1.a ;
wire \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.u1.b ;
wire \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.u1.cin ;
wire \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.u1.cout ;
wire \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.u1.s ;
wire [1:0] \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.u2.a ;
wire [1:0] \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.u2.b ;
wire \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.u2.cin ;
wire \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.u2.cout ;
wire [1:0] \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.u2.s ;
wire \add_4ns_4ns_4_2_1_U1.ce ;
wire \add_4ns_4ns_4_2_1_U1.clk ;
wire [3:0] \add_4ns_4ns_4_2_1_U1.din0 ;
wire [3:0] \add_4ns_4ns_4_2_1_U1.din1 ;
wire [3:0] \add_4ns_4ns_4_2_1_U1.dout ;
wire \add_4ns_4ns_4_2_1_U1.reset ;
wire [3:0] \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.a ;
wire [3:0] \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.ain_s0 ;
wire [3:0] \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.b ;
wire [3:0] \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.bin_s0 ;
wire \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.ce ;
wire \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.clk ;
wire \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.facout_s1 ;
wire \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.facout_s2 ;
wire [1:0] \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.fas_s1 ;
wire [1:0] \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.fas_s2 ;
wire \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.reset ;
wire [3:0] \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.s ;
wire [1:0] \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.u1.a ;
wire [1:0] \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.u1.b ;
wire \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.u1.cin ;
wire \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.u1.cout ;
wire [1:0] \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.u1.s ;
wire [1:0] \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.u2.a ;
wire [1:0] \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.u2.b ;
wire \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.u2.cin ;
wire \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.u2.cout ;
wire [1:0] \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.u2.s ;
wire \add_4ns_4s_4_2_1_U11.ce ;
wire \add_4ns_4s_4_2_1_U11.clk ;
wire [3:0] \add_4ns_4s_4_2_1_U11.din0 ;
wire [3:0] \add_4ns_4s_4_2_1_U11.din1 ;
wire [3:0] \add_4ns_4s_4_2_1_U11.dout ;
wire \add_4ns_4s_4_2_1_U11.reset ;
wire [3:0] \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.a ;
wire [3:0] \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.ain_s0 ;
wire [3:0] \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.b ;
wire [3:0] \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.bin_s0 ;
wire \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.ce ;
wire \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.clk ;
wire \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.facout_s1 ;
wire \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.facout_s2 ;
wire [1:0] \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.fas_s1 ;
wire [1:0] \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.fas_s2 ;
wire \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.reset ;
wire [3:0] \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.s ;
wire [1:0] \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.u1.a ;
wire [1:0] \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.u1.b ;
wire \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.u1.cin ;
wire \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.u1.cout ;
wire [1:0] \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.u1.s ;
wire [1:0] \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.u2.a ;
wire [1:0] \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.u2.b ;
wire \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.u2.cin ;
wire \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.u2.cout ;
wire [1:0] \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.u2.s ;
wire \add_5s_5ns_5_2_1_U16.ce ;
wire \add_5s_5ns_5_2_1_U16.clk ;
wire [4:0] \add_5s_5ns_5_2_1_U16.din0 ;
wire [4:0] \add_5s_5ns_5_2_1_U16.din1 ;
wire [4:0] \add_5s_5ns_5_2_1_U16.dout ;
wire \add_5s_5ns_5_2_1_U16.reset ;
wire [4:0] \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.a ;
wire [4:0] \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.ain_s0 ;
wire [4:0] \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.b ;
wire [4:0] \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.bin_s0 ;
wire \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.ce ;
wire \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.clk ;
wire \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.facout_s1 ;
wire \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.facout_s2 ;
wire [1:0] \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.fas_s1 ;
wire [2:0] \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.fas_s2 ;
wire \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.reset ;
wire [4:0] \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.s ;
wire [1:0] \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.u1.a ;
wire [1:0] \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.u1.b ;
wire \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.u1.cin ;
wire \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.u1.cout ;
wire [1:0] \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.u1.s ;
wire [2:0] \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.u2.a ;
wire [2:0] \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.u2.b ;
wire \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.u2.cin ;
wire \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.u2.cout ;
wire [2:0] \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.u2.s ;
wire \add_9ns_9s_9_2_1_U2.ce ;
wire \add_9ns_9s_9_2_1_U2.clk ;
wire [8:0] \add_9ns_9s_9_2_1_U2.din0 ;
wire [8:0] \add_9ns_9s_9_2_1_U2.din1 ;
wire [8:0] \add_9ns_9s_9_2_1_U2.dout ;
wire \add_9ns_9s_9_2_1_U2.reset ;
wire [8:0] \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.a ;
wire [8:0] \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.ain_s0 ;
wire [8:0] \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.b ;
wire [8:0] \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.bin_s0 ;
wire \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.ce ;
wire \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.clk ;
wire \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.facout_s1 ;
wire \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.facout_s2 ;
wire [3:0] \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.fas_s1 ;
wire [4:0] \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.fas_s2 ;
wire \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.reset ;
wire [8:0] \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.s ;
wire [3:0] \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.u1.a ;
wire [3:0] \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.u1.b ;
wire \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.u1.cin ;
wire \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.u1.cout ;
wire [3:0] \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.u1.s ;
wire [4:0] \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.u2.a ;
wire [4:0] \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.u2.b ;
wire \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.u2.cin ;
wire \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.u2.cout ;
wire [4:0] \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.u2.s ;
wire and_ln781_1_fu_320_p2;
wire and_ln781_fu_324_p2;
wire and_ln785_1_fu_448_p2;
wire and_ln785_fu_439_p2;
wire and_ln786_1_fu_340_p2;
wire and_ln786_fu_345_p2;
wire ap_CS_fsm_state1;
wire ap_CS_fsm_state10;
wire ap_CS_fsm_state11;
wire ap_CS_fsm_state12;
wire ap_CS_fsm_state13;
wire ap_CS_fsm_state14;
wire ap_CS_fsm_state15;
wire ap_CS_fsm_state16;
wire ap_CS_fsm_state17;
wire ap_CS_fsm_state18;
wire ap_CS_fsm_state19;
wire ap_CS_fsm_state2;
wire ap_CS_fsm_state20;
wire ap_CS_fsm_state21;
wire ap_CS_fsm_state22;
wire ap_CS_fsm_state23;
wire ap_CS_fsm_state3;
wire ap_CS_fsm_state4;
wire ap_CS_fsm_state5;
wire ap_CS_fsm_state6;
wire ap_CS_fsm_state7;
wire ap_CS_fsm_state8;
wire ap_CS_fsm_state9;
wire [22:0] ap_NS_fsm;
wire ap_clk;
wire ap_done;
wire ap_idle;
wire ap_ready;
wire ap_rst;
wire ap_start;
wire deleted_zeros_fu_298_p2;
wire [3:0] grp_fu_235_p0;
wire [3:0] grp_fu_235_p1;
wire [3:0] grp_fu_235_p2;
wire [8:0] grp_fu_293_p1;
wire [8:0] grp_fu_293_p2;
wire [16:0] grp_fu_376_p0;
wire [16:0] grp_fu_376_p1;
wire [16:0] grp_fu_376_p2;
wire [1:0] grp_fu_420_p2;
wire [12:0] grp_fu_478_p2;
wire [4:0] grp_fu_495_p2;
wire [1:0] grp_fu_593_p2;
wire [13:0] grp_fu_613_p0;
wire [13:0] grp_fu_613_p1;
wire [13:0] grp_fu_613_p2;
wire [2:0] grp_fu_619_p0;
wire [2:0] grp_fu_619_p1;
wire [2:0] grp_fu_619_p2;
wire [13:0] grp_fu_654_p2;
wire [3:0] grp_fu_661_p0;
wire [3:0] grp_fu_661_p1;
wire [3:0] grp_fu_661_p2;
wire [13:0] grp_fu_670_p0;
wire [13:0] grp_fu_670_p2;
wire [14:0] grp_fu_694_p0;
wire [14:0] grp_fu_694_p1;
wire [14:0] grp_fu_694_p2;
wire [14:0] grp_fu_717_p0;
wire [14:0] grp_fu_717_p1;
wire [14:0] grp_fu_717_p2;
wire [17:0] grp_fu_740_p0;
wire [17:0] grp_fu_740_p1;
wire [17:0] grp_fu_740_p2;
wire [4:0] grp_fu_746_p0;
wire [4:0] grp_fu_746_p1;
wire [4:0] grp_fu_746_p2;
wire [17:0] grp_fu_755_p0;
wire [17:0] grp_fu_755_p2;
wire icmp_ln851_1_fu_473_p2;
wire icmp_ln851_2_fu_253_p2;
wire icmp_ln851_3_fu_588_p2;
wire icmp_ln851_fu_199_p2;
wire neg_src_fu_335_p2;
wire [15:0] op_0;
wire op_1;
wire [3:0] op_12;
wire op_13;
wire [1:0] op_14;
wire [1:0] op_16;
wire [3:0] op_17;
wire [7:0] op_2;
wire op_3;
wire [31:0] op_30;
wire op_30_ap_vld;
wire [3:0] op_6_V_fu_453_p3;
wire [3:0] op_9;
wire or_ln340_1_fu_408_p2;
wire or_ln340_fu_403_p2;
wire or_ln778_fu_285_p2;
wire or_ln780_fu_315_p2;
wire or_ln785_1_fu_443_p2;
wire or_ln785_fu_387_p2;
wire overflow_fu_397_p2;
wire p_Result_1_fu_536_p3;
wire p_Result_2_fu_569_p3;
wire [7:0] p_Result_3_fu_187_p1;
wire [7:0] p_Result_4_fu_215_p1;
wire p_Result_s_fu_625_p3;
wire [7:0] p_Val2_2_fu_205_p1;
wire p_Val2_s_fu_675_p1;
wire [1:0] p_Val2_s_fu_675_p3;
wire [1:0] ret_V_18_fu_548_p3;
wire [12:0] ret_V_20_fu_581_p3;
wire [1:0] ret_V_22_fu_637_p3;
wire [4:0] ret_V_23_fu_520_p2;
wire ret_V_9_fu_483_p2;
wire [4:0] rhs_2_fu_512_p3;
wire [4:0] rhs_fu_364_p3;
wire select_ln1192_fu_267_p0;
wire [8:0] select_ln1192_fu_267_p3;
wire [3:0] select_ln340_fu_413_p3;
wire [1:0] select_ln353_fu_506_p3;
wire select_ln69_fu_644_p0;
wire [7:0] select_ln69_fu_644_p3;
wire select_ln703_fu_466_p0;
wire [4:0] select_ln703_fu_466_p3;
wire [1:0] select_ln831_fu_459_p3;
wire [12:0] select_ln850_1_fu_576_p3;
wire [1:0] select_ln850_3_fu_632_p3;
wire [1:0] select_ln850_6_fu_500_p3;
wire [1:0] select_ln850_fu_543_p3;
wire [15:0] sext_ln69_2_fu_730_p1;
wire [4:0] sext_ln703_2_fu_492_p1;
wire [7:0] sext_ln703_fu_290_p0;
wire \sub_5ns_5s_5_2_1_U6.ce ;
wire \sub_5ns_5s_5_2_1_U6.clk ;
wire [4:0] \sub_5ns_5s_5_2_1_U6.din0 ;
wire [4:0] \sub_5ns_5s_5_2_1_U6.din1 ;
wire [4:0] \sub_5ns_5s_5_2_1_U6.dout ;
wire \sub_5ns_5s_5_2_1_U6.reset ;
wire [4:0] \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.a ;
wire [4:0] \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.ain_s0 ;
wire [4:0] \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.b ;
wire [4:0] \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.bin_s0 ;
wire \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.ce ;
wire \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.clk ;
wire \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.facout_s1 ;
wire \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.facout_s2 ;
wire [1:0] \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.fas_s1 ;
wire [2:0] \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.fas_s2 ;
wire \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.reset ;
wire [4:0] \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.s ;
wire [1:0] \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.u1.a ;
wire [1:0] \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.u1.b ;
wire \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.u1.cin ;
wire \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.u1.cout ;
wire [1:0] \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.u1.s ;
wire [2:0] \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.u2.a ;
wire [2:0] \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.u2.b ;
wire \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.u2.cin ;
wire \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.u2.cout ;
wire [2:0] \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.u2.s ;
wire [7:0] tmp_6_fu_223_p1;
wire tmp_6_fu_223_p3;
wire [7:0] tmp_9_fu_302_p1;
wire tmp_9_fu_302_p3;
wire [7:0] trunc_ln1192_fu_195_p0;
wire [6:0] trunc_ln1192_fu_195_p1;
wire [7:0] trunc_ln851_1_fu_249_p0;
wire [6:0] trunc_ln851_1_fu_249_p1;
wire [2:0] trunc_ln851_2_fu_565_p1;
wire [3:0] trunc_ln851_fu_435_p1;
wire xor_ln416_fu_275_p2;
wire xor_ln778_fu_280_p2;
wire xor_ln780_fu_309_p2;
wire xor_ln781_fu_329_p2;
wire xor_ln785_1_fu_392_p2;
wire xor_ln785_fu_382_p2;
wire [1:0] zext_ln831_fu_488_p1;


assign _046_ = _049_ & ap_CS_fsm[6];
assign _047_ = _050_ & ap_CS_fsm[0];
assign _048_ = ap_start & ap_CS_fsm[0];
assign and_ln781_1_fu_320_p2 = xor_ln416_reg_839 & Range2_all_ones_reg_800;
assign and_ln781_fu_324_p2 = p_Result_4_reg_789 & and_ln781_1_fu_320_p2;
assign and_ln785_1_fu_448_p2 = or_ln785_1_fu_443_p2 & and_ln786_reg_867;
assign and_ln785_fu_439_p2 = xor_ln416_reg_839 & deleted_zeros_reg_856;
assign and_ln786_1_fu_340_p2 = p_Result_5_reg_820 & or_ln780_fu_315_p2;
assign and_ln786_fu_345_p2 = and_ln786_1_fu_340_p2 & Range2_all_ones_reg_800;
assign neg_src_fu_335_p2 = xor_ln781_fu_329_p2 & p_Result_3_reg_771;
assign overflow_fu_397_p2 = xor_ln785_1_fu_392_p2 & or_ln785_fu_387_p2;
assign ret_V_23_fu_520_p2 = { op_6_V_reg_917[3], op_6_V_reg_917 } & { select_ln353_fu_506_p3, 3'h0 };
assign xor_ln780_fu_309_p2 = ~ op_2[7];
assign xor_ln781_fu_329_p2 = ~ and_ln781_fu_324_p2;
assign xor_ln785_fu_382_p2 = ~ deleted_zeros_reg_856;
assign xor_ln785_1_fu_392_p2 = ~ p_Result_3_reg_771;
assign xor_ln778_fu_280_p2 = ~ p_Result_4_reg_789;
assign ret_V_9_fu_483_p2 = ~ Range2_all_ones_reg_800;
assign xor_ln416_fu_275_p2 = ~ p_Result_5_reg_820;
assign _049_ = ~ icmp_ln851_reg_779;
assign _050_ = ~ ap_start;
assign _051_ = ! trunc_ln851_reg_912;
assign _052_ = ! op_2[6:0];
assign _053_ = ! trunc_ln851_2_reg_975;
always @(posedge \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.clk )
\add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.bin_s1  <= _055_;
always @(posedge \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.clk )
\add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.ain_s1  <= _054_;
always @(posedge \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.clk )
\add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.sum_s1  <= _057_;
always @(posedge \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.clk )
\add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.carry_s1  <= _056_;
assign _055_ = \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.ce  ? \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.b [12:6] : \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.bin_s1 ;
assign _054_ = \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.ce  ? \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.a [12:6] : \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.ain_s1 ;
assign _056_ = \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.ce  ? \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.facout_s1  : \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.carry_s1 ;
assign _057_ = \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.ce  ? \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.fas_s1  : \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.sum_s1 ;
assign _058_ = \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.u1.a  + \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.u1.b ;
assign { \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.u1.cout , \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.u1.s  } = _058_ + \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.u1.cin ;
assign _059_ = \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.u2.a  + \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.u2.b ;
assign { \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.u2.cout , \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.u2.s  } = _059_ + \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.u2.cin ;
always @(posedge \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.clk )
\add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.bin_s1  <= _061_;
always @(posedge \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.clk )
\add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.ain_s1  <= _060_;
always @(posedge \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.clk )
\add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.sum_s1  <= _063_;
always @(posedge \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.clk )
\add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.carry_s1  <= _062_;
assign _061_ = \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.ce  ? \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.b [13:7] : \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.bin_s1 ;
assign _060_ = \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.ce  ? \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.a [13:7] : \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.ain_s1 ;
assign _062_ = \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.ce  ? \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.facout_s1  : \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.carry_s1 ;
assign _063_ = \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.ce  ? \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.fas_s1  : \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.sum_s1 ;
assign _064_ = \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.u1.a  + \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.u1.b ;
assign { \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.u1.cout , \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.u1.s  } = _064_ + \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.u1.cin ;
assign _065_ = \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.u2.a  + \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.u2.b ;
assign { \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.u2.cout , \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.u2.s  } = _065_ + \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.u2.cin ;
always @(posedge \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.clk )
\add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.bin_s1  <= _067_;
always @(posedge \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.clk )
\add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.ain_s1  <= _066_;
always @(posedge \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.clk )
\add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.sum_s1  <= _069_;
always @(posedge \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.clk )
\add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.carry_s1  <= _068_;
assign _067_ = \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.ce  ? \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.b [13:7] : \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.bin_s1 ;
assign _066_ = \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.ce  ? \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.a [13:7] : \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.ain_s1 ;
assign _068_ = \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.ce  ? \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.facout_s1  : \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.carry_s1 ;
assign _069_ = \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.ce  ? \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.fas_s1  : \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.sum_s1 ;
assign _070_ = \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.u1.a  + \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.u1.b ;
assign { \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.u1.cout , \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.u1.s  } = _070_ + \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.u1.cin ;
assign _071_ = \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.u2.a  + \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.u2.b ;
assign { \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.u2.cout , \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.u2.s  } = _071_ + \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.u2.cin ;
always @(posedge \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.clk )
\add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.bin_s1  <= _073_;
always @(posedge \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.clk )
\add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.ain_s1  <= _072_;
always @(posedge \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.clk )
\add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.sum_s1  <= _075_;
always @(posedge \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.clk )
\add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.carry_s1  <= _074_;
assign _073_ = \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.ce  ? \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.b [13:7] : \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.bin_s1 ;
assign _072_ = \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.ce  ? \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.a [13:7] : \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.ain_s1 ;
assign _074_ = \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.ce  ? \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.facout_s1  : \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.carry_s1 ;
assign _075_ = \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.ce  ? \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.fas_s1  : \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.sum_s1 ;
assign _076_ = \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.u1.a  + \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.u1.b ;
assign { \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.u1.cout , \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.u1.s  } = _076_ + \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.u1.cin ;
assign _077_ = \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.u2.a  + \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.u2.b ;
assign { \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.u2.cout , \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.u2.s  } = _077_ + \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.u2.cin ;
always @(posedge \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.clk )
\add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.bin_s1  <= _079_;
always @(posedge \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.clk )
\add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.ain_s1  <= _078_;
always @(posedge \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.clk )
\add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.sum_s1  <= _081_;
always @(posedge \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.clk )
\add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.carry_s1  <= _080_;
assign _079_ = \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.ce  ? \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.b [14:7] : \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.bin_s1 ;
assign _078_ = \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.ce  ? \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.a [14:7] : \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.ain_s1 ;
assign _080_ = \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.ce  ? \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.facout_s1  : \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.carry_s1 ;
assign _081_ = \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.ce  ? \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.fas_s1  : \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.sum_s1 ;
assign _082_ = \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.u1.a  + \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.u1.b ;
assign { \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.u1.cout , \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.u1.s  } = _082_ + \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.u1.cin ;
assign _083_ = \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.u2.a  + \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.u2.b ;
assign { \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.u2.cout , \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.u2.s  } = _083_ + \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.u2.cin ;
always @(posedge \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.clk )
\add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.bin_s1  <= _085_;
always @(posedge \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.clk )
\add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.ain_s1  <= _084_;
always @(posedge \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.clk )
\add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.sum_s1  <= _087_;
always @(posedge \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.clk )
\add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.carry_s1  <= _086_;
assign _085_ = \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.ce  ? \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.b [14:7] : \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.bin_s1 ;
assign _084_ = \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.ce  ? \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.a [14:7] : \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.ain_s1 ;
assign _086_ = \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.ce  ? \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.facout_s1  : \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.carry_s1 ;
assign _087_ = \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.ce  ? \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.fas_s1  : \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.sum_s1 ;
assign _088_ = \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.u1.a  + \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.u1.b ;
assign { \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.u1.cout , \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.u1.s  } = _088_ + \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.u1.cin ;
assign _089_ = \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.u2.a  + \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.u2.b ;
assign { \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.u2.cout , \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.u2.s  } = _089_ + \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.u2.cin ;
always @(posedge \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.clk )
\add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.bin_s1  <= _091_;
always @(posedge \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.clk )
\add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.ain_s1  <= _090_;
always @(posedge \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.clk )
\add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.sum_s1  <= _093_;
always @(posedge \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.clk )
\add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.carry_s1  <= _092_;
assign _091_ = \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.ce  ? \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.b [16:8] : \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.bin_s1 ;
assign _090_ = \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.ce  ? \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.a [16:8] : \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.ain_s1 ;
assign _092_ = \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.ce  ? \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.facout_s1  : \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.carry_s1 ;
assign _093_ = \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.ce  ? \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.fas_s1  : \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.sum_s1 ;
assign _094_ = \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.u1.a  + \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.u1.b ;
assign { \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.u1.cout , \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.u1.s  } = _094_ + \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.u1.cin ;
assign _095_ = \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.u2.a  + \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.u2.b ;
assign { \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.u2.cout , \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.u2.s  } = _095_ + \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.u2.cin ;
always @(posedge \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.clk )
\add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.bin_s1  <= _097_;
always @(posedge \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.clk )
\add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.ain_s1  <= _096_;
always @(posedge \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.clk )
\add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.sum_s1  <= _099_;
always @(posedge \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.clk )
\add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.carry_s1  <= _098_;
assign _097_ = \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.ce  ? \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.b [17:9] : \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.bin_s1 ;
assign _096_ = \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.ce  ? \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.a [17:9] : \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.ain_s1 ;
assign _098_ = \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.ce  ? \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.facout_s1  : \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.carry_s1 ;
assign _099_ = \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.ce  ? \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.fas_s1  : \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.sum_s1 ;
assign _100_ = \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.u1.a  + \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.u1.b ;
assign { \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.u1.cout , \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.u1.s  } = _100_ + \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.u1.cin ;
assign _101_ = \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.u2.a  + \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.u2.b ;
assign { \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.u2.cout , \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.u2.s  } = _101_ + \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.u2.cin ;
always @(posedge \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.clk )
\add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.bin_s1  <= _103_;
always @(posedge \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.clk )
\add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.ain_s1  <= _102_;
always @(posedge \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.clk )
\add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.sum_s1  <= _105_;
always @(posedge \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.clk )
\add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.carry_s1  <= _104_;
assign _103_ = \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.ce  ? \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.b [17:9] : \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.bin_s1 ;
assign _102_ = \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.ce  ? \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.a [17:9] : \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.ain_s1 ;
assign _104_ = \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.ce  ? \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.facout_s1  : \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.carry_s1 ;
assign _105_ = \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.ce  ? \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.fas_s1  : \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.sum_s1 ;
assign _106_ = \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.u1.a  + \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.u1.b ;
assign { \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.u1.cout , \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.u1.s  } = _106_ + \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.u1.cin ;
assign _107_ = \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.u2.a  + \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.u2.b ;
assign { \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.u2.cout , \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.u2.s  } = _107_ + \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.u2.cin ;
always @(posedge \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.clk )
\add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.bin_s1  <= _109_;
always @(posedge \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.clk )
\add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.ain_s1  <= _108_;
always @(posedge \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.clk )
\add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.sum_s1  <= _111_;
always @(posedge \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.clk )
\add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.carry_s1  <= _110_;
assign _109_ = \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.ce  ? \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.b [1] : \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.bin_s1 ;
assign _108_ = \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.ce  ? \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.a [1] : \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.ain_s1 ;
assign _110_ = \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.ce  ? \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.facout_s1  : \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.carry_s1 ;
assign _111_ = \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.ce  ? \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.fas_s1  : \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.sum_s1 ;
assign _112_ = \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.u1.a  + \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.u1.b ;
assign { \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.u1.cout , \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.u1.s  } = _112_ + \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.u1.cin ;
assign _113_ = \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.u2.a  + \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.u2.b ;
assign { \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.u2.cout , \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.u2.s  } = _113_ + \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.u2.cin ;
always @(posedge \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.clk )
\add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.bin_s1  <= _115_;
always @(posedge \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.clk )
\add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.ain_s1  <= _114_;
always @(posedge \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.clk )
\add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.sum_s1  <= _117_;
always @(posedge \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.clk )
\add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.carry_s1  <= _116_;
assign _115_ = \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.ce  ? \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.b [1] : \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.bin_s1 ;
assign _114_ = \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.ce  ? \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.a [1] : \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.ain_s1 ;
assign _116_ = \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.ce  ? \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.facout_s1  : \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.carry_s1 ;
assign _117_ = \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.ce  ? \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.fas_s1  : \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.sum_s1 ;
assign _118_ = \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.u1.a  + \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.u1.b ;
assign { \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.u1.cout , \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.u1.s  } = _118_ + \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.u1.cin ;
assign _119_ = \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.u2.a  + \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.u2.b ;
assign { \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.u2.cout , \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.u2.s  } = _119_ + \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.u2.cin ;
always @(posedge \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.clk )
\add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.bin_s1  <= _121_;
always @(posedge \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.clk )
\add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.ain_s1  <= _120_;
always @(posedge \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.clk )
\add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.sum_s1  <= _123_;
always @(posedge \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.clk )
\add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.carry_s1  <= _122_;
assign _121_ = \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.ce  ? \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.b [2:1] : \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.bin_s1 ;
assign _120_ = \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.ce  ? \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.a [2:1] : \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.ain_s1 ;
assign _122_ = \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.ce  ? \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.facout_s1  : \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.carry_s1 ;
assign _123_ = \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.ce  ? \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.fas_s1  : \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.sum_s1 ;
assign _124_ = \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.u1.a  + \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.u1.b ;
assign { \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.u1.cout , \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.u1.s  } = _124_ + \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.u1.cin ;
assign _125_ = \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.u2.a  + \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.u2.b ;
assign { \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.u2.cout , \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.u2.s  } = _125_ + \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.u2.cin ;
always @(posedge \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.clk )
\add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.bin_s1  <= _127_;
always @(posedge \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.clk )
\add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.ain_s1  <= _126_;
always @(posedge \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.clk )
\add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.sum_s1  <= _129_;
always @(posedge \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.clk )
\add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.carry_s1  <= _128_;
assign _127_ = \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.ce  ? \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.b [3:2] : \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.bin_s1 ;
assign _126_ = \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.ce  ? \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.a [3:2] : \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.ain_s1 ;
assign _128_ = \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.ce  ? \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.facout_s1  : \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.carry_s1 ;
assign _129_ = \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.ce  ? \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.fas_s1  : \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.sum_s1 ;
assign _130_ = \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.u1.a  + \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.u1.b ;
assign { \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.u1.cout , \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.u1.s  } = _130_ + \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.u1.cin ;
assign _131_ = \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.u2.a  + \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.u2.b ;
assign { \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.u2.cout , \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.u2.s  } = _131_ + \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.u2.cin ;
always @(posedge \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.clk )
\add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.bin_s1  <= _133_;
always @(posedge \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.clk )
\add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.ain_s1  <= _132_;
always @(posedge \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.clk )
\add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.sum_s1  <= _135_;
always @(posedge \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.clk )
\add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.carry_s1  <= _134_;
assign _133_ = \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.ce  ? \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.b [3:2] : \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.bin_s1 ;
assign _132_ = \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.ce  ? \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.a [3:2] : \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.ain_s1 ;
assign _134_ = \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.ce  ? \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.facout_s1  : \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.carry_s1 ;
assign _135_ = \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.ce  ? \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.fas_s1  : \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.sum_s1 ;
assign _136_ = \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.u1.a  + \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.u1.b ;
assign { \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.u1.cout , \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.u1.s  } = _136_ + \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.u1.cin ;
assign _137_ = \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.u2.a  + \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.u2.b ;
assign { \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.u2.cout , \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.u2.s  } = _137_ + \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.u2.cin ;
always @(posedge \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.clk )
\add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.bin_s1  <= _139_;
always @(posedge \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.clk )
\add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.ain_s1  <= _138_;
always @(posedge \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.clk )
\add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.sum_s1  <= _141_;
always @(posedge \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.clk )
\add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.carry_s1  <= _140_;
assign _139_ = \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.ce  ? \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.b [4:2] : \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.bin_s1 ;
assign _138_ = \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.ce  ? \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.a [4:2] : \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.ain_s1 ;
assign _140_ = \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.ce  ? \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.facout_s1  : \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.carry_s1 ;
assign _141_ = \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.ce  ? \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.fas_s1  : \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.sum_s1 ;
assign _142_ = \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.u1.a  + \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.u1.b ;
assign { \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.u1.cout , \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.u1.s  } = _142_ + \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.u1.cin ;
assign _143_ = \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.u2.a  + \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.u2.b ;
assign { \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.u2.cout , \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.u2.s  } = _143_ + \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.u2.cin ;
always @(posedge \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.clk )
\add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.bin_s1  <= _145_;
always @(posedge \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.clk )
\add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.ain_s1  <= _144_;
always @(posedge \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.clk )
\add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.sum_s1  <= _147_;
always @(posedge \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.clk )
\add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.carry_s1  <= _146_;
assign _145_ = \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.ce  ? \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.b [8:4] : \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.bin_s1 ;
assign _144_ = \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.ce  ? \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.a [8:4] : \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.ain_s1 ;
assign _146_ = \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.ce  ? \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.facout_s1  : \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.carry_s1 ;
assign _147_ = \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.ce  ? \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.fas_s1  : \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.sum_s1 ;
assign _148_ = \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.u1.a  + \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.u1.b ;
assign { \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.u1.cout , \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.u1.s  } = _148_ + \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.u1.cin ;
assign _149_ = \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.u2.a  + \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.u2.b ;
assign { \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.u2.cout , \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.u2.s  } = _149_ + \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.u2.cin ;
assign \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.bin_s0  = ~ \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.b ;
always @(posedge \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.clk )
\sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.bin_s1  <= _151_;
always @(posedge \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.clk )
\sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.ain_s1  <= _150_;
always @(posedge \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.clk )
\sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.sum_s1  <= _153_;
always @(posedge \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.clk )
\sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.carry_s1  <= _152_;
assign _151_ = \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.ce  ? \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.bin_s0 [4:2] : \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.bin_s1 ;
assign _150_ = \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.ce  ? \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.a [4:2] : \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.ain_s1 ;
assign _152_ = \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.ce  ? \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.facout_s1  : \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.carry_s1 ;
assign _153_ = \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.ce  ? \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.fas_s1  : \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.sum_s1 ;
assign _154_ = \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.u1.a  + \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.u1.b ;
assign { \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.u1.cout , \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.u1.s  } = _154_ + \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.u1.cin ;
assign _155_ = \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.u2.a  + \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.u2.b ;
assign { \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.u2.cout , \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.u2.s  } = _155_ + \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.u2.cin ;
assign or_ln340_1_fu_408_p2 = or_ln340_fu_403_p2 | neg_src_reg_862;
assign or_ln340_fu_403_p2 = overflow_fu_397_p2 | and_ln786_reg_867;
assign or_ln778_fu_285_p2 = xor_ln778_fu_280_p2 | p_Result_5_reg_820;
assign or_ln780_fu_315_p2 = xor_ln780_fu_309_p2 | or_ln778_reg_845;
assign or_ln785_1_fu_443_p2 = p_Result_3_reg_771 | and_ln785_fu_439_p2;
assign or_ln785_fu_387_p2 = xor_ln785_fu_382_p2 | p_Result_5_reg_820;
always @(posedge ap_clk)
select_ln1192_reg_834[6:0] <= 7'h00;
always @(posedge ap_clk)
select_ln703_reg_928[2:0] <= 3'h0;
always @(posedge ap_clk)
select_ln69_reg_1020[13:8] <= 6'h00;
always @(posedge ap_clk)
ret_V_2_reg_933 <= _032_;
always @(posedge ap_clk)
ret_V_24_reg_1090 <= _031_;
always @(posedge ap_clk)
ret_V_17_reg_873 <= _025_;
always @(posedge ap_clk)
ret_V_reg_878 <= _035_;
always @(posedge ap_clk)
select_ln340_reg_895 <= _037_;
always @(posedge ap_clk)
ret_V_12_reg_995 <= _024_;
always @(posedge ap_clk)
ret_V_18_reg_953 <= _026_;
always @(posedge ap_clk)
ret_V_6_reg_958 <= _034_;
always @(posedge ap_clk)
ret_V_21_reg_963 <= _029_;
always @(posedge ap_clk)
ret_V_11_reg_968 <= _023_;
always @(posedge ap_clk)
trunc_ln851_2_reg_975 <= _042_;
always @(posedge ap_clk)
p_Val2_3_reg_814 <= _022_;
always @(posedge ap_clk)
p_Result_5_reg_820 <= _021_;
always @(posedge ap_clk)
select_ln1192_reg_834[8:7] <= _036_;
always @(posedge ap_clk)
xor_ln416_reg_839 <= _044_;
always @(posedge ap_clk)
or_ln778_reg_845 <= _018_;
always @(posedge ap_clk)
ret_V_19_reg_900 <= _027_;
always @(posedge ap_clk)
ret_V_4_reg_905 <= _033_;
always @(posedge ap_clk)
trunc_ln851_reg_912 <= _043_;
always @(posedge ap_clk)
op_6_V_reg_917 <= _017_;
always @(posedge ap_clk)
select_ln831_reg_922 <= _040_;
always @(posedge ap_clk)
select_ln703_reg_928[4:3] <= _039_;
always @(posedge ap_clk)
op_26_V_reg_1075 <= _016_;
always @(posedge ap_clk)
op_25_V_reg_1060 <= _015_;
always @(posedge ap_clk)
ret_V_20_reg_980 <= _028_;
always @(posedge ap_clk)
icmp_ln851_3_reg_985 <= _012_;
always @(posedge ap_clk)
icmp_ln851_1_reg_938 <= _010_;
always @(posedge ap_clk)
tmp_reg_948 <= _041_;
always @(posedge ap_clk)
deleted_zeros_reg_856 <= _009_;
always @(posedge ap_clk)
neg_src_reg_862 <= _014_;
always @(posedge ap_clk)
and_ln786_reg_867 <= _007_;
always @(posedge ap_clk)
add_ln69_5_reg_1115 <= _004_;
always @(posedge ap_clk)
add_ln69_7_reg_1120 <= _005_;
always @(posedge ap_clk)
ret_V_22_reg_1015 <= _030_;
always @(posedge ap_clk)
select_ln69_reg_1020[7:0] <= _038_;
always @(posedge ap_clk)
add_ln69_reg_1025 <= _006_;
always @(posedge ap_clk)
add_ln69_2_reg_1030 <= _002_;
always @(posedge ap_clk)
add_ln69_1_reg_1045 <= _001_;
always @(posedge ap_clk)
add_ln69_3_reg_1050 <= _003_;
always @(posedge ap_clk)
p_Result_3_reg_771 <= _019_;
always @(posedge ap_clk)
icmp_ln851_reg_779 <= _013_;
always @(posedge ap_clk)
p_Result_4_reg_789 <= _020_;
always @(posedge ap_clk)
Range2_all_ones_reg_800 <= _000_;
always @(posedge ap_clk)
icmp_ln851_2_reg_809 <= _011_;
always @(posedge ap_clk)
ap_CS_fsm <= _008_;
assign _045_ = _048_ ? 2'h2 : 2'h1;
assign _156_ = ap_CS_fsm == 1'h1;
function [22:0] _464_;
input [22:0] a;
input [528:0] b;
input [22:0] s;
case (s)
23'b00000000000000000000001:
_464_ = b[22:0];
23'b00000000000000000000010:
_464_ = b[45:23];
23'b00000000000000000000100:
_464_ = b[68:46];
23'b00000000000000000001000:
_464_ = b[91:69];
23'b00000000000000000010000:
_464_ = b[114:92];
23'b00000000000000000100000:
_464_ = b[137:115];
23'b00000000000000001000000:
_464_ = b[160:138];
23'b00000000000000010000000:
_464_ = b[183:161];
23'b00000000000000100000000:
_464_ = b[206:184];
23'b00000000000001000000000:
_464_ = b[229:207];
23'b00000000000010000000000:
_464_ = b[252:230];
23'b00000000000100000000000:
_464_ = b[275:253];
23'b00000000001000000000000:
_464_ = b[298:276];
23'b00000000010000000000000:
_464_ = b[321:299];
23'b00000000100000000000000:
_464_ = b[344:322];
23'b00000001000000000000000:
_464_ = b[367:345];
23'b00000010000000000000000:
_464_ = b[390:368];
23'b00000100000000000000000:
_464_ = b[413:391];
23'b00001000000000000000000:
_464_ = b[436:414];
23'b00010000000000000000000:
_464_ = b[459:437];
23'b00100000000000000000000:
_464_ = b[482:460];
23'b01000000000000000000000:
_464_ = b[505:483];
23'b10000000000000000000000:
_464_ = b[528:506];
23'b00000000000000000000000:
_464_ = a;
default:
_464_ = 23'bx;
endcase
endfunction
assign ap_NS_fsm = _464_(23'hxxxxxx, { 21'h000000, _045_, 506'h0000020000080000200000800002000008000020000080000200000800002000008000020000080000200000800002000008000020000080000200000000001 }, { _156_, _178_, _177_, _176_, _175_, _174_, _173_, _172_, _171_, _170_, _169_, _168_, _167_, _166_, _165_, _164_, _163_, _162_, _161_, _160_, _159_, _158_, _157_ });
assign _157_ = ap_CS_fsm == 23'h400000;
assign _158_ = ap_CS_fsm == 22'h200000;
assign _159_ = ap_CS_fsm == 21'h100000;
assign _160_ = ap_CS_fsm == 20'h80000;
assign _161_ = ap_CS_fsm == 19'h40000;
assign _162_ = ap_CS_fsm == 18'h20000;
assign _163_ = ap_CS_fsm == 17'h10000;
assign _164_ = ap_CS_fsm == 16'h8000;
assign _165_ = ap_CS_fsm == 15'h4000;
assign _166_ = ap_CS_fsm == 14'h2000;
assign _167_ = ap_CS_fsm == 13'h1000;
assign _168_ = ap_CS_fsm == 12'h800;
assign _169_ = ap_CS_fsm == 11'h400;
assign _170_ = ap_CS_fsm == 10'h200;
assign _171_ = ap_CS_fsm == 9'h100;
assign _172_ = ap_CS_fsm == 8'h80;
assign _173_ = ap_CS_fsm == 7'h40;
assign _174_ = ap_CS_fsm == 6'h20;
assign _175_ = ap_CS_fsm == 5'h10;
assign _176_ = ap_CS_fsm == 4'h8;
assign _177_ = ap_CS_fsm == 3'h4;
assign _178_ = ap_CS_fsm == 2'h2;
assign op_30_ap_vld = ap_CS_fsm[22] ? 1'h1 : 1'h0;
assign ap_idle = _047_ ? 1'h1 : 1'h0;
assign _032_ = _046_ ? grp_fu_420_p2 : ret_V_2_reg_933;
assign _031_ = ap_CS_fsm[18] ? grp_fu_717_p2 : ret_V_24_reg_1090;
assign _037_ = ap_CS_fsm[4] ? select_ln340_fu_413_p3 : select_ln340_reg_895;
assign _035_ = ap_CS_fsm[4] ? grp_fu_293_p2[8:7] : ret_V_reg_878;
assign _025_ = ap_CS_fsm[4] ? grp_fu_293_p2 : ret_V_17_reg_873;
assign _024_ = ap_CS_fsm[9] ? grp_fu_593_p2 : ret_V_12_reg_995;
assign _042_ = ap_CS_fsm[7] ? grp_fu_495_p2[2:0] : trunc_ln851_2_reg_975;
assign _023_ = ap_CS_fsm[7] ? grp_fu_495_p2[4:3] : ret_V_11_reg_968;
assign _029_ = ap_CS_fsm[7] ? grp_fu_495_p2 : ret_V_21_reg_963;
assign _034_ = ap_CS_fsm[7] ? grp_fu_478_p2 : ret_V_6_reg_958;
assign _026_ = ap_CS_fsm[7] ? ret_V_18_fu_548_p3 : ret_V_18_reg_953;
assign _021_ = ap_CS_fsm[1] ? grp_fu_235_p2[3] : p_Result_5_reg_820;
assign _022_ = ap_CS_fsm[1] ? grp_fu_235_p2 : p_Val2_3_reg_814;
assign _018_ = ap_CS_fsm[2] ? or_ln778_fu_285_p2 : or_ln778_reg_845;
assign _044_ = ap_CS_fsm[2] ? xor_ln416_fu_275_p2 : xor_ln416_reg_839;
assign _036_ = ap_CS_fsm[2] ? select_ln1192_fu_267_p3[8:7] : select_ln1192_reg_834[8:7];
assign _039_ = ap_CS_fsm[5] ? select_ln703_fu_466_p3[4:3] : select_ln703_reg_928[4:3];
assign _040_ = ap_CS_fsm[5] ? select_ln831_fu_459_p3 : select_ln831_reg_922;
assign _017_ = ap_CS_fsm[5] ? op_6_V_fu_453_p3 : op_6_V_reg_917;
assign _043_ = ap_CS_fsm[5] ? grp_fu_376_p2[3:0] : trunc_ln851_reg_912;
assign _033_ = ap_CS_fsm[5] ? grp_fu_376_p2[16:4] : ret_V_4_reg_905;
assign _027_ = ap_CS_fsm[5] ? grp_fu_376_p2 : ret_V_19_reg_900;
assign _016_ = ap_CS_fsm[16] ? grp_fu_694_p2[14:1] : op_26_V_reg_1075;
assign _015_ = ap_CS_fsm[14] ? grp_fu_670_p2 : op_25_V_reg_1060;
assign _012_ = ap_CS_fsm[8] ? icmp_ln851_3_fu_588_p2 : icmp_ln851_3_reg_985;
assign _028_ = ap_CS_fsm[8] ? ret_V_20_fu_581_p3 : ret_V_20_reg_980;
assign _041_ = ap_CS_fsm[6] ? ret_V_23_fu_520_p2[4:3] : tmp_reg_948;
assign _010_ = ap_CS_fsm[6] ? icmp_ln851_1_fu_473_p2 : icmp_ln851_1_reg_938;
assign _007_ = ap_CS_fsm[3] ? and_ln786_fu_345_p2 : and_ln786_reg_867;
assign _014_ = ap_CS_fsm[3] ? neg_src_fu_335_p2 : neg_src_reg_862;
assign _009_ = ap_CS_fsm[3] ? deleted_zeros_fu_298_p2 : deleted_zeros_reg_856;
assign _005_ = ap_CS_fsm[20] ? grp_fu_746_p2 : add_ln69_7_reg_1120;
assign _004_ = ap_CS_fsm[20] ? grp_fu_740_p2 : add_ln69_5_reg_1115;
assign _002_ = ap_CS_fsm[10] ? grp_fu_619_p2 : add_ln69_2_reg_1030;
assign _006_ = ap_CS_fsm[10] ? grp_fu_613_p2 : add_ln69_reg_1025;
assign _038_ = ap_CS_fsm[10] ? select_ln69_fu_644_p3 : select_ln69_reg_1020[7:0];
assign _030_ = ap_CS_fsm[10] ? ret_V_22_fu_637_p3 : ret_V_22_reg_1015;
assign _003_ = ap_CS_fsm[12] ? grp_fu_661_p2 : add_ln69_3_reg_1050;
assign _001_ = ap_CS_fsm[12] ? grp_fu_654_p2 : add_ln69_1_reg_1045;
assign _011_ = ap_CS_fsm[0] ? icmp_ln851_2_fu_253_p2 : icmp_ln851_2_reg_809;
assign _000_ = ap_CS_fsm[0] ? op_2[7] : Range2_all_ones_reg_800;
assign _020_ = ap_CS_fsm[0] ? op_2[7] : p_Result_4_reg_789;
assign _013_ = ap_CS_fsm[0] ? icmp_ln851_2_fu_253_p2 : icmp_ln851_reg_779;
assign _019_ = ap_CS_fsm[0] ? op_2[7] : p_Result_3_reg_771;
assign _008_ = ap_rst ? 23'h000001 : ap_NS_fsm;
assign icmp_ln851_1_fu_473_p2 = _051_ ? 1'h1 : 1'h0;
assign icmp_ln851_2_fu_253_p2 = _052_ ? 1'h1 : 1'h0;
assign icmp_ln851_3_fu_588_p2 = _053_ ? 1'h1 : 1'h0;
assign op_6_V_fu_453_p3 = and_ln785_1_fu_448_p2 ? p_Val2_3_reg_814 : select_ln340_reg_895;
assign ret_V_18_fu_548_p3 = ret_V_17_reg_873[8] ? select_ln850_fu_543_p3 : ret_V_reg_878;
assign ret_V_20_fu_581_p3 = ret_V_19_reg_900[16] ? select_ln850_1_fu_576_p3 : ret_V_4_reg_905;
assign ret_V_22_fu_637_p3 = ret_V_21_reg_963[4] ? select_ln850_3_fu_632_p3 : ret_V_11_reg_968;
assign select_ln1192_fu_267_p3 = op_3 ? 9'h180 : 9'h000;
assign select_ln340_fu_413_p3 = or_ln340_1_fu_408_p2 ? 4'h0 : p_Val2_3_reg_814;
assign select_ln353_fu_506_p3 = p_Result_3_reg_771 ? select_ln850_6_fu_500_p3 : select_ln831_reg_922;
assign select_ln69_fu_644_p3 = op_3 ? 8'hff : 8'h00;
assign select_ln703_fu_466_p3 = op_3 ? 5'h18 : 5'h00;
assign select_ln831_fu_459_p3 = Range2_all_ones_reg_800 ? 2'h3 : 2'h0;
assign select_ln850_1_fu_576_p3 = icmp_ln851_1_reg_938 ? ret_V_4_reg_905 : ret_V_6_reg_958;
assign select_ln850_3_fu_632_p3 = icmp_ln851_3_reg_985 ? ret_V_11_reg_968 : ret_V_12_reg_995;
assign select_ln850_6_fu_500_p3 = icmp_ln851_2_reg_809 ? select_ln831_reg_922 : { 1'h0, ret_V_9_fu_483_p2 };
assign select_ln850_fu_543_p3 = icmp_ln851_reg_779 ? ret_V_reg_878 : ret_V_2_reg_933;
assign deleted_zeros_fu_298_p2 = or_ln778_reg_845 ^ Range2_all_ones_reg_800;
assign Range2_all_ones_fu_241_p1 = op_2;
assign ap_CS_fsm_state1 = ap_CS_fsm[0];
assign ap_CS_fsm_state10 = ap_CS_fsm[9];
assign ap_CS_fsm_state11 = ap_CS_fsm[10];
assign ap_CS_fsm_state12 = ap_CS_fsm[11];
assign ap_CS_fsm_state13 = ap_CS_fsm[12];
assign ap_CS_fsm_state14 = ap_CS_fsm[13];
assign ap_CS_fsm_state15 = ap_CS_fsm[14];
assign ap_CS_fsm_state16 = ap_CS_fsm[15];
assign ap_CS_fsm_state17 = ap_CS_fsm[16];
assign ap_CS_fsm_state18 = ap_CS_fsm[17];
assign ap_CS_fsm_state19 = ap_CS_fsm[18];
assign ap_CS_fsm_state2 = ap_CS_fsm[1];
assign ap_CS_fsm_state20 = ap_CS_fsm[19];
assign ap_CS_fsm_state21 = ap_CS_fsm[20];
assign ap_CS_fsm_state22 = ap_CS_fsm[21];
assign ap_CS_fsm_state23 = ap_CS_fsm[22];
assign ap_CS_fsm_state3 = ap_CS_fsm[2];
assign ap_CS_fsm_state4 = ap_CS_fsm[3];
assign ap_CS_fsm_state5 = ap_CS_fsm[4];
assign ap_CS_fsm_state6 = ap_CS_fsm[5];
assign ap_CS_fsm_state7 = ap_CS_fsm[6];
assign ap_CS_fsm_state8 = ap_CS_fsm[7];
assign ap_CS_fsm_state9 = ap_CS_fsm[8];
assign ap_done = op_30_ap_vld;
assign ap_ready = op_30_ap_vld;
assign grp_fu_235_p0 = { 3'h0, op_2[3] };
assign grp_fu_235_p1 = op_2[7:4];
assign grp_fu_293_p1 = { op_2[7], op_2 };
assign grp_fu_376_p0 = { op_9[3], op_9[3], op_9[3], op_9[3], op_9[3], op_9[3], op_9[3], op_9[3], op_9[3], op_9[3], op_9[3], op_9[3], op_9, 1'h0 };
assign grp_fu_376_p1 = { op_0[15], op_0 };
assign grp_fu_613_p0 = { ret_V_20_reg_980[12], ret_V_20_reg_980 };
assign grp_fu_613_p1 = { 10'h000, op_12 };
assign grp_fu_619_p0 = { 1'h0, op_14 };
assign grp_fu_619_p1 = { 2'h0, op_13 };
assign grp_fu_661_p0 = { 1'h0, add_ln69_2_reg_1030 };
assign grp_fu_661_p1 = { ret_V_22_reg_1015[1], ret_V_22_reg_1015[1], ret_V_22_reg_1015 };
assign grp_fu_670_p0 = { add_ln69_3_reg_1050[3], add_ln69_3_reg_1050[3], add_ln69_3_reg_1050[3], add_ln69_3_reg_1050[3], add_ln69_3_reg_1050[3], add_ln69_3_reg_1050[3], add_ln69_3_reg_1050[3], add_ln69_3_reg_1050[3], add_ln69_3_reg_1050[3], add_ln69_3_reg_1050[3], add_ln69_3_reg_1050 };
assign grp_fu_694_p0 = { op_25_V_reg_1060, 1'h0 };
assign grp_fu_694_p1 = { op_1, op_1, op_1, op_1, op_1, op_1, op_1, op_1, op_1, op_1, op_1, op_1, op_1, op_1, 1'h0 };
assign grp_fu_717_p0 = { op_26_V_reg_1075[13], op_26_V_reg_1075 };
assign grp_fu_717_p1 = { op_16[1], op_16[1], op_16[1], op_16[1], op_16[1], op_16[1], op_16[1], op_16[1], op_16[1], op_16[1], op_16[1], op_16[1], op_16[1], op_16 };
assign grp_fu_740_p0 = { ret_V_24_reg_1090[14], ret_V_24_reg_1090[14], ret_V_24_reg_1090[14], ret_V_24_reg_1090 };
assign grp_fu_740_p1 = { 2'h0, ret_V_18_reg_953[1], ret_V_18_reg_953[1], ret_V_18_reg_953[1], ret_V_18_reg_953[1], ret_V_18_reg_953[1], ret_V_18_reg_953[1], ret_V_18_reg_953[1], ret_V_18_reg_953[1], ret_V_18_reg_953[1], ret_V_18_reg_953[1], ret_V_18_reg_953[1], ret_V_18_reg_953[1], ret_V_18_reg_953[1], ret_V_18_reg_953[1], ret_V_18_reg_953 };
assign grp_fu_746_p0 = { op_17[3], op_17 };
assign grp_fu_746_p1 = { 3'h0, tmp_reg_948 };
assign grp_fu_755_p0 = { add_ln69_7_reg_1120[4], add_ln69_7_reg_1120[4], add_ln69_7_reg_1120[4], add_ln69_7_reg_1120[4], add_ln69_7_reg_1120[4], add_ln69_7_reg_1120[4], add_ln69_7_reg_1120[4], add_ln69_7_reg_1120[4], add_ln69_7_reg_1120[4], add_ln69_7_reg_1120[4], add_ln69_7_reg_1120[4], add_ln69_7_reg_1120[4], add_ln69_7_reg_1120[4], add_ln69_7_reg_1120 };
assign icmp_ln851_fu_199_p2 = icmp_ln851_2_fu_253_p2;
assign op_30 = { grp_fu_755_p2[17], grp_fu_755_p2[17], grp_fu_755_p2[17], grp_fu_755_p2[17], grp_fu_755_p2[17], grp_fu_755_p2[17], grp_fu_755_p2[17], grp_fu_755_p2[17], grp_fu_755_p2[17], grp_fu_755_p2[17], grp_fu_755_p2[17], grp_fu_755_p2[17], grp_fu_755_p2[17], grp_fu_755_p2[17], grp_fu_755_p2 };
assign p_Result_1_fu_536_p3 = ret_V_17_reg_873[8];
assign p_Result_2_fu_569_p3 = ret_V_19_reg_900[16];
assign p_Result_3_fu_187_p1 = op_2;
assign p_Result_4_fu_215_p1 = op_2;
assign p_Result_s_fu_625_p3 = ret_V_21_reg_963[4];
assign p_Val2_2_fu_205_p1 = op_2;
assign p_Val2_s_fu_675_p1 = op_1;
assign p_Val2_s_fu_675_p3 = { op_1, 1'h0 };
assign rhs_2_fu_512_p3 = { select_ln353_fu_506_p3, 3'h0 };
assign rhs_fu_364_p3 = { op_9, 1'h0 };
assign select_ln1192_fu_267_p0 = op_3;
assign select_ln69_fu_644_p0 = op_3;
assign select_ln703_fu_466_p0 = op_3;
assign sext_ln69_2_fu_730_p1 = { ret_V_18_reg_953[1], ret_V_18_reg_953[1], ret_V_18_reg_953[1], ret_V_18_reg_953[1], ret_V_18_reg_953[1], ret_V_18_reg_953[1], ret_V_18_reg_953[1], ret_V_18_reg_953[1], ret_V_18_reg_953[1], ret_V_18_reg_953[1], ret_V_18_reg_953[1], ret_V_18_reg_953[1], ret_V_18_reg_953[1], ret_V_18_reg_953[1], ret_V_18_reg_953 };
assign sext_ln703_2_fu_492_p1 = { op_6_V_reg_917[3], op_6_V_reg_917 };
assign sext_ln703_fu_290_p0 = op_2;
assign tmp_6_fu_223_p1 = op_2;
assign tmp_6_fu_223_p3 = op_2[3];
assign tmp_9_fu_302_p1 = op_2;
assign tmp_9_fu_302_p3 = op_2[7];
assign trunc_ln1192_fu_195_p0 = op_2;
assign trunc_ln1192_fu_195_p1 = op_2[6:0];
assign trunc_ln851_1_fu_249_p0 = op_2;
assign trunc_ln851_1_fu_249_p1 = op_2[6:0];
assign trunc_ln851_2_fu_565_p1 = grp_fu_495_p2[2:0];
assign trunc_ln851_fu_435_p1 = grp_fu_376_p2[3:0];
assign zext_ln831_fu_488_p1 = { 1'h0, ret_V_9_fu_483_p2 };
assign \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.ain_s0  = \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.a ;
assign \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.s  = { \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.fas_s2 , \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.sum_s1  };
assign \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.u2.a  = \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.ain_s1 ;
assign \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.u2.b  = \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.bin_s1 ;
assign \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.u2.cin  = \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.carry_s1 ;
assign \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.facout_s2  = \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.u2.cout ;
assign \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.fas_s2  = \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.u2.s ;
assign \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.u1.a  = \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.a [1:0];
assign \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.u1.b  = \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.bin_s0 [1:0];
assign \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.u1.cin  = 1'h1;
assign \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.facout_s1  = \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.u1.cout ;
assign \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.fas_s1  = \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.u1.s ;
assign \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.a  = \sub_5ns_5s_5_2_1_U6.din0 ;
assign \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.b  = \sub_5ns_5s_5_2_1_U6.din1 ;
assign \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.ce  = \sub_5ns_5s_5_2_1_U6.ce ;
assign \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.clk  = \sub_5ns_5s_5_2_1_U6.clk ;
assign \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.reset  = \sub_5ns_5s_5_2_1_U6.reset ;
assign \sub_5ns_5s_5_2_1_U6.dout  = \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.s ;
assign \sub_5ns_5s_5_2_1_U6.ce  = 1'h1;
assign \sub_5ns_5s_5_2_1_U6.clk  = ap_clk;
assign \sub_5ns_5s_5_2_1_U6.din0  = select_ln703_reg_928;
assign \sub_5ns_5s_5_2_1_U6.din1  = { op_6_V_reg_917[3], op_6_V_reg_917 };
assign grp_fu_495_p2 = \sub_5ns_5s_5_2_1_U6.dout ;
assign \sub_5ns_5s_5_2_1_U6.reset  = ap_rst;
assign \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.ain_s0  = \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.a ;
assign \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.bin_s0  = \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.b ;
assign \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.s  = { \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.fas_s2 , \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.sum_s1  };
assign \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.u2.a  = \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.ain_s1 ;
assign \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.u2.b  = \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.bin_s1 ;
assign \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.u2.cin  = \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.carry_s1 ;
assign \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.facout_s2  = \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.u2.cout ;
assign \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.fas_s2  = \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.u2.s ;
assign \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.u1.a  = \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.a [3:0];
assign \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.u1.b  = \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.b [3:0];
assign \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.u1.cin  = 1'h0;
assign \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.facout_s1  = \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.u1.cout ;
assign \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.fas_s1  = \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.u1.s ;
assign \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.a  = \add_9ns_9s_9_2_1_U2.din0 ;
assign \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.b  = \add_9ns_9s_9_2_1_U2.din1 ;
assign \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.ce  = \add_9ns_9s_9_2_1_U2.ce ;
assign \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.clk  = \add_9ns_9s_9_2_1_U2.clk ;
assign \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.reset  = \add_9ns_9s_9_2_1_U2.reset ;
assign \add_9ns_9s_9_2_1_U2.dout  = \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.s ;
assign \add_9ns_9s_9_2_1_U2.ce  = 1'h1;
assign \add_9ns_9s_9_2_1_U2.clk  = ap_clk;
assign \add_9ns_9s_9_2_1_U2.din0  = select_ln1192_reg_834;
assign \add_9ns_9s_9_2_1_U2.din1  = { op_2[7], op_2 };
assign grp_fu_293_p2 = \add_9ns_9s_9_2_1_U2.dout ;
assign \add_9ns_9s_9_2_1_U2.reset  = ap_rst;
assign \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.ain_s0  = \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.a ;
assign \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.bin_s0  = \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.b ;
assign \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.s  = { \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.fas_s2 , \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.sum_s1  };
assign \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.u2.a  = \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.ain_s1 ;
assign \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.u2.b  = \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.bin_s1 ;
assign \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.u2.cin  = \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.carry_s1 ;
assign \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.facout_s2  = \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.u2.cout ;
assign \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.fas_s2  = \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.u2.s ;
assign \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.u1.a  = \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.a [1:0];
assign \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.u1.b  = \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.b [1:0];
assign \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.u1.cin  = 1'h0;
assign \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.facout_s1  = \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.u1.cout ;
assign \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.fas_s1  = \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.u1.s ;
assign \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.a  = \add_5s_5ns_5_2_1_U16.din0 ;
assign \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.b  = \add_5s_5ns_5_2_1_U16.din1 ;
assign \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.ce  = \add_5s_5ns_5_2_1_U16.ce ;
assign \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.clk  = \add_5s_5ns_5_2_1_U16.clk ;
assign \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.reset  = \add_5s_5ns_5_2_1_U16.reset ;
assign \add_5s_5ns_5_2_1_U16.dout  = \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.s ;
assign \add_5s_5ns_5_2_1_U16.ce  = 1'h1;
assign \add_5s_5ns_5_2_1_U16.clk  = ap_clk;
assign \add_5s_5ns_5_2_1_U16.din0  = { op_17[3], op_17 };
assign \add_5s_5ns_5_2_1_U16.din1  = { 3'h0, tmp_reg_948 };
assign grp_fu_746_p2 = \add_5s_5ns_5_2_1_U16.dout ;
assign \add_5s_5ns_5_2_1_U16.reset  = ap_rst;
assign \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.ain_s0  = \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.a ;
assign \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.bin_s0  = \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.b ;
assign \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.s  = { \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.fas_s2 , \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.sum_s1  };
assign \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.u2.a  = \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.ain_s1 ;
assign \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.u2.b  = \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.bin_s1 ;
assign \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.u2.cin  = \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.carry_s1 ;
assign \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.facout_s2  = \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.u2.cout ;
assign \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.fas_s2  = \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.u2.s ;
assign \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.u1.a  = \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.a [1:0];
assign \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.u1.b  = \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.b [1:0];
assign \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.u1.cin  = 1'h0;
assign \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.facout_s1  = \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.u1.cout ;
assign \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.fas_s1  = \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.u1.s ;
assign \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.a  = \add_4ns_4s_4_2_1_U11.din0 ;
assign \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.b  = \add_4ns_4s_4_2_1_U11.din1 ;
assign \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.ce  = \add_4ns_4s_4_2_1_U11.ce ;
assign \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.clk  = \add_4ns_4s_4_2_1_U11.clk ;
assign \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.reset  = \add_4ns_4s_4_2_1_U11.reset ;
assign \add_4ns_4s_4_2_1_U11.dout  = \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.s ;
assign \add_4ns_4s_4_2_1_U11.ce  = 1'h1;
assign \add_4ns_4s_4_2_1_U11.clk  = ap_clk;
assign \add_4ns_4s_4_2_1_U11.din0  = { 1'h0, add_ln69_2_reg_1030 };
assign \add_4ns_4s_4_2_1_U11.din1  = { ret_V_22_reg_1015[1], ret_V_22_reg_1015[1], ret_V_22_reg_1015 };
assign grp_fu_661_p2 = \add_4ns_4s_4_2_1_U11.dout ;
assign \add_4ns_4s_4_2_1_U11.reset  = ap_rst;
assign \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.ain_s0  = \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.a ;
assign \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.bin_s0  = \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.b ;
assign \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.s  = { \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.fas_s2 , \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.sum_s1  };
assign \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.u2.a  = \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.ain_s1 ;
assign \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.u2.b  = \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.bin_s1 ;
assign \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.u2.cin  = \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.carry_s1 ;
assign \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.facout_s2  = \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.u2.cout ;
assign \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.fas_s2  = \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.u2.s ;
assign \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.u1.a  = \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.a [1:0];
assign \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.u1.b  = \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.b [1:0];
assign \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.u1.cin  = 1'h0;
assign \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.facout_s1  = \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.u1.cout ;
assign \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.fas_s1  = \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.u1.s ;
assign \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.a  = \add_4ns_4ns_4_2_1_U1.din0 ;
assign \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.b  = \add_4ns_4ns_4_2_1_U1.din1 ;
assign \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.ce  = \add_4ns_4ns_4_2_1_U1.ce ;
assign \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.clk  = \add_4ns_4ns_4_2_1_U1.clk ;
assign \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.reset  = \add_4ns_4ns_4_2_1_U1.reset ;
assign \add_4ns_4ns_4_2_1_U1.dout  = \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.s ;
assign \add_4ns_4ns_4_2_1_U1.ce  = 1'h1;
assign \add_4ns_4ns_4_2_1_U1.clk  = ap_clk;
assign \add_4ns_4ns_4_2_1_U1.din0  = { 3'h0, op_2[3] };
assign \add_4ns_4ns_4_2_1_U1.din1  = op_2[7:4];
assign grp_fu_235_p2 = \add_4ns_4ns_4_2_1_U1.dout ;
assign \add_4ns_4ns_4_2_1_U1.reset  = ap_rst;
assign \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.ain_s0  = \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.a ;
assign \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.bin_s0  = \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.b ;
assign \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.s  = { \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.fas_s2 , \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.sum_s1  };
assign \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.u2.a  = \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.ain_s1 ;
assign \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.u2.b  = \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.bin_s1 ;
assign \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.u2.cin  = \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.carry_s1 ;
assign \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.facout_s2  = \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.u2.cout ;
assign \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.fas_s2  = \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.u2.s ;
assign \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.u1.a  = \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.a [0];
assign \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.u1.b  = \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.b [0];
assign \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.u1.cin  = 1'h0;
assign \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.facout_s1  = \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.u1.cout ;
assign \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.fas_s1  = \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.u1.s ;
assign \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.a  = \add_3ns_3ns_3_2_1_U9.din0 ;
assign \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.b  = \add_3ns_3ns_3_2_1_U9.din1 ;
assign \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.ce  = \add_3ns_3ns_3_2_1_U9.ce ;
assign \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.clk  = \add_3ns_3ns_3_2_1_U9.clk ;
assign \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.reset  = \add_3ns_3ns_3_2_1_U9.reset ;
assign \add_3ns_3ns_3_2_1_U9.dout  = \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.s ;
assign \add_3ns_3ns_3_2_1_U9.ce  = 1'h1;
assign \add_3ns_3ns_3_2_1_U9.clk  = ap_clk;
assign \add_3ns_3ns_3_2_1_U9.din0  = { 1'h0, op_14 };
assign \add_3ns_3ns_3_2_1_U9.din1  = { 2'h0, op_13 };
assign grp_fu_619_p2 = \add_3ns_3ns_3_2_1_U9.dout ;
assign \add_3ns_3ns_3_2_1_U9.reset  = ap_rst;
assign \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.ain_s0  = \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.a ;
assign \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.bin_s0  = \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.b ;
assign \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.s  = { \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.fas_s2 , \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.sum_s1  };
assign \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.u2.a  = \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.ain_s1 ;
assign \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.u2.b  = \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.bin_s1 ;
assign \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.u2.cin  = \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.carry_s1 ;
assign \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.facout_s2  = \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.u2.cout ;
assign \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.fas_s2  = \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.u2.s ;
assign \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.u1.a  = \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.a [0];
assign \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.u1.b  = \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.b [0];
assign \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.u1.cin  = 1'h0;
assign \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.facout_s1  = \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.u1.cout ;
assign \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.fas_s1  = \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.u1.s ;
assign \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.a  = \add_2ns_2ns_2_2_1_U7.din0 ;
assign \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.b  = \add_2ns_2ns_2_2_1_U7.din1 ;
assign \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.ce  = \add_2ns_2ns_2_2_1_U7.ce ;
assign \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.clk  = \add_2ns_2ns_2_2_1_U7.clk ;
assign \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.reset  = \add_2ns_2ns_2_2_1_U7.reset ;
assign \add_2ns_2ns_2_2_1_U7.dout  = \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.s ;
assign \add_2ns_2ns_2_2_1_U7.ce  = 1'h1;
assign \add_2ns_2ns_2_2_1_U7.clk  = ap_clk;
assign \add_2ns_2ns_2_2_1_U7.din0  = ret_V_11_reg_968;
assign \add_2ns_2ns_2_2_1_U7.din1  = 2'h1;
assign grp_fu_593_p2 = \add_2ns_2ns_2_2_1_U7.dout ;
assign \add_2ns_2ns_2_2_1_U7.reset  = ap_rst;
assign \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.ain_s0  = \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.a ;
assign \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.bin_s0  = \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.b ;
assign \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.s  = { \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.fas_s2 , \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.sum_s1  };
assign \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.u2.a  = \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.ain_s1 ;
assign \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.u2.b  = \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.bin_s1 ;
assign \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.u2.cin  = \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.carry_s1 ;
assign \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.facout_s2  = \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.u2.cout ;
assign \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.fas_s2  = \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.u2.s ;
assign \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.u1.a  = \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.a [0];
assign \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.u1.b  = \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.b [0];
assign \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.u1.cin  = 1'h0;
assign \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.facout_s1  = \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.u1.cout ;
assign \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.fas_s1  = \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.u1.s ;
assign \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.a  = \add_2ns_2ns_2_2_1_U4.din0 ;
assign \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.b  = \add_2ns_2ns_2_2_1_U4.din1 ;
assign \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.ce  = \add_2ns_2ns_2_2_1_U4.ce ;
assign \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.clk  = \add_2ns_2ns_2_2_1_U4.clk ;
assign \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.reset  = \add_2ns_2ns_2_2_1_U4.reset ;
assign \add_2ns_2ns_2_2_1_U4.dout  = \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.s ;
assign \add_2ns_2ns_2_2_1_U4.ce  = 1'h1;
assign \add_2ns_2ns_2_2_1_U4.clk  = ap_clk;
assign \add_2ns_2ns_2_2_1_U4.din0  = ret_V_reg_878;
assign \add_2ns_2ns_2_2_1_U4.din1  = 2'h1;
assign grp_fu_420_p2 = \add_2ns_2ns_2_2_1_U4.dout ;
assign \add_2ns_2ns_2_2_1_U4.reset  = ap_rst;
assign \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.ain_s0  = \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.a ;
assign \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.bin_s0  = \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.b ;
assign \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.s  = { \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.fas_s2 , \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.sum_s1  };
assign \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.u2.a  = \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.ain_s1 ;
assign \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.u2.b  = \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.bin_s1 ;
assign \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.u2.cin  = \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.carry_s1 ;
assign \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.facout_s2  = \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.u2.cout ;
assign \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.fas_s2  = \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.u2.s ;
assign \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.u1.a  = \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.a [8:0];
assign \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.u1.b  = \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.b [8:0];
assign \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.u1.cin  = 1'h0;
assign \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.facout_s1  = \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.u1.cout ;
assign \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.fas_s1  = \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.u1.s ;
assign \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.a  = \add_18s_18ns_18_2_1_U17.din0 ;
assign \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.b  = \add_18s_18ns_18_2_1_U17.din1 ;
assign \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.ce  = \add_18s_18ns_18_2_1_U17.ce ;
assign \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.clk  = \add_18s_18ns_18_2_1_U17.clk ;
assign \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.reset  = \add_18s_18ns_18_2_1_U17.reset ;
assign \add_18s_18ns_18_2_1_U17.dout  = \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.s ;
assign \add_18s_18ns_18_2_1_U17.ce  = 1'h1;
assign \add_18s_18ns_18_2_1_U17.clk  = ap_clk;
assign \add_18s_18ns_18_2_1_U17.din0  = { add_ln69_7_reg_1120[4], add_ln69_7_reg_1120[4], add_ln69_7_reg_1120[4], add_ln69_7_reg_1120[4], add_ln69_7_reg_1120[4], add_ln69_7_reg_1120[4], add_ln69_7_reg_1120[4], add_ln69_7_reg_1120[4], add_ln69_7_reg_1120[4], add_ln69_7_reg_1120[4], add_ln69_7_reg_1120[4], add_ln69_7_reg_1120[4], add_ln69_7_reg_1120[4], add_ln69_7_reg_1120 };
assign \add_18s_18ns_18_2_1_U17.din1  = add_ln69_5_reg_1115;
assign grp_fu_755_p2 = \add_18s_18ns_18_2_1_U17.dout ;
assign \add_18s_18ns_18_2_1_U17.reset  = ap_rst;
assign \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.ain_s0  = \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.a ;
assign \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.bin_s0  = \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.b ;
assign \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.s  = { \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.fas_s2 , \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.sum_s1  };
assign \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.u2.a  = \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.ain_s1 ;
assign \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.u2.b  = \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.bin_s1 ;
assign \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.u2.cin  = \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.carry_s1 ;
assign \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.facout_s2  = \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.u2.cout ;
assign \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.fas_s2  = \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.u2.s ;
assign \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.u1.a  = \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.a [8:0];
assign \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.u1.b  = \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.b [8:0];
assign \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.u1.cin  = 1'h0;
assign \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.facout_s1  = \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.u1.cout ;
assign \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.fas_s1  = \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.u1.s ;
assign \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.a  = \add_18s_18ns_18_2_1_U15.din0 ;
assign \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.b  = \add_18s_18ns_18_2_1_U15.din1 ;
assign \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.ce  = \add_18s_18ns_18_2_1_U15.ce ;
assign \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.clk  = \add_18s_18ns_18_2_1_U15.clk ;
assign \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.reset  = \add_18s_18ns_18_2_1_U15.reset ;
assign \add_18s_18ns_18_2_1_U15.dout  = \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.s ;
assign \add_18s_18ns_18_2_1_U15.ce  = 1'h1;
assign \add_18s_18ns_18_2_1_U15.clk  = ap_clk;
assign \add_18s_18ns_18_2_1_U15.din0  = { ret_V_24_reg_1090[14], ret_V_24_reg_1090[14], ret_V_24_reg_1090[14], ret_V_24_reg_1090 };
assign \add_18s_18ns_18_2_1_U15.din1  = { 2'h0, ret_V_18_reg_953[1], ret_V_18_reg_953[1], ret_V_18_reg_953[1], ret_V_18_reg_953[1], ret_V_18_reg_953[1], ret_V_18_reg_953[1], ret_V_18_reg_953[1], ret_V_18_reg_953[1], ret_V_18_reg_953[1], ret_V_18_reg_953[1], ret_V_18_reg_953[1], ret_V_18_reg_953[1], ret_V_18_reg_953[1], ret_V_18_reg_953[1], ret_V_18_reg_953 };
assign grp_fu_740_p2 = \add_18s_18ns_18_2_1_U15.dout ;
assign \add_18s_18ns_18_2_1_U15.reset  = ap_rst;
assign \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.ain_s0  = \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.a ;
assign \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.bin_s0  = \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.b ;
assign \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.s  = { \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.fas_s2 , \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.sum_s1  };
assign \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.u2.a  = \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.ain_s1 ;
assign \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.u2.b  = \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.bin_s1 ;
assign \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.u2.cin  = \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.carry_s1 ;
assign \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.facout_s2  = \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.u2.cout ;
assign \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.fas_s2  = \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.u2.s ;
assign \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.u1.a  = \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.a [7:0];
assign \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.u1.b  = \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.b [7:0];
assign \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.u1.cin  = 1'h0;
assign \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.facout_s1  = \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.u1.cout ;
assign \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.fas_s1  = \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.u1.s ;
assign \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.a  = \add_17s_17s_17_2_1_U3.din0 ;
assign \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.b  = \add_17s_17s_17_2_1_U3.din1 ;
assign \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.ce  = \add_17s_17s_17_2_1_U3.ce ;
assign \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.clk  = \add_17s_17s_17_2_1_U3.clk ;
assign \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.reset  = \add_17s_17s_17_2_1_U3.reset ;
assign \add_17s_17s_17_2_1_U3.dout  = \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.s ;
assign \add_17s_17s_17_2_1_U3.ce  = 1'h1;
assign \add_17s_17s_17_2_1_U3.clk  = ap_clk;
assign \add_17s_17s_17_2_1_U3.din0  = { op_9[3], op_9[3], op_9[3], op_9[3], op_9[3], op_9[3], op_9[3], op_9[3], op_9[3], op_9[3], op_9[3], op_9[3], op_9, 1'h0 };
assign \add_17s_17s_17_2_1_U3.din1  = { op_0[15], op_0 };
assign grp_fu_376_p2 = \add_17s_17s_17_2_1_U3.dout ;
assign \add_17s_17s_17_2_1_U3.reset  = ap_rst;
assign \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.ain_s0  = \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.a ;
assign \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.bin_s0  = \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.b ;
assign \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.s  = { \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.fas_s2 , \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.sum_s1  };
assign \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.u2.a  = \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.ain_s1 ;
assign \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.u2.b  = \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.bin_s1 ;
assign \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.u2.cin  = \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.carry_s1 ;
assign \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.facout_s2  = \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.u2.cout ;
assign \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.fas_s2  = \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.u2.s ;
assign \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.u1.a  = \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.a [6:0];
assign \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.u1.b  = \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.b [6:0];
assign \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.u1.cin  = 1'h0;
assign \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.facout_s1  = \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.u1.cout ;
assign \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.fas_s1  = \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.u1.s ;
assign \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.a  = \add_15s_15s_15_2_1_U14.din0 ;
assign \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.b  = \add_15s_15s_15_2_1_U14.din1 ;
assign \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.ce  = \add_15s_15s_15_2_1_U14.ce ;
assign \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.clk  = \add_15s_15s_15_2_1_U14.clk ;
assign \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.reset  = \add_15s_15s_15_2_1_U14.reset ;
assign \add_15s_15s_15_2_1_U14.dout  = \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.s ;
assign \add_15s_15s_15_2_1_U14.ce  = 1'h1;
assign \add_15s_15s_15_2_1_U14.clk  = ap_clk;
assign \add_15s_15s_15_2_1_U14.din0  = { op_26_V_reg_1075[13], op_26_V_reg_1075 };
assign \add_15s_15s_15_2_1_U14.din1  = { op_16[1], op_16[1], op_16[1], op_16[1], op_16[1], op_16[1], op_16[1], op_16[1], op_16[1], op_16[1], op_16[1], op_16[1], op_16[1], op_16 };
assign grp_fu_717_p2 = \add_15s_15s_15_2_1_U14.dout ;
assign \add_15s_15s_15_2_1_U14.reset  = ap_rst;
assign \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.ain_s0  = \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.a ;
assign \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.bin_s0  = \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.b ;
assign \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.s  = { \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.fas_s2 , \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.sum_s1  };
assign \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.u2.a  = \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.ain_s1 ;
assign \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.u2.b  = \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.bin_s1 ;
assign \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.u2.cin  = \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.carry_s1 ;
assign \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.facout_s2  = \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.u2.cout ;
assign \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.fas_s2  = \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.u2.s ;
assign \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.u1.a  = \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.a [6:0];
assign \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.u1.b  = \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.b [6:0];
assign \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.u1.cin  = 1'h0;
assign \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.facout_s1  = \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.u1.cout ;
assign \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.fas_s1  = \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.u1.s ;
assign \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.a  = \add_15ns_15s_15_2_1_U13.din0 ;
assign \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.b  = \add_15ns_15s_15_2_1_U13.din1 ;
assign \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.ce  = \add_15ns_15s_15_2_1_U13.ce ;
assign \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.clk  = \add_15ns_15s_15_2_1_U13.clk ;
assign \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.reset  = \add_15ns_15s_15_2_1_U13.reset ;
assign \add_15ns_15s_15_2_1_U13.dout  = \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.s ;
assign \add_15ns_15s_15_2_1_U13.ce  = 1'h1;
assign \add_15ns_15s_15_2_1_U13.clk  = ap_clk;
assign \add_15ns_15s_15_2_1_U13.din0  = { op_25_V_reg_1060, 1'h0 };
assign \add_15ns_15s_15_2_1_U13.din1  = { op_1, op_1, op_1, op_1, op_1, op_1, op_1, op_1, op_1, op_1, op_1, op_1, op_1, op_1, 1'h0 };
assign grp_fu_694_p2 = \add_15ns_15s_15_2_1_U13.dout ;
assign \add_15ns_15s_15_2_1_U13.reset  = ap_rst;
assign \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.ain_s0  = \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.a ;
assign \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.bin_s0  = \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.b ;
assign \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.s  = { \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.fas_s2 , \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.sum_s1  };
assign \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.u2.a  = \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.ain_s1 ;
assign \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.u2.b  = \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.bin_s1 ;
assign \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.u2.cin  = \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.carry_s1 ;
assign \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.facout_s2  = \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.u2.cout ;
assign \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.fas_s2  = \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.u2.s ;
assign \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.u1.a  = \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.a [6:0];
assign \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.u1.b  = \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.b [6:0];
assign \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.u1.cin  = 1'h0;
assign \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.facout_s1  = \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.u1.cout ;
assign \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.fas_s1  = \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.u1.s ;
assign \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.a  = \add_14s_14ns_14_2_1_U8.din0 ;
assign \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.b  = \add_14s_14ns_14_2_1_U8.din1 ;
assign \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.ce  = \add_14s_14ns_14_2_1_U8.ce ;
assign \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.clk  = \add_14s_14ns_14_2_1_U8.clk ;
assign \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.reset  = \add_14s_14ns_14_2_1_U8.reset ;
assign \add_14s_14ns_14_2_1_U8.dout  = \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.s ;
assign \add_14s_14ns_14_2_1_U8.ce  = 1'h1;
assign \add_14s_14ns_14_2_1_U8.clk  = ap_clk;
assign \add_14s_14ns_14_2_1_U8.din0  = { ret_V_20_reg_980[12], ret_V_20_reg_980 };
assign \add_14s_14ns_14_2_1_U8.din1  = { 10'h000, op_12 };
assign grp_fu_613_p2 = \add_14s_14ns_14_2_1_U8.dout ;
assign \add_14s_14ns_14_2_1_U8.reset  = ap_rst;
assign \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.ain_s0  = \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.a ;
assign \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.bin_s0  = \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.b ;
assign \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.s  = { \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.fas_s2 , \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.sum_s1  };
assign \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.u2.a  = \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.ain_s1 ;
assign \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.u2.b  = \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.bin_s1 ;
assign \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.u2.cin  = \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.carry_s1 ;
assign \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.facout_s2  = \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.u2.cout ;
assign \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.fas_s2  = \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.u2.s ;
assign \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.u1.a  = \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.a [6:0];
assign \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.u1.b  = \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.b [6:0];
assign \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.u1.cin  = 1'h0;
assign \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.facout_s1  = \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.u1.cout ;
assign \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.fas_s1  = \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.u1.s ;
assign \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.a  = \add_14s_14ns_14_2_1_U12.din0 ;
assign \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.b  = \add_14s_14ns_14_2_1_U12.din1 ;
assign \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.ce  = \add_14s_14ns_14_2_1_U12.ce ;
assign \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.clk  = \add_14s_14ns_14_2_1_U12.clk ;
assign \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.reset  = \add_14s_14ns_14_2_1_U12.reset ;
assign \add_14s_14ns_14_2_1_U12.dout  = \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.s ;
assign \add_14s_14ns_14_2_1_U12.ce  = 1'h1;
assign \add_14s_14ns_14_2_1_U12.clk  = ap_clk;
assign \add_14s_14ns_14_2_1_U12.din0  = { add_ln69_3_reg_1050[3], add_ln69_3_reg_1050[3], add_ln69_3_reg_1050[3], add_ln69_3_reg_1050[3], add_ln69_3_reg_1050[3], add_ln69_3_reg_1050[3], add_ln69_3_reg_1050[3], add_ln69_3_reg_1050[3], add_ln69_3_reg_1050[3], add_ln69_3_reg_1050[3], add_ln69_3_reg_1050 };
assign \add_14s_14ns_14_2_1_U12.din1  = add_ln69_1_reg_1045;
assign grp_fu_670_p2 = \add_14s_14ns_14_2_1_U12.dout ;
assign \add_14s_14ns_14_2_1_U12.reset  = ap_rst;
assign \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.ain_s0  = \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.a ;
assign \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.bin_s0  = \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.b ;
assign \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.s  = { \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.fas_s2 , \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.sum_s1  };
assign \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.u2.a  = \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.ain_s1 ;
assign \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.u2.b  = \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.bin_s1 ;
assign \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.u2.cin  = \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.carry_s1 ;
assign \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.facout_s2  = \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.u2.cout ;
assign \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.fas_s2  = \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.u2.s ;
assign \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.u1.a  = \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.a [6:0];
assign \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.u1.b  = \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.b [6:0];
assign \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.u1.cin  = 1'h0;
assign \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.facout_s1  = \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.u1.cout ;
assign \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.fas_s1  = \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.u1.s ;
assign \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.a  = \add_14ns_14ns_14_2_1_U10.din0 ;
assign \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.b  = \add_14ns_14ns_14_2_1_U10.din1 ;
assign \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.ce  = \add_14ns_14ns_14_2_1_U10.ce ;
assign \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.clk  = \add_14ns_14ns_14_2_1_U10.clk ;
assign \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.reset  = \add_14ns_14ns_14_2_1_U10.reset ;
assign \add_14ns_14ns_14_2_1_U10.dout  = \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.s ;
assign \add_14ns_14ns_14_2_1_U10.ce  = 1'h1;
assign \add_14ns_14ns_14_2_1_U10.clk  = ap_clk;
assign \add_14ns_14ns_14_2_1_U10.din0  = add_ln69_reg_1025;
assign \add_14ns_14ns_14_2_1_U10.din1  = select_ln69_reg_1020;
assign grp_fu_654_p2 = \add_14ns_14ns_14_2_1_U10.dout ;
assign \add_14ns_14ns_14_2_1_U10.reset  = ap_rst;
assign \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.ain_s0  = \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.a ;
assign \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.bin_s0  = \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.b ;
assign \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.s  = { \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.fas_s2 , \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.sum_s1  };
assign \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.u2.a  = \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.ain_s1 ;
assign \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.u2.b  = \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.bin_s1 ;
assign \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.u2.cin  = \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.carry_s1 ;
assign \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.facout_s2  = \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.u2.cout ;
assign \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.fas_s2  = \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.u2.s ;
assign \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.u1.a  = \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.a [5:0];
assign \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.u1.b  = \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.b [5:0];
assign \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.u1.cin  = 1'h0;
assign \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.facout_s1  = \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.u1.cout ;
assign \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.fas_s1  = \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.u1.s ;
assign \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.a  = \add_13ns_13ns_13_2_1_U5.din0 ;
assign \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.b  = \add_13ns_13ns_13_2_1_U5.din1 ;
assign \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.ce  = \add_13ns_13ns_13_2_1_U5.ce ;
assign \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.clk  = \add_13ns_13ns_13_2_1_U5.clk ;
assign \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.reset  = \add_13ns_13ns_13_2_1_U5.reset ;
assign \add_13ns_13ns_13_2_1_U5.dout  = \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.s ;
assign \add_13ns_13ns_13_2_1_U5.ce  = 1'h1;
assign \add_13ns_13ns_13_2_1_U5.clk  = ap_clk;
assign \add_13ns_13ns_13_2_1_U5.din0  = ret_V_4_reg_905;
assign \add_13ns_13ns_13_2_1_U5.din1  = 13'h0001;
assign grp_fu_478_p2 = \add_13ns_13ns_13_2_1_U5.dout ;
assign \add_13ns_13ns_13_2_1_U5.reset  = ap_rst;
endmodule


// Machine B:
// Processed by function `add_clk_enable_signal` in `verilog_tricks.py`.
// Processed by function `remove_reset_signal` in `verilog_tricks.py`.
module top_B (
  ap_clk,
  ap_start,
  ap_done,
  ap_idle,
  ap_ready,
  op_0,
  op_1,
  op_2,
  op_3,
  op_9,
  op_12,
  op_13,
  op_14,
  op_16,
  op_17,
  op_30,
  op_30_ap_vld,
clk_enable
);
input clk_enable;


input ap_clk;
wire ap_rst;
assign ap_rst = op_30_ap_vld;
input ap_start;
input [15:0] op_0;
input op_1;
input [3:0] op_12;
input op_13;
input [1:0] op_14;
input [1:0] op_16;
input [3:0] op_17;
input [7:0] op_2;
input op_3;
input [3:0] op_9;
output ap_done;
output ap_idle;
output ap_ready;
output [31:0] op_30;
output op_30_ap_vld;


reg Range2_all_ones_reg_800;
reg [6:0] \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.ain_s1 ;
reg [6:0] \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.bin_s1 ;
reg \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.carry_s1 ;
reg [5:0] \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.sum_s1 ;
reg [6:0] \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.ain_s1 ;
reg [6:0] \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.bin_s1 ;
reg \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.carry_s1 ;
reg [6:0] \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.sum_s1 ;
reg [6:0] \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.ain_s1 ;
reg [6:0] \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.bin_s1 ;
reg \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.carry_s1 ;
reg [6:0] \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.sum_s1 ;
reg [6:0] \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.ain_s1 ;
reg [6:0] \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.bin_s1 ;
reg \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.carry_s1 ;
reg [6:0] \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.sum_s1 ;
reg [7:0] \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.ain_s1 ;
reg [7:0] \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.bin_s1 ;
reg \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.carry_s1 ;
reg [6:0] \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.sum_s1 ;
reg [7:0] \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.ain_s1 ;
reg [7:0] \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.bin_s1 ;
reg \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.carry_s1 ;
reg [6:0] \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.sum_s1 ;
reg [8:0] \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.ain_s1 ;
reg [8:0] \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.bin_s1 ;
reg \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.carry_s1 ;
reg [7:0] \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.sum_s1 ;
reg [8:0] \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.ain_s1 ;
reg [8:0] \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.bin_s1 ;
reg \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.carry_s1 ;
reg [8:0] \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.sum_s1 ;
reg [8:0] \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.ain_s1 ;
reg [8:0] \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.bin_s1 ;
reg \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.carry_s1 ;
reg [8:0] \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.sum_s1 ;
reg \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.ain_s1 ;
reg \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.bin_s1 ;
reg \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.carry_s1 ;
reg \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.sum_s1 ;
reg \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.ain_s1 ;
reg \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.bin_s1 ;
reg \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.carry_s1 ;
reg \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.sum_s1 ;
reg [1:0] \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.ain_s1 ;
reg [1:0] \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.bin_s1 ;
reg \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.carry_s1 ;
reg \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.sum_s1 ;
reg [1:0] \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.ain_s1 ;
reg [1:0] \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.bin_s1 ;
reg \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.carry_s1 ;
reg [1:0] \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.sum_s1 ;
reg [1:0] \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.ain_s1 ;
reg [1:0] \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.bin_s1 ;
reg \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.carry_s1 ;
reg [1:0] \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.sum_s1 ;
reg [2:0] \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.ain_s1 ;
reg [2:0] \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.bin_s1 ;
reg \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.carry_s1 ;
reg [1:0] \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.sum_s1 ;
reg [4:0] \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.ain_s1 ;
reg [4:0] \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.bin_s1 ;
reg \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.carry_s1 ;
reg [3:0] \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.sum_s1 ;
reg [13:0] add_ln69_1_reg_1045;
reg [2:0] add_ln69_2_reg_1030;
reg [3:0] add_ln69_3_reg_1050;
reg [17:0] add_ln69_5_reg_1115;
reg [4:0] add_ln69_7_reg_1120;
reg [13:0] add_ln69_reg_1025;
reg and_ln786_reg_867;
reg [22:0] ap_CS_fsm = 23'h000001;
reg deleted_zeros_reg_856;
reg icmp_ln851_1_reg_938;
reg icmp_ln851_2_reg_809;
reg icmp_ln851_3_reg_985;
reg icmp_ln851_reg_779;
reg neg_src_reg_862;
reg [13:0] op_25_V_reg_1060;
reg [13:0] op_26_V_reg_1075;
reg [3:0] op_6_V_reg_917;
reg or_ln778_reg_845;
reg p_Result_3_reg_771;
reg p_Result_4_reg_789;
reg p_Result_5_reg_820;
reg [3:0] p_Val2_3_reg_814;
reg [1:0] ret_V_11_reg_968;
reg [1:0] ret_V_12_reg_995;
reg [8:0] ret_V_17_reg_873;
reg [1:0] ret_V_18_reg_953;
reg [16:0] ret_V_19_reg_900;
reg [12:0] ret_V_20_reg_980;
reg [4:0] ret_V_21_reg_963;
reg [1:0] ret_V_22_reg_1015;
reg [14:0] ret_V_24_reg_1090;
reg [1:0] ret_V_2_reg_933;
reg [12:0] ret_V_4_reg_905;
reg [12:0] ret_V_6_reg_958;
reg [1:0] ret_V_reg_878;
reg [8:0] select_ln1192_reg_834;
reg [3:0] select_ln340_reg_895;
reg [13:0] select_ln69_reg_1020;
reg [4:0] select_ln703_reg_928;
reg [1:0] select_ln831_reg_922;
reg [2:0] \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.ain_s1 ;
reg [2:0] \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.bin_s1 ;
reg \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.carry_s1 ;
reg [1:0] \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.sum_s1 ;
reg [1:0] tmp_reg_948;
reg [2:0] trunc_ln851_2_reg_975;
reg [3:0] trunc_ln851_reg_912;
reg xor_ln416_reg_839;
wire _000_;
wire [13:0] _001_;
wire [2:0] _002_;
wire [3:0] _003_;
wire [17:0] _004_;
wire [4:0] _005_;
wire [13:0] _006_;
wire _007_;
wire [22:0] _008_;
wire _009_;
wire _010_;
wire _011_;
wire _012_;
wire _013_;
wire _014_;
wire [13:0] _015_;
wire [13:0] _016_;
wire [3:0] _017_;
wire _018_;
wire _019_;
wire _020_;
wire _021_;
wire [3:0] _022_;
wire [1:0] _023_;
wire [1:0] _024_;
wire [8:0] _025_;
wire [1:0] _026_;
wire [16:0] _027_;
wire [12:0] _028_;
wire [4:0] _029_;
wire [1:0] _030_;
wire [14:0] _031_;
wire [1:0] _032_;
wire [12:0] _033_;
wire [12:0] _034_;
wire [1:0] _035_;
wire [1:0] _036_;
wire [3:0] _037_;
wire [7:0] _038_;
wire [1:0] _039_;
wire [1:0] _040_;
wire [1:0] _041_;
wire [2:0] _042_;
wire [3:0] _043_;
wire _044_;
wire [1:0] _045_;
wire _046_;
wire _047_;
wire _048_;
wire _049_;
wire _050_;
wire _051_;
wire _052_;
wire _053_;
wire [6:0] _054_;
wire [6:0] _055_;
wire _056_;
wire [5:0] _057_;
wire [6:0] _058_;
wire [7:0] _059_;
wire [6:0] _060_;
wire [6:0] _061_;
wire _062_;
wire [6:0] _063_;
wire [7:0] _064_;
wire [7:0] _065_;
wire [6:0] _066_;
wire [6:0] _067_;
wire _068_;
wire [6:0] _069_;
wire [7:0] _070_;
wire [7:0] _071_;
wire [6:0] _072_;
wire [6:0] _073_;
wire _074_;
wire [6:0] _075_;
wire [7:0] _076_;
wire [7:0] _077_;
wire [7:0] _078_;
wire [7:0] _079_;
wire _080_;
wire [6:0] _081_;
wire [7:0] _082_;
wire [8:0] _083_;
wire [7:0] _084_;
wire [7:0] _085_;
wire _086_;
wire [6:0] _087_;
wire [7:0] _088_;
wire [8:0] _089_;
wire [8:0] _090_;
wire [8:0] _091_;
wire _092_;
wire [7:0] _093_;
wire [8:0] _094_;
wire [9:0] _095_;
wire [8:0] _096_;
wire [8:0] _097_;
wire _098_;
wire [8:0] _099_;
wire [9:0] _100_;
wire [9:0] _101_;
wire [8:0] _102_;
wire [8:0] _103_;
wire _104_;
wire [8:0] _105_;
wire [9:0] _106_;
wire [9:0] _107_;
wire _108_;
wire _109_;
wire _110_;
wire _111_;
wire [1:0] _112_;
wire [1:0] _113_;
wire _114_;
wire _115_;
wire _116_;
wire _117_;
wire [1:0] _118_;
wire [1:0] _119_;
wire [1:0] _120_;
wire [1:0] _121_;
wire _122_;
wire _123_;
wire [1:0] _124_;
wire [2:0] _125_;
wire [1:0] _126_;
wire [1:0] _127_;
wire _128_;
wire [1:0] _129_;
wire [2:0] _130_;
wire [2:0] _131_;
wire [1:0] _132_;
wire [1:0] _133_;
wire _134_;
wire [1:0] _135_;
wire [2:0] _136_;
wire [2:0] _137_;
wire [2:0] _138_;
wire [2:0] _139_;
wire _140_;
wire [1:0] _141_;
wire [2:0] _142_;
wire [3:0] _143_;
wire [4:0] _144_;
wire [4:0] _145_;
wire _146_;
wire [3:0] _147_;
wire [4:0] _148_;
wire [5:0] _149_;
wire [2:0] _150_;
wire [2:0] _151_;
wire _152_;
wire [1:0] _153_;
wire [2:0] _154_;
wire [3:0] _155_;
wire _156_;
wire _157_;
wire _158_;
wire _159_;
wire _160_;
wire _161_;
wire _162_;
wire _163_;
wire _164_;
wire _165_;
wire _166_;
wire _167_;
wire _168_;
wire _169_;
wire _170_;
wire _171_;
wire _172_;
wire _173_;
wire _174_;
wire _175_;
wire _176_;
wire _177_;
wire _178_;
wire [7:0] Range2_all_ones_fu_241_p1;
wire \add_13ns_13ns_13_2_1_U5.ce ;
wire \add_13ns_13ns_13_2_1_U5.clk ;
wire [12:0] \add_13ns_13ns_13_2_1_U5.din0 ;
wire [12:0] \add_13ns_13ns_13_2_1_U5.din1 ;
wire [12:0] \add_13ns_13ns_13_2_1_U5.dout ;
wire \add_13ns_13ns_13_2_1_U5.reset ;
wire [12:0] \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.a ;
wire [12:0] \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.ain_s0 ;
wire [12:0] \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.b ;
wire [12:0] \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.bin_s0 ;
wire \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.ce ;
wire \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.clk ;
wire \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.facout_s1 ;
wire \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.facout_s2 ;
wire [5:0] \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.fas_s1 ;
wire [6:0] \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.fas_s2 ;
wire \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.reset ;
wire [12:0] \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.s ;
wire [5:0] \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.u1.a ;
wire [5:0] \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.u1.b ;
wire \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.u1.cin ;
wire \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.u1.cout ;
wire [5:0] \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.u1.s ;
wire [6:0] \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.u2.a ;
wire [6:0] \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.u2.b ;
wire \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.u2.cin ;
wire \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.u2.cout ;
wire [6:0] \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.u2.s ;
wire \add_14ns_14ns_14_2_1_U10.ce ;
wire \add_14ns_14ns_14_2_1_U10.clk ;
wire [13:0] \add_14ns_14ns_14_2_1_U10.din0 ;
wire [13:0] \add_14ns_14ns_14_2_1_U10.din1 ;
wire [13:0] \add_14ns_14ns_14_2_1_U10.dout ;
wire \add_14ns_14ns_14_2_1_U10.reset ;
wire [13:0] \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.a ;
wire [13:0] \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.ain_s0 ;
wire [13:0] \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.b ;
wire [13:0] \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.bin_s0 ;
wire \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.ce ;
wire \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.clk ;
wire \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.facout_s1 ;
wire \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.facout_s2 ;
wire [6:0] \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.fas_s1 ;
wire [6:0] \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.fas_s2 ;
wire \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.reset ;
wire [13:0] \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.s ;
wire [6:0] \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.u1.a ;
wire [6:0] \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.u1.b ;
wire \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.u1.cin ;
wire \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.u1.cout ;
wire [6:0] \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.u1.s ;
wire [6:0] \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.u2.a ;
wire [6:0] \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.u2.b ;
wire \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.u2.cin ;
wire \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.u2.cout ;
wire [6:0] \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.u2.s ;
wire \add_14s_14ns_14_2_1_U12.ce ;
wire \add_14s_14ns_14_2_1_U12.clk ;
wire [13:0] \add_14s_14ns_14_2_1_U12.din0 ;
wire [13:0] \add_14s_14ns_14_2_1_U12.din1 ;
wire [13:0] \add_14s_14ns_14_2_1_U12.dout ;
wire \add_14s_14ns_14_2_1_U12.reset ;
wire [13:0] \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.a ;
wire [13:0] \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.ain_s0 ;
wire [13:0] \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.b ;
wire [13:0] \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.bin_s0 ;
wire \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.ce ;
wire \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.clk ;
wire \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.facout_s1 ;
wire \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.facout_s2 ;
wire [6:0] \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.fas_s1 ;
wire [6:0] \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.fas_s2 ;
wire \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.reset ;
wire [13:0] \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.s ;
wire [6:0] \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.u1.a ;
wire [6:0] \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.u1.b ;
wire \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.u1.cin ;
wire \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.u1.cout ;
wire [6:0] \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.u1.s ;
wire [6:0] \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.u2.a ;
wire [6:0] \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.u2.b ;
wire \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.u2.cin ;
wire \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.u2.cout ;
wire [6:0] \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.u2.s ;
wire \add_14s_14ns_14_2_1_U8.ce ;
wire \add_14s_14ns_14_2_1_U8.clk ;
wire [13:0] \add_14s_14ns_14_2_1_U8.din0 ;
wire [13:0] \add_14s_14ns_14_2_1_U8.din1 ;
wire [13:0] \add_14s_14ns_14_2_1_U8.dout ;
wire \add_14s_14ns_14_2_1_U8.reset ;
wire [13:0] \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.a ;
wire [13:0] \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.ain_s0 ;
wire [13:0] \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.b ;
wire [13:0] \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.bin_s0 ;
wire \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.ce ;
wire \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.clk ;
wire \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.facout_s1 ;
wire \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.facout_s2 ;
wire [6:0] \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.fas_s1 ;
wire [6:0] \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.fas_s2 ;
wire \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.reset ;
wire [13:0] \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.s ;
wire [6:0] \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.u1.a ;
wire [6:0] \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.u1.b ;
wire \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.u1.cin ;
wire \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.u1.cout ;
wire [6:0] \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.u1.s ;
wire [6:0] \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.u2.a ;
wire [6:0] \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.u2.b ;
wire \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.u2.cin ;
wire \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.u2.cout ;
wire [6:0] \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.u2.s ;
wire \add_15ns_15s_15_2_1_U13.ce ;
wire \add_15ns_15s_15_2_1_U13.clk ;
wire [14:0] \add_15ns_15s_15_2_1_U13.din0 ;
wire [14:0] \add_15ns_15s_15_2_1_U13.din1 ;
wire [14:0] \add_15ns_15s_15_2_1_U13.dout ;
wire \add_15ns_15s_15_2_1_U13.reset ;
wire [14:0] \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.a ;
wire [14:0] \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.ain_s0 ;
wire [14:0] \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.b ;
wire [14:0] \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.bin_s0 ;
wire \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.ce ;
wire \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.clk ;
wire \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.facout_s1 ;
wire \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.facout_s2 ;
wire [6:0] \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.fas_s1 ;
wire [7:0] \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.fas_s2 ;
wire \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.reset ;
wire [14:0] \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.s ;
wire [6:0] \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.u1.a ;
wire [6:0] \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.u1.b ;
wire \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.u1.cin ;
wire \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.u1.cout ;
wire [6:0] \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.u1.s ;
wire [7:0] \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.u2.a ;
wire [7:0] \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.u2.b ;
wire \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.u2.cin ;
wire \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.u2.cout ;
wire [7:0] \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.u2.s ;
wire \add_15s_15s_15_2_1_U14.ce ;
wire \add_15s_15s_15_2_1_U14.clk ;
wire [14:0] \add_15s_15s_15_2_1_U14.din0 ;
wire [14:0] \add_15s_15s_15_2_1_U14.din1 ;
wire [14:0] \add_15s_15s_15_2_1_U14.dout ;
wire \add_15s_15s_15_2_1_U14.reset ;
wire [14:0] \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.a ;
wire [14:0] \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.ain_s0 ;
wire [14:0] \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.b ;
wire [14:0] \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.bin_s0 ;
wire \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.ce ;
wire \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.clk ;
wire \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.facout_s1 ;
wire \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.facout_s2 ;
wire [6:0] \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.fas_s1 ;
wire [7:0] \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.fas_s2 ;
wire \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.reset ;
wire [14:0] \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.s ;
wire [6:0] \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.u1.a ;
wire [6:0] \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.u1.b ;
wire \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.u1.cin ;
wire \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.u1.cout ;
wire [6:0] \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.u1.s ;
wire [7:0] \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.u2.a ;
wire [7:0] \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.u2.b ;
wire \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.u2.cin ;
wire \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.u2.cout ;
wire [7:0] \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.u2.s ;
wire \add_17s_17s_17_2_1_U3.ce ;
wire \add_17s_17s_17_2_1_U3.clk ;
wire [16:0] \add_17s_17s_17_2_1_U3.din0 ;
wire [16:0] \add_17s_17s_17_2_1_U3.din1 ;
wire [16:0] \add_17s_17s_17_2_1_U3.dout ;
wire \add_17s_17s_17_2_1_U3.reset ;
wire [16:0] \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.a ;
wire [16:0] \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.ain_s0 ;
wire [16:0] \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.b ;
wire [16:0] \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.bin_s0 ;
wire \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.ce ;
wire \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.clk ;
wire \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.facout_s1 ;
wire \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.facout_s2 ;
wire [7:0] \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.fas_s1 ;
wire [8:0] \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.fas_s2 ;
wire \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.reset ;
wire [16:0] \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.s ;
wire [7:0] \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.u1.a ;
wire [7:0] \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.u1.b ;
wire \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.u1.cin ;
wire \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.u1.cout ;
wire [7:0] \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.u1.s ;
wire [8:0] \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.u2.a ;
wire [8:0] \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.u2.b ;
wire \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.u2.cin ;
wire \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.u2.cout ;
wire [8:0] \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.u2.s ;
wire \add_18s_18ns_18_2_1_U15.ce ;
wire \add_18s_18ns_18_2_1_U15.clk ;
wire [17:0] \add_18s_18ns_18_2_1_U15.din0 ;
wire [17:0] \add_18s_18ns_18_2_1_U15.din1 ;
wire [17:0] \add_18s_18ns_18_2_1_U15.dout ;
wire \add_18s_18ns_18_2_1_U15.reset ;
wire [17:0] \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.a ;
wire [17:0] \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.ain_s0 ;
wire [17:0] \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.b ;
wire [17:0] \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.bin_s0 ;
wire \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.ce ;
wire \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.clk ;
wire \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.facout_s1 ;
wire \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.facout_s2 ;
wire [8:0] \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.fas_s1 ;
wire [8:0] \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.fas_s2 ;
wire \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.reset ;
wire [17:0] \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.s ;
wire [8:0] \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.u1.a ;
wire [8:0] \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.u1.b ;
wire \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.u1.cin ;
wire \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.u1.cout ;
wire [8:0] \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.u1.s ;
wire [8:0] \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.u2.a ;
wire [8:0] \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.u2.b ;
wire \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.u2.cin ;
wire \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.u2.cout ;
wire [8:0] \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.u2.s ;
wire \add_18s_18ns_18_2_1_U17.ce ;
wire \add_18s_18ns_18_2_1_U17.clk ;
wire [17:0] \add_18s_18ns_18_2_1_U17.din0 ;
wire [17:0] \add_18s_18ns_18_2_1_U17.din1 ;
wire [17:0] \add_18s_18ns_18_2_1_U17.dout ;
wire \add_18s_18ns_18_2_1_U17.reset ;
wire [17:0] \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.a ;
wire [17:0] \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.ain_s0 ;
wire [17:0] \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.b ;
wire [17:0] \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.bin_s0 ;
wire \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.ce ;
wire \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.clk ;
wire \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.facout_s1 ;
wire \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.facout_s2 ;
wire [8:0] \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.fas_s1 ;
wire [8:0] \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.fas_s2 ;
wire \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.reset ;
wire [17:0] \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.s ;
wire [8:0] \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.u1.a ;
wire [8:0] \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.u1.b ;
wire \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.u1.cin ;
wire \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.u1.cout ;
wire [8:0] \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.u1.s ;
wire [8:0] \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.u2.a ;
wire [8:0] \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.u2.b ;
wire \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.u2.cin ;
wire \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.u2.cout ;
wire [8:0] \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.u2.s ;
wire \add_2ns_2ns_2_2_1_U4.ce ;
wire \add_2ns_2ns_2_2_1_U4.clk ;
wire [1:0] \add_2ns_2ns_2_2_1_U4.din0 ;
wire [1:0] \add_2ns_2ns_2_2_1_U4.din1 ;
wire [1:0] \add_2ns_2ns_2_2_1_U4.dout ;
wire \add_2ns_2ns_2_2_1_U4.reset ;
wire [1:0] \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.a ;
wire [1:0] \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.ain_s0 ;
wire [1:0] \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.b ;
wire [1:0] \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.bin_s0 ;
wire \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.ce ;
wire \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.clk ;
wire \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.facout_s1 ;
wire \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.facout_s2 ;
wire \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.fas_s1 ;
wire \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.fas_s2 ;
wire \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.reset ;
wire [1:0] \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.s ;
wire \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.u1.a ;
wire \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.u1.b ;
wire \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.u1.cin ;
wire \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.u1.cout ;
wire \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.u1.s ;
wire \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.u2.a ;
wire \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.u2.b ;
wire \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.u2.cin ;
wire \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.u2.cout ;
wire \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.u2.s ;
wire \add_2ns_2ns_2_2_1_U7.ce ;
wire \add_2ns_2ns_2_2_1_U7.clk ;
wire [1:0] \add_2ns_2ns_2_2_1_U7.din0 ;
wire [1:0] \add_2ns_2ns_2_2_1_U7.din1 ;
wire [1:0] \add_2ns_2ns_2_2_1_U7.dout ;
wire \add_2ns_2ns_2_2_1_U7.reset ;
wire [1:0] \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.a ;
wire [1:0] \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.ain_s0 ;
wire [1:0] \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.b ;
wire [1:0] \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.bin_s0 ;
wire \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.ce ;
wire \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.clk ;
wire \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.facout_s1 ;
wire \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.facout_s2 ;
wire \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.fas_s1 ;
wire \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.fas_s2 ;
wire \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.reset ;
wire [1:0] \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.s ;
wire \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.u1.a ;
wire \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.u1.b ;
wire \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.u1.cin ;
wire \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.u1.cout ;
wire \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.u1.s ;
wire \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.u2.a ;
wire \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.u2.b ;
wire \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.u2.cin ;
wire \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.u2.cout ;
wire \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.u2.s ;
wire \add_3ns_3ns_3_2_1_U9.ce ;
wire \add_3ns_3ns_3_2_1_U9.clk ;
wire [2:0] \add_3ns_3ns_3_2_1_U9.din0 ;
wire [2:0] \add_3ns_3ns_3_2_1_U9.din1 ;
wire [2:0] \add_3ns_3ns_3_2_1_U9.dout ;
wire \add_3ns_3ns_3_2_1_U9.reset ;
wire [2:0] \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.a ;
wire [2:0] \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.ain_s0 ;
wire [2:0] \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.b ;
wire [2:0] \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.bin_s0 ;
wire \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.ce ;
wire \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.clk ;
wire \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.facout_s1 ;
wire \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.facout_s2 ;
wire \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.fas_s1 ;
wire [1:0] \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.fas_s2 ;
wire \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.reset ;
wire [2:0] \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.s ;
wire \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.u1.a ;
wire \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.u1.b ;
wire \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.u1.cin ;
wire \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.u1.cout ;
wire \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.u1.s ;
wire [1:0] \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.u2.a ;
wire [1:0] \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.u2.b ;
wire \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.u2.cin ;
wire \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.u2.cout ;
wire [1:0] \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.u2.s ;
wire \add_4ns_4ns_4_2_1_U1.ce ;
wire \add_4ns_4ns_4_2_1_U1.clk ;
wire [3:0] \add_4ns_4ns_4_2_1_U1.din0 ;
wire [3:0] \add_4ns_4ns_4_2_1_U1.din1 ;
wire [3:0] \add_4ns_4ns_4_2_1_U1.dout ;
wire \add_4ns_4ns_4_2_1_U1.reset ;
wire [3:0] \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.a ;
wire [3:0] \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.ain_s0 ;
wire [3:0] \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.b ;
wire [3:0] \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.bin_s0 ;
wire \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.ce ;
wire \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.clk ;
wire \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.facout_s1 ;
wire \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.facout_s2 ;
wire [1:0] \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.fas_s1 ;
wire [1:0] \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.fas_s2 ;
wire \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.reset ;
wire [3:0] \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.s ;
wire [1:0] \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.u1.a ;
wire [1:0] \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.u1.b ;
wire \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.u1.cin ;
wire \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.u1.cout ;
wire [1:0] \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.u1.s ;
wire [1:0] \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.u2.a ;
wire [1:0] \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.u2.b ;
wire \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.u2.cin ;
wire \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.u2.cout ;
wire [1:0] \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.u2.s ;
wire \add_4ns_4s_4_2_1_U11.ce ;
wire \add_4ns_4s_4_2_1_U11.clk ;
wire [3:0] \add_4ns_4s_4_2_1_U11.din0 ;
wire [3:0] \add_4ns_4s_4_2_1_U11.din1 ;
wire [3:0] \add_4ns_4s_4_2_1_U11.dout ;
wire \add_4ns_4s_4_2_1_U11.reset ;
wire [3:0] \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.a ;
wire [3:0] \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.ain_s0 ;
wire [3:0] \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.b ;
wire [3:0] \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.bin_s0 ;
wire \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.ce ;
wire \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.clk ;
wire \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.facout_s1 ;
wire \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.facout_s2 ;
wire [1:0] \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.fas_s1 ;
wire [1:0] \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.fas_s2 ;
wire \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.reset ;
wire [3:0] \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.s ;
wire [1:0] \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.u1.a ;
wire [1:0] \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.u1.b ;
wire \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.u1.cin ;
wire \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.u1.cout ;
wire [1:0] \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.u1.s ;
wire [1:0] \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.u2.a ;
wire [1:0] \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.u2.b ;
wire \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.u2.cin ;
wire \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.u2.cout ;
wire [1:0] \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.u2.s ;
wire \add_5s_5ns_5_2_1_U16.ce ;
wire \add_5s_5ns_5_2_1_U16.clk ;
wire [4:0] \add_5s_5ns_5_2_1_U16.din0 ;
wire [4:0] \add_5s_5ns_5_2_1_U16.din1 ;
wire [4:0] \add_5s_5ns_5_2_1_U16.dout ;
wire \add_5s_5ns_5_2_1_U16.reset ;
wire [4:0] \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.a ;
wire [4:0] \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.ain_s0 ;
wire [4:0] \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.b ;
wire [4:0] \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.bin_s0 ;
wire \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.ce ;
wire \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.clk ;
wire \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.facout_s1 ;
wire \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.facout_s2 ;
wire [1:0] \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.fas_s1 ;
wire [2:0] \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.fas_s2 ;
wire \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.reset ;
wire [4:0] \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.s ;
wire [1:0] \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.u1.a ;
wire [1:0] \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.u1.b ;
wire \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.u1.cin ;
wire \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.u1.cout ;
wire [1:0] \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.u1.s ;
wire [2:0] \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.u2.a ;
wire [2:0] \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.u2.b ;
wire \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.u2.cin ;
wire \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.u2.cout ;
wire [2:0] \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.u2.s ;
wire \add_9ns_9s_9_2_1_U2.ce ;
wire \add_9ns_9s_9_2_1_U2.clk ;
wire [8:0] \add_9ns_9s_9_2_1_U2.din0 ;
wire [8:0] \add_9ns_9s_9_2_1_U2.din1 ;
wire [8:0] \add_9ns_9s_9_2_1_U2.dout ;
wire \add_9ns_9s_9_2_1_U2.reset ;
wire [8:0] \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.a ;
wire [8:0] \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.ain_s0 ;
wire [8:0] \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.b ;
wire [8:0] \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.bin_s0 ;
wire \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.ce ;
wire \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.clk ;
wire \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.facout_s1 ;
wire \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.facout_s2 ;
wire [3:0] \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.fas_s1 ;
wire [4:0] \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.fas_s2 ;
wire \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.reset ;
wire [8:0] \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.s ;
wire [3:0] \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.u1.a ;
wire [3:0] \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.u1.b ;
wire \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.u1.cin ;
wire \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.u1.cout ;
wire [3:0] \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.u1.s ;
wire [4:0] \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.u2.a ;
wire [4:0] \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.u2.b ;
wire \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.u2.cin ;
wire \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.u2.cout ;
wire [4:0] \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.u2.s ;
wire and_ln781_1_fu_320_p2;
wire and_ln781_fu_324_p2;
wire and_ln785_1_fu_448_p2;
wire and_ln785_fu_439_p2;
wire and_ln786_1_fu_340_p2;
wire and_ln786_fu_345_p2;
wire ap_CS_fsm_state1;
wire ap_CS_fsm_state10;
wire ap_CS_fsm_state11;
wire ap_CS_fsm_state12;
wire ap_CS_fsm_state13;
wire ap_CS_fsm_state14;
wire ap_CS_fsm_state15;
wire ap_CS_fsm_state16;
wire ap_CS_fsm_state17;
wire ap_CS_fsm_state18;
wire ap_CS_fsm_state19;
wire ap_CS_fsm_state2;
wire ap_CS_fsm_state20;
wire ap_CS_fsm_state21;
wire ap_CS_fsm_state22;
wire ap_CS_fsm_state23;
wire ap_CS_fsm_state3;
wire ap_CS_fsm_state4;
wire ap_CS_fsm_state5;
wire ap_CS_fsm_state6;
wire ap_CS_fsm_state7;
wire ap_CS_fsm_state8;
wire ap_CS_fsm_state9;
wire [22:0] ap_NS_fsm;
wire ap_clk;
wire ap_done;
wire ap_idle;
wire ap_ready;
wire ap_rst;
wire ap_start;
wire deleted_zeros_fu_298_p2;
wire [3:0] grp_fu_235_p0;
wire [3:0] grp_fu_235_p1;
wire [3:0] grp_fu_235_p2;
wire [8:0] grp_fu_293_p1;
wire [8:0] grp_fu_293_p2;
wire [16:0] grp_fu_376_p0;
wire [16:0] grp_fu_376_p1;
wire [16:0] grp_fu_376_p2;
wire [1:0] grp_fu_420_p2;
wire [12:0] grp_fu_478_p2;
wire [4:0] grp_fu_495_p2;
wire [1:0] grp_fu_593_p2;
wire [13:0] grp_fu_613_p0;
wire [13:0] grp_fu_613_p1;
wire [13:0] grp_fu_613_p2;
wire [2:0] grp_fu_619_p0;
wire [2:0] grp_fu_619_p1;
wire [2:0] grp_fu_619_p2;
wire [13:0] grp_fu_654_p2;
wire [3:0] grp_fu_661_p0;
wire [3:0] grp_fu_661_p1;
wire [3:0] grp_fu_661_p2;
wire [13:0] grp_fu_670_p0;
wire [13:0] grp_fu_670_p2;
wire [14:0] grp_fu_694_p0;
wire [14:0] grp_fu_694_p1;
wire [14:0] grp_fu_694_p2;
wire [14:0] grp_fu_717_p0;
wire [14:0] grp_fu_717_p1;
wire [14:0] grp_fu_717_p2;
wire [17:0] grp_fu_740_p0;
wire [17:0] grp_fu_740_p1;
wire [17:0] grp_fu_740_p2;
wire [4:0] grp_fu_746_p0;
wire [4:0] grp_fu_746_p1;
wire [4:0] grp_fu_746_p2;
wire [17:0] grp_fu_755_p0;
wire [17:0] grp_fu_755_p2;
wire icmp_ln851_1_fu_473_p2;
wire icmp_ln851_2_fu_253_p2;
wire icmp_ln851_3_fu_588_p2;
wire icmp_ln851_fu_199_p2;
wire neg_src_fu_335_p2;
wire [15:0] op_0;
wire op_1;
wire [3:0] op_12;
wire op_13;
wire [1:0] op_14;
wire [1:0] op_16;
wire [3:0] op_17;
wire [7:0] op_2;
wire op_3;
wire [31:0] op_30;
wire op_30_ap_vld;
wire [3:0] op_6_V_fu_453_p3;
wire [3:0] op_9;
wire or_ln340_1_fu_408_p2;
wire or_ln340_fu_403_p2;
wire or_ln778_fu_285_p2;
wire or_ln780_fu_315_p2;
wire or_ln785_1_fu_443_p2;
wire or_ln785_fu_387_p2;
wire overflow_fu_397_p2;
wire p_Result_1_fu_536_p3;
wire p_Result_2_fu_569_p3;
wire [7:0] p_Result_3_fu_187_p1;
wire [7:0] p_Result_4_fu_215_p1;
wire p_Result_s_fu_625_p3;
wire [7:0] p_Val2_2_fu_205_p1;
wire p_Val2_s_fu_675_p1;
wire [1:0] p_Val2_s_fu_675_p3;
wire [1:0] ret_V_18_fu_548_p3;
wire [12:0] ret_V_20_fu_581_p3;
wire [1:0] ret_V_22_fu_637_p3;
wire [4:0] ret_V_23_fu_520_p2;
wire ret_V_9_fu_483_p2;
wire [4:0] rhs_2_fu_512_p3;
wire [4:0] rhs_fu_364_p3;
wire select_ln1192_fu_267_p0;
wire [8:0] select_ln1192_fu_267_p3;
wire [3:0] select_ln340_fu_413_p3;
wire [1:0] select_ln353_fu_506_p3;
wire select_ln69_fu_644_p0;
wire [7:0] select_ln69_fu_644_p3;
wire select_ln703_fu_466_p0;
wire [4:0] select_ln703_fu_466_p3;
wire [1:0] select_ln831_fu_459_p3;
wire [12:0] select_ln850_1_fu_576_p3;
wire [1:0] select_ln850_3_fu_632_p3;
wire [1:0] select_ln850_6_fu_500_p3;
wire [1:0] select_ln850_fu_543_p3;
wire [15:0] sext_ln69_2_fu_730_p1;
wire [4:0] sext_ln703_2_fu_492_p1;
wire [7:0] sext_ln703_fu_290_p0;
wire \sub_5ns_5s_5_2_1_U6.ce ;
wire \sub_5ns_5s_5_2_1_U6.clk ;
wire [4:0] \sub_5ns_5s_5_2_1_U6.din0 ;
wire [4:0] \sub_5ns_5s_5_2_1_U6.din1 ;
wire [4:0] \sub_5ns_5s_5_2_1_U6.dout ;
wire \sub_5ns_5s_5_2_1_U6.reset ;
wire [4:0] \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.a ;
wire [4:0] \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.ain_s0 ;
wire [4:0] \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.b ;
wire [4:0] \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.bin_s0 ;
wire \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.ce ;
wire \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.clk ;
wire \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.facout_s1 ;
wire \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.facout_s2 ;
wire [1:0] \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.fas_s1 ;
wire [2:0] \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.fas_s2 ;
wire \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.reset ;
wire [4:0] \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.s ;
wire [1:0] \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.u1.a ;
wire [1:0] \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.u1.b ;
wire \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.u1.cin ;
wire \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.u1.cout ;
wire [1:0] \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.u1.s ;
wire [2:0] \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.u2.a ;
wire [2:0] \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.u2.b ;
wire \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.u2.cin ;
wire \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.u2.cout ;
wire [2:0] \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.u2.s ;
wire [7:0] tmp_6_fu_223_p1;
wire tmp_6_fu_223_p3;
wire [7:0] tmp_9_fu_302_p1;
wire tmp_9_fu_302_p3;
wire [7:0] trunc_ln1192_fu_195_p0;
wire [6:0] trunc_ln1192_fu_195_p1;
wire [7:0] trunc_ln851_1_fu_249_p0;
wire [6:0] trunc_ln851_1_fu_249_p1;
wire [2:0] trunc_ln851_2_fu_565_p1;
wire [3:0] trunc_ln851_fu_435_p1;
wire xor_ln416_fu_275_p2;
wire xor_ln778_fu_280_p2;
wire xor_ln780_fu_309_p2;
wire xor_ln781_fu_329_p2;
wire xor_ln785_1_fu_392_p2;
wire xor_ln785_fu_382_p2;
wire [1:0] zext_ln831_fu_488_p1;


assign _046_ = _049_ & ap_CS_fsm[6];
assign _047_ = _050_ & ap_CS_fsm[0];
assign _048_ = ap_start & ap_CS_fsm[0];
assign and_ln781_1_fu_320_p2 = xor_ln416_reg_839 & Range2_all_ones_reg_800;
assign and_ln781_fu_324_p2 = p_Result_4_reg_789 & and_ln781_1_fu_320_p2;
assign and_ln785_1_fu_448_p2 = or_ln785_1_fu_443_p2 & and_ln786_reg_867;
assign and_ln785_fu_439_p2 = xor_ln416_reg_839 & deleted_zeros_reg_856;
assign and_ln786_1_fu_340_p2 = p_Result_5_reg_820 & or_ln780_fu_315_p2;
assign and_ln786_fu_345_p2 = and_ln786_1_fu_340_p2 & Range2_all_ones_reg_800;
assign neg_src_fu_335_p2 = xor_ln781_fu_329_p2 & p_Result_3_reg_771;
assign overflow_fu_397_p2 = xor_ln785_1_fu_392_p2 & or_ln785_fu_387_p2;
assign ret_V_23_fu_520_p2 = { op_6_V_reg_917[3], op_6_V_reg_917 } & { select_ln353_fu_506_p3, 3'h0 };
assign xor_ln780_fu_309_p2 = ~ op_2[7];
assign xor_ln781_fu_329_p2 = ~ and_ln781_fu_324_p2;
assign xor_ln785_fu_382_p2 = ~ deleted_zeros_reg_856;
assign xor_ln785_1_fu_392_p2 = ~ p_Result_3_reg_771;
assign xor_ln778_fu_280_p2 = ~ p_Result_4_reg_789;
assign ret_V_9_fu_483_p2 = ~ Range2_all_ones_reg_800;
assign xor_ln416_fu_275_p2 = ~ p_Result_5_reg_820;
assign _049_ = ~ icmp_ln851_reg_779;
assign _050_ = ~ ap_start;
assign _051_ = ! trunc_ln851_reg_912;
assign _052_ = ! op_2[6:0];
assign _053_ = ! trunc_ln851_2_reg_975;
always @(posedge \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.clk )
\add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.bin_s1  <= _055_;
always @(posedge \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.clk )
\add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.ain_s1  <= _054_;
always @(posedge \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.clk )
\add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.sum_s1  <= _057_;
always @(posedge \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.clk )
\add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.carry_s1  <= _056_;
assign _055_ = \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.ce  ? \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.b [12:6] : \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.bin_s1 ;
assign _054_ = \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.ce  ? \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.a [12:6] : \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.ain_s1 ;
assign _056_ = \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.ce  ? \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.facout_s1  : \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.carry_s1 ;
assign _057_ = \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.ce  ? \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.fas_s1  : \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.sum_s1 ;
assign _058_ = \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.u1.a  + \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.u1.b ;
assign { \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.u1.cout , \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.u1.s  } = _058_ + \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.u1.cin ;
assign _059_ = \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.u2.a  + \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.u2.b ;
assign { \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.u2.cout , \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.u2.s  } = _059_ + \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.u2.cin ;
always @(posedge \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.clk )
\add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.bin_s1  <= _061_;
always @(posedge \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.clk )
\add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.ain_s1  <= _060_;
always @(posedge \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.clk )
\add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.sum_s1  <= _063_;
always @(posedge \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.clk )
\add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.carry_s1  <= _062_;
assign _061_ = \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.ce  ? \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.b [13:7] : \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.bin_s1 ;
assign _060_ = \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.ce  ? \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.a [13:7] : \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.ain_s1 ;
assign _062_ = \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.ce  ? \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.facout_s1  : \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.carry_s1 ;
assign _063_ = \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.ce  ? \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.fas_s1  : \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.sum_s1 ;
assign _064_ = \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.u1.a  + \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.u1.b ;
assign { \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.u1.cout , \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.u1.s  } = _064_ + \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.u1.cin ;
assign _065_ = \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.u2.a  + \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.u2.b ;
assign { \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.u2.cout , \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.u2.s  } = _065_ + \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.u2.cin ;
always @(posedge \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.clk )
\add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.bin_s1  <= _067_;
always @(posedge \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.clk )
\add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.ain_s1  <= _066_;
always @(posedge \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.clk )
\add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.sum_s1  <= _069_;
always @(posedge \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.clk )
\add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.carry_s1  <= _068_;
assign _067_ = \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.ce  ? \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.b [13:7] : \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.bin_s1 ;
assign _066_ = \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.ce  ? \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.a [13:7] : \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.ain_s1 ;
assign _068_ = \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.ce  ? \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.facout_s1  : \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.carry_s1 ;
assign _069_ = \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.ce  ? \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.fas_s1  : \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.sum_s1 ;
assign _070_ = \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.u1.a  + \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.u1.b ;
assign { \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.u1.cout , \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.u1.s  } = _070_ + \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.u1.cin ;
assign _071_ = \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.u2.a  + \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.u2.b ;
assign { \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.u2.cout , \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.u2.s  } = _071_ + \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.u2.cin ;
always @(posedge \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.clk )
\add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.bin_s1  <= _073_;
always @(posedge \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.clk )
\add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.ain_s1  <= _072_;
always @(posedge \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.clk )
\add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.sum_s1  <= _075_;
always @(posedge \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.clk )
\add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.carry_s1  <= _074_;
assign _073_ = \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.ce  ? \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.b [13:7] : \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.bin_s1 ;
assign _072_ = \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.ce  ? \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.a [13:7] : \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.ain_s1 ;
assign _074_ = \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.ce  ? \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.facout_s1  : \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.carry_s1 ;
assign _075_ = \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.ce  ? \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.fas_s1  : \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.sum_s1 ;
assign _076_ = \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.u1.a  + \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.u1.b ;
assign { \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.u1.cout , \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.u1.s  } = _076_ + \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.u1.cin ;
assign _077_ = \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.u2.a  + \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.u2.b ;
assign { \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.u2.cout , \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.u2.s  } = _077_ + \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.u2.cin ;
always @(posedge \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.clk )
\add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.bin_s1  <= _079_;
always @(posedge \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.clk )
\add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.ain_s1  <= _078_;
always @(posedge \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.clk )
\add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.sum_s1  <= _081_;
always @(posedge \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.clk )
\add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.carry_s1  <= _080_;
assign _079_ = \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.ce  ? \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.b [14:7] : \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.bin_s1 ;
assign _078_ = \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.ce  ? \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.a [14:7] : \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.ain_s1 ;
assign _080_ = \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.ce  ? \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.facout_s1  : \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.carry_s1 ;
assign _081_ = \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.ce  ? \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.fas_s1  : \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.sum_s1 ;
assign _082_ = \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.u1.a  + \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.u1.b ;
assign { \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.u1.cout , \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.u1.s  } = _082_ + \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.u1.cin ;
assign _083_ = \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.u2.a  + \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.u2.b ;
assign { \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.u2.cout , \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.u2.s  } = _083_ + \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.u2.cin ;
always @(posedge \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.clk )
\add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.bin_s1  <= _085_;
always @(posedge \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.clk )
\add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.ain_s1  <= _084_;
always @(posedge \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.clk )
\add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.sum_s1  <= _087_;
always @(posedge \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.clk )
\add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.carry_s1  <= _086_;
assign _085_ = \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.ce  ? \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.b [14:7] : \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.bin_s1 ;
assign _084_ = \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.ce  ? \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.a [14:7] : \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.ain_s1 ;
assign _086_ = \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.ce  ? \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.facout_s1  : \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.carry_s1 ;
assign _087_ = \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.ce  ? \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.fas_s1  : \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.sum_s1 ;
assign _088_ = \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.u1.a  + \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.u1.b ;
assign { \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.u1.cout , \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.u1.s  } = _088_ + \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.u1.cin ;
assign _089_ = \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.u2.a  + \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.u2.b ;
assign { \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.u2.cout , \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.u2.s  } = _089_ + \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.u2.cin ;
always @(posedge \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.clk )
\add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.bin_s1  <= _091_;
always @(posedge \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.clk )
\add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.ain_s1  <= _090_;
always @(posedge \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.clk )
\add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.sum_s1  <= _093_;
always @(posedge \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.clk )
\add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.carry_s1  <= _092_;
assign _091_ = \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.ce  ? \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.b [16:8] : \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.bin_s1 ;
assign _090_ = \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.ce  ? \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.a [16:8] : \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.ain_s1 ;
assign _092_ = \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.ce  ? \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.facout_s1  : \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.carry_s1 ;
assign _093_ = \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.ce  ? \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.fas_s1  : \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.sum_s1 ;
assign _094_ = \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.u1.a  + \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.u1.b ;
assign { \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.u1.cout , \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.u1.s  } = _094_ + \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.u1.cin ;
assign _095_ = \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.u2.a  + \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.u2.b ;
assign { \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.u2.cout , \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.u2.s  } = _095_ + \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.u2.cin ;
always @(posedge \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.clk )
\add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.bin_s1  <= _097_;
always @(posedge \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.clk )
\add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.ain_s1  <= _096_;
always @(posedge \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.clk )
\add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.sum_s1  <= _099_;
always @(posedge \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.clk )
\add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.carry_s1  <= _098_;
assign _097_ = \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.ce  ? \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.b [17:9] : \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.bin_s1 ;
assign _096_ = \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.ce  ? \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.a [17:9] : \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.ain_s1 ;
assign _098_ = \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.ce  ? \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.facout_s1  : \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.carry_s1 ;
assign _099_ = \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.ce  ? \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.fas_s1  : \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.sum_s1 ;
assign _100_ = \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.u1.a  + \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.u1.b ;
assign { \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.u1.cout , \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.u1.s  } = _100_ + \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.u1.cin ;
assign _101_ = \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.u2.a  + \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.u2.b ;
assign { \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.u2.cout , \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.u2.s  } = _101_ + \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.u2.cin ;
always @(posedge \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.clk )
\add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.bin_s1  <= _103_;
always @(posedge \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.clk )
\add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.ain_s1  <= _102_;
always @(posedge \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.clk )
\add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.sum_s1  <= _105_;
always @(posedge \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.clk )
\add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.carry_s1  <= _104_;
assign _103_ = \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.ce  ? \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.b [17:9] : \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.bin_s1 ;
assign _102_ = \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.ce  ? \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.a [17:9] : \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.ain_s1 ;
assign _104_ = \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.ce  ? \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.facout_s1  : \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.carry_s1 ;
assign _105_ = \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.ce  ? \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.fas_s1  : \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.sum_s1 ;
assign _106_ = \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.u1.a  + \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.u1.b ;
assign { \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.u1.cout , \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.u1.s  } = _106_ + \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.u1.cin ;
assign _107_ = \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.u2.a  + \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.u2.b ;
assign { \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.u2.cout , \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.u2.s  } = _107_ + \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.u2.cin ;
always @(posedge \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.clk )
\add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.bin_s1  <= _109_;
always @(posedge \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.clk )
\add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.ain_s1  <= _108_;
always @(posedge \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.clk )
\add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.sum_s1  <= _111_;
always @(posedge \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.clk )
\add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.carry_s1  <= _110_;
assign _109_ = \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.ce  ? \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.b [1] : \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.bin_s1 ;
assign _108_ = \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.ce  ? \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.a [1] : \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.ain_s1 ;
assign _110_ = \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.ce  ? \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.facout_s1  : \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.carry_s1 ;
assign _111_ = \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.ce  ? \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.fas_s1  : \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.sum_s1 ;
assign _112_ = \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.u1.a  + \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.u1.b ;
assign { \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.u1.cout , \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.u1.s  } = _112_ + \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.u1.cin ;
assign _113_ = \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.u2.a  + \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.u2.b ;
assign { \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.u2.cout , \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.u2.s  } = _113_ + \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.u2.cin ;
always @(posedge \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.clk )
\add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.bin_s1  <= _115_;
always @(posedge \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.clk )
\add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.ain_s1  <= _114_;
always @(posedge \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.clk )
\add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.sum_s1  <= _117_;
always @(posedge \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.clk )
\add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.carry_s1  <= _116_;
assign _115_ = \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.ce  ? \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.b [1] : \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.bin_s1 ;
assign _114_ = \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.ce  ? \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.a [1] : \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.ain_s1 ;
assign _116_ = \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.ce  ? \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.facout_s1  : \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.carry_s1 ;
assign _117_ = \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.ce  ? \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.fas_s1  : \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.sum_s1 ;
assign _118_ = \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.u1.a  + \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.u1.b ;
assign { \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.u1.cout , \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.u1.s  } = _118_ + \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.u1.cin ;
assign _119_ = \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.u2.a  + \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.u2.b ;
assign { \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.u2.cout , \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.u2.s  } = _119_ + \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.u2.cin ;
always @(posedge \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.clk )
\add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.bin_s1  <= _121_;
always @(posedge \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.clk )
\add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.ain_s1  <= _120_;
always @(posedge \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.clk )
\add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.sum_s1  <= _123_;
always @(posedge \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.clk )
\add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.carry_s1  <= _122_;
assign _121_ = \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.ce  ? \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.b [2:1] : \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.bin_s1 ;
assign _120_ = \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.ce  ? \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.a [2:1] : \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.ain_s1 ;
assign _122_ = \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.ce  ? \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.facout_s1  : \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.carry_s1 ;
assign _123_ = \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.ce  ? \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.fas_s1  : \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.sum_s1 ;
assign _124_ = \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.u1.a  + \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.u1.b ;
assign { \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.u1.cout , \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.u1.s  } = _124_ + \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.u1.cin ;
assign _125_ = \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.u2.a  + \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.u2.b ;
assign { \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.u2.cout , \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.u2.s  } = _125_ + \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.u2.cin ;
always @(posedge \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.clk )
\add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.bin_s1  <= _127_;
always @(posedge \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.clk )
\add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.ain_s1  <= _126_;
always @(posedge \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.clk )
\add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.sum_s1  <= _129_;
always @(posedge \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.clk )
\add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.carry_s1  <= _128_;
assign _127_ = \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.ce  ? \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.b [3:2] : \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.bin_s1 ;
assign _126_ = \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.ce  ? \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.a [3:2] : \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.ain_s1 ;
assign _128_ = \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.ce  ? \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.facout_s1  : \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.carry_s1 ;
assign _129_ = \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.ce  ? \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.fas_s1  : \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.sum_s1 ;
assign _130_ = \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.u1.a  + \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.u1.b ;
assign { \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.u1.cout , \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.u1.s  } = _130_ + \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.u1.cin ;
assign _131_ = \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.u2.a  + \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.u2.b ;
assign { \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.u2.cout , \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.u2.s  } = _131_ + \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.u2.cin ;
always @(posedge \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.clk )
\add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.bin_s1  <= _133_;
always @(posedge \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.clk )
\add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.ain_s1  <= _132_;
always @(posedge \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.clk )
\add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.sum_s1  <= _135_;
always @(posedge \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.clk )
\add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.carry_s1  <= _134_;
assign _133_ = \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.ce  ? \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.b [3:2] : \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.bin_s1 ;
assign _132_ = \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.ce  ? \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.a [3:2] : \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.ain_s1 ;
assign _134_ = \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.ce  ? \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.facout_s1  : \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.carry_s1 ;
assign _135_ = \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.ce  ? \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.fas_s1  : \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.sum_s1 ;
assign _136_ = \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.u1.a  + \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.u1.b ;
assign { \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.u1.cout , \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.u1.s  } = _136_ + \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.u1.cin ;
assign _137_ = \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.u2.a  + \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.u2.b ;
assign { \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.u2.cout , \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.u2.s  } = _137_ + \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.u2.cin ;
always @(posedge \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.clk )
\add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.bin_s1  <= _139_;
always @(posedge \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.clk )
\add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.ain_s1  <= _138_;
always @(posedge \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.clk )
\add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.sum_s1  <= _141_;
always @(posedge \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.clk )
\add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.carry_s1  <= _140_;
assign _139_ = \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.ce  ? \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.b [4:2] : \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.bin_s1 ;
assign _138_ = \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.ce  ? \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.a [4:2] : \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.ain_s1 ;
assign _140_ = \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.ce  ? \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.facout_s1  : \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.carry_s1 ;
assign _141_ = \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.ce  ? \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.fas_s1  : \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.sum_s1 ;
assign _142_ = \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.u1.a  + \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.u1.b ;
assign { \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.u1.cout , \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.u1.s  } = _142_ + \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.u1.cin ;
assign _143_ = \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.u2.a  + \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.u2.b ;
assign { \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.u2.cout , \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.u2.s  } = _143_ + \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.u2.cin ;
always @(posedge \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.clk )
\add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.bin_s1  <= _145_;
always @(posedge \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.clk )
\add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.ain_s1  <= _144_;
always @(posedge \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.clk )
\add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.sum_s1  <= _147_;
always @(posedge \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.clk )
\add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.carry_s1  <= _146_;
assign _145_ = \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.ce  ? \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.b [8:4] : \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.bin_s1 ;
assign _144_ = \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.ce  ? \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.a [8:4] : \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.ain_s1 ;
assign _146_ = \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.ce  ? \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.facout_s1  : \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.carry_s1 ;
assign _147_ = \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.ce  ? \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.fas_s1  : \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.sum_s1 ;
assign _148_ = \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.u1.a  + \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.u1.b ;
assign { \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.u1.cout , \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.u1.s  } = _148_ + \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.u1.cin ;
assign _149_ = \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.u2.a  + \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.u2.b ;
assign { \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.u2.cout , \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.u2.s  } = _149_ + \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.u2.cin ;
assign \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.bin_s0  = ~ \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.b ;
always @(posedge \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.clk )
\sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.bin_s1  <= _151_;
always @(posedge \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.clk )
\sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.ain_s1  <= _150_;
always @(posedge \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.clk )
\sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.sum_s1  <= _153_;
always @(posedge \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.clk )
\sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.carry_s1  <= _152_;
assign _151_ = \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.ce  ? \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.bin_s0 [4:2] : \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.bin_s1 ;
assign _150_ = \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.ce  ? \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.a [4:2] : \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.ain_s1 ;
assign _152_ = \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.ce  ? \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.facout_s1  : \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.carry_s1 ;
assign _153_ = \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.ce  ? \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.fas_s1  : \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.sum_s1 ;
assign _154_ = \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.u1.a  + \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.u1.b ;
assign { \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.u1.cout , \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.u1.s  } = _154_ + \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.u1.cin ;
assign _155_ = \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.u2.a  + \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.u2.b ;
assign { \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.u2.cout , \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.u2.s  } = _155_ + \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.u2.cin ;
assign or_ln340_1_fu_408_p2 = or_ln340_fu_403_p2 | neg_src_reg_862;
assign or_ln340_fu_403_p2 = overflow_fu_397_p2 | and_ln786_reg_867;
assign or_ln778_fu_285_p2 = xor_ln778_fu_280_p2 | p_Result_5_reg_820;
assign or_ln780_fu_315_p2 = xor_ln780_fu_309_p2 | or_ln778_reg_845;
assign or_ln785_1_fu_443_p2 = p_Result_3_reg_771 | and_ln785_fu_439_p2;
assign or_ln785_fu_387_p2 = xor_ln785_fu_382_p2 | p_Result_5_reg_820;
always @(posedge ap_clk)
select_ln1192_reg_834[6:0] <= 7'h00;
always @(posedge ap_clk)
select_ln703_reg_928[2:0] <= 3'h0;
always @(posedge ap_clk)
select_ln69_reg_1020[13:8] <= 6'h00;
always @(posedge ap_clk)
ret_V_2_reg_933 <= _032_;
always @(posedge ap_clk)
ret_V_24_reg_1090 <= _031_;
always @(posedge ap_clk)
ret_V_17_reg_873 <= _025_;
always @(posedge ap_clk)
ret_V_reg_878 <= _035_;
always @(posedge ap_clk)
select_ln340_reg_895 <= _037_;
always @(posedge ap_clk)
ret_V_12_reg_995 <= _024_;
always @(posedge ap_clk)
ret_V_18_reg_953 <= _026_;
always @(posedge ap_clk)
ret_V_6_reg_958 <= _034_;
always @(posedge ap_clk)
ret_V_21_reg_963 <= _029_;
always @(posedge ap_clk)
ret_V_11_reg_968 <= _023_;
always @(posedge ap_clk)
trunc_ln851_2_reg_975 <= _042_;
always @(posedge ap_clk)
p_Val2_3_reg_814 <= _022_;
always @(posedge ap_clk)
p_Result_5_reg_820 <= _021_;
always @(posedge ap_clk)
select_ln1192_reg_834[8:7] <= _036_;
always @(posedge ap_clk)
xor_ln416_reg_839 <= _044_;
always @(posedge ap_clk)
or_ln778_reg_845 <= _018_;
always @(posedge ap_clk)
ret_V_19_reg_900 <= _027_;
always @(posedge ap_clk)
ret_V_4_reg_905 <= _033_;
always @(posedge ap_clk)
trunc_ln851_reg_912 <= _043_;
always @(posedge ap_clk)
op_6_V_reg_917 <= _017_;
always @(posedge ap_clk)
select_ln831_reg_922 <= _040_;
always @(posedge ap_clk)
select_ln703_reg_928[4:3] <= _039_;
always @(posedge ap_clk)
op_26_V_reg_1075 <= _016_;
always @(posedge ap_clk)
op_25_V_reg_1060 <= _015_;
always @(posedge ap_clk)
ret_V_20_reg_980 <= _028_;
always @(posedge ap_clk)
icmp_ln851_3_reg_985 <= _012_;
always @(posedge ap_clk)
icmp_ln851_1_reg_938 <= _010_;
always @(posedge ap_clk)
tmp_reg_948 <= _041_;
always @(posedge ap_clk)
deleted_zeros_reg_856 <= _009_;
always @(posedge ap_clk)
neg_src_reg_862 <= _014_;
always @(posedge ap_clk)
and_ln786_reg_867 <= _007_;
always @(posedge ap_clk)
add_ln69_5_reg_1115 <= _004_;
always @(posedge ap_clk)
add_ln69_7_reg_1120 <= _005_;
always @(posedge ap_clk)
ret_V_22_reg_1015 <= _030_;
always @(posedge ap_clk)
select_ln69_reg_1020[7:0] <= _038_;
always @(posedge ap_clk)
add_ln69_reg_1025 <= _006_;
always @(posedge ap_clk)
add_ln69_2_reg_1030 <= _002_;
always @(posedge ap_clk)
add_ln69_1_reg_1045 <= _001_;
always @(posedge ap_clk)
add_ln69_3_reg_1050 <= _003_;
always @(posedge ap_clk)
p_Result_3_reg_771 <= _019_;
always @(posedge ap_clk)
icmp_ln851_reg_779 <= _013_;
always @(posedge ap_clk)
p_Result_4_reg_789 <= _020_;
always @(posedge ap_clk)
Range2_all_ones_reg_800 <= _000_;
always @(posedge ap_clk)
icmp_ln851_2_reg_809 <= _011_;
always @(posedge ap_clk)
ap_CS_fsm <= _008_;
assign _045_ = _048_ ? 2'h2 : 2'h1;
assign _156_ = ap_CS_fsm == 1'h1;
function [22:0] _464_;
input [22:0] a;
input [528:0] b;
input [22:0] s;
case (s)
23'b00000000000000000000001:
_464_ = b[22:0];
23'b00000000000000000000010:
_464_ = b[45:23];
23'b00000000000000000000100:
_464_ = b[68:46];
23'b00000000000000000001000:
_464_ = b[91:69];
23'b00000000000000000010000:
_464_ = b[114:92];
23'b00000000000000000100000:
_464_ = b[137:115];
23'b00000000000000001000000:
_464_ = b[160:138];
23'b00000000000000010000000:
_464_ = b[183:161];
23'b00000000000000100000000:
_464_ = b[206:184];
23'b00000000000001000000000:
_464_ = b[229:207];
23'b00000000000010000000000:
_464_ = b[252:230];
23'b00000000000100000000000:
_464_ = b[275:253];
23'b00000000001000000000000:
_464_ = b[298:276];
23'b00000000010000000000000:
_464_ = b[321:299];
23'b00000000100000000000000:
_464_ = b[344:322];
23'b00000001000000000000000:
_464_ = b[367:345];
23'b00000010000000000000000:
_464_ = b[390:368];
23'b00000100000000000000000:
_464_ = b[413:391];
23'b00001000000000000000000:
_464_ = b[436:414];
23'b00010000000000000000000:
_464_ = b[459:437];
23'b00100000000000000000000:
_464_ = b[482:460];
23'b01000000000000000000000:
_464_ = b[505:483];
23'b10000000000000000000000:
_464_ = b[528:506];
23'b00000000000000000000000:
_464_ = a;
default:
_464_ = 23'bx;
endcase
endfunction
assign ap_NS_fsm = _464_(23'hxxxxxx, { 21'h000000, _045_, 506'h0000020000080000200000800002000008000020000080000200000800002000008000020000080000200000800002000008000020000080000200000000001 }, { _156_, _178_, _177_, _176_, _175_, _174_, _173_, _172_, _171_, _170_, _169_, _168_, _167_, _166_, _165_, _164_, _163_, _162_, _161_, _160_, _159_, _158_, _157_ });
assign _157_ = ap_CS_fsm == 23'h400000;
assign _158_ = ap_CS_fsm == 22'h200000;
assign _159_ = ap_CS_fsm == 21'h100000;
assign _160_ = ap_CS_fsm == 20'h80000;
assign _161_ = ap_CS_fsm == 19'h40000;
assign _162_ = ap_CS_fsm == 18'h20000;
assign _163_ = ap_CS_fsm == 17'h10000;
assign _164_ = ap_CS_fsm == 16'h8000;
assign _165_ = ap_CS_fsm == 15'h4000;
assign _166_ = ap_CS_fsm == 14'h2000;
assign _167_ = ap_CS_fsm == 13'h1000;
assign _168_ = ap_CS_fsm == 12'h800;
assign _169_ = ap_CS_fsm == 11'h400;
assign _170_ = ap_CS_fsm == 10'h200;
assign _171_ = ap_CS_fsm == 9'h100;
assign _172_ = ap_CS_fsm == 8'h80;
assign _173_ = ap_CS_fsm == 7'h40;
assign _174_ = ap_CS_fsm == 6'h20;
assign _175_ = ap_CS_fsm == 5'h10;
assign _176_ = ap_CS_fsm == 4'h8;
assign _177_ = ap_CS_fsm == 3'h4;
assign _178_ = ap_CS_fsm == 2'h2;
assign op_30_ap_vld = ap_CS_fsm[22] ? 1'h1 : 1'h0;
assign ap_idle = _047_ ? 1'h1 : 1'h0;
assign _032_ = _046_ ? grp_fu_420_p2 : ret_V_2_reg_933;
assign _031_ = ap_CS_fsm[18] ? grp_fu_717_p2 : ret_V_24_reg_1090;
assign _037_ = ap_CS_fsm[4] ? select_ln340_fu_413_p3 : select_ln340_reg_895;
assign _035_ = ap_CS_fsm[4] ? grp_fu_293_p2[8:7] : ret_V_reg_878;
assign _025_ = ap_CS_fsm[4] ? grp_fu_293_p2 : ret_V_17_reg_873;
assign _024_ = ap_CS_fsm[9] ? grp_fu_593_p2 : ret_V_12_reg_995;
assign _042_ = ap_CS_fsm[7] ? grp_fu_495_p2[2:0] : trunc_ln851_2_reg_975;
assign _023_ = ap_CS_fsm[7] ? grp_fu_495_p2[4:3] : ret_V_11_reg_968;
assign _029_ = ap_CS_fsm[7] ? grp_fu_495_p2 : ret_V_21_reg_963;
assign _034_ = ap_CS_fsm[7] ? grp_fu_478_p2 : ret_V_6_reg_958;
assign _026_ = ap_CS_fsm[7] ? ret_V_18_fu_548_p3 : ret_V_18_reg_953;
assign _021_ = ap_CS_fsm[1] ? grp_fu_235_p2[3] : p_Result_5_reg_820;
assign _022_ = ap_CS_fsm[1] ? grp_fu_235_p2 : p_Val2_3_reg_814;
assign _018_ = ap_CS_fsm[2] ? or_ln778_fu_285_p2 : or_ln778_reg_845;
assign _044_ = ap_CS_fsm[2] ? xor_ln416_fu_275_p2 : xor_ln416_reg_839;
assign _036_ = ap_CS_fsm[2] ? select_ln1192_fu_267_p3[8:7] : select_ln1192_reg_834[8:7];
assign _039_ = ap_CS_fsm[5] ? select_ln703_fu_466_p3[4:3] : select_ln703_reg_928[4:3];
assign _040_ = ap_CS_fsm[5] ? select_ln831_fu_459_p3 : select_ln831_reg_922;
assign _017_ = ap_CS_fsm[5] ? op_6_V_fu_453_p3 : op_6_V_reg_917;
assign _043_ = ap_CS_fsm[5] ? grp_fu_376_p2[3:0] : trunc_ln851_reg_912;
assign _033_ = ap_CS_fsm[5] ? grp_fu_376_p2[16:4] : ret_V_4_reg_905;
assign _027_ = ap_CS_fsm[5] ? grp_fu_376_p2 : ret_V_19_reg_900;
assign _016_ = ap_CS_fsm[16] ? grp_fu_694_p2[14:1] : op_26_V_reg_1075;
assign _015_ = ap_CS_fsm[14] ? grp_fu_670_p2 : op_25_V_reg_1060;
assign _012_ = ap_CS_fsm[8] ? icmp_ln851_3_fu_588_p2 : icmp_ln851_3_reg_985;
assign _028_ = ap_CS_fsm[8] ? ret_V_20_fu_581_p3 : ret_V_20_reg_980;
assign _041_ = ap_CS_fsm[6] ? ret_V_23_fu_520_p2[4:3] : tmp_reg_948;
assign _010_ = ap_CS_fsm[6] ? icmp_ln851_1_fu_473_p2 : icmp_ln851_1_reg_938;
assign _007_ = ap_CS_fsm[3] ? and_ln786_fu_345_p2 : and_ln786_reg_867;
assign _014_ = ap_CS_fsm[3] ? neg_src_fu_335_p2 : neg_src_reg_862;
assign _009_ = ap_CS_fsm[3] ? deleted_zeros_fu_298_p2 : deleted_zeros_reg_856;
assign _005_ = ap_CS_fsm[20] ? grp_fu_746_p2 : add_ln69_7_reg_1120;
assign _004_ = ap_CS_fsm[20] ? grp_fu_740_p2 : add_ln69_5_reg_1115;
assign _002_ = ap_CS_fsm[10] ? grp_fu_619_p2 : add_ln69_2_reg_1030;
assign _006_ = ap_CS_fsm[10] ? grp_fu_613_p2 : add_ln69_reg_1025;
assign _038_ = ap_CS_fsm[10] ? select_ln69_fu_644_p3 : select_ln69_reg_1020[7:0];
assign _030_ = ap_CS_fsm[10] ? ret_V_22_fu_637_p3 : ret_V_22_reg_1015;
assign _003_ = ap_CS_fsm[12] ? grp_fu_661_p2 : add_ln69_3_reg_1050;
assign _001_ = ap_CS_fsm[12] ? grp_fu_654_p2 : add_ln69_1_reg_1045;
assign _011_ = ap_CS_fsm[0] ? icmp_ln851_2_fu_253_p2 : icmp_ln851_2_reg_809;
assign _000_ = ap_CS_fsm[0] ? op_2[7] : Range2_all_ones_reg_800;
assign _020_ = ap_CS_fsm[0] ? op_2[7] : p_Result_4_reg_789;
assign _013_ = ap_CS_fsm[0] ? icmp_ln851_2_fu_253_p2 : icmp_ln851_reg_779;
assign _019_ = ap_CS_fsm[0] ? op_2[7] : p_Result_3_reg_771;
assign _008_ = ap_rst ? 23'h000001 : ap_NS_fsm;
assign icmp_ln851_1_fu_473_p2 = _051_ ? 1'h1 : 1'h0;
assign icmp_ln851_2_fu_253_p2 = _052_ ? 1'h1 : 1'h0;
assign icmp_ln851_3_fu_588_p2 = _053_ ? 1'h1 : 1'h0;
assign op_6_V_fu_453_p3 = and_ln785_1_fu_448_p2 ? p_Val2_3_reg_814 : select_ln340_reg_895;
assign ret_V_18_fu_548_p3 = ret_V_17_reg_873[8] ? select_ln850_fu_543_p3 : ret_V_reg_878;
assign ret_V_20_fu_581_p3 = ret_V_19_reg_900[16] ? select_ln850_1_fu_576_p3 : ret_V_4_reg_905;
assign ret_V_22_fu_637_p3 = ret_V_21_reg_963[4] ? select_ln850_3_fu_632_p3 : ret_V_11_reg_968;
assign select_ln1192_fu_267_p3 = op_3 ? 9'h180 : 9'h000;
assign select_ln340_fu_413_p3 = or_ln340_1_fu_408_p2 ? 4'h0 : p_Val2_3_reg_814;
assign select_ln353_fu_506_p3 = p_Result_3_reg_771 ? select_ln850_6_fu_500_p3 : select_ln831_reg_922;
assign select_ln69_fu_644_p3 = op_3 ? 8'hff : 8'h00;
assign select_ln703_fu_466_p3 = op_3 ? 5'h18 : 5'h00;
assign select_ln831_fu_459_p3 = Range2_all_ones_reg_800 ? 2'h3 : 2'h0;
assign select_ln850_1_fu_576_p3 = icmp_ln851_1_reg_938 ? ret_V_4_reg_905 : ret_V_6_reg_958;
assign select_ln850_3_fu_632_p3 = icmp_ln851_3_reg_985 ? ret_V_11_reg_968 : ret_V_12_reg_995;
assign select_ln850_6_fu_500_p3 = icmp_ln851_2_reg_809 ? select_ln831_reg_922 : { 1'h0, ret_V_9_fu_483_p2 };
assign select_ln850_fu_543_p3 = icmp_ln851_reg_779 ? ret_V_reg_878 : ret_V_2_reg_933;
assign deleted_zeros_fu_298_p2 = or_ln778_reg_845 ^ Range2_all_ones_reg_800;
assign Range2_all_ones_fu_241_p1 = op_2;
assign ap_CS_fsm_state1 = ap_CS_fsm[0];
assign ap_CS_fsm_state10 = ap_CS_fsm[9];
assign ap_CS_fsm_state11 = ap_CS_fsm[10];
assign ap_CS_fsm_state12 = ap_CS_fsm[11];
assign ap_CS_fsm_state13 = ap_CS_fsm[12];
assign ap_CS_fsm_state14 = ap_CS_fsm[13];
assign ap_CS_fsm_state15 = ap_CS_fsm[14];
assign ap_CS_fsm_state16 = ap_CS_fsm[15];
assign ap_CS_fsm_state17 = ap_CS_fsm[16];
assign ap_CS_fsm_state18 = ap_CS_fsm[17];
assign ap_CS_fsm_state19 = ap_CS_fsm[18];
assign ap_CS_fsm_state2 = ap_CS_fsm[1];
assign ap_CS_fsm_state20 = ap_CS_fsm[19];
assign ap_CS_fsm_state21 = ap_CS_fsm[20];
assign ap_CS_fsm_state22 = ap_CS_fsm[21];
assign ap_CS_fsm_state23 = ap_CS_fsm[22];
assign ap_CS_fsm_state3 = ap_CS_fsm[2];
assign ap_CS_fsm_state4 = ap_CS_fsm[3];
assign ap_CS_fsm_state5 = ap_CS_fsm[4];
assign ap_CS_fsm_state6 = ap_CS_fsm[5];
assign ap_CS_fsm_state7 = ap_CS_fsm[6];
assign ap_CS_fsm_state8 = ap_CS_fsm[7];
assign ap_CS_fsm_state9 = ap_CS_fsm[8];
assign ap_done = op_30_ap_vld;
assign ap_ready = op_30_ap_vld;
assign grp_fu_235_p0 = { 3'h0, op_2[3] };
assign grp_fu_235_p1 = op_2[7:4];
assign grp_fu_293_p1 = { op_2[7], op_2 };
assign grp_fu_376_p0 = { op_9[3], op_9[3], op_9[3], op_9[3], op_9[3], op_9[3], op_9[3], op_9[3], op_9[3], op_9[3], op_9[3], op_9[3], op_9, 1'h0 };
assign grp_fu_376_p1 = { op_0[15], op_0 };
assign grp_fu_613_p0 = { ret_V_20_reg_980[12], ret_V_20_reg_980 };
assign grp_fu_613_p1 = { 10'h000, op_12 };
assign grp_fu_619_p0 = { 1'h0, op_14 };
assign grp_fu_619_p1 = { 2'h0, op_13 };
assign grp_fu_661_p0 = { 1'h0, add_ln69_2_reg_1030 };
assign grp_fu_661_p1 = { ret_V_22_reg_1015[1], ret_V_22_reg_1015[1], ret_V_22_reg_1015 };
assign grp_fu_670_p0 = { add_ln69_3_reg_1050[3], add_ln69_3_reg_1050[3], add_ln69_3_reg_1050[3], add_ln69_3_reg_1050[3], add_ln69_3_reg_1050[3], add_ln69_3_reg_1050[3], add_ln69_3_reg_1050[3], add_ln69_3_reg_1050[3], add_ln69_3_reg_1050[3], add_ln69_3_reg_1050[3], add_ln69_3_reg_1050 };
assign grp_fu_694_p0 = { op_25_V_reg_1060, 1'h0 };
assign grp_fu_694_p1 = { op_1, op_1, op_1, op_1, op_1, op_1, op_1, op_1, op_1, op_1, op_1, op_1, op_1, op_1, 1'h0 };
assign grp_fu_717_p0 = { op_26_V_reg_1075[13], op_26_V_reg_1075 };
assign grp_fu_717_p1 = { op_16[1], op_16[1], op_16[1], op_16[1], op_16[1], op_16[1], op_16[1], op_16[1], op_16[1], op_16[1], op_16[1], op_16[1], op_16[1], op_16 };
assign grp_fu_740_p0 = { ret_V_24_reg_1090[14], ret_V_24_reg_1090[14], ret_V_24_reg_1090[14], ret_V_24_reg_1090 };
assign grp_fu_740_p1 = { 2'h0, ret_V_18_reg_953[1], ret_V_18_reg_953[1], ret_V_18_reg_953[1], ret_V_18_reg_953[1], ret_V_18_reg_953[1], ret_V_18_reg_953[1], ret_V_18_reg_953[1], ret_V_18_reg_953[1], ret_V_18_reg_953[1], ret_V_18_reg_953[1], ret_V_18_reg_953[1], ret_V_18_reg_953[1], ret_V_18_reg_953[1], ret_V_18_reg_953[1], ret_V_18_reg_953 };
assign grp_fu_746_p0 = { op_17[3], op_17 };
assign grp_fu_746_p1 = { 3'h0, tmp_reg_948 };
assign grp_fu_755_p0 = { add_ln69_7_reg_1120[4], add_ln69_7_reg_1120[4], add_ln69_7_reg_1120[4], add_ln69_7_reg_1120[4], add_ln69_7_reg_1120[4], add_ln69_7_reg_1120[4], add_ln69_7_reg_1120[4], add_ln69_7_reg_1120[4], add_ln69_7_reg_1120[4], add_ln69_7_reg_1120[4], add_ln69_7_reg_1120[4], add_ln69_7_reg_1120[4], add_ln69_7_reg_1120[4], add_ln69_7_reg_1120 };
assign icmp_ln851_fu_199_p2 = icmp_ln851_2_fu_253_p2;
assign op_30 = { grp_fu_755_p2[17], grp_fu_755_p2[17], grp_fu_755_p2[17], grp_fu_755_p2[17], grp_fu_755_p2[17], grp_fu_755_p2[17], grp_fu_755_p2[17], grp_fu_755_p2[17], grp_fu_755_p2[17], grp_fu_755_p2[17], grp_fu_755_p2[17], grp_fu_755_p2[17], grp_fu_755_p2[17], grp_fu_755_p2[17], grp_fu_755_p2 };
assign p_Result_1_fu_536_p3 = ret_V_17_reg_873[8];
assign p_Result_2_fu_569_p3 = ret_V_19_reg_900[16];
assign p_Result_3_fu_187_p1 = op_2;
assign p_Result_4_fu_215_p1 = op_2;
assign p_Result_s_fu_625_p3 = ret_V_21_reg_963[4];
assign p_Val2_2_fu_205_p1 = op_2;
assign p_Val2_s_fu_675_p1 = op_1;
assign p_Val2_s_fu_675_p3 = { op_1, 1'h0 };
assign rhs_2_fu_512_p3 = { select_ln353_fu_506_p3, 3'h0 };
assign rhs_fu_364_p3 = { op_9, 1'h0 };
assign select_ln1192_fu_267_p0 = op_3;
assign select_ln69_fu_644_p0 = op_3;
assign select_ln703_fu_466_p0 = op_3;
assign sext_ln69_2_fu_730_p1 = { ret_V_18_reg_953[1], ret_V_18_reg_953[1], ret_V_18_reg_953[1], ret_V_18_reg_953[1], ret_V_18_reg_953[1], ret_V_18_reg_953[1], ret_V_18_reg_953[1], ret_V_18_reg_953[1], ret_V_18_reg_953[1], ret_V_18_reg_953[1], ret_V_18_reg_953[1], ret_V_18_reg_953[1], ret_V_18_reg_953[1], ret_V_18_reg_953[1], ret_V_18_reg_953 };
assign sext_ln703_2_fu_492_p1 = { op_6_V_reg_917[3], op_6_V_reg_917 };
assign sext_ln703_fu_290_p0 = op_2;
assign tmp_6_fu_223_p1 = op_2;
assign tmp_6_fu_223_p3 = op_2[3];
assign tmp_9_fu_302_p1 = op_2;
assign tmp_9_fu_302_p3 = op_2[7];
assign trunc_ln1192_fu_195_p0 = op_2;
assign trunc_ln1192_fu_195_p1 = op_2[6:0];
assign trunc_ln851_1_fu_249_p0 = op_2;
assign trunc_ln851_1_fu_249_p1 = op_2[6:0];
assign trunc_ln851_2_fu_565_p1 = grp_fu_495_p2[2:0];
assign trunc_ln851_fu_435_p1 = grp_fu_376_p2[3:0];
assign zext_ln831_fu_488_p1 = { 1'h0, ret_V_9_fu_483_p2 };
assign \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.ain_s0  = \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.a ;
assign \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.s  = { \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.fas_s2 , \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.sum_s1  };
assign \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.u2.a  = \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.ain_s1 ;
assign \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.u2.b  = \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.bin_s1 ;
assign \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.u2.cin  = \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.carry_s1 ;
assign \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.facout_s2  = \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.u2.cout ;
assign \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.fas_s2  = \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.u2.s ;
assign \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.u1.a  = \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.a [1:0];
assign \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.u1.b  = \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.bin_s0 [1:0];
assign \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.u1.cin  = 1'h1;
assign \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.facout_s1  = \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.u1.cout ;
assign \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.fas_s1  = \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.u1.s ;
assign \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.a  = \sub_5ns_5s_5_2_1_U6.din0 ;
assign \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.b  = \sub_5ns_5s_5_2_1_U6.din1 ;
assign \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.ce  = \sub_5ns_5s_5_2_1_U6.ce ;
assign \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.clk  = \sub_5ns_5s_5_2_1_U6.clk ;
assign \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.reset  = \sub_5ns_5s_5_2_1_U6.reset ;
assign \sub_5ns_5s_5_2_1_U6.dout  = \sub_5ns_5s_5_2_1_U6.top_sub_5ns_5s_5_2_1_Adder_5_U.s ;
assign \sub_5ns_5s_5_2_1_U6.ce  = 1'h1;
assign \sub_5ns_5s_5_2_1_U6.clk  = ap_clk;
assign \sub_5ns_5s_5_2_1_U6.din0  = select_ln703_reg_928;
assign \sub_5ns_5s_5_2_1_U6.din1  = { op_6_V_reg_917[3], op_6_V_reg_917 };
assign grp_fu_495_p2 = \sub_5ns_5s_5_2_1_U6.dout ;
assign \sub_5ns_5s_5_2_1_U6.reset  = ap_rst;
assign \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.ain_s0  = \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.a ;
assign \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.bin_s0  = \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.b ;
assign \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.s  = { \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.fas_s2 , \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.sum_s1  };
assign \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.u2.a  = \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.ain_s1 ;
assign \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.u2.b  = \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.bin_s1 ;
assign \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.u2.cin  = \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.carry_s1 ;
assign \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.facout_s2  = \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.u2.cout ;
assign \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.fas_s2  = \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.u2.s ;
assign \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.u1.a  = \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.a [3:0];
assign \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.u1.b  = \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.b [3:0];
assign \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.u1.cin  = 1'h0;
assign \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.facout_s1  = \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.u1.cout ;
assign \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.fas_s1  = \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.u1.s ;
assign \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.a  = \add_9ns_9s_9_2_1_U2.din0 ;
assign \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.b  = \add_9ns_9s_9_2_1_U2.din1 ;
assign \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.ce  = \add_9ns_9s_9_2_1_U2.ce ;
assign \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.clk  = \add_9ns_9s_9_2_1_U2.clk ;
assign \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.reset  = \add_9ns_9s_9_2_1_U2.reset ;
assign \add_9ns_9s_9_2_1_U2.dout  = \add_9ns_9s_9_2_1_U2.top_add_9ns_9s_9_2_1_Adder_1_U.s ;
assign \add_9ns_9s_9_2_1_U2.ce  = 1'h1;
assign \add_9ns_9s_9_2_1_U2.clk  = ap_clk;
assign \add_9ns_9s_9_2_1_U2.din0  = select_ln1192_reg_834;
assign \add_9ns_9s_9_2_1_U2.din1  = { op_2[7], op_2 };
assign grp_fu_293_p2 = \add_9ns_9s_9_2_1_U2.dout ;
assign \add_9ns_9s_9_2_1_U2.reset  = ap_rst;
assign \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.ain_s0  = \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.a ;
assign \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.bin_s0  = \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.b ;
assign \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.s  = { \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.fas_s2 , \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.sum_s1  };
assign \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.u2.a  = \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.ain_s1 ;
assign \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.u2.b  = \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.bin_s1 ;
assign \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.u2.cin  = \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.carry_s1 ;
assign \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.facout_s2  = \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.u2.cout ;
assign \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.fas_s2  = \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.u2.s ;
assign \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.u1.a  = \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.a [1:0];
assign \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.u1.b  = \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.b [1:0];
assign \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.u1.cin  = 1'h0;
assign \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.facout_s1  = \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.u1.cout ;
assign \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.fas_s1  = \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.u1.s ;
assign \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.a  = \add_5s_5ns_5_2_1_U16.din0 ;
assign \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.b  = \add_5s_5ns_5_2_1_U16.din1 ;
assign \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.ce  = \add_5s_5ns_5_2_1_U16.ce ;
assign \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.clk  = \add_5s_5ns_5_2_1_U16.clk ;
assign \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.reset  = \add_5s_5ns_5_2_1_U16.reset ;
assign \add_5s_5ns_5_2_1_U16.dout  = \add_5s_5ns_5_2_1_U16.top_add_5s_5ns_5_2_1_Adder_13_U.s ;
assign \add_5s_5ns_5_2_1_U16.ce  = 1'h1;
assign \add_5s_5ns_5_2_1_U16.clk  = ap_clk;
assign \add_5s_5ns_5_2_1_U16.din0  = { op_17[3], op_17 };
assign \add_5s_5ns_5_2_1_U16.din1  = { 3'h0, tmp_reg_948 };
assign grp_fu_746_p2 = \add_5s_5ns_5_2_1_U16.dout ;
assign \add_5s_5ns_5_2_1_U16.reset  = ap_rst;
assign \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.ain_s0  = \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.a ;
assign \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.bin_s0  = \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.b ;
assign \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.s  = { \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.fas_s2 , \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.sum_s1  };
assign \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.u2.a  = \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.ain_s1 ;
assign \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.u2.b  = \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.bin_s1 ;
assign \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.u2.cin  = \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.carry_s1 ;
assign \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.facout_s2  = \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.u2.cout ;
assign \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.fas_s2  = \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.u2.s ;
assign \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.u1.a  = \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.a [1:0];
assign \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.u1.b  = \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.b [1:0];
assign \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.u1.cin  = 1'h0;
assign \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.facout_s1  = \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.u1.cout ;
assign \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.fas_s1  = \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.u1.s ;
assign \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.a  = \add_4ns_4s_4_2_1_U11.din0 ;
assign \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.b  = \add_4ns_4s_4_2_1_U11.din1 ;
assign \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.ce  = \add_4ns_4s_4_2_1_U11.ce ;
assign \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.clk  = \add_4ns_4s_4_2_1_U11.clk ;
assign \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.reset  = \add_4ns_4s_4_2_1_U11.reset ;
assign \add_4ns_4s_4_2_1_U11.dout  = \add_4ns_4s_4_2_1_U11.top_add_4ns_4s_4_2_1_Adder_9_U.s ;
assign \add_4ns_4s_4_2_1_U11.ce  = 1'h1;
assign \add_4ns_4s_4_2_1_U11.clk  = ap_clk;
assign \add_4ns_4s_4_2_1_U11.din0  = { 1'h0, add_ln69_2_reg_1030 };
assign \add_4ns_4s_4_2_1_U11.din1  = { ret_V_22_reg_1015[1], ret_V_22_reg_1015[1], ret_V_22_reg_1015 };
assign grp_fu_661_p2 = \add_4ns_4s_4_2_1_U11.dout ;
assign \add_4ns_4s_4_2_1_U11.reset  = ap_rst;
assign \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.ain_s0  = \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.a ;
assign \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.bin_s0  = \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.b ;
assign \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.s  = { \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.fas_s2 , \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.sum_s1  };
assign \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.u2.a  = \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.ain_s1 ;
assign \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.u2.b  = \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.bin_s1 ;
assign \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.u2.cin  = \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.carry_s1 ;
assign \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.facout_s2  = \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.u2.cout ;
assign \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.fas_s2  = \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.u2.s ;
assign \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.u1.a  = \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.a [1:0];
assign \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.u1.b  = \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.b [1:0];
assign \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.u1.cin  = 1'h0;
assign \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.facout_s1  = \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.u1.cout ;
assign \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.fas_s1  = \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.u1.s ;
assign \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.a  = \add_4ns_4ns_4_2_1_U1.din0 ;
assign \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.b  = \add_4ns_4ns_4_2_1_U1.din1 ;
assign \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.ce  = \add_4ns_4ns_4_2_1_U1.ce ;
assign \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.clk  = \add_4ns_4ns_4_2_1_U1.clk ;
assign \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.reset  = \add_4ns_4ns_4_2_1_U1.reset ;
assign \add_4ns_4ns_4_2_1_U1.dout  = \add_4ns_4ns_4_2_1_U1.top_add_4ns_4ns_4_2_1_Adder_0_U.s ;
assign \add_4ns_4ns_4_2_1_U1.ce  = 1'h1;
assign \add_4ns_4ns_4_2_1_U1.clk  = ap_clk;
assign \add_4ns_4ns_4_2_1_U1.din0  = { 3'h0, op_2[3] };
assign \add_4ns_4ns_4_2_1_U1.din1  = op_2[7:4];
assign grp_fu_235_p2 = \add_4ns_4ns_4_2_1_U1.dout ;
assign \add_4ns_4ns_4_2_1_U1.reset  = ap_rst;
assign \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.ain_s0  = \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.a ;
assign \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.bin_s0  = \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.b ;
assign \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.s  = { \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.fas_s2 , \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.sum_s1  };
assign \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.u2.a  = \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.ain_s1 ;
assign \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.u2.b  = \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.bin_s1 ;
assign \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.u2.cin  = \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.carry_s1 ;
assign \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.facout_s2  = \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.u2.cout ;
assign \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.fas_s2  = \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.u2.s ;
assign \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.u1.a  = \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.a [0];
assign \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.u1.b  = \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.b [0];
assign \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.u1.cin  = 1'h0;
assign \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.facout_s1  = \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.u1.cout ;
assign \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.fas_s1  = \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.u1.s ;
assign \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.a  = \add_3ns_3ns_3_2_1_U9.din0 ;
assign \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.b  = \add_3ns_3ns_3_2_1_U9.din1 ;
assign \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.ce  = \add_3ns_3ns_3_2_1_U9.ce ;
assign \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.clk  = \add_3ns_3ns_3_2_1_U9.clk ;
assign \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.reset  = \add_3ns_3ns_3_2_1_U9.reset ;
assign \add_3ns_3ns_3_2_1_U9.dout  = \add_3ns_3ns_3_2_1_U9.top_add_3ns_3ns_3_2_1_Adder_7_U.s ;
assign \add_3ns_3ns_3_2_1_U9.ce  = 1'h1;
assign \add_3ns_3ns_3_2_1_U9.clk  = ap_clk;
assign \add_3ns_3ns_3_2_1_U9.din0  = { 1'h0, op_14 };
assign \add_3ns_3ns_3_2_1_U9.din1  = { 2'h0, op_13 };
assign grp_fu_619_p2 = \add_3ns_3ns_3_2_1_U9.dout ;
assign \add_3ns_3ns_3_2_1_U9.reset  = ap_rst;
assign \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.ain_s0  = \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.a ;
assign \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.bin_s0  = \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.b ;
assign \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.s  = { \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.fas_s2 , \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.sum_s1  };
assign \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.u2.a  = \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.ain_s1 ;
assign \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.u2.b  = \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.bin_s1 ;
assign \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.u2.cin  = \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.carry_s1 ;
assign \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.facout_s2  = \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.u2.cout ;
assign \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.fas_s2  = \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.u2.s ;
assign \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.u1.a  = \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.a [0];
assign \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.u1.b  = \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.b [0];
assign \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.u1.cin  = 1'h0;
assign \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.facout_s1  = \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.u1.cout ;
assign \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.fas_s1  = \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.u1.s ;
assign \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.a  = \add_2ns_2ns_2_2_1_U7.din0 ;
assign \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.b  = \add_2ns_2ns_2_2_1_U7.din1 ;
assign \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.ce  = \add_2ns_2ns_2_2_1_U7.ce ;
assign \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.clk  = \add_2ns_2ns_2_2_1_U7.clk ;
assign \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.reset  = \add_2ns_2ns_2_2_1_U7.reset ;
assign \add_2ns_2ns_2_2_1_U7.dout  = \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_3_U.s ;
assign \add_2ns_2ns_2_2_1_U7.ce  = 1'h1;
assign \add_2ns_2ns_2_2_1_U7.clk  = ap_clk;
assign \add_2ns_2ns_2_2_1_U7.din0  = ret_V_11_reg_968;
assign \add_2ns_2ns_2_2_1_U7.din1  = 2'h1;
assign grp_fu_593_p2 = \add_2ns_2ns_2_2_1_U7.dout ;
assign \add_2ns_2ns_2_2_1_U7.reset  = ap_rst;
assign \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.ain_s0  = \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.a ;
assign \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.bin_s0  = \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.b ;
assign \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.s  = { \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.fas_s2 , \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.sum_s1  };
assign \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.u2.a  = \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.ain_s1 ;
assign \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.u2.b  = \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.bin_s1 ;
assign \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.u2.cin  = \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.carry_s1 ;
assign \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.facout_s2  = \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.u2.cout ;
assign \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.fas_s2  = \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.u2.s ;
assign \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.u1.a  = \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.a [0];
assign \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.u1.b  = \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.b [0];
assign \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.u1.cin  = 1'h0;
assign \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.facout_s1  = \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.u1.cout ;
assign \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.fas_s1  = \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.u1.s ;
assign \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.a  = \add_2ns_2ns_2_2_1_U4.din0 ;
assign \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.b  = \add_2ns_2ns_2_2_1_U4.din1 ;
assign \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.ce  = \add_2ns_2ns_2_2_1_U4.ce ;
assign \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.clk  = \add_2ns_2ns_2_2_1_U4.clk ;
assign \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.reset  = \add_2ns_2ns_2_2_1_U4.reset ;
assign \add_2ns_2ns_2_2_1_U4.dout  = \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_3_U.s ;
assign \add_2ns_2ns_2_2_1_U4.ce  = 1'h1;
assign \add_2ns_2ns_2_2_1_U4.clk  = ap_clk;
assign \add_2ns_2ns_2_2_1_U4.din0  = ret_V_reg_878;
assign \add_2ns_2ns_2_2_1_U4.din1  = 2'h1;
assign grp_fu_420_p2 = \add_2ns_2ns_2_2_1_U4.dout ;
assign \add_2ns_2ns_2_2_1_U4.reset  = ap_rst;
assign \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.ain_s0  = \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.a ;
assign \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.bin_s0  = \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.b ;
assign \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.s  = { \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.fas_s2 , \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.sum_s1  };
assign \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.u2.a  = \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.ain_s1 ;
assign \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.u2.b  = \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.bin_s1 ;
assign \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.u2.cin  = \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.carry_s1 ;
assign \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.facout_s2  = \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.u2.cout ;
assign \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.fas_s2  = \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.u2.s ;
assign \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.u1.a  = \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.a [8:0];
assign \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.u1.b  = \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.b [8:0];
assign \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.u1.cin  = 1'h0;
assign \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.facout_s1  = \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.u1.cout ;
assign \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.fas_s1  = \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.u1.s ;
assign \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.a  = \add_18s_18ns_18_2_1_U17.din0 ;
assign \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.b  = \add_18s_18ns_18_2_1_U17.din1 ;
assign \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.ce  = \add_18s_18ns_18_2_1_U17.ce ;
assign \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.clk  = \add_18s_18ns_18_2_1_U17.clk ;
assign \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.reset  = \add_18s_18ns_18_2_1_U17.reset ;
assign \add_18s_18ns_18_2_1_U17.dout  = \add_18s_18ns_18_2_1_U17.top_add_18s_18ns_18_2_1_Adder_12_U.s ;
assign \add_18s_18ns_18_2_1_U17.ce  = 1'h1;
assign \add_18s_18ns_18_2_1_U17.clk  = ap_clk;
assign \add_18s_18ns_18_2_1_U17.din0  = { add_ln69_7_reg_1120[4], add_ln69_7_reg_1120[4], add_ln69_7_reg_1120[4], add_ln69_7_reg_1120[4], add_ln69_7_reg_1120[4], add_ln69_7_reg_1120[4], add_ln69_7_reg_1120[4], add_ln69_7_reg_1120[4], add_ln69_7_reg_1120[4], add_ln69_7_reg_1120[4], add_ln69_7_reg_1120[4], add_ln69_7_reg_1120[4], add_ln69_7_reg_1120[4], add_ln69_7_reg_1120 };
assign \add_18s_18ns_18_2_1_U17.din1  = add_ln69_5_reg_1115;
assign grp_fu_755_p2 = \add_18s_18ns_18_2_1_U17.dout ;
assign \add_18s_18ns_18_2_1_U17.reset  = ap_rst;
assign \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.ain_s0  = \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.a ;
assign \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.bin_s0  = \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.b ;
assign \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.s  = { \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.fas_s2 , \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.sum_s1  };
assign \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.u2.a  = \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.ain_s1 ;
assign \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.u2.b  = \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.bin_s1 ;
assign \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.u2.cin  = \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.carry_s1 ;
assign \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.facout_s2  = \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.u2.cout ;
assign \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.fas_s2  = \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.u2.s ;
assign \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.u1.a  = \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.a [8:0];
assign \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.u1.b  = \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.b [8:0];
assign \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.u1.cin  = 1'h0;
assign \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.facout_s1  = \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.u1.cout ;
assign \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.fas_s1  = \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.u1.s ;
assign \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.a  = \add_18s_18ns_18_2_1_U15.din0 ;
assign \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.b  = \add_18s_18ns_18_2_1_U15.din1 ;
assign \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.ce  = \add_18s_18ns_18_2_1_U15.ce ;
assign \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.clk  = \add_18s_18ns_18_2_1_U15.clk ;
assign \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.reset  = \add_18s_18ns_18_2_1_U15.reset ;
assign \add_18s_18ns_18_2_1_U15.dout  = \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_12_U.s ;
assign \add_18s_18ns_18_2_1_U15.ce  = 1'h1;
assign \add_18s_18ns_18_2_1_U15.clk  = ap_clk;
assign \add_18s_18ns_18_2_1_U15.din0  = { ret_V_24_reg_1090[14], ret_V_24_reg_1090[14], ret_V_24_reg_1090[14], ret_V_24_reg_1090 };
assign \add_18s_18ns_18_2_1_U15.din1  = { 2'h0, ret_V_18_reg_953[1], ret_V_18_reg_953[1], ret_V_18_reg_953[1], ret_V_18_reg_953[1], ret_V_18_reg_953[1], ret_V_18_reg_953[1], ret_V_18_reg_953[1], ret_V_18_reg_953[1], ret_V_18_reg_953[1], ret_V_18_reg_953[1], ret_V_18_reg_953[1], ret_V_18_reg_953[1], ret_V_18_reg_953[1], ret_V_18_reg_953[1], ret_V_18_reg_953 };
assign grp_fu_740_p2 = \add_18s_18ns_18_2_1_U15.dout ;
assign \add_18s_18ns_18_2_1_U15.reset  = ap_rst;
assign \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.ain_s0  = \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.a ;
assign \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.bin_s0  = \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.b ;
assign \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.s  = { \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.fas_s2 , \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.sum_s1  };
assign \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.u2.a  = \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.ain_s1 ;
assign \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.u2.b  = \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.bin_s1 ;
assign \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.u2.cin  = \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.carry_s1 ;
assign \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.facout_s2  = \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.u2.cout ;
assign \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.fas_s2  = \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.u2.s ;
assign \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.u1.a  = \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.a [7:0];
assign \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.u1.b  = \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.b [7:0];
assign \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.u1.cin  = 1'h0;
assign \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.facout_s1  = \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.u1.cout ;
assign \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.fas_s1  = \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.u1.s ;
assign \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.a  = \add_17s_17s_17_2_1_U3.din0 ;
assign \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.b  = \add_17s_17s_17_2_1_U3.din1 ;
assign \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.ce  = \add_17s_17s_17_2_1_U3.ce ;
assign \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.clk  = \add_17s_17s_17_2_1_U3.clk ;
assign \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.reset  = \add_17s_17s_17_2_1_U3.reset ;
assign \add_17s_17s_17_2_1_U3.dout  = \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.s ;
assign \add_17s_17s_17_2_1_U3.ce  = 1'h1;
assign \add_17s_17s_17_2_1_U3.clk  = ap_clk;
assign \add_17s_17s_17_2_1_U3.din0  = { op_9[3], op_9[3], op_9[3], op_9[3], op_9[3], op_9[3], op_9[3], op_9[3], op_9[3], op_9[3], op_9[3], op_9[3], op_9, 1'h0 };
assign \add_17s_17s_17_2_1_U3.din1  = { op_0[15], op_0 };
assign grp_fu_376_p2 = \add_17s_17s_17_2_1_U3.dout ;
assign \add_17s_17s_17_2_1_U3.reset  = ap_rst;
assign \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.ain_s0  = \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.a ;
assign \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.bin_s0  = \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.b ;
assign \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.s  = { \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.fas_s2 , \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.sum_s1  };
assign \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.u2.a  = \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.ain_s1 ;
assign \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.u2.b  = \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.bin_s1 ;
assign \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.u2.cin  = \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.carry_s1 ;
assign \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.facout_s2  = \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.u2.cout ;
assign \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.fas_s2  = \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.u2.s ;
assign \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.u1.a  = \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.a [6:0];
assign \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.u1.b  = \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.b [6:0];
assign \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.u1.cin  = 1'h0;
assign \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.facout_s1  = \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.u1.cout ;
assign \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.fas_s1  = \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.u1.s ;
assign \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.a  = \add_15s_15s_15_2_1_U14.din0 ;
assign \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.b  = \add_15s_15s_15_2_1_U14.din1 ;
assign \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.ce  = \add_15s_15s_15_2_1_U14.ce ;
assign \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.clk  = \add_15s_15s_15_2_1_U14.clk ;
assign \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.reset  = \add_15s_15s_15_2_1_U14.reset ;
assign \add_15s_15s_15_2_1_U14.dout  = \add_15s_15s_15_2_1_U14.top_add_15s_15s_15_2_1_Adder_11_U.s ;
assign \add_15s_15s_15_2_1_U14.ce  = 1'h1;
assign \add_15s_15s_15_2_1_U14.clk  = ap_clk;
assign \add_15s_15s_15_2_1_U14.din0  = { op_26_V_reg_1075[13], op_26_V_reg_1075 };
assign \add_15s_15s_15_2_1_U14.din1  = { op_16[1], op_16[1], op_16[1], op_16[1], op_16[1], op_16[1], op_16[1], op_16[1], op_16[1], op_16[1], op_16[1], op_16[1], op_16[1], op_16 };
assign grp_fu_717_p2 = \add_15s_15s_15_2_1_U14.dout ;
assign \add_15s_15s_15_2_1_U14.reset  = ap_rst;
assign \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.ain_s0  = \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.a ;
assign \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.bin_s0  = \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.b ;
assign \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.s  = { \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.fas_s2 , \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.sum_s1  };
assign \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.u2.a  = \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.ain_s1 ;
assign \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.u2.b  = \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.bin_s1 ;
assign \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.u2.cin  = \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.carry_s1 ;
assign \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.facout_s2  = \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.u2.cout ;
assign \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.fas_s2  = \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.u2.s ;
assign \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.u1.a  = \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.a [6:0];
assign \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.u1.b  = \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.b [6:0];
assign \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.u1.cin  = 1'h0;
assign \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.facout_s1  = \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.u1.cout ;
assign \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.fas_s1  = \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.u1.s ;
assign \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.a  = \add_15ns_15s_15_2_1_U13.din0 ;
assign \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.b  = \add_15ns_15s_15_2_1_U13.din1 ;
assign \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.ce  = \add_15ns_15s_15_2_1_U13.ce ;
assign \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.clk  = \add_15ns_15s_15_2_1_U13.clk ;
assign \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.reset  = \add_15ns_15s_15_2_1_U13.reset ;
assign \add_15ns_15s_15_2_1_U13.dout  = \add_15ns_15s_15_2_1_U13.top_add_15ns_15s_15_2_1_Adder_10_U.s ;
assign \add_15ns_15s_15_2_1_U13.ce  = 1'h1;
assign \add_15ns_15s_15_2_1_U13.clk  = ap_clk;
assign \add_15ns_15s_15_2_1_U13.din0  = { op_25_V_reg_1060, 1'h0 };
assign \add_15ns_15s_15_2_1_U13.din1  = { op_1, op_1, op_1, op_1, op_1, op_1, op_1, op_1, op_1, op_1, op_1, op_1, op_1, op_1, 1'h0 };
assign grp_fu_694_p2 = \add_15ns_15s_15_2_1_U13.dout ;
assign \add_15ns_15s_15_2_1_U13.reset  = ap_rst;
assign \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.ain_s0  = \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.a ;
assign \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.bin_s0  = \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.b ;
assign \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.s  = { \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.fas_s2 , \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.sum_s1  };
assign \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.u2.a  = \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.ain_s1 ;
assign \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.u2.b  = \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.bin_s1 ;
assign \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.u2.cin  = \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.carry_s1 ;
assign \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.facout_s2  = \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.u2.cout ;
assign \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.fas_s2  = \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.u2.s ;
assign \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.u1.a  = \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.a [6:0];
assign \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.u1.b  = \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.b [6:0];
assign \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.u1.cin  = 1'h0;
assign \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.facout_s1  = \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.u1.cout ;
assign \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.fas_s1  = \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.u1.s ;
assign \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.a  = \add_14s_14ns_14_2_1_U8.din0 ;
assign \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.b  = \add_14s_14ns_14_2_1_U8.din1 ;
assign \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.ce  = \add_14s_14ns_14_2_1_U8.ce ;
assign \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.clk  = \add_14s_14ns_14_2_1_U8.clk ;
assign \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.reset  = \add_14s_14ns_14_2_1_U8.reset ;
assign \add_14s_14ns_14_2_1_U8.dout  = \add_14s_14ns_14_2_1_U8.top_add_14s_14ns_14_2_1_Adder_6_U.s ;
assign \add_14s_14ns_14_2_1_U8.ce  = 1'h1;
assign \add_14s_14ns_14_2_1_U8.clk  = ap_clk;
assign \add_14s_14ns_14_2_1_U8.din0  = { ret_V_20_reg_980[12], ret_V_20_reg_980 };
assign \add_14s_14ns_14_2_1_U8.din1  = { 10'h000, op_12 };
assign grp_fu_613_p2 = \add_14s_14ns_14_2_1_U8.dout ;
assign \add_14s_14ns_14_2_1_U8.reset  = ap_rst;
assign \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.ain_s0  = \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.a ;
assign \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.bin_s0  = \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.b ;
assign \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.s  = { \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.fas_s2 , \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.sum_s1  };
assign \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.u2.a  = \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.ain_s1 ;
assign \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.u2.b  = \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.bin_s1 ;
assign \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.u2.cin  = \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.carry_s1 ;
assign \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.facout_s2  = \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.u2.cout ;
assign \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.fas_s2  = \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.u2.s ;
assign \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.u1.a  = \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.a [6:0];
assign \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.u1.b  = \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.b [6:0];
assign \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.u1.cin  = 1'h0;
assign \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.facout_s1  = \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.u1.cout ;
assign \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.fas_s1  = \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.u1.s ;
assign \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.a  = \add_14s_14ns_14_2_1_U12.din0 ;
assign \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.b  = \add_14s_14ns_14_2_1_U12.din1 ;
assign \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.ce  = \add_14s_14ns_14_2_1_U12.ce ;
assign \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.clk  = \add_14s_14ns_14_2_1_U12.clk ;
assign \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.reset  = \add_14s_14ns_14_2_1_U12.reset ;
assign \add_14s_14ns_14_2_1_U12.dout  = \add_14s_14ns_14_2_1_U12.top_add_14s_14ns_14_2_1_Adder_6_U.s ;
assign \add_14s_14ns_14_2_1_U12.ce  = 1'h1;
assign \add_14s_14ns_14_2_1_U12.clk  = ap_clk;
assign \add_14s_14ns_14_2_1_U12.din0  = { add_ln69_3_reg_1050[3], add_ln69_3_reg_1050[3], add_ln69_3_reg_1050[3], add_ln69_3_reg_1050[3], add_ln69_3_reg_1050[3], add_ln69_3_reg_1050[3], add_ln69_3_reg_1050[3], add_ln69_3_reg_1050[3], add_ln69_3_reg_1050[3], add_ln69_3_reg_1050[3], add_ln69_3_reg_1050 };
assign \add_14s_14ns_14_2_1_U12.din1  = add_ln69_1_reg_1045;
assign grp_fu_670_p2 = \add_14s_14ns_14_2_1_U12.dout ;
assign \add_14s_14ns_14_2_1_U12.reset  = ap_rst;
assign \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.ain_s0  = \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.a ;
assign \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.bin_s0  = \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.b ;
assign \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.s  = { \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.fas_s2 , \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.sum_s1  };
assign \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.u2.a  = \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.ain_s1 ;
assign \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.u2.b  = \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.bin_s1 ;
assign \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.u2.cin  = \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.carry_s1 ;
assign \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.facout_s2  = \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.u2.cout ;
assign \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.fas_s2  = \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.u2.s ;
assign \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.u1.a  = \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.a [6:0];
assign \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.u1.b  = \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.b [6:0];
assign \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.u1.cin  = 1'h0;
assign \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.facout_s1  = \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.u1.cout ;
assign \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.fas_s1  = \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.u1.s ;
assign \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.a  = \add_14ns_14ns_14_2_1_U10.din0 ;
assign \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.b  = \add_14ns_14ns_14_2_1_U10.din1 ;
assign \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.ce  = \add_14ns_14ns_14_2_1_U10.ce ;
assign \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.clk  = \add_14ns_14ns_14_2_1_U10.clk ;
assign \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.reset  = \add_14ns_14ns_14_2_1_U10.reset ;
assign \add_14ns_14ns_14_2_1_U10.dout  = \add_14ns_14ns_14_2_1_U10.top_add_14ns_14ns_14_2_1_Adder_8_U.s ;
assign \add_14ns_14ns_14_2_1_U10.ce  = 1'h1;
assign \add_14ns_14ns_14_2_1_U10.clk  = ap_clk;
assign \add_14ns_14ns_14_2_1_U10.din0  = add_ln69_reg_1025;
assign \add_14ns_14ns_14_2_1_U10.din1  = select_ln69_reg_1020;
assign grp_fu_654_p2 = \add_14ns_14ns_14_2_1_U10.dout ;
assign \add_14ns_14ns_14_2_1_U10.reset  = ap_rst;
assign \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.ain_s0  = \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.a ;
assign \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.bin_s0  = \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.b ;
assign \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.s  = { \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.fas_s2 , \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.sum_s1  };
assign \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.u2.a  = \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.ain_s1 ;
assign \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.u2.b  = \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.bin_s1 ;
assign \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.u2.cin  = \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.carry_s1 ;
assign \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.facout_s2  = \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.u2.cout ;
assign \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.fas_s2  = \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.u2.s ;
assign \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.u1.a  = \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.a [5:0];
assign \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.u1.b  = \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.b [5:0];
assign \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.u1.cin  = 1'h0;
assign \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.facout_s1  = \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.u1.cout ;
assign \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.fas_s1  = \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.u1.s ;
assign \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.a  = \add_13ns_13ns_13_2_1_U5.din0 ;
assign \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.b  = \add_13ns_13ns_13_2_1_U5.din1 ;
assign \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.ce  = \add_13ns_13ns_13_2_1_U5.ce ;
assign \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.clk  = \add_13ns_13ns_13_2_1_U5.clk ;
assign \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.reset  = \add_13ns_13ns_13_2_1_U5.reset ;
assign \add_13ns_13ns_13_2_1_U5.dout  = \add_13ns_13ns_13_2_1_U5.top_add_13ns_13ns_13_2_1_Adder_4_U.s ;
assign \add_13ns_13ns_13_2_1_U5.ce  = 1'h1;
assign \add_13ns_13ns_13_2_1_U5.clk  = ap_clk;
assign \add_13ns_13ns_13_2_1_U5.din0  = ret_V_4_reg_905;
assign \add_13ns_13ns_13_2_1_U5.din1  = 13'h0001;
assign grp_fu_478_p2 = \add_13ns_13ns_13_2_1_U5.dout ;
assign \add_13ns_13ns_13_2_1_U5.reset  = ap_rst;
endmodule


// Product machine:
module top_A_times_top_B (ap_start, op_0, op_1, op_12, op_13, op_14, op_16, op_17, op_2, op_3, op_9, ap_clk, unsafe_signal);
input ap_start;
input [15:0] op_0;
input op_1;
input [3:0] op_12;
input op_13;
input [1:0] op_14;
input [1:0] op_16;
input [3:0] op_17;
input [7:0] op_2;
input op_3;
input [3:0] op_9;
input ap_clk;
output unsafe_signal;
reg _setup;
initial _setup = 1'b0;
always @ (posedge ap_clk) _setup <= 1'b1;
reg ap_start_internal;
always @ (posedge ap_clk) if (!_setup) ap_start_internal <= ap_start;
reg [15:0] op_0_internal;
always @ (posedge ap_clk) if (!_setup) op_0_internal <= op_0;
reg op_1_internal;
always @ (posedge ap_clk) if (!_setup) op_1_internal <= op_1;
reg [3:0] op_12_internal;
always @ (posedge ap_clk) if (!_setup) op_12_internal <= op_12;
reg op_13_internal;
always @ (posedge ap_clk) if (!_setup) op_13_internal <= op_13;
reg [1:0] op_14_internal;
always @ (posedge ap_clk) if (!_setup) op_14_internal <= op_14;
reg [1:0] op_16_internal;
always @ (posedge ap_clk) if (!_setup) op_16_internal <= op_16;
reg [3:0] op_17_internal;
always @ (posedge ap_clk) if (!_setup) op_17_internal <= op_17;
reg [7:0] op_2_internal;
always @ (posedge ap_clk) if (!_setup) op_2_internal <= op_2;
reg op_3_internal;
always @ (posedge ap_clk) if (!_setup) op_3_internal <= op_3;
reg [3:0] op_9_internal;
always @ (posedge ap_clk) if (!_setup) op_9_internal <= op_9;
wire ap_done_A;
wire ap_done_B;
wire ap_done_eq;
assign ap_done_eq = ap_done_A == ap_done_B;
wire ap_idle_A;
wire ap_idle_B;
wire ap_idle_eq;
assign ap_idle_eq = ap_idle_A == ap_idle_B;
wire ap_ready_A;
wire ap_ready_B;
wire ap_ready_eq;
assign ap_ready_eq = ap_ready_A == ap_ready_B;
wire [31:0] op_30_A;
wire [31:0] op_30_B;
wire op_30_eq;
assign op_30_eq = op_30_A == op_30_B;
wire op_30_ap_vld_A;
wire op_30_ap_vld_B;
wire clk_enable_A;
wire clk_enable_B;
assign clk_enable_A = _setup & (~op_30_ap_vld_A | op_30_ap_vld_B);
assign clk_enable_B = _setup;
wire divergent;
assign divergent = ~(ap_done_eq & ap_idle_eq & ap_ready_eq & op_30_eq);
assign unsafe_signal = op_30_ap_vld_A & op_30_ap_vld_B & divergent;
top_A instance_A (
    .ap_clk(ap_clk),
    .clk_enable(clk_enable_A),
    .ap_start(ap_start_internal),
    .op_0(op_0_internal),
    .op_1(op_1_internal),
    .op_12(op_12_internal),
    .op_13(op_13_internal),
    .op_14(op_14_internal),
    .op_16(op_16_internal),
    .op_17(op_17_internal),
    .op_2(op_2_internal),
    .op_3(op_3_internal),
    .op_9(op_9_internal),
    .ap_done(ap_done_A),
    .ap_idle(ap_idle_A),
    .ap_ready(ap_ready_A),
    .op_30(op_30_A),
    .op_30_ap_vld(op_30_ap_vld_A)
);
top_B instance_B (
    .ap_clk(ap_clk),
    .clk_enable(clk_enable_B),
    .ap_start(ap_start_internal),
    .op_0(op_0_internal),
    .op_1(op_1_internal),
    .op_12(op_12_internal),
    .op_13(op_13_internal),
    .op_14(op_14_internal),
    .op_16(op_16_internal),
    .op_17(op_17_internal),
    .op_2(op_2_internal),
    .op_3(op_3_internal),
    .op_9(op_9_internal),
    .ap_done(ap_done_B),
    .ap_idle(ap_idle_B),
    .ap_ready(ap_ready_B),
    .op_30(op_30_B),
    .op_30_ap_vld(op_30_ap_vld_B)
);
endmodule
