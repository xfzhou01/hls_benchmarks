// Processed by function `construct_kairos` in `verilog_tricks.py`.
// Machine A:
// Processed by function `add_clk_enable_signal` in `verilog_tricks.py`.
// Processed by function `remove_reset_signal` in `verilog_tricks.py`.
module top_A (
  ap_clk,
  ap_start,
  ap_done,
  ap_idle,
  ap_ready,
  op_0,
  op_1,
  op_2,
  op_5,
  op_6,
  op_7,
  op_9,
  op_13,
  op_19,
  op_28,
  op_28_ap_vld,
clk_enable
);
input clk_enable;


input ap_clk;
wire ap_rst;
assign ap_rst = op_28_ap_vld;
input ap_start;
input op_0;
input [31:0] op_1;
input [1:0] op_13;
input [7:0] op_19;
input [3:0] op_2;
input [1:0] op_5;
input [31:0] op_6;
input [3:0] op_7;
input [1:0] op_9;
output ap_done;
output ap_idle;
output ap_ready;
output [31:0] op_28;
output op_28_ap_vld;


reg Range1_all_ones_1_reg_2195;
reg Range1_all_ones_2_reg_2325;
reg Range1_all_ones_reg_1789;
reg Range1_all_zeros_1_reg_2202;
reg Range1_all_zeros_2_reg_2332;
reg Range1_all_zeros_reg_1796;
reg Range2_all_ones_1_reg_2190;
reg Range2_all_ones_reg_1784;
reg [12:0] \add_25ns_25ns_25_2_1_U6.top_add_25ns_25ns_25_2_1_Adder_3_U.ain_s1 ;
reg [12:0] \add_25ns_25ns_25_2_1_U6.top_add_25ns_25ns_25_2_1_Adder_3_U.bin_s1 ;
reg \add_25ns_25ns_25_2_1_U6.top_add_25ns_25ns_25_2_1_Adder_3_U.carry_s1 ;
reg [11:0] \add_25ns_25ns_25_2_1_U6.top_add_25ns_25ns_25_2_1_Adder_3_U.sum_s1 ;
reg [12:0] \add_26ns_26ns_26_2_1_U5.top_add_26ns_26ns_26_2_1_Adder_2_U.ain_s1 ;
reg [12:0] \add_26ns_26ns_26_2_1_U5.top_add_26ns_26ns_26_2_1_Adder_2_U.bin_s1 ;
reg \add_26ns_26ns_26_2_1_U5.top_add_26ns_26ns_26_2_1_Adder_2_U.carry_s1 ;
reg [12:0] \add_26ns_26ns_26_2_1_U5.top_add_26ns_26ns_26_2_1_Adder_2_U.sum_s1 ;
reg \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_1_U.ain_s1 ;
reg \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_1_U.bin_s1 ;
reg \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_1_U.carry_s1 ;
reg \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_1_U.sum_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_17_U.ain_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_17_U.bin_s1 ;
reg \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_17_U.carry_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_17_U.sum_s1 ;
reg [15:0] \add_32s_32ns_32_2_1_U24.top_add_32s_32ns_32_2_1_Adder_19_U.ain_s1 ;
reg [15:0] \add_32s_32ns_32_2_1_U24.top_add_32s_32ns_32_2_1_Adder_19_U.bin_s1 ;
reg \add_32s_32ns_32_2_1_U24.top_add_32s_32ns_32_2_1_Adder_19_U.carry_s1 ;
reg [15:0] \add_32s_32ns_32_2_1_U24.top_add_32s_32ns_32_2_1_Adder_19_U.sum_s1 ;
reg [16:0] \add_33s_33s_33_2_1_U8.top_add_33s_33s_33_2_1_Adder_5_U.ain_s1 ;
reg [16:0] \add_33s_33s_33_2_1_U8.top_add_33s_33s_33_2_1_Adder_5_U.bin_s1 ;
reg \add_33s_33s_33_2_1_U8.top_add_33s_33s_33_2_1_Adder_5_U.carry_s1 ;
reg [15:0] \add_33s_33s_33_2_1_U8.top_add_33s_33s_33_2_1_Adder_5_U.sum_s1 ;
reg [19:0] \add_39s_39s_39_2_1_U21.top_add_39s_39s_39_2_1_Adder_16_U.ain_s1 ;
reg [19:0] \add_39s_39s_39_2_1_U21.top_add_39s_39s_39_2_1_Adder_16_U.bin_s1 ;
reg \add_39s_39s_39_2_1_U21.top_add_39s_39s_39_2_1_Adder_16_U.carry_s1 ;
reg [18:0] \add_39s_39s_39_2_1_U21.top_add_39s_39s_39_2_1_Adder_16_U.sum_s1 ;
reg [1:0] \add_3s_3ns_3_2_1_U11.top_add_3s_3ns_3_2_1_Adder_8_U.ain_s1 ;
reg [1:0] \add_3s_3ns_3_2_1_U11.top_add_3s_3ns_3_2_1_Adder_8_U.bin_s1 ;
reg \add_3s_3ns_3_2_1_U11.top_add_3s_3ns_3_2_1_Adder_8_U.carry_s1 ;
reg \add_3s_3ns_3_2_1_U11.top_add_3s_3ns_3_2_1_Adder_8_U.sum_s1 ;
reg [1:0] \add_4ns_4ns_4_2_1_U12.top_add_4ns_4ns_4_2_1_Adder_9_U.ain_s1 ;
reg [1:0] \add_4ns_4ns_4_2_1_U12.top_add_4ns_4ns_4_2_1_Adder_9_U.bin_s1 ;
reg \add_4ns_4ns_4_2_1_U12.top_add_4ns_4ns_4_2_1_Adder_9_U.carry_s1 ;
reg [1:0] \add_4ns_4ns_4_2_1_U12.top_add_4ns_4ns_4_2_1_Adder_9_U.sum_s1 ;
reg [1:0] \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_9_U.ain_s1 ;
reg [1:0] \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_9_U.bin_s1 ;
reg \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_9_U.carry_s1 ;
reg [1:0] \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_9_U.sum_s1 ;
reg [1:0] \add_4ns_4ns_4_2_1_U15.top_add_4ns_4ns_4_2_1_Adder_9_U.ain_s1 ;
reg [1:0] \add_4ns_4ns_4_2_1_U15.top_add_4ns_4ns_4_2_1_Adder_9_U.bin_s1 ;
reg \add_4ns_4ns_4_2_1_U15.top_add_4ns_4ns_4_2_1_Adder_9_U.carry_s1 ;
reg [1:0] \add_4ns_4ns_4_2_1_U15.top_add_4ns_4ns_4_2_1_Adder_9_U.sum_s1 ;
reg [1:0] \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_10_U.ain_s1 ;
reg [1:0] \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_10_U.bin_s1 ;
reg \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_10_U.carry_s1 ;
reg [1:0] \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_10_U.sum_s1 ;
reg [1:0] \add_4s_4ns_4_2_1_U16.top_add_4s_4ns_4_2_1_Adder_11_U.ain_s1 ;
reg [1:0] \add_4s_4ns_4_2_1_U16.top_add_4s_4ns_4_2_1_Adder_11_U.bin_s1 ;
reg \add_4s_4ns_4_2_1_U16.top_add_4s_4ns_4_2_1_Adder_11_U.carry_s1 ;
reg [1:0] \add_4s_4ns_4_2_1_U16.top_add_4s_4ns_4_2_1_Adder_11_U.sum_s1 ;
reg [2:0] \add_5ns_5s_5_2_1_U18.top_add_5ns_5s_5_2_1_Adder_13_U.ain_s1 ;
reg [2:0] \add_5ns_5s_5_2_1_U18.top_add_5ns_5s_5_2_1_Adder_13_U.bin_s1 ;
reg \add_5ns_5s_5_2_1_U18.top_add_5ns_5s_5_2_1_Adder_13_U.carry_s1 ;
reg [1:0] \add_5ns_5s_5_2_1_U18.top_add_5ns_5s_5_2_1_Adder_13_U.sum_s1 ;
reg [2:0] \add_5s_5s_5_2_1_U17.top_add_5s_5s_5_2_1_Adder_12_U.ain_s1 ;
reg [2:0] \add_5s_5s_5_2_1_U17.top_add_5s_5s_5_2_1_Adder_12_U.bin_s1 ;
reg \add_5s_5s_5_2_1_U17.top_add_5s_5s_5_2_1_Adder_12_U.carry_s1 ;
reg [1:0] \add_5s_5s_5_2_1_U17.top_add_5s_5s_5_2_1_Adder_12_U.sum_s1 ;
reg [2:0] \add_6ns_6s_6_2_1_U20.top_add_6ns_6s_6_2_1_Adder_15_U.ain_s1 ;
reg [2:0] \add_6ns_6s_6_2_1_U20.top_add_6ns_6s_6_2_1_Adder_15_U.bin_s1 ;
reg \add_6ns_6s_6_2_1_U20.top_add_6ns_6s_6_2_1_Adder_15_U.carry_s1 ;
reg [2:0] \add_6ns_6s_6_2_1_U20.top_add_6ns_6s_6_2_1_Adder_15_U.sum_s1 ;
reg [2:0] \add_6s_6s_6_2_1_U19.top_add_6s_6s_6_2_1_Adder_14_U.ain_s1 ;
reg [2:0] \add_6s_6s_6_2_1_U19.top_add_6s_6s_6_2_1_Adder_14_U.bin_s1 ;
reg \add_6s_6s_6_2_1_U19.top_add_6s_6s_6_2_1_Adder_14_U.carry_s1 ;
reg [2:0] \add_6s_6s_6_2_1_U19.top_add_6s_6s_6_2_1_Adder_14_U.sum_s1 ;
reg [3:0] \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_4_U.ain_s1 ;
reg [3:0] \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_4_U.bin_s1 ;
reg \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_4_U.carry_s1 ;
reg [3:0] \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_4_U.sum_s1 ;
reg [4:0] \add_9s_9ns_9_2_1_U3.top_add_9s_9ns_9_2_1_Adder_0_U.ain_s1 ;
reg [4:0] \add_9s_9ns_9_2_1_U3.top_add_9s_9ns_9_2_1_Adder_0_U.bin_s1 ;
reg \add_9s_9ns_9_2_1_U3.top_add_9s_9ns_9_2_1_Adder_0_U.carry_s1 ;
reg [3:0] \add_9s_9ns_9_2_1_U3.top_add_9s_9ns_9_2_1_Adder_0_U.sum_s1 ;
reg [4:0] \add_9s_9s_9_2_1_U23.top_add_9s_9s_9_2_1_Adder_18_U.ain_s1 ;
reg [4:0] \add_9s_9s_9_2_1_U23.top_add_9s_9s_9_2_1_Adder_18_U.bin_s1 ;
reg \add_9s_9s_9_2_1_U23.top_add_9s_9s_9_2_1_Adder_18_U.carry_s1 ;
reg [3:0] \add_9s_9s_9_2_1_U23.top_add_9s_9s_9_2_1_Adder_18_U.sum_s1 ;
reg [25:0] add_ln1192_1_reg_1927;
reg [24:0] add_ln1192_2_reg_1932;
reg [31:0] add_ln691_3_reg_2455;
reg [3:0] add_ln691_reg_2337;
reg [8:0] add_ln69_3_reg_2470;
reg [4:0] add_ln69_reg_2373;
reg and_ln408_reg_2234;
reg and_ln412_reg_1959;
reg and_ln414_reg_1811;
reg and_ln785_1_reg_2007;
reg and_ln786_1_reg_2228;
reg and_ln786_3_reg_2363;
reg and_ln786_reg_1982;
reg [31:0] ap_CS_fsm = 32'd1;
reg carry_1_reg_1952;
reg carry_3_reg_2183;
reg carry_5_reg_2318;
reg deleted_zeros_1_reg_2222;
reg deleted_zeros_reg_1970;
reg [24:0] empty_reg_1750;
reg icmp_ln414_reg_1773;
reg icmp_ln768_reg_1732;
reg icmp_ln785_reg_1869;
reg icmp_ln786_1_reg_1874;
reg icmp_ln786_2_reg_1737;
reg icmp_ln786_reg_1916;
reg icmp_ln790_reg_1879;
reg icmp_ln851_1_reg_2217;
reg icmp_ln851_2_reg_2378;
reg icmp_ln851_reg_2212;
reg [3:0] \mul_4s_4s_4_7_1_U1.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.a_reg0 ;
reg [3:0] \mul_4s_4s_4_7_1_U1.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.b_reg0 ;
reg [3:0] \mul_4s_4s_4_7_1_U1.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.buff0 ;
reg [3:0] \mul_4s_4s_4_7_1_U1.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.buff1 ;
reg [3:0] \mul_4s_4s_4_7_1_U1.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.buff2 ;
reg [3:0] \mul_4s_4s_4_7_1_U1.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.buff3 ;
reg [3:0] \mul_4s_4s_4_7_1_U1.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.buff4 ;
reg [3:0] \mul_4s_4s_8_7_1_U2.top_mul_4s_4s_8_7_1_Mul_DSP_1_U.a_reg0 ;
reg [3:0] \mul_4s_4s_8_7_1_U2.top_mul_4s_4s_8_7_1_Mul_DSP_1_U.b_reg0 ;
reg [7:0] \mul_4s_4s_8_7_1_U2.top_mul_4s_4s_8_7_1_Mul_DSP_1_U.buff0 ;
reg [7:0] \mul_4s_4s_8_7_1_U2.top_mul_4s_4s_8_7_1_Mul_DSP_1_U.buff1 ;
reg [7:0] \mul_4s_4s_8_7_1_U2.top_mul_4s_4s_8_7_1_Mul_DSP_1_U.buff2 ;
reg [7:0] \mul_4s_4s_8_7_1_U2.top_mul_4s_4s_8_7_1_Mul_DSP_1_U.buff3 ;
reg [7:0] \mul_4s_4s_8_7_1_U2.top_mul_4s_4s_8_7_1_Mul_DSP_1_U.buff4 ;
reg [1:0] op_12_V_reg_2172;
reg [3:0] op_15_V_reg_2393;
reg [3:0] op_16_V_reg_1705;
reg [7:0] op_17_V_reg_2313;
reg [4:0] op_23_V_reg_2398;
reg [5:0] op_25_V_reg_2423;
reg [3:0] op_3_V_reg_1816;
reg [7:0] op_4_V_reg_1693;
reg [7:0] op_8_V_reg_1964;
reg or_ln340_3_reg_2259;
reg or_ln340_reg_2001;
reg or_ln384_2_reg_2383;
reg or_ln384_reg_1947;
reg overflow_3_reg_1995;
reg overflow_4_reg_2357;
reg overflow_reg_1910;
reg p_Result_29_reg_1826;
reg [1:0] p_Result_2_reg_2132;
reg p_Result_30_reg_1755;
reg p_Result_31_reg_1768;
reg p_Result_32_reg_1893;
reg p_Result_33_reg_1778;
reg p_Result_34_reg_2080;
reg p_Result_36_reg_1942;
reg p_Result_37_reg_2033;
reg p_Result_38_reg_1720;
reg p_Result_39_reg_1698;
reg p_Result_40_reg_2111;
reg p_Result_41_reg_2122;
reg p_Result_43_reg_2299;
reg [6:0] p_Result_5_reg_2093;
reg [7:0] p_Result_6_reg_2098;
reg [7:0] p_Result_8_reg_1726;
reg [4:0] p_Result_s_reg_1838;
reg [3:0] p_Val2_12_reg_2117;
reg [3:0] p_Val2_13_reg_2294;
reg [1:0] p_Val2_2_reg_1763;
reg [1:0] p_Val2_3_reg_1884;
reg [7:0] p_Val2_7_reg_1937;
reg [7:0] p_Val2_8_reg_2027;
reg r_1_reg_2207;
reg r_reg_1806;
reg [3:0] ret_V_10_reg_2254;
reg [2:0] ret_V_15_reg_2178;
reg [10:0] ret_V_17_reg_2104;
reg [3:0] ret_V_18_reg_2269;
reg [3:0] ret_V_19_reg_2368;
reg [31:0] ret_V_20_cast_reg_2443;
reg [8:0] ret_V_20_reg_2138;
reg [3:0] ret_V_21_reg_2279;
reg [31:0] ret_V_22_reg_2155;
reg [3:0] ret_V_23_reg_2284;
reg [5:0] ret_V_24_reg_2413;
reg [38:0] ret_V_25_reg_2438;
reg [31:0] ret_V_26_reg_2465;
reg [3:0] ret_V_7_cast_reg_2160;
reg [3:0] ret_V_7_reg_2249;
reg [3:0] ret_V_reg_2143;
reg [7:0] ret_reg_1821;
reg [23:0] rhs_3_reg_2060;
reg sel_tmp11_reg_2070;
reg [7:0] select_ln340_1_reg_2289;
reg [1:0] select_ln340_reg_2065;
reg [2:0] select_ln703_reg_2012;
reg [3:0] sext_ln850_reg_2306;
reg [5:0] \sub_11ns_11s_11_2_1_U9.top_sub_11ns_11s_11_2_1_Adder_6_U.ain_s1 ;
reg [5:0] \sub_11ns_11s_11_2_1_U9.top_sub_11ns_11s_11_2_1_Adder_6_U.bin_s1 ;
reg \sub_11ns_11s_11_2_1_U9.top_sub_11ns_11s_11_2_1_Adder_6_U.carry_s1 ;
reg [4:0] \sub_11ns_11s_11_2_1_U9.top_sub_11ns_11s_11_2_1_Adder_6_U.sum_s1 ;
reg [4:0] \sub_9s_9s_9_2_1_U10.top_sub_9s_9s_9_2_1_Adder_7_U.ain_s1 ;
reg [4:0] \sub_9s_9s_9_2_1_U10.top_sub_9s_9s_9_2_1_Adder_7_U.bin_s1 ;
reg \sub_9s_9s_9_2_1_U10.top_sub_9s_9s_9_2_1_Adder_7_U.carry_s1 ;
reg [3:0] \sub_9s_9s_9_2_1_U10.top_sub_9s_9s_9_2_1_Adder_7_U.sum_s1 ;
reg [2:0] tmp_5_reg_2274;
reg tmp_reg_1832;
reg [25:0] trunc_ln1192_2_reg_1801;
reg [2:0] trunc_ln1192_3_reg_1864;
reg [1:0] trunc_ln1192_reg_1859;
reg trunc_ln703_reg_1854;
reg [3:0] trunc_ln718_1_reg_2127;
reg [1:0] trunc_ln790_reg_1844;
reg [4:0] trunc_ln851_1_reg_2150;
reg [22:0] trunc_ln851_2_reg_2167;
reg [5:0] trunc_ln851_3_reg_2352;
reg xor_ln416_1_reg_2087;
reg xor_ln416_reg_1921;
reg xor_ln785_2_reg_1976;
wire _0000_;
wire _0001_;
wire _0002_;
wire _0003_;
wire _0004_;
wire _0005_;
wire _0006_;
wire _0007_;
wire [25:0] _0008_;
wire [24:0] _0009_;
wire [31:0] _0010_;
wire [3:0] _0011_;
wire [8:0] _0012_;
wire [4:0] _0013_;
wire _0014_;
wire _0015_;
wire _0016_;
wire _0017_;
wire _0018_;
wire _0019_;
wire _0020_;
wire [31:0] _0021_;
wire _0022_;
wire _0023_;
wire _0024_;
wire _0025_;
wire _0026_;
wire [24:0] _0027_;
wire _0028_;
wire _0029_;
wire _0030_;
wire _0031_;
wire _0032_;
wire _0033_;
wire _0034_;
wire _0035_;
wire _0036_;
wire _0037_;
wire [1:0] _0038_;
wire [3:0] _0039_;
wire [3:0] _0040_;
wire [7:0] _0041_;
wire [4:0] _0042_;
wire [5:0] _0043_;
wire [3:0] _0044_;
wire [7:0] _0045_;
wire [7:0] _0046_;
wire _0047_;
wire _0048_;
wire _0049_;
wire _0050_;
wire _0051_;
wire _0052_;
wire _0053_;
wire _0054_;
wire [1:0] _0055_;
wire _0056_;
wire _0057_;
wire _0058_;
wire _0059_;
wire _0060_;
wire _0061_;
wire _0062_;
wire _0063_;
wire _0064_;
wire _0065_;
wire _0066_;
wire _0067_;
wire [6:0] _0068_;
wire [7:0] _0069_;
wire [7:0] _0070_;
wire [4:0] _0071_;
wire [3:0] _0072_;
wire [3:0] _0073_;
wire [1:0] _0074_;
wire [1:0] _0075_;
wire [7:0] _0076_;
wire [7:0] _0077_;
wire _0078_;
wire _0079_;
wire [3:0] _0080_;
wire [2:0] _0081_;
wire [10:0] _0082_;
wire [3:0] _0083_;
wire [3:0] _0084_;
wire [31:0] _0085_;
wire [8:0] _0086_;
wire [3:0] _0087_;
wire [31:0] _0088_;
wire [3:0] _0089_;
wire [5:0] _0090_;
wire [38:0] _0091_;
wire [31:0] _0092_;
wire [3:0] _0093_;
wire [3:0] _0094_;
wire [3:0] _0095_;
wire [7:0] _0096_;
wire [1:0] _0097_;
wire _0098_;
wire [7:0] _0099_;
wire [1:0] _0100_;
wire [2:0] _0101_;
wire [3:0] _0102_;
wire [2:0] _0103_;
wire _0104_;
wire [25:0] _0105_;
wire [2:0] _0106_;
wire [1:0] _0107_;
wire _0108_;
wire [3:0] _0109_;
wire [1:0] _0110_;
wire [4:0] _0111_;
wire [22:0] _0112_;
wire [5:0] _0113_;
wire _0114_;
wire _0115_;
wire _0116_;
wire [1:0] _0117_;
wire _0118_;
wire _0119_;
wire _0120_;
wire _0121_;
wire _0122_;
wire _0123_;
wire _0124_;
wire _0125_;
wire _0126_;
wire _0127_;
wire _0128_;
wire _0129_;
wire _0130_;
wire _0131_;
wire _0132_;
wire _0133_;
wire _0134_;
wire _0135_;
wire [12:0] _0136_;
wire [12:0] _0137_;
wire _0138_;
wire [11:0] _0139_;
wire [12:0] _0140_;
wire [13:0] _0141_;
wire [12:0] _0142_;
wire [12:0] _0143_;
wire _0144_;
wire [12:0] _0145_;
wire [13:0] _0146_;
wire [13:0] _0147_;
wire _0148_;
wire _0149_;
wire _0150_;
wire _0151_;
wire [1:0] _0152_;
wire [1:0] _0153_;
wire [15:0] _0154_;
wire [15:0] _0155_;
wire _0156_;
wire [15:0] _0157_;
wire [16:0] _0158_;
wire [16:0] _0159_;
wire [15:0] _0160_;
wire [15:0] _0161_;
wire _0162_;
wire [15:0] _0163_;
wire [16:0] _0164_;
wire [16:0] _0165_;
wire [16:0] _0166_;
wire [16:0] _0167_;
wire _0168_;
wire [15:0] _0169_;
wire [16:0] _0170_;
wire [17:0] _0171_;
wire [19:0] _0172_;
wire [19:0] _0173_;
wire _0174_;
wire [18:0] _0175_;
wire [19:0] _0176_;
wire [20:0] _0177_;
wire [1:0] _0178_;
wire [1:0] _0179_;
wire _0180_;
wire _0181_;
wire [1:0] _0182_;
wire [2:0] _0183_;
wire [1:0] _0184_;
wire [1:0] _0185_;
wire _0186_;
wire [1:0] _0187_;
wire [2:0] _0188_;
wire [2:0] _0189_;
wire [1:0] _0190_;
wire [1:0] _0191_;
wire _0192_;
wire [1:0] _0193_;
wire [2:0] _0194_;
wire [2:0] _0195_;
wire [1:0] _0196_;
wire [1:0] _0197_;
wire _0198_;
wire [1:0] _0199_;
wire [2:0] _0200_;
wire [2:0] _0201_;
wire [1:0] _0202_;
wire [1:0] _0203_;
wire _0204_;
wire [1:0] _0205_;
wire [2:0] _0206_;
wire [2:0] _0207_;
wire [1:0] _0208_;
wire [1:0] _0209_;
wire _0210_;
wire [1:0] _0211_;
wire [2:0] _0212_;
wire [2:0] _0213_;
wire [2:0] _0214_;
wire [2:0] _0215_;
wire _0216_;
wire [1:0] _0217_;
wire [2:0] _0218_;
wire [3:0] _0219_;
wire [2:0] _0220_;
wire [2:0] _0221_;
wire _0222_;
wire [1:0] _0223_;
wire [2:0] _0224_;
wire [3:0] _0225_;
wire [2:0] _0226_;
wire [2:0] _0227_;
wire _0228_;
wire [2:0] _0229_;
wire [3:0] _0230_;
wire [3:0] _0231_;
wire [2:0] _0232_;
wire [2:0] _0233_;
wire _0234_;
wire [2:0] _0235_;
wire [3:0] _0236_;
wire [3:0] _0237_;
wire [3:0] _0238_;
wire [3:0] _0239_;
wire _0240_;
wire [3:0] _0241_;
wire [4:0] _0242_;
wire [4:0] _0243_;
wire [4:0] _0244_;
wire [4:0] _0245_;
wire _0246_;
wire [3:0] _0247_;
wire [4:0] _0248_;
wire [5:0] _0249_;
wire [4:0] _0250_;
wire [4:0] _0251_;
wire _0252_;
wire [3:0] _0253_;
wire [4:0] _0254_;
wire [5:0] _0255_;
wire [3:0] _0256_;
wire [3:0] _0257_;
wire [3:0] _0258_;
wire [3:0] _0259_;
wire [3:0] _0260_;
wire [3:0] _0261_;
wire [3:0] _0262_;
wire [3:0] _0263_;
wire [3:0] _0264_;
wire [7:0] _0265_;
wire [7:0] _0266_;
wire [7:0] _0267_;
wire [7:0] _0268_;
wire [7:0] _0269_;
wire [5:0] _0270_;
wire [5:0] _0271_;
wire _0272_;
wire [4:0] _0273_;
wire [5:0] _0274_;
wire [6:0] _0275_;
wire [4:0] _0276_;
wire [4:0] _0277_;
wire _0278_;
wire [3:0] _0279_;
wire [4:0] _0280_;
wire [5:0] _0281_;
wire _0282_;
wire _0283_;
wire _0284_;
wire _0285_;
wire _0286_;
wire _0287_;
wire _0288_;
wire _0289_;
wire _0290_;
wire _0291_;
wire _0292_;
wire _0293_;
wire _0294_;
wire _0295_;
wire _0296_;
wire _0297_;
wire _0298_;
wire _0299_;
wire _0300_;
wire _0301_;
wire _0302_;
wire _0303_;
wire _0304_;
wire _0305_;
wire _0306_;
wire _0307_;
wire _0308_;
wire _0309_;
wire _0310_;
wire _0311_;
wire _0312_;
wire _0313_;
wire _0314_;
wire _0315_;
wire _0316_;
wire _0317_;
wire _0318_;
wire _0319_;
wire _0320_;
wire _0321_;
wire Range1_all_ones_1_fu_1158_p2;
wire Range1_all_ones_2_fu_1411_p2;
wire Range1_all_ones_fu_455_p2;
wire Range1_all_zeros_1_fu_1163_p2;
wire Range1_all_zeros_2_fu_1416_p2;
wire Range1_all_zeros_fu_461_p2;
wire Range2_all_ones_1_fu_1153_p2;
wire Range2_all_ones_2_fu_1438_p3;
wire Range2_all_ones_fu_439_p2;
wire \add_25ns_25ns_25_2_1_U6.ce ;
wire \add_25ns_25ns_25_2_1_U6.clk ;
wire [24:0] \add_25ns_25ns_25_2_1_U6.din0 ;
wire [24:0] \add_25ns_25ns_25_2_1_U6.din1 ;
wire [24:0] \add_25ns_25ns_25_2_1_U6.dout ;
wire \add_25ns_25ns_25_2_1_U6.reset ;
wire [24:0] \add_25ns_25ns_25_2_1_U6.top_add_25ns_25ns_25_2_1_Adder_3_U.a ;
wire [24:0] \add_25ns_25ns_25_2_1_U6.top_add_25ns_25ns_25_2_1_Adder_3_U.ain_s0 ;
wire [24:0] \add_25ns_25ns_25_2_1_U6.top_add_25ns_25ns_25_2_1_Adder_3_U.b ;
wire [24:0] \add_25ns_25ns_25_2_1_U6.top_add_25ns_25ns_25_2_1_Adder_3_U.bin_s0 ;
wire \add_25ns_25ns_25_2_1_U6.top_add_25ns_25ns_25_2_1_Adder_3_U.ce ;
wire \add_25ns_25ns_25_2_1_U6.top_add_25ns_25ns_25_2_1_Adder_3_U.clk ;
wire \add_25ns_25ns_25_2_1_U6.top_add_25ns_25ns_25_2_1_Adder_3_U.facout_s1 ;
wire \add_25ns_25ns_25_2_1_U6.top_add_25ns_25ns_25_2_1_Adder_3_U.facout_s2 ;
wire [11:0] \add_25ns_25ns_25_2_1_U6.top_add_25ns_25ns_25_2_1_Adder_3_U.fas_s1 ;
wire [12:0] \add_25ns_25ns_25_2_1_U6.top_add_25ns_25ns_25_2_1_Adder_3_U.fas_s2 ;
wire \add_25ns_25ns_25_2_1_U6.top_add_25ns_25ns_25_2_1_Adder_3_U.reset ;
wire [24:0] \add_25ns_25ns_25_2_1_U6.top_add_25ns_25ns_25_2_1_Adder_3_U.s ;
wire [11:0] \add_25ns_25ns_25_2_1_U6.top_add_25ns_25ns_25_2_1_Adder_3_U.u1.a ;
wire [11:0] \add_25ns_25ns_25_2_1_U6.top_add_25ns_25ns_25_2_1_Adder_3_U.u1.b ;
wire \add_25ns_25ns_25_2_1_U6.top_add_25ns_25ns_25_2_1_Adder_3_U.u1.cin ;
wire \add_25ns_25ns_25_2_1_U6.top_add_25ns_25ns_25_2_1_Adder_3_U.u1.cout ;
wire [11:0] \add_25ns_25ns_25_2_1_U6.top_add_25ns_25ns_25_2_1_Adder_3_U.u1.s ;
wire [12:0] \add_25ns_25ns_25_2_1_U6.top_add_25ns_25ns_25_2_1_Adder_3_U.u2.a ;
wire [12:0] \add_25ns_25ns_25_2_1_U6.top_add_25ns_25ns_25_2_1_Adder_3_U.u2.b ;
wire \add_25ns_25ns_25_2_1_U6.top_add_25ns_25ns_25_2_1_Adder_3_U.u2.cin ;
wire \add_25ns_25ns_25_2_1_U6.top_add_25ns_25ns_25_2_1_Adder_3_U.u2.cout ;
wire [12:0] \add_25ns_25ns_25_2_1_U6.top_add_25ns_25ns_25_2_1_Adder_3_U.u2.s ;
wire \add_26ns_26ns_26_2_1_U5.ce ;
wire \add_26ns_26ns_26_2_1_U5.clk ;
wire [25:0] \add_26ns_26ns_26_2_1_U5.din0 ;
wire [25:0] \add_26ns_26ns_26_2_1_U5.din1 ;
wire [25:0] \add_26ns_26ns_26_2_1_U5.dout ;
wire \add_26ns_26ns_26_2_1_U5.reset ;
wire [25:0] \add_26ns_26ns_26_2_1_U5.top_add_26ns_26ns_26_2_1_Adder_2_U.a ;
wire [25:0] \add_26ns_26ns_26_2_1_U5.top_add_26ns_26ns_26_2_1_Adder_2_U.ain_s0 ;
wire [25:0] \add_26ns_26ns_26_2_1_U5.top_add_26ns_26ns_26_2_1_Adder_2_U.b ;
wire [25:0] \add_26ns_26ns_26_2_1_U5.top_add_26ns_26ns_26_2_1_Adder_2_U.bin_s0 ;
wire \add_26ns_26ns_26_2_1_U5.top_add_26ns_26ns_26_2_1_Adder_2_U.ce ;
wire \add_26ns_26ns_26_2_1_U5.top_add_26ns_26ns_26_2_1_Adder_2_U.clk ;
wire \add_26ns_26ns_26_2_1_U5.top_add_26ns_26ns_26_2_1_Adder_2_U.facout_s1 ;
wire \add_26ns_26ns_26_2_1_U5.top_add_26ns_26ns_26_2_1_Adder_2_U.facout_s2 ;
wire [12:0] \add_26ns_26ns_26_2_1_U5.top_add_26ns_26ns_26_2_1_Adder_2_U.fas_s1 ;
wire [12:0] \add_26ns_26ns_26_2_1_U5.top_add_26ns_26ns_26_2_1_Adder_2_U.fas_s2 ;
wire \add_26ns_26ns_26_2_1_U5.top_add_26ns_26ns_26_2_1_Adder_2_U.reset ;
wire [25:0] \add_26ns_26ns_26_2_1_U5.top_add_26ns_26ns_26_2_1_Adder_2_U.s ;
wire [12:0] \add_26ns_26ns_26_2_1_U5.top_add_26ns_26ns_26_2_1_Adder_2_U.u1.a ;
wire [12:0] \add_26ns_26ns_26_2_1_U5.top_add_26ns_26ns_26_2_1_Adder_2_U.u1.b ;
wire \add_26ns_26ns_26_2_1_U5.top_add_26ns_26ns_26_2_1_Adder_2_U.u1.cin ;
wire \add_26ns_26ns_26_2_1_U5.top_add_26ns_26ns_26_2_1_Adder_2_U.u1.cout ;
wire [12:0] \add_26ns_26ns_26_2_1_U5.top_add_26ns_26ns_26_2_1_Adder_2_U.u1.s ;
wire [12:0] \add_26ns_26ns_26_2_1_U5.top_add_26ns_26ns_26_2_1_Adder_2_U.u2.a ;
wire [12:0] \add_26ns_26ns_26_2_1_U5.top_add_26ns_26ns_26_2_1_Adder_2_U.u2.b ;
wire \add_26ns_26ns_26_2_1_U5.top_add_26ns_26ns_26_2_1_Adder_2_U.u2.cin ;
wire \add_26ns_26ns_26_2_1_U5.top_add_26ns_26ns_26_2_1_Adder_2_U.u2.cout ;
wire [12:0] \add_26ns_26ns_26_2_1_U5.top_add_26ns_26ns_26_2_1_Adder_2_U.u2.s ;
wire \add_2ns_2ns_2_2_1_U4.ce ;
wire \add_2ns_2ns_2_2_1_U4.clk ;
wire [1:0] \add_2ns_2ns_2_2_1_U4.din0 ;
wire [1:0] \add_2ns_2ns_2_2_1_U4.din1 ;
wire [1:0] \add_2ns_2ns_2_2_1_U4.dout ;
wire \add_2ns_2ns_2_2_1_U4.reset ;
wire [1:0] \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_1_U.a ;
wire [1:0] \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_1_U.ain_s0 ;
wire [1:0] \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_1_U.b ;
wire [1:0] \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_1_U.bin_s0 ;
wire \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_1_U.ce ;
wire \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_1_U.clk ;
wire \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_1_U.facout_s1 ;
wire \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_1_U.facout_s2 ;
wire \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_1_U.fas_s1 ;
wire \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_1_U.fas_s2 ;
wire \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_1_U.reset ;
wire [1:0] \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_1_U.s ;
wire \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.a ;
wire \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.b ;
wire \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.cin ;
wire \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.cout ;
wire \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.s ;
wire \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.a ;
wire \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.b ;
wire \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.cin ;
wire \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.cout ;
wire \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.s ;
wire \add_32ns_32ns_32_2_1_U22.ce ;
wire \add_32ns_32ns_32_2_1_U22.clk ;
wire [31:0] \add_32ns_32ns_32_2_1_U22.din0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U22.din1 ;
wire [31:0] \add_32ns_32ns_32_2_1_U22.dout ;
wire \add_32ns_32ns_32_2_1_U22.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_17_U.a ;
wire [31:0] \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_17_U.ain_s0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_17_U.b ;
wire [31:0] \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_17_U.bin_s0 ;
wire \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_17_U.ce ;
wire \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_17_U.clk ;
wire \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_17_U.facout_s1 ;
wire \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_17_U.facout_s2 ;
wire [15:0] \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_17_U.fas_s1 ;
wire [15:0] \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_17_U.fas_s2 ;
wire \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_17_U.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_17_U.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_17_U.u1.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_17_U.u1.b ;
wire \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_17_U.u1.cin ;
wire \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_17_U.u1.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_17_U.u1.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_17_U.u2.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_17_U.u2.b ;
wire \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_17_U.u2.cin ;
wire \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_17_U.u2.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_17_U.u2.s ;
wire \add_32s_32ns_32_2_1_U24.ce ;
wire \add_32s_32ns_32_2_1_U24.clk ;
wire [31:0] \add_32s_32ns_32_2_1_U24.din0 ;
wire [31:0] \add_32s_32ns_32_2_1_U24.din1 ;
wire [31:0] \add_32s_32ns_32_2_1_U24.dout ;
wire \add_32s_32ns_32_2_1_U24.reset ;
wire [31:0] \add_32s_32ns_32_2_1_U24.top_add_32s_32ns_32_2_1_Adder_19_U.a ;
wire [31:0] \add_32s_32ns_32_2_1_U24.top_add_32s_32ns_32_2_1_Adder_19_U.ain_s0 ;
wire [31:0] \add_32s_32ns_32_2_1_U24.top_add_32s_32ns_32_2_1_Adder_19_U.b ;
wire [31:0] \add_32s_32ns_32_2_1_U24.top_add_32s_32ns_32_2_1_Adder_19_U.bin_s0 ;
wire \add_32s_32ns_32_2_1_U24.top_add_32s_32ns_32_2_1_Adder_19_U.ce ;
wire \add_32s_32ns_32_2_1_U24.top_add_32s_32ns_32_2_1_Adder_19_U.clk ;
wire \add_32s_32ns_32_2_1_U24.top_add_32s_32ns_32_2_1_Adder_19_U.facout_s1 ;
wire \add_32s_32ns_32_2_1_U24.top_add_32s_32ns_32_2_1_Adder_19_U.facout_s2 ;
wire [15:0] \add_32s_32ns_32_2_1_U24.top_add_32s_32ns_32_2_1_Adder_19_U.fas_s1 ;
wire [15:0] \add_32s_32ns_32_2_1_U24.top_add_32s_32ns_32_2_1_Adder_19_U.fas_s2 ;
wire \add_32s_32ns_32_2_1_U24.top_add_32s_32ns_32_2_1_Adder_19_U.reset ;
wire [31:0] \add_32s_32ns_32_2_1_U24.top_add_32s_32ns_32_2_1_Adder_19_U.s ;
wire [15:0] \add_32s_32ns_32_2_1_U24.top_add_32s_32ns_32_2_1_Adder_19_U.u1.a ;
wire [15:0] \add_32s_32ns_32_2_1_U24.top_add_32s_32ns_32_2_1_Adder_19_U.u1.b ;
wire \add_32s_32ns_32_2_1_U24.top_add_32s_32ns_32_2_1_Adder_19_U.u1.cin ;
wire \add_32s_32ns_32_2_1_U24.top_add_32s_32ns_32_2_1_Adder_19_U.u1.cout ;
wire [15:0] \add_32s_32ns_32_2_1_U24.top_add_32s_32ns_32_2_1_Adder_19_U.u1.s ;
wire [15:0] \add_32s_32ns_32_2_1_U24.top_add_32s_32ns_32_2_1_Adder_19_U.u2.a ;
wire [15:0] \add_32s_32ns_32_2_1_U24.top_add_32s_32ns_32_2_1_Adder_19_U.u2.b ;
wire \add_32s_32ns_32_2_1_U24.top_add_32s_32ns_32_2_1_Adder_19_U.u2.cin ;
wire \add_32s_32ns_32_2_1_U24.top_add_32s_32ns_32_2_1_Adder_19_U.u2.cout ;
wire [15:0] \add_32s_32ns_32_2_1_U24.top_add_32s_32ns_32_2_1_Adder_19_U.u2.s ;
wire \add_33s_33s_33_2_1_U8.ce ;
wire \add_33s_33s_33_2_1_U8.clk ;
wire [32:0] \add_33s_33s_33_2_1_U8.din0 ;
wire [32:0] \add_33s_33s_33_2_1_U8.din1 ;
wire [32:0] \add_33s_33s_33_2_1_U8.dout ;
wire \add_33s_33s_33_2_1_U8.reset ;
wire [32:0] \add_33s_33s_33_2_1_U8.top_add_33s_33s_33_2_1_Adder_5_U.a ;
wire [32:0] \add_33s_33s_33_2_1_U8.top_add_33s_33s_33_2_1_Adder_5_U.ain_s0 ;
wire [32:0] \add_33s_33s_33_2_1_U8.top_add_33s_33s_33_2_1_Adder_5_U.b ;
wire [32:0] \add_33s_33s_33_2_1_U8.top_add_33s_33s_33_2_1_Adder_5_U.bin_s0 ;
wire \add_33s_33s_33_2_1_U8.top_add_33s_33s_33_2_1_Adder_5_U.ce ;
wire \add_33s_33s_33_2_1_U8.top_add_33s_33s_33_2_1_Adder_5_U.clk ;
wire \add_33s_33s_33_2_1_U8.top_add_33s_33s_33_2_1_Adder_5_U.facout_s1 ;
wire \add_33s_33s_33_2_1_U8.top_add_33s_33s_33_2_1_Adder_5_U.facout_s2 ;
wire [15:0] \add_33s_33s_33_2_1_U8.top_add_33s_33s_33_2_1_Adder_5_U.fas_s1 ;
wire [16:0] \add_33s_33s_33_2_1_U8.top_add_33s_33s_33_2_1_Adder_5_U.fas_s2 ;
wire \add_33s_33s_33_2_1_U8.top_add_33s_33s_33_2_1_Adder_5_U.reset ;
wire [32:0] \add_33s_33s_33_2_1_U8.top_add_33s_33s_33_2_1_Adder_5_U.s ;
wire [15:0] \add_33s_33s_33_2_1_U8.top_add_33s_33s_33_2_1_Adder_5_U.u1.a ;
wire [15:0] \add_33s_33s_33_2_1_U8.top_add_33s_33s_33_2_1_Adder_5_U.u1.b ;
wire \add_33s_33s_33_2_1_U8.top_add_33s_33s_33_2_1_Adder_5_U.u1.cin ;
wire \add_33s_33s_33_2_1_U8.top_add_33s_33s_33_2_1_Adder_5_U.u1.cout ;
wire [15:0] \add_33s_33s_33_2_1_U8.top_add_33s_33s_33_2_1_Adder_5_U.u1.s ;
wire [16:0] \add_33s_33s_33_2_1_U8.top_add_33s_33s_33_2_1_Adder_5_U.u2.a ;
wire [16:0] \add_33s_33s_33_2_1_U8.top_add_33s_33s_33_2_1_Adder_5_U.u2.b ;
wire \add_33s_33s_33_2_1_U8.top_add_33s_33s_33_2_1_Adder_5_U.u2.cin ;
wire \add_33s_33s_33_2_1_U8.top_add_33s_33s_33_2_1_Adder_5_U.u2.cout ;
wire [16:0] \add_33s_33s_33_2_1_U8.top_add_33s_33s_33_2_1_Adder_5_U.u2.s ;
wire \add_39s_39s_39_2_1_U21.ce ;
wire \add_39s_39s_39_2_1_U21.clk ;
wire [38:0] \add_39s_39s_39_2_1_U21.din0 ;
wire [38:0] \add_39s_39s_39_2_1_U21.din1 ;
wire [38:0] \add_39s_39s_39_2_1_U21.dout ;
wire \add_39s_39s_39_2_1_U21.reset ;
wire [38:0] \add_39s_39s_39_2_1_U21.top_add_39s_39s_39_2_1_Adder_16_U.a ;
wire [38:0] \add_39s_39s_39_2_1_U21.top_add_39s_39s_39_2_1_Adder_16_U.ain_s0 ;
wire [38:0] \add_39s_39s_39_2_1_U21.top_add_39s_39s_39_2_1_Adder_16_U.b ;
wire [38:0] \add_39s_39s_39_2_1_U21.top_add_39s_39s_39_2_1_Adder_16_U.bin_s0 ;
wire \add_39s_39s_39_2_1_U21.top_add_39s_39s_39_2_1_Adder_16_U.ce ;
wire \add_39s_39s_39_2_1_U21.top_add_39s_39s_39_2_1_Adder_16_U.clk ;
wire \add_39s_39s_39_2_1_U21.top_add_39s_39s_39_2_1_Adder_16_U.facout_s1 ;
wire \add_39s_39s_39_2_1_U21.top_add_39s_39s_39_2_1_Adder_16_U.facout_s2 ;
wire [18:0] \add_39s_39s_39_2_1_U21.top_add_39s_39s_39_2_1_Adder_16_U.fas_s1 ;
wire [19:0] \add_39s_39s_39_2_1_U21.top_add_39s_39s_39_2_1_Adder_16_U.fas_s2 ;
wire \add_39s_39s_39_2_1_U21.top_add_39s_39s_39_2_1_Adder_16_U.reset ;
wire [38:0] \add_39s_39s_39_2_1_U21.top_add_39s_39s_39_2_1_Adder_16_U.s ;
wire [18:0] \add_39s_39s_39_2_1_U21.top_add_39s_39s_39_2_1_Adder_16_U.u1.a ;
wire [18:0] \add_39s_39s_39_2_1_U21.top_add_39s_39s_39_2_1_Adder_16_U.u1.b ;
wire \add_39s_39s_39_2_1_U21.top_add_39s_39s_39_2_1_Adder_16_U.u1.cin ;
wire \add_39s_39s_39_2_1_U21.top_add_39s_39s_39_2_1_Adder_16_U.u1.cout ;
wire [18:0] \add_39s_39s_39_2_1_U21.top_add_39s_39s_39_2_1_Adder_16_U.u1.s ;
wire [19:0] \add_39s_39s_39_2_1_U21.top_add_39s_39s_39_2_1_Adder_16_U.u2.a ;
wire [19:0] \add_39s_39s_39_2_1_U21.top_add_39s_39s_39_2_1_Adder_16_U.u2.b ;
wire \add_39s_39s_39_2_1_U21.top_add_39s_39s_39_2_1_Adder_16_U.u2.cin ;
wire \add_39s_39s_39_2_1_U21.top_add_39s_39s_39_2_1_Adder_16_U.u2.cout ;
wire [19:0] \add_39s_39s_39_2_1_U21.top_add_39s_39s_39_2_1_Adder_16_U.u2.s ;
wire \add_3s_3ns_3_2_1_U11.ce ;
wire \add_3s_3ns_3_2_1_U11.clk ;
wire [2:0] \add_3s_3ns_3_2_1_U11.din0 ;
wire [2:0] \add_3s_3ns_3_2_1_U11.din1 ;
wire [2:0] \add_3s_3ns_3_2_1_U11.dout ;
wire \add_3s_3ns_3_2_1_U11.reset ;
wire [2:0] \add_3s_3ns_3_2_1_U11.top_add_3s_3ns_3_2_1_Adder_8_U.a ;
wire [2:0] \add_3s_3ns_3_2_1_U11.top_add_3s_3ns_3_2_1_Adder_8_U.ain_s0 ;
wire [2:0] \add_3s_3ns_3_2_1_U11.top_add_3s_3ns_3_2_1_Adder_8_U.b ;
wire [2:0] \add_3s_3ns_3_2_1_U11.top_add_3s_3ns_3_2_1_Adder_8_U.bin_s0 ;
wire \add_3s_3ns_3_2_1_U11.top_add_3s_3ns_3_2_1_Adder_8_U.ce ;
wire \add_3s_3ns_3_2_1_U11.top_add_3s_3ns_3_2_1_Adder_8_U.clk ;
wire \add_3s_3ns_3_2_1_U11.top_add_3s_3ns_3_2_1_Adder_8_U.facout_s1 ;
wire \add_3s_3ns_3_2_1_U11.top_add_3s_3ns_3_2_1_Adder_8_U.facout_s2 ;
wire \add_3s_3ns_3_2_1_U11.top_add_3s_3ns_3_2_1_Adder_8_U.fas_s1 ;
wire [1:0] \add_3s_3ns_3_2_1_U11.top_add_3s_3ns_3_2_1_Adder_8_U.fas_s2 ;
wire \add_3s_3ns_3_2_1_U11.top_add_3s_3ns_3_2_1_Adder_8_U.reset ;
wire [2:0] \add_3s_3ns_3_2_1_U11.top_add_3s_3ns_3_2_1_Adder_8_U.s ;
wire \add_3s_3ns_3_2_1_U11.top_add_3s_3ns_3_2_1_Adder_8_U.u1.a ;
wire \add_3s_3ns_3_2_1_U11.top_add_3s_3ns_3_2_1_Adder_8_U.u1.b ;
wire \add_3s_3ns_3_2_1_U11.top_add_3s_3ns_3_2_1_Adder_8_U.u1.cin ;
wire \add_3s_3ns_3_2_1_U11.top_add_3s_3ns_3_2_1_Adder_8_U.u1.cout ;
wire \add_3s_3ns_3_2_1_U11.top_add_3s_3ns_3_2_1_Adder_8_U.u1.s ;
wire [1:0] \add_3s_3ns_3_2_1_U11.top_add_3s_3ns_3_2_1_Adder_8_U.u2.a ;
wire [1:0] \add_3s_3ns_3_2_1_U11.top_add_3s_3ns_3_2_1_Adder_8_U.u2.b ;
wire \add_3s_3ns_3_2_1_U11.top_add_3s_3ns_3_2_1_Adder_8_U.u2.cin ;
wire \add_3s_3ns_3_2_1_U11.top_add_3s_3ns_3_2_1_Adder_8_U.u2.cout ;
wire [1:0] \add_3s_3ns_3_2_1_U11.top_add_3s_3ns_3_2_1_Adder_8_U.u2.s ;
wire \add_4ns_4ns_4_2_1_U12.ce ;
wire \add_4ns_4ns_4_2_1_U12.clk ;
wire [3:0] \add_4ns_4ns_4_2_1_U12.din0 ;
wire [3:0] \add_4ns_4ns_4_2_1_U12.din1 ;
wire [3:0] \add_4ns_4ns_4_2_1_U12.dout ;
wire \add_4ns_4ns_4_2_1_U12.reset ;
wire [3:0] \add_4ns_4ns_4_2_1_U12.top_add_4ns_4ns_4_2_1_Adder_9_U.a ;
wire [3:0] \add_4ns_4ns_4_2_1_U12.top_add_4ns_4ns_4_2_1_Adder_9_U.ain_s0 ;
wire [3:0] \add_4ns_4ns_4_2_1_U12.top_add_4ns_4ns_4_2_1_Adder_9_U.b ;
wire [3:0] \add_4ns_4ns_4_2_1_U12.top_add_4ns_4ns_4_2_1_Adder_9_U.bin_s0 ;
wire \add_4ns_4ns_4_2_1_U12.top_add_4ns_4ns_4_2_1_Adder_9_U.ce ;
wire \add_4ns_4ns_4_2_1_U12.top_add_4ns_4ns_4_2_1_Adder_9_U.clk ;
wire \add_4ns_4ns_4_2_1_U12.top_add_4ns_4ns_4_2_1_Adder_9_U.facout_s1 ;
wire \add_4ns_4ns_4_2_1_U12.top_add_4ns_4ns_4_2_1_Adder_9_U.facout_s2 ;
wire [1:0] \add_4ns_4ns_4_2_1_U12.top_add_4ns_4ns_4_2_1_Adder_9_U.fas_s1 ;
wire [1:0] \add_4ns_4ns_4_2_1_U12.top_add_4ns_4ns_4_2_1_Adder_9_U.fas_s2 ;
wire \add_4ns_4ns_4_2_1_U12.top_add_4ns_4ns_4_2_1_Adder_9_U.reset ;
wire [3:0] \add_4ns_4ns_4_2_1_U12.top_add_4ns_4ns_4_2_1_Adder_9_U.s ;
wire [1:0] \add_4ns_4ns_4_2_1_U12.top_add_4ns_4ns_4_2_1_Adder_9_U.u1.a ;
wire [1:0] \add_4ns_4ns_4_2_1_U12.top_add_4ns_4ns_4_2_1_Adder_9_U.u1.b ;
wire \add_4ns_4ns_4_2_1_U12.top_add_4ns_4ns_4_2_1_Adder_9_U.u1.cin ;
wire \add_4ns_4ns_4_2_1_U12.top_add_4ns_4ns_4_2_1_Adder_9_U.u1.cout ;
wire [1:0] \add_4ns_4ns_4_2_1_U12.top_add_4ns_4ns_4_2_1_Adder_9_U.u1.s ;
wire [1:0] \add_4ns_4ns_4_2_1_U12.top_add_4ns_4ns_4_2_1_Adder_9_U.u2.a ;
wire [1:0] \add_4ns_4ns_4_2_1_U12.top_add_4ns_4ns_4_2_1_Adder_9_U.u2.b ;
wire \add_4ns_4ns_4_2_1_U12.top_add_4ns_4ns_4_2_1_Adder_9_U.u2.cin ;
wire \add_4ns_4ns_4_2_1_U12.top_add_4ns_4ns_4_2_1_Adder_9_U.u2.cout ;
wire [1:0] \add_4ns_4ns_4_2_1_U12.top_add_4ns_4ns_4_2_1_Adder_9_U.u2.s ;
wire \add_4ns_4ns_4_2_1_U13.ce ;
wire \add_4ns_4ns_4_2_1_U13.clk ;
wire [3:0] \add_4ns_4ns_4_2_1_U13.din0 ;
wire [3:0] \add_4ns_4ns_4_2_1_U13.din1 ;
wire [3:0] \add_4ns_4ns_4_2_1_U13.dout ;
wire \add_4ns_4ns_4_2_1_U13.reset ;
wire [3:0] \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_9_U.a ;
wire [3:0] \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_9_U.ain_s0 ;
wire [3:0] \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_9_U.b ;
wire [3:0] \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_9_U.bin_s0 ;
wire \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_9_U.ce ;
wire \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_9_U.clk ;
wire \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_9_U.facout_s1 ;
wire \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_9_U.facout_s2 ;
wire [1:0] \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_9_U.fas_s1 ;
wire [1:0] \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_9_U.fas_s2 ;
wire \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_9_U.reset ;
wire [3:0] \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_9_U.s ;
wire [1:0] \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_9_U.u1.a ;
wire [1:0] \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_9_U.u1.b ;
wire \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_9_U.u1.cin ;
wire \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_9_U.u1.cout ;
wire [1:0] \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_9_U.u1.s ;
wire [1:0] \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_9_U.u2.a ;
wire [1:0] \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_9_U.u2.b ;
wire \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_9_U.u2.cin ;
wire \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_9_U.u2.cout ;
wire [1:0] \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_9_U.u2.s ;
wire \add_4ns_4ns_4_2_1_U15.ce ;
wire \add_4ns_4ns_4_2_1_U15.clk ;
wire [3:0] \add_4ns_4ns_4_2_1_U15.din0 ;
wire [3:0] \add_4ns_4ns_4_2_1_U15.din1 ;
wire [3:0] \add_4ns_4ns_4_2_1_U15.dout ;
wire \add_4ns_4ns_4_2_1_U15.reset ;
wire [3:0] \add_4ns_4ns_4_2_1_U15.top_add_4ns_4ns_4_2_1_Adder_9_U.a ;
wire [3:0] \add_4ns_4ns_4_2_1_U15.top_add_4ns_4ns_4_2_1_Adder_9_U.ain_s0 ;
wire [3:0] \add_4ns_4ns_4_2_1_U15.top_add_4ns_4ns_4_2_1_Adder_9_U.b ;
wire [3:0] \add_4ns_4ns_4_2_1_U15.top_add_4ns_4ns_4_2_1_Adder_9_U.bin_s0 ;
wire \add_4ns_4ns_4_2_1_U15.top_add_4ns_4ns_4_2_1_Adder_9_U.ce ;
wire \add_4ns_4ns_4_2_1_U15.top_add_4ns_4ns_4_2_1_Adder_9_U.clk ;
wire \add_4ns_4ns_4_2_1_U15.top_add_4ns_4ns_4_2_1_Adder_9_U.facout_s1 ;
wire \add_4ns_4ns_4_2_1_U15.top_add_4ns_4ns_4_2_1_Adder_9_U.facout_s2 ;
wire [1:0] \add_4ns_4ns_4_2_1_U15.top_add_4ns_4ns_4_2_1_Adder_9_U.fas_s1 ;
wire [1:0] \add_4ns_4ns_4_2_1_U15.top_add_4ns_4ns_4_2_1_Adder_9_U.fas_s2 ;
wire \add_4ns_4ns_4_2_1_U15.top_add_4ns_4ns_4_2_1_Adder_9_U.reset ;
wire [3:0] \add_4ns_4ns_4_2_1_U15.top_add_4ns_4ns_4_2_1_Adder_9_U.s ;
wire [1:0] \add_4ns_4ns_4_2_1_U15.top_add_4ns_4ns_4_2_1_Adder_9_U.u1.a ;
wire [1:0] \add_4ns_4ns_4_2_1_U15.top_add_4ns_4ns_4_2_1_Adder_9_U.u1.b ;
wire \add_4ns_4ns_4_2_1_U15.top_add_4ns_4ns_4_2_1_Adder_9_U.u1.cin ;
wire \add_4ns_4ns_4_2_1_U15.top_add_4ns_4ns_4_2_1_Adder_9_U.u1.cout ;
wire [1:0] \add_4ns_4ns_4_2_1_U15.top_add_4ns_4ns_4_2_1_Adder_9_U.u1.s ;
wire [1:0] \add_4ns_4ns_4_2_1_U15.top_add_4ns_4ns_4_2_1_Adder_9_U.u2.a ;
wire [1:0] \add_4ns_4ns_4_2_1_U15.top_add_4ns_4ns_4_2_1_Adder_9_U.u2.b ;
wire \add_4ns_4ns_4_2_1_U15.top_add_4ns_4ns_4_2_1_Adder_9_U.u2.cin ;
wire \add_4ns_4ns_4_2_1_U15.top_add_4ns_4ns_4_2_1_Adder_9_U.u2.cout ;
wire [1:0] \add_4ns_4ns_4_2_1_U15.top_add_4ns_4ns_4_2_1_Adder_9_U.u2.s ;
wire \add_4ns_4s_4_2_1_U14.ce ;
wire \add_4ns_4s_4_2_1_U14.clk ;
wire [3:0] \add_4ns_4s_4_2_1_U14.din0 ;
wire [3:0] \add_4ns_4s_4_2_1_U14.din1 ;
wire [3:0] \add_4ns_4s_4_2_1_U14.dout ;
wire \add_4ns_4s_4_2_1_U14.reset ;
wire [3:0] \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_10_U.a ;
wire [3:0] \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_10_U.ain_s0 ;
wire [3:0] \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_10_U.b ;
wire [3:0] \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_10_U.bin_s0 ;
wire \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_10_U.ce ;
wire \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_10_U.clk ;
wire \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_10_U.facout_s1 ;
wire \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_10_U.facout_s2 ;
wire [1:0] \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_10_U.fas_s1 ;
wire [1:0] \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_10_U.fas_s2 ;
wire \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_10_U.reset ;
wire [3:0] \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_10_U.s ;
wire [1:0] \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_10_U.u1.a ;
wire [1:0] \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_10_U.u1.b ;
wire \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_10_U.u1.cin ;
wire \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_10_U.u1.cout ;
wire [1:0] \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_10_U.u1.s ;
wire [1:0] \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_10_U.u2.a ;
wire [1:0] \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_10_U.u2.b ;
wire \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_10_U.u2.cin ;
wire \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_10_U.u2.cout ;
wire [1:0] \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_10_U.u2.s ;
wire \add_4s_4ns_4_2_1_U16.ce ;
wire \add_4s_4ns_4_2_1_U16.clk ;
wire [3:0] \add_4s_4ns_4_2_1_U16.din0 ;
wire [3:0] \add_4s_4ns_4_2_1_U16.din1 ;
wire [3:0] \add_4s_4ns_4_2_1_U16.dout ;
wire \add_4s_4ns_4_2_1_U16.reset ;
wire [3:0] \add_4s_4ns_4_2_1_U16.top_add_4s_4ns_4_2_1_Adder_11_U.a ;
wire [3:0] \add_4s_4ns_4_2_1_U16.top_add_4s_4ns_4_2_1_Adder_11_U.ain_s0 ;
wire [3:0] \add_4s_4ns_4_2_1_U16.top_add_4s_4ns_4_2_1_Adder_11_U.b ;
wire [3:0] \add_4s_4ns_4_2_1_U16.top_add_4s_4ns_4_2_1_Adder_11_U.bin_s0 ;
wire \add_4s_4ns_4_2_1_U16.top_add_4s_4ns_4_2_1_Adder_11_U.ce ;
wire \add_4s_4ns_4_2_1_U16.top_add_4s_4ns_4_2_1_Adder_11_U.clk ;
wire \add_4s_4ns_4_2_1_U16.top_add_4s_4ns_4_2_1_Adder_11_U.facout_s1 ;
wire \add_4s_4ns_4_2_1_U16.top_add_4s_4ns_4_2_1_Adder_11_U.facout_s2 ;
wire [1:0] \add_4s_4ns_4_2_1_U16.top_add_4s_4ns_4_2_1_Adder_11_U.fas_s1 ;
wire [1:0] \add_4s_4ns_4_2_1_U16.top_add_4s_4ns_4_2_1_Adder_11_U.fas_s2 ;
wire \add_4s_4ns_4_2_1_U16.top_add_4s_4ns_4_2_1_Adder_11_U.reset ;
wire [3:0] \add_4s_4ns_4_2_1_U16.top_add_4s_4ns_4_2_1_Adder_11_U.s ;
wire [1:0] \add_4s_4ns_4_2_1_U16.top_add_4s_4ns_4_2_1_Adder_11_U.u1.a ;
wire [1:0] \add_4s_4ns_4_2_1_U16.top_add_4s_4ns_4_2_1_Adder_11_U.u1.b ;
wire \add_4s_4ns_4_2_1_U16.top_add_4s_4ns_4_2_1_Adder_11_U.u1.cin ;
wire \add_4s_4ns_4_2_1_U16.top_add_4s_4ns_4_2_1_Adder_11_U.u1.cout ;
wire [1:0] \add_4s_4ns_4_2_1_U16.top_add_4s_4ns_4_2_1_Adder_11_U.u1.s ;
wire [1:0] \add_4s_4ns_4_2_1_U16.top_add_4s_4ns_4_2_1_Adder_11_U.u2.a ;
wire [1:0] \add_4s_4ns_4_2_1_U16.top_add_4s_4ns_4_2_1_Adder_11_U.u2.b ;
wire \add_4s_4ns_4_2_1_U16.top_add_4s_4ns_4_2_1_Adder_11_U.u2.cin ;
wire \add_4s_4ns_4_2_1_U16.top_add_4s_4ns_4_2_1_Adder_11_U.u2.cout ;
wire [1:0] \add_4s_4ns_4_2_1_U16.top_add_4s_4ns_4_2_1_Adder_11_U.u2.s ;
wire \add_5ns_5s_5_2_1_U18.ce ;
wire \add_5ns_5s_5_2_1_U18.clk ;
wire [4:0] \add_5ns_5s_5_2_1_U18.din0 ;
wire [4:0] \add_5ns_5s_5_2_1_U18.din1 ;
wire [4:0] \add_5ns_5s_5_2_1_U18.dout ;
wire \add_5ns_5s_5_2_1_U18.reset ;
wire [4:0] \add_5ns_5s_5_2_1_U18.top_add_5ns_5s_5_2_1_Adder_13_U.a ;
wire [4:0] \add_5ns_5s_5_2_1_U18.top_add_5ns_5s_5_2_1_Adder_13_U.ain_s0 ;
wire [4:0] \add_5ns_5s_5_2_1_U18.top_add_5ns_5s_5_2_1_Adder_13_U.b ;
wire [4:0] \add_5ns_5s_5_2_1_U18.top_add_5ns_5s_5_2_1_Adder_13_U.bin_s0 ;
wire \add_5ns_5s_5_2_1_U18.top_add_5ns_5s_5_2_1_Adder_13_U.ce ;
wire \add_5ns_5s_5_2_1_U18.top_add_5ns_5s_5_2_1_Adder_13_U.clk ;
wire \add_5ns_5s_5_2_1_U18.top_add_5ns_5s_5_2_1_Adder_13_U.facout_s1 ;
wire \add_5ns_5s_5_2_1_U18.top_add_5ns_5s_5_2_1_Adder_13_U.facout_s2 ;
wire [1:0] \add_5ns_5s_5_2_1_U18.top_add_5ns_5s_5_2_1_Adder_13_U.fas_s1 ;
wire [2:0] \add_5ns_5s_5_2_1_U18.top_add_5ns_5s_5_2_1_Adder_13_U.fas_s2 ;
wire \add_5ns_5s_5_2_1_U18.top_add_5ns_5s_5_2_1_Adder_13_U.reset ;
wire [4:0] \add_5ns_5s_5_2_1_U18.top_add_5ns_5s_5_2_1_Adder_13_U.s ;
wire [1:0] \add_5ns_5s_5_2_1_U18.top_add_5ns_5s_5_2_1_Adder_13_U.u1.a ;
wire [1:0] \add_5ns_5s_5_2_1_U18.top_add_5ns_5s_5_2_1_Adder_13_U.u1.b ;
wire \add_5ns_5s_5_2_1_U18.top_add_5ns_5s_5_2_1_Adder_13_U.u1.cin ;
wire \add_5ns_5s_5_2_1_U18.top_add_5ns_5s_5_2_1_Adder_13_U.u1.cout ;
wire [1:0] \add_5ns_5s_5_2_1_U18.top_add_5ns_5s_5_2_1_Adder_13_U.u1.s ;
wire [2:0] \add_5ns_5s_5_2_1_U18.top_add_5ns_5s_5_2_1_Adder_13_U.u2.a ;
wire [2:0] \add_5ns_5s_5_2_1_U18.top_add_5ns_5s_5_2_1_Adder_13_U.u2.b ;
wire \add_5ns_5s_5_2_1_U18.top_add_5ns_5s_5_2_1_Adder_13_U.u2.cin ;
wire \add_5ns_5s_5_2_1_U18.top_add_5ns_5s_5_2_1_Adder_13_U.u2.cout ;
wire [2:0] \add_5ns_5s_5_2_1_U18.top_add_5ns_5s_5_2_1_Adder_13_U.u2.s ;
wire \add_5s_5s_5_2_1_U17.ce ;
wire \add_5s_5s_5_2_1_U17.clk ;
wire [4:0] \add_5s_5s_5_2_1_U17.din0 ;
wire [4:0] \add_5s_5s_5_2_1_U17.din1 ;
wire [4:0] \add_5s_5s_5_2_1_U17.dout ;
wire \add_5s_5s_5_2_1_U17.reset ;
wire [4:0] \add_5s_5s_5_2_1_U17.top_add_5s_5s_5_2_1_Adder_12_U.a ;
wire [4:0] \add_5s_5s_5_2_1_U17.top_add_5s_5s_5_2_1_Adder_12_U.ain_s0 ;
wire [4:0] \add_5s_5s_5_2_1_U17.top_add_5s_5s_5_2_1_Adder_12_U.b ;
wire [4:0] \add_5s_5s_5_2_1_U17.top_add_5s_5s_5_2_1_Adder_12_U.bin_s0 ;
wire \add_5s_5s_5_2_1_U17.top_add_5s_5s_5_2_1_Adder_12_U.ce ;
wire \add_5s_5s_5_2_1_U17.top_add_5s_5s_5_2_1_Adder_12_U.clk ;
wire \add_5s_5s_5_2_1_U17.top_add_5s_5s_5_2_1_Adder_12_U.facout_s1 ;
wire \add_5s_5s_5_2_1_U17.top_add_5s_5s_5_2_1_Adder_12_U.facout_s2 ;
wire [1:0] \add_5s_5s_5_2_1_U17.top_add_5s_5s_5_2_1_Adder_12_U.fas_s1 ;
wire [2:0] \add_5s_5s_5_2_1_U17.top_add_5s_5s_5_2_1_Adder_12_U.fas_s2 ;
wire \add_5s_5s_5_2_1_U17.top_add_5s_5s_5_2_1_Adder_12_U.reset ;
wire [4:0] \add_5s_5s_5_2_1_U17.top_add_5s_5s_5_2_1_Adder_12_U.s ;
wire [1:0] \add_5s_5s_5_2_1_U17.top_add_5s_5s_5_2_1_Adder_12_U.u1.a ;
wire [1:0] \add_5s_5s_5_2_1_U17.top_add_5s_5s_5_2_1_Adder_12_U.u1.b ;
wire \add_5s_5s_5_2_1_U17.top_add_5s_5s_5_2_1_Adder_12_U.u1.cin ;
wire \add_5s_5s_5_2_1_U17.top_add_5s_5s_5_2_1_Adder_12_U.u1.cout ;
wire [1:0] \add_5s_5s_5_2_1_U17.top_add_5s_5s_5_2_1_Adder_12_U.u1.s ;
wire [2:0] \add_5s_5s_5_2_1_U17.top_add_5s_5s_5_2_1_Adder_12_U.u2.a ;
wire [2:0] \add_5s_5s_5_2_1_U17.top_add_5s_5s_5_2_1_Adder_12_U.u2.b ;
wire \add_5s_5s_5_2_1_U17.top_add_5s_5s_5_2_1_Adder_12_U.u2.cin ;
wire \add_5s_5s_5_2_1_U17.top_add_5s_5s_5_2_1_Adder_12_U.u2.cout ;
wire [2:0] \add_5s_5s_5_2_1_U17.top_add_5s_5s_5_2_1_Adder_12_U.u2.s ;
wire \add_6ns_6s_6_2_1_U20.ce ;
wire \add_6ns_6s_6_2_1_U20.clk ;
wire [5:0] \add_6ns_6s_6_2_1_U20.din0 ;
wire [5:0] \add_6ns_6s_6_2_1_U20.din1 ;
wire [5:0] \add_6ns_6s_6_2_1_U20.dout ;
wire \add_6ns_6s_6_2_1_U20.reset ;
wire [5:0] \add_6ns_6s_6_2_1_U20.top_add_6ns_6s_6_2_1_Adder_15_U.a ;
wire [5:0] \add_6ns_6s_6_2_1_U20.top_add_6ns_6s_6_2_1_Adder_15_U.ain_s0 ;
wire [5:0] \add_6ns_6s_6_2_1_U20.top_add_6ns_6s_6_2_1_Adder_15_U.b ;
wire [5:0] \add_6ns_6s_6_2_1_U20.top_add_6ns_6s_6_2_1_Adder_15_U.bin_s0 ;
wire \add_6ns_6s_6_2_1_U20.top_add_6ns_6s_6_2_1_Adder_15_U.ce ;
wire \add_6ns_6s_6_2_1_U20.top_add_6ns_6s_6_2_1_Adder_15_U.clk ;
wire \add_6ns_6s_6_2_1_U20.top_add_6ns_6s_6_2_1_Adder_15_U.facout_s1 ;
wire \add_6ns_6s_6_2_1_U20.top_add_6ns_6s_6_2_1_Adder_15_U.facout_s2 ;
wire [2:0] \add_6ns_6s_6_2_1_U20.top_add_6ns_6s_6_2_1_Adder_15_U.fas_s1 ;
wire [2:0] \add_6ns_6s_6_2_1_U20.top_add_6ns_6s_6_2_1_Adder_15_U.fas_s2 ;
wire \add_6ns_6s_6_2_1_U20.top_add_6ns_6s_6_2_1_Adder_15_U.reset ;
wire [5:0] \add_6ns_6s_6_2_1_U20.top_add_6ns_6s_6_2_1_Adder_15_U.s ;
wire [2:0] \add_6ns_6s_6_2_1_U20.top_add_6ns_6s_6_2_1_Adder_15_U.u1.a ;
wire [2:0] \add_6ns_6s_6_2_1_U20.top_add_6ns_6s_6_2_1_Adder_15_U.u1.b ;
wire \add_6ns_6s_6_2_1_U20.top_add_6ns_6s_6_2_1_Adder_15_U.u1.cin ;
wire \add_6ns_6s_6_2_1_U20.top_add_6ns_6s_6_2_1_Adder_15_U.u1.cout ;
wire [2:0] \add_6ns_6s_6_2_1_U20.top_add_6ns_6s_6_2_1_Adder_15_U.u1.s ;
wire [2:0] \add_6ns_6s_6_2_1_U20.top_add_6ns_6s_6_2_1_Adder_15_U.u2.a ;
wire [2:0] \add_6ns_6s_6_2_1_U20.top_add_6ns_6s_6_2_1_Adder_15_U.u2.b ;
wire \add_6ns_6s_6_2_1_U20.top_add_6ns_6s_6_2_1_Adder_15_U.u2.cin ;
wire \add_6ns_6s_6_2_1_U20.top_add_6ns_6s_6_2_1_Adder_15_U.u2.cout ;
wire [2:0] \add_6ns_6s_6_2_1_U20.top_add_6ns_6s_6_2_1_Adder_15_U.u2.s ;
wire \add_6s_6s_6_2_1_U19.ce ;
wire \add_6s_6s_6_2_1_U19.clk ;
wire [5:0] \add_6s_6s_6_2_1_U19.din0 ;
wire [5:0] \add_6s_6s_6_2_1_U19.din1 ;
wire [5:0] \add_6s_6s_6_2_1_U19.dout ;
wire \add_6s_6s_6_2_1_U19.reset ;
wire [5:0] \add_6s_6s_6_2_1_U19.top_add_6s_6s_6_2_1_Adder_14_U.a ;
wire [5:0] \add_6s_6s_6_2_1_U19.top_add_6s_6s_6_2_1_Adder_14_U.ain_s0 ;
wire [5:0] \add_6s_6s_6_2_1_U19.top_add_6s_6s_6_2_1_Adder_14_U.b ;
wire [5:0] \add_6s_6s_6_2_1_U19.top_add_6s_6s_6_2_1_Adder_14_U.bin_s0 ;
wire \add_6s_6s_6_2_1_U19.top_add_6s_6s_6_2_1_Adder_14_U.ce ;
wire \add_6s_6s_6_2_1_U19.top_add_6s_6s_6_2_1_Adder_14_U.clk ;
wire \add_6s_6s_6_2_1_U19.top_add_6s_6s_6_2_1_Adder_14_U.facout_s1 ;
wire \add_6s_6s_6_2_1_U19.top_add_6s_6s_6_2_1_Adder_14_U.facout_s2 ;
wire [2:0] \add_6s_6s_6_2_1_U19.top_add_6s_6s_6_2_1_Adder_14_U.fas_s1 ;
wire [2:0] \add_6s_6s_6_2_1_U19.top_add_6s_6s_6_2_1_Adder_14_U.fas_s2 ;
wire \add_6s_6s_6_2_1_U19.top_add_6s_6s_6_2_1_Adder_14_U.reset ;
wire [5:0] \add_6s_6s_6_2_1_U19.top_add_6s_6s_6_2_1_Adder_14_U.s ;
wire [2:0] \add_6s_6s_6_2_1_U19.top_add_6s_6s_6_2_1_Adder_14_U.u1.a ;
wire [2:0] \add_6s_6s_6_2_1_U19.top_add_6s_6s_6_2_1_Adder_14_U.u1.b ;
wire \add_6s_6s_6_2_1_U19.top_add_6s_6s_6_2_1_Adder_14_U.u1.cin ;
wire \add_6s_6s_6_2_1_U19.top_add_6s_6s_6_2_1_Adder_14_U.u1.cout ;
wire [2:0] \add_6s_6s_6_2_1_U19.top_add_6s_6s_6_2_1_Adder_14_U.u1.s ;
wire [2:0] \add_6s_6s_6_2_1_U19.top_add_6s_6s_6_2_1_Adder_14_U.u2.a ;
wire [2:0] \add_6s_6s_6_2_1_U19.top_add_6s_6s_6_2_1_Adder_14_U.u2.b ;
wire \add_6s_6s_6_2_1_U19.top_add_6s_6s_6_2_1_Adder_14_U.u2.cin ;
wire \add_6s_6s_6_2_1_U19.top_add_6s_6s_6_2_1_Adder_14_U.u2.cout ;
wire [2:0] \add_6s_6s_6_2_1_U19.top_add_6s_6s_6_2_1_Adder_14_U.u2.s ;
wire \add_8ns_8ns_8_2_1_U7.ce ;
wire \add_8ns_8ns_8_2_1_U7.clk ;
wire [7:0] \add_8ns_8ns_8_2_1_U7.din0 ;
wire [7:0] \add_8ns_8ns_8_2_1_U7.din1 ;
wire [7:0] \add_8ns_8ns_8_2_1_U7.dout ;
wire \add_8ns_8ns_8_2_1_U7.reset ;
wire [7:0] \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_4_U.a ;
wire [7:0] \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_4_U.ain_s0 ;
wire [7:0] \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_4_U.b ;
wire [7:0] \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_4_U.bin_s0 ;
wire \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_4_U.ce ;
wire \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_4_U.clk ;
wire \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_4_U.facout_s1 ;
wire \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_4_U.facout_s2 ;
wire [3:0] \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_4_U.fas_s1 ;
wire [3:0] \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_4_U.fas_s2 ;
wire \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_4_U.reset ;
wire [7:0] \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_4_U.s ;
wire [3:0] \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_4_U.u1.a ;
wire [3:0] \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_4_U.u1.b ;
wire \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_4_U.u1.cin ;
wire \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_4_U.u1.cout ;
wire [3:0] \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_4_U.u1.s ;
wire [3:0] \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_4_U.u2.a ;
wire [3:0] \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_4_U.u2.b ;
wire \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_4_U.u2.cin ;
wire \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_4_U.u2.cout ;
wire [3:0] \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_4_U.u2.s ;
wire \add_9s_9ns_9_2_1_U3.ce ;
wire \add_9s_9ns_9_2_1_U3.clk ;
wire [8:0] \add_9s_9ns_9_2_1_U3.din0 ;
wire [8:0] \add_9s_9ns_9_2_1_U3.din1 ;
wire [8:0] \add_9s_9ns_9_2_1_U3.dout ;
wire \add_9s_9ns_9_2_1_U3.reset ;
wire [8:0] \add_9s_9ns_9_2_1_U3.top_add_9s_9ns_9_2_1_Adder_0_U.a ;
wire [8:0] \add_9s_9ns_9_2_1_U3.top_add_9s_9ns_9_2_1_Adder_0_U.ain_s0 ;
wire [8:0] \add_9s_9ns_9_2_1_U3.top_add_9s_9ns_9_2_1_Adder_0_U.b ;
wire [8:0] \add_9s_9ns_9_2_1_U3.top_add_9s_9ns_9_2_1_Adder_0_U.bin_s0 ;
wire \add_9s_9ns_9_2_1_U3.top_add_9s_9ns_9_2_1_Adder_0_U.ce ;
wire \add_9s_9ns_9_2_1_U3.top_add_9s_9ns_9_2_1_Adder_0_U.clk ;
wire \add_9s_9ns_9_2_1_U3.top_add_9s_9ns_9_2_1_Adder_0_U.facout_s1 ;
wire \add_9s_9ns_9_2_1_U3.top_add_9s_9ns_9_2_1_Adder_0_U.facout_s2 ;
wire [3:0] \add_9s_9ns_9_2_1_U3.top_add_9s_9ns_9_2_1_Adder_0_U.fas_s1 ;
wire [4:0] \add_9s_9ns_9_2_1_U3.top_add_9s_9ns_9_2_1_Adder_0_U.fas_s2 ;
wire \add_9s_9ns_9_2_1_U3.top_add_9s_9ns_9_2_1_Adder_0_U.reset ;
wire [8:0] \add_9s_9ns_9_2_1_U3.top_add_9s_9ns_9_2_1_Adder_0_U.s ;
wire [3:0] \add_9s_9ns_9_2_1_U3.top_add_9s_9ns_9_2_1_Adder_0_U.u1.a ;
wire [3:0] \add_9s_9ns_9_2_1_U3.top_add_9s_9ns_9_2_1_Adder_0_U.u1.b ;
wire \add_9s_9ns_9_2_1_U3.top_add_9s_9ns_9_2_1_Adder_0_U.u1.cin ;
wire \add_9s_9ns_9_2_1_U3.top_add_9s_9ns_9_2_1_Adder_0_U.u1.cout ;
wire [3:0] \add_9s_9ns_9_2_1_U3.top_add_9s_9ns_9_2_1_Adder_0_U.u1.s ;
wire [4:0] \add_9s_9ns_9_2_1_U3.top_add_9s_9ns_9_2_1_Adder_0_U.u2.a ;
wire [4:0] \add_9s_9ns_9_2_1_U3.top_add_9s_9ns_9_2_1_Adder_0_U.u2.b ;
wire \add_9s_9ns_9_2_1_U3.top_add_9s_9ns_9_2_1_Adder_0_U.u2.cin ;
wire \add_9s_9ns_9_2_1_U3.top_add_9s_9ns_9_2_1_Adder_0_U.u2.cout ;
wire [4:0] \add_9s_9ns_9_2_1_U3.top_add_9s_9ns_9_2_1_Adder_0_U.u2.s ;
wire \add_9s_9s_9_2_1_U23.ce ;
wire \add_9s_9s_9_2_1_U23.clk ;
wire [8:0] \add_9s_9s_9_2_1_U23.din0 ;
wire [8:0] \add_9s_9s_9_2_1_U23.din1 ;
wire [8:0] \add_9s_9s_9_2_1_U23.dout ;
wire \add_9s_9s_9_2_1_U23.reset ;
wire [8:0] \add_9s_9s_9_2_1_U23.top_add_9s_9s_9_2_1_Adder_18_U.a ;
wire [8:0] \add_9s_9s_9_2_1_U23.top_add_9s_9s_9_2_1_Adder_18_U.ain_s0 ;
wire [8:0] \add_9s_9s_9_2_1_U23.top_add_9s_9s_9_2_1_Adder_18_U.b ;
wire [8:0] \add_9s_9s_9_2_1_U23.top_add_9s_9s_9_2_1_Adder_18_U.bin_s0 ;
wire \add_9s_9s_9_2_1_U23.top_add_9s_9s_9_2_1_Adder_18_U.ce ;
wire \add_9s_9s_9_2_1_U23.top_add_9s_9s_9_2_1_Adder_18_U.clk ;
wire \add_9s_9s_9_2_1_U23.top_add_9s_9s_9_2_1_Adder_18_U.facout_s1 ;
wire \add_9s_9s_9_2_1_U23.top_add_9s_9s_9_2_1_Adder_18_U.facout_s2 ;
wire [3:0] \add_9s_9s_9_2_1_U23.top_add_9s_9s_9_2_1_Adder_18_U.fas_s1 ;
wire [4:0] \add_9s_9s_9_2_1_U23.top_add_9s_9s_9_2_1_Adder_18_U.fas_s2 ;
wire \add_9s_9s_9_2_1_U23.top_add_9s_9s_9_2_1_Adder_18_U.reset ;
wire [8:0] \add_9s_9s_9_2_1_U23.top_add_9s_9s_9_2_1_Adder_18_U.s ;
wire [3:0] \add_9s_9s_9_2_1_U23.top_add_9s_9s_9_2_1_Adder_18_U.u1.a ;
wire [3:0] \add_9s_9s_9_2_1_U23.top_add_9s_9s_9_2_1_Adder_18_U.u1.b ;
wire \add_9s_9s_9_2_1_U23.top_add_9s_9s_9_2_1_Adder_18_U.u1.cin ;
wire \add_9s_9s_9_2_1_U23.top_add_9s_9s_9_2_1_Adder_18_U.u1.cout ;
wire [3:0] \add_9s_9s_9_2_1_U23.top_add_9s_9s_9_2_1_Adder_18_U.u1.s ;
wire [4:0] \add_9s_9s_9_2_1_U23.top_add_9s_9s_9_2_1_Adder_18_U.u2.a ;
wire [4:0] \add_9s_9s_9_2_1_U23.top_add_9s_9s_9_2_1_Adder_18_U.u2.b ;
wire \add_9s_9s_9_2_1_U23.top_add_9s_9s_9_2_1_Adder_18_U.u2.cin ;
wire \add_9s_9s_9_2_1_U23.top_add_9s_9s_9_2_1_Adder_18_U.u2.cout ;
wire [4:0] \add_9s_9s_9_2_1_U23.top_add_9s_9s_9_2_1_Adder_18_U.u2.s ;
wire and_ln340_fu_1003_p2;
wire and_ln408_fu_1227_p2;
wire and_ln412_fu_687_p2;
wire and_ln414_fu_481_p2;
wire and_ln780_1_fu_1211_p2;
wire and_ln780_2_fu_1463_p2;
wire and_ln780_fu_722_p2;
wire and_ln781_1_fu_1329_p2;
wire and_ln781_2_fu_1530_p2;
wire and_ln781_fu_766_p2;
wire and_ln785_1_fu_811_p2;
wire and_ln785_2_fu_994_p2;
wire and_ln785_4_fu_1373_p2;
wire and_ln785_5_fu_1382_p2;
wire and_ln785_fu_802_p2;
wire and_ln786_1_fu_1222_p2;
wire and_ln786_3_fu_1497_p2;
wire and_ln786_fu_738_p2;
wire [7:0] and_ln_fu_599_p3;
wire ap_CS_fsm_state1;
wire ap_CS_fsm_state10;
wire ap_CS_fsm_state11;
wire ap_CS_fsm_state12;
wire ap_CS_fsm_state13;
wire ap_CS_fsm_state14;
wire ap_CS_fsm_state15;
wire ap_CS_fsm_state16;
wire ap_CS_fsm_state17;
wire ap_CS_fsm_state18;
wire ap_CS_fsm_state19;
wire ap_CS_fsm_state2;
wire ap_CS_fsm_state20;
wire ap_CS_fsm_state21;
wire ap_CS_fsm_state22;
wire ap_CS_fsm_state23;
wire ap_CS_fsm_state24;
wire ap_CS_fsm_state25;
wire ap_CS_fsm_state26;
wire ap_CS_fsm_state27;
wire ap_CS_fsm_state28;
wire ap_CS_fsm_state29;
wire ap_CS_fsm_state3;
wire ap_CS_fsm_state30;
wire ap_CS_fsm_state31;
wire ap_CS_fsm_state32;
wire ap_CS_fsm_state4;
wire ap_CS_fsm_state5;
wire ap_CS_fsm_state6;
wire ap_CS_fsm_state7;
wire ap_CS_fsm_state8;
wire ap_CS_fsm_state9;
wire [31:0] ap_NS_fsm;
wire ap_clk;
wire ap_done;
wire ap_idle;
wire ap_ready;
wire ap_rst;
wire ap_start;
wire carry_1_fu_664_p2;
wire carry_3_fu_1149_p2;
wire carry_5_fu_1405_p2;
wire deleted_ones_1_fu_1216_p3;
wire deleted_ones_2_fu_1469_p3;
wire deleted_ones_fu_727_p3;
wire deleted_zeros_1_fu_1193_p3;
wire deleted_zeros_2_fu_1445_p3;
wire deleted_zeros_fu_712_p3;
wire [31:0] empty_fu_381_p0;
wire [24:0] empty_fu_381_p1;
wire [2:0] grp_fu_1024_p0;
wire [2:0] grp_fu_1024_p2;
wire [3:0] grp_fu_1178_p2;
wire [3:0] grp_fu_1188_p2;
wire [3:0] grp_fu_1241_p0;
wire [3:0] grp_fu_1241_p1;
wire [3:0] grp_fu_1241_p2;
wire [3:0] grp_fu_1276_p1;
wire [3:0] grp_fu_1276_p2;
wire [3:0] grp_fu_1367_p0;
wire [3:0] grp_fu_1367_p2;
wire [4:0] grp_fu_1428_p0;
wire [4:0] grp_fu_1428_p1;
wire [4:0] grp_fu_1428_p2;
wire [4:0] grp_fu_1558_p1;
wire [4:0] grp_fu_1558_p2;
wire [5:0] grp_fu_1582_p0;
wire [5:0] grp_fu_1582_p1;
wire [5:0] grp_fu_1582_p2;
wire [5:0] grp_fu_1591_p1;
wire [5:0] grp_fu_1591_p2;
wire [38:0] grp_fu_1610_p0;
wire [38:0] grp_fu_1610_p1;
wire [38:0] grp_fu_1610_p2;
wire [31:0] grp_fu_1626_p2;
wire [8:0] grp_fu_1638_p0;
wire [8:0] grp_fu_1638_p1;
wire [8:0] grp_fu_1638_p2;
wire [31:0] grp_fu_1666_p0;
wire [31:0] grp_fu_1666_p2;
wire [3:0] grp_fu_279_p2;
wire [3:0] grp_fu_307_p0;
wire [3:0] grp_fu_307_p1;
wire [7:0] grp_fu_307_p2;
wire [8:0] grp_fu_347_p0;
wire [8:0] grp_fu_347_p1;
wire [8:0] grp_fu_347_p2;
wire [1:0] grp_fu_518_p1;
wire [1:0] grp_fu_518_p2;
wire [25:0] grp_fu_589_p0;
wire [25:0] grp_fu_589_p2;
wire [24:0] grp_fu_594_p0;
wire [24:0] grp_fu_594_p2;
wire [7:0] grp_fu_746_p1;
wire [7:0] grp_fu_746_p2;
wire [32:0] grp_fu_838_p0;
wire [32:0] grp_fu_838_p1;
wire [32:0] grp_fu_838_p2;
wire [10:0] grp_fu_894_p0;
wire [10:0] grp_fu_894_p1;
wire [10:0] grp_fu_894_p2;
wire [8:0] grp_fu_914_p0;
wire [8:0] grp_fu_914_p1;
wire [8:0] grp_fu_914_p2;
wire icmp_ln414_fu_415_p2;
wire icmp_ln768_fu_371_p2;
wire icmp_ln785_fu_543_p2;
wire icmp_ln786_1_fu_549_p2;
wire icmp_ln786_2_fu_376_p2;
wire icmp_ln786_fu_616_p2;
wire icmp_ln790_fu_561_p2;
wire icmp_ln851_1_fu_1183_p2;
wire icmp_ln851_2_fu_1525_p2;
wire icmp_ln851_fu_1173_p2;
wire [26:0] lhs_V_1_fu_824_p3;
wire [8:0] lhs_V_3_fu_879_p3;
wire \mul_4s_4s_4_7_1_U1.ce ;
wire \mul_4s_4s_4_7_1_U1.clk ;
wire [3:0] \mul_4s_4s_4_7_1_U1.din0 ;
wire [3:0] \mul_4s_4s_4_7_1_U1.din1 ;
wire [3:0] \mul_4s_4s_4_7_1_U1.dout ;
wire \mul_4s_4s_4_7_1_U1.reset ;
wire [3:0] \mul_4s_4s_4_7_1_U1.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.a ;
wire [3:0] \mul_4s_4s_4_7_1_U1.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.b ;
wire \mul_4s_4s_4_7_1_U1.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.ce ;
wire \mul_4s_4s_4_7_1_U1.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.clk ;
wire [3:0] \mul_4s_4s_4_7_1_U1.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.p ;
wire [3:0] \mul_4s_4s_4_7_1_U1.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.tmp_product ;
wire \mul_4s_4s_8_7_1_U2.ce ;
wire \mul_4s_4s_8_7_1_U2.clk ;
wire [3:0] \mul_4s_4s_8_7_1_U2.din0 ;
wire [3:0] \mul_4s_4s_8_7_1_U2.din1 ;
wire [7:0] \mul_4s_4s_8_7_1_U2.dout ;
wire \mul_4s_4s_8_7_1_U2.reset ;
wire [3:0] \mul_4s_4s_8_7_1_U2.top_mul_4s_4s_8_7_1_Mul_DSP_1_U.a ;
wire [3:0] \mul_4s_4s_8_7_1_U2.top_mul_4s_4s_8_7_1_Mul_DSP_1_U.b ;
wire \mul_4s_4s_8_7_1_U2.top_mul_4s_4s_8_7_1_Mul_DSP_1_U.ce ;
wire \mul_4s_4s_8_7_1_U2.top_mul_4s_4s_8_7_1_Mul_DSP_1_U.clk ;
wire [7:0] \mul_4s_4s_8_7_1_U2.top_mul_4s_4s_8_7_1_Mul_DSP_1_U.p ;
wire [7:0] \mul_4s_4s_8_7_1_U2.top_mul_4s_4s_8_7_1_Mul_DSP_1_U.tmp_product ;
wire neg_src_7_fu_1339_p2;
wire neg_src_fu_776_p2;
wire op_0;
wire [31:0] op_1;
wire [1:0] op_12_V_fu_1143_p3;
wire [1:0] op_13;
wire [3:0] op_15_V_fu_1570_p3;
wire [3:0] op_16_V_fu_335_p2;
wire [7:0] op_17_V_fu_1387_p3;
wire [7:0] op_19;
wire [3:0] op_2;
wire [31:0] op_28;
wire op_28_ap_vld;
wire [7:0] op_4_V_fu_301_p2;
wire [1:0] op_5;
wire [31:0] op_6;
wire [3:0] op_7;
wire [7:0] op_8_V_fu_705_p3;
wire [1:0] op_9;
wire or_ln340_1_fu_983_p2;
wire or_ln340_2_fu_1008_p2;
wire or_ln340_3_fu_1268_p2;
wire or_ln340_4_fu_1344_p2;
wire or_ln340_fu_796_p2;
wire or_ln384_1_fu_874_p2;
wire or_ln384_2_fu_1550_p2;
wire or_ln384_fu_659_p2;
wire or_ln412_fu_682_p2;
wire or_ln731_fu_317_p2;
wire [3:0] or_ln760_fu_329_p1;
wire [3:0] or_ln760_fu_329_p2;
wire or_ln785_1_fu_1252_p2;
wire or_ln785_2_fu_751_p2;
wire or_ln785_3_fu_1481_p2;
wire or_ln785_4_fu_806_p2;
wire or_ln785_5_fu_1377_p2;
wire or_ln785_fu_786_p2;
wire or_ln786_1_fu_1534_p2;
wire or_ln786_fu_864_p2;
wire or_ln788_1_fu_649_p2;
wire or_ln788_fu_645_p2;
wire [7:0] or_ln_fu_535_p4;
wire overflow_1_fu_791_p2;
wire overflow_2_fu_1262_p2;
wire overflow_3_fu_760_p2;
wire overflow_4_fu_1491_p2;
wire overflow_fu_611_p2;
wire [1:0] p_Result_12_fu_974_p4;
wire p_Result_17_fu_668_p3;
wire [31:0] p_Result_1_fu_429_p1;
wire [6:0] p_Result_1_fu_429_p4;
wire p_Result_25_fu_1502_p3;
wire p_Result_26_fu_1291_p3;
wire p_Result_27_fu_1310_p3;
wire p_Result_28_fu_1644_p3;
wire [31:0] p_Result_30_fu_385_p1;
wire [31:0] p_Result_31_fu_403_p1;
wire [31:0] p_Result_33_fu_421_p1;
wire [31:0] p_Result_35_fu_675_p1;
wire p_Result_35_fu_675_p3;
wire p_Result_39_fu_323_p2;
wire [31:0] p_Result_3_fu_445_p1;
wire [7:0] p_Result_3_fu_445_p4;
wire p_Result_42_fu_1393_p3;
wire [6:0] p_Result_s_20_fu_554_p3;
wire [1:0] p_Val2_10_fu_852_p3;
wire [7:0] p_Val2_1_fu_693_p2;
wire [31:0] p_Val2_2_fu_393_p1;
wire p_Val2_4_fu_969_p2;
wire r_1_fu_1168_p2;
wire r_fu_475_p2;
wire [3:0] ret_V_19_fu_1518_p3;
wire [3:0] ret_V_21_fu_1303_p3;
wire [31:0] ret_V_22_fu_1119_p1;
wire [31:0] ret_V_22_fu_1119_p2;
wire [3:0] ret_V_23_fu_1322_p3;
wire [31:0] ret_V_26_fu_1656_p3;
wire [23:0] rhs_3_fu_935_p3;
wire [6:0] rhs_fu_903_p3;
wire sel_tmp11_fu_1014_p2;
wire [7:0] select_ln340_1_fu_1349_p3;
wire [1:0] select_ln340_fu_987_p3;
wire [3:0] select_ln384_2_fu_1563_p3;
wire [1:0] select_ln384_4_fu_920_p3;
wire [1:0] select_ln384_5_fu_927_p3;
wire [7:0] select_ln384_fu_698_p3;
wire [2:0] select_ln703_fu_816_p3;
wire [1:0] select_ln785_fu_1138_p3;
wire [3:0] select_ln850_1_fu_1298_p3;
wire [3:0] select_ln850_2_fu_1317_p3;
wire [31:0] select_ln850_3_fu_1651_p3;
wire [3:0] select_ln850_fu_1512_p3;
wire [31:0] sext_ln1195_fu_1116_p1;
wire [3:0] sext_ln69_fu_289_p0;
wire [7:0] sext_ln69_fu_289_p1;
wire [31:0] sext_ln703_1_fu_835_p0;
wire [3:0] sext_ln850_fu_1364_p1;
wire \sub_11ns_11s_11_2_1_U9.ce ;
wire \sub_11ns_11s_11_2_1_U9.clk ;
wire [10:0] \sub_11ns_11s_11_2_1_U9.din0 ;
wire [10:0] \sub_11ns_11s_11_2_1_U9.din1 ;
wire [10:0] \sub_11ns_11s_11_2_1_U9.dout ;
wire \sub_11ns_11s_11_2_1_U9.reset ;
wire [10:0] \sub_11ns_11s_11_2_1_U9.top_sub_11ns_11s_11_2_1_Adder_6_U.a ;
wire [10:0] \sub_11ns_11s_11_2_1_U9.top_sub_11ns_11s_11_2_1_Adder_6_U.ain_s0 ;
wire [10:0] \sub_11ns_11s_11_2_1_U9.top_sub_11ns_11s_11_2_1_Adder_6_U.b ;
wire [10:0] \sub_11ns_11s_11_2_1_U9.top_sub_11ns_11s_11_2_1_Adder_6_U.bin_s0 ;
wire \sub_11ns_11s_11_2_1_U9.top_sub_11ns_11s_11_2_1_Adder_6_U.ce ;
wire \sub_11ns_11s_11_2_1_U9.top_sub_11ns_11s_11_2_1_Adder_6_U.clk ;
wire \sub_11ns_11s_11_2_1_U9.top_sub_11ns_11s_11_2_1_Adder_6_U.facout_s1 ;
wire \sub_11ns_11s_11_2_1_U9.top_sub_11ns_11s_11_2_1_Adder_6_U.facout_s2 ;
wire [4:0] \sub_11ns_11s_11_2_1_U9.top_sub_11ns_11s_11_2_1_Adder_6_U.fas_s1 ;
wire [5:0] \sub_11ns_11s_11_2_1_U9.top_sub_11ns_11s_11_2_1_Adder_6_U.fas_s2 ;
wire \sub_11ns_11s_11_2_1_U9.top_sub_11ns_11s_11_2_1_Adder_6_U.reset ;
wire [10:0] \sub_11ns_11s_11_2_1_U9.top_sub_11ns_11s_11_2_1_Adder_6_U.s ;
wire [4:0] \sub_11ns_11s_11_2_1_U9.top_sub_11ns_11s_11_2_1_Adder_6_U.u1.a ;
wire [4:0] \sub_11ns_11s_11_2_1_U9.top_sub_11ns_11s_11_2_1_Adder_6_U.u1.b ;
wire \sub_11ns_11s_11_2_1_U9.top_sub_11ns_11s_11_2_1_Adder_6_U.u1.cin ;
wire \sub_11ns_11s_11_2_1_U9.top_sub_11ns_11s_11_2_1_Adder_6_U.u1.cout ;
wire [4:0] \sub_11ns_11s_11_2_1_U9.top_sub_11ns_11s_11_2_1_Adder_6_U.u1.s ;
wire [5:0] \sub_11ns_11s_11_2_1_U9.top_sub_11ns_11s_11_2_1_Adder_6_U.u2.a ;
wire [5:0] \sub_11ns_11s_11_2_1_U9.top_sub_11ns_11s_11_2_1_Adder_6_U.u2.b ;
wire \sub_11ns_11s_11_2_1_U9.top_sub_11ns_11s_11_2_1_Adder_6_U.u2.cin ;
wire \sub_11ns_11s_11_2_1_U9.top_sub_11ns_11s_11_2_1_Adder_6_U.u2.cout ;
wire [5:0] \sub_11ns_11s_11_2_1_U9.top_sub_11ns_11s_11_2_1_Adder_6_U.u2.s ;
wire \sub_9s_9s_9_2_1_U10.ce ;
wire \sub_9s_9s_9_2_1_U10.clk ;
wire [8:0] \sub_9s_9s_9_2_1_U10.din0 ;
wire [8:0] \sub_9s_9s_9_2_1_U10.din1 ;
wire [8:0] \sub_9s_9s_9_2_1_U10.dout ;
wire \sub_9s_9s_9_2_1_U10.reset ;
wire [8:0] \sub_9s_9s_9_2_1_U10.top_sub_9s_9s_9_2_1_Adder_7_U.a ;
wire [8:0] \sub_9s_9s_9_2_1_U10.top_sub_9s_9s_9_2_1_Adder_7_U.ain_s0 ;
wire [8:0] \sub_9s_9s_9_2_1_U10.top_sub_9s_9s_9_2_1_Adder_7_U.b ;
wire [8:0] \sub_9s_9s_9_2_1_U10.top_sub_9s_9s_9_2_1_Adder_7_U.bin_s0 ;
wire \sub_9s_9s_9_2_1_U10.top_sub_9s_9s_9_2_1_Adder_7_U.ce ;
wire \sub_9s_9s_9_2_1_U10.top_sub_9s_9s_9_2_1_Adder_7_U.clk ;
wire \sub_9s_9s_9_2_1_U10.top_sub_9s_9s_9_2_1_Adder_7_U.facout_s1 ;
wire \sub_9s_9s_9_2_1_U10.top_sub_9s_9s_9_2_1_Adder_7_U.facout_s2 ;
wire [3:0] \sub_9s_9s_9_2_1_U10.top_sub_9s_9s_9_2_1_Adder_7_U.fas_s1 ;
wire [4:0] \sub_9s_9s_9_2_1_U10.top_sub_9s_9s_9_2_1_Adder_7_U.fas_s2 ;
wire \sub_9s_9s_9_2_1_U10.top_sub_9s_9s_9_2_1_Adder_7_U.reset ;
wire [8:0] \sub_9s_9s_9_2_1_U10.top_sub_9s_9s_9_2_1_Adder_7_U.s ;
wire [3:0] \sub_9s_9s_9_2_1_U10.top_sub_9s_9s_9_2_1_Adder_7_U.u1.a ;
wire [3:0] \sub_9s_9s_9_2_1_U10.top_sub_9s_9s_9_2_1_Adder_7_U.u1.b ;
wire \sub_9s_9s_9_2_1_U10.top_sub_9s_9s_9_2_1_Adder_7_U.u1.cin ;
wire \sub_9s_9s_9_2_1_U10.top_sub_9s_9s_9_2_1_Adder_7_U.u1.cout ;
wire [3:0] \sub_9s_9s_9_2_1_U10.top_sub_9s_9s_9_2_1_Adder_7_U.u1.s ;
wire [4:0] \sub_9s_9s_9_2_1_U10.top_sub_9s_9s_9_2_1_Adder_7_U.u2.a ;
wire [4:0] \sub_9s_9s_9_2_1_U10.top_sub_9s_9s_9_2_1_Adder_7_U.u2.b ;
wire \sub_9s_9s_9_2_1_U10.top_sub_9s_9s_9_2_1_Adder_7_U.u2.cin ;
wire \sub_9s_9s_9_2_1_U10.top_sub_9s_9s_9_2_1_Adder_7_U.u2.cout ;
wire [4:0] \sub_9s_9s_9_2_1_U10.top_sub_9s_9s_9_2_1_Adder_7_U.u2.s ;
wire tmp_14_fu_1198_p3;
wire tmp_21_fu_1450_p3;
wire [11:0] tmp_25_fu_1599_p3;
wire [31:0] tmp_6_fu_943_p1;
wire tmp_6_fu_943_p3;
wire tmp_7_fu_950_p3;
wire [31:0] trunc_ln1192_2_fu_467_p0;
wire [25:0] trunc_ln1192_2_fu_467_p1;
wire [2:0] trunc_ln1192_3_fu_531_p1;
wire [1:0] trunc_ln1192_fu_527_p1;
wire [31:0] trunc_ln414_fu_411_p0;
wire [21:0] trunc_ln414_fu_411_p1;
wire [7:0] trunc_ln69_1_fu_285_p1;
wire trunc_ln69_2_fu_293_p1;
wire [3:0] trunc_ln69_3_fu_297_p0;
wire trunc_ln69_3_fu_297_p1;
wire [3:0] trunc_ln69_fu_275_p1;
wire trunc_ln703_fu_523_p1;
wire [3:0] trunc_ln718_1_fu_1088_p1;
wire [31:0] trunc_ln718_fu_471_p0;
wire [15:0] trunc_ln718_fu_471_p1;
wire trunc_ln731_fu_313_p1;
wire [1:0] trunc_ln790_fu_511_p1;
wire [4:0] trunc_ln851_1_fu_1112_p1;
wire [22:0] trunc_ln851_2_fu_1134_p1;
wire [5:0] trunc_ln851_3_fu_1434_p1;
wire trunc_ln851_fu_1509_p1;
wire underflow_3_fu_869_p2;
wire underflow_4_fu_1545_p2;
wire underflow_fu_654_p2;
wire xor_ln365_1_fu_963_p2;
wire xor_ln365_fu_957_p2;
wire xor_ln416_1_fu_1037_p2;
wire xor_ln416_2_fu_1400_p2;
wire xor_ln416_fu_622_p2;
wire xor_ln780_1_fu_1205_p2;
wire xor_ln780_2_fu_1457_p2;
wire xor_ln780_fu_717_p2;
wire xor_ln781_1_fu_1333_p2;
wire xor_ln781_fu_770_p2;
wire xor_ln785_1_fu_781_p2;
wire xor_ln785_2_fu_733_p2;
wire xor_ln785_3_fu_1247_p2;
wire xor_ln785_4_fu_1257_p2;
wire xor_ln785_5_fu_755_p2;
wire xor_ln785_6_fu_1475_p2;
wire xor_ln785_7_fu_1486_p2;
wire xor_ln785_fu_606_p2;
wire xor_ln786_1_fu_998_p2;
wire xor_ln786_2_fu_1539_p2;
wire xor_ln786_fu_859_p2;


assign _0118_ = icmp_ln851_2_reg_2378 & ap_CS_fsm[28];
assign _0119_ = _0122_ & ap_CS_fsm[12];
assign _0120_ = _0123_ & ap_CS_fsm[0];
assign _0121_ = ap_start & ap_CS_fsm[0];
assign and_ln340_fu_1003_p2 = xor_ln786_1_fu_998_p2 & or_ln340_reg_2001;
assign and_ln408_fu_1227_p2 = r_1_reg_2207 & p_Result_41_reg_2122;
assign and_ln412_fu_687_p2 = op_6[16] & or_ln412_fu_682_p2;
assign and_ln414_fu_481_p2 = p_Result_30_reg_1755 & icmp_ln414_reg_1773;
assign and_ln780_1_fu_1211_p2 = xor_ln780_1_fu_1205_p2 & Range2_all_ones_1_reg_2190;
assign and_ln780_2_fu_1463_p2 = xor_ln780_2_fu_1457_p2 & ret_V_17_reg_2104[10];
assign and_ln780_fu_722_p2 = xor_ln780_fu_717_p2 & Range2_all_ones_reg_1784;
assign and_ln781_1_fu_1329_p2 = carry_3_reg_2183 & Range1_all_ones_1_reg_2195;
assign and_ln781_2_fu_1530_p2 = carry_5_reg_2318 & Range1_all_ones_2_reg_2325;
assign and_ln781_fu_766_p2 = carry_1_reg_1952 & Range1_all_ones_reg_1789;
assign and_ln785_1_fu_811_p2 = or_ln785_4_fu_806_p2 & and_ln786_reg_1982;
assign and_ln785_2_fu_994_p2 = xor_ln785_2_reg_1976 & and_ln786_reg_1982;
assign and_ln785_4_fu_1373_p2 = xor_ln416_1_reg_2087 & deleted_zeros_1_reg_2222;
assign and_ln785_5_fu_1382_p2 = or_ln785_5_fu_1377_p2 & and_ln786_1_reg_2228;
assign and_ln785_fu_802_p2 = xor_ln416_reg_1921 & deleted_zeros_reg_1970;
assign and_ln786_1_fu_1222_p2 = p_Result_37_reg_2033 & deleted_ones_1_fu_1216_p3;
assign and_ln786_3_fu_1497_p2 = p_Result_43_reg_2299 & deleted_ones_2_fu_1469_p3;
assign and_ln786_fu_738_p2 = p_Result_32_reg_1893 & deleted_ones_fu_727_p3;
assign carry_1_fu_664_p2 = xor_ln416_reg_1921 & p_Result_31_reg_1768;
assign carry_3_fu_1149_p2 = xor_ln416_1_reg_2087 & p_Result_36_reg_1942;
assign carry_5_fu_1405_p2 = xor_ln416_2_fu_1400_p2 & ret_V_17_reg_2104[8];
assign neg_src_7_fu_1339_p2 = xor_ln781_1_fu_1333_p2 & p_Result_34_reg_2080;
assign neg_src_fu_776_p2 = xor_ln781_fu_770_p2 & p_Result_30_reg_1755;
assign overflow_1_fu_791_p2 = xor_ln785_2_reg_1976 & or_ln785_fu_786_p2;
assign overflow_2_fu_1262_p2 = xor_ln785_4_fu_1257_p2 & or_ln785_1_fu_1252_p2;
assign overflow_3_fu_760_p2 = xor_ln785_5_fu_755_p2 & or_ln785_2_fu_751_p2;
assign overflow_4_fu_1491_p2 = xor_ln785_7_fu_1486_p2 & or_ln785_3_fu_1481_p2;
assign overflow_fu_611_p2 = xor_ln785_fu_606_p2 & icmp_ln785_reg_1869;
assign sel_tmp11_fu_1014_p2 = xor_ln365_1_fu_963_p2 & or_ln340_2_fu_1008_p2;
assign underflow_3_fu_869_p2 = p_Result_38_reg_1720 & or_ln786_fu_864_p2;
assign underflow_4_fu_1545_p2 = xor_ln786_2_fu_1539_p2 & p_Result_40_reg_2111;
assign underflow_fu_654_p2 = p_Result_29_reg_1826 & or_ln788_1_fu_649_p2;
assign xor_ln786_1_fu_998_p2 = ~ and_ln786_reg_1982;
assign xor_ln780_1_fu_1205_p2 = ~ add_ln1192_1_reg_1927[25];
assign xor_ln780_2_fu_1457_p2 = ~ ret_V_17_reg_2104[9];
assign xor_ln780_fu_717_p2 = ~ p_Result_33_reg_1778;
assign xor_ln416_2_fu_1400_p2 = ~ p_Result_43_reg_2299;
assign xor_ln781_1_fu_1333_p2 = ~ and_ln781_1_fu_1329_p2;
assign xor_ln781_fu_770_p2 = ~ and_ln781_fu_766_p2;
assign xor_ln785_3_fu_1247_p2 = ~ deleted_zeros_1_reg_2222;
assign xor_ln785_4_fu_1257_p2 = ~ p_Result_34_reg_2080;
assign xor_ln785_1_fu_781_p2 = ~ deleted_zeros_reg_1970;
assign xor_ln786_fu_859_p2 = ~ p_Result_39_reg_1698;
assign xor_ln786_2_fu_1539_p2 = ~ or_ln786_1_fu_1534_p2;
assign xor_ln785_6_fu_1475_p2 = ~ deleted_zeros_2_fu_1445_p3;
assign xor_ln785_5_fu_755_p2 = ~ p_Result_38_reg_1720;
assign xor_ln785_7_fu_1486_p2 = ~ p_Result_40_reg_2111;
assign xor_ln785_fu_606_p2 = ~ p_Result_29_reg_1826;
assign xor_ln365_1_fu_963_p2 = ~ xor_ln365_fu_957_p2;
assign xor_ln416_1_fu_1037_p2 = ~ p_Result_37_reg_2033;
assign xor_ln416_fu_622_p2 = ~ p_Result_32_reg_1893;
assign xor_ln785_2_fu_733_p2 = ~ p_Result_30_reg_1755;
assign op_16_V_fu_335_p2 = ~ or_ln760_fu_329_p2;
assign p_Val2_4_fu_969_p2 = ~ p_Val2_3_reg_1884[0];
assign _0122_ = ~ and_ln785_1_reg_2007;
assign _0123_ = ~ ap_start;
assign _0124_ = p_Result_6_reg_2098 == 8'hff;
assign _0125_ = p_Result_2_reg_2132 == 2'h3;
assign _0126_ = op_6[31:24] == 8'hff;
assign _0127_ = ! p_Result_6_reg_2098;
assign _0128_ = ! p_Result_2_reg_2132;
assign _0129_ = ! op_6[31:24];
assign _0130_ = p_Result_5_reg_2093 == 7'h7f;
assign _0131_ = op_6[31:25] == 7'h7f;
assign _0132_ = ! { tmp_reg_1832, 7'h00 };
assign _0133_ = ! { trunc_ln790_reg_1844, 5'h00 };
assign _0134_ = ! trunc_ln851_2_reg_2167;
assign _0135_ = ! trunc_ln851_1_reg_2150;
always @(posedge \add_25ns_25ns_25_2_1_U6.top_add_25ns_25ns_25_2_1_Adder_3_U.clk )
\add_25ns_25ns_25_2_1_U6.top_add_25ns_25ns_25_2_1_Adder_3_U.bin_s1  <= _0137_;
always @(posedge \add_25ns_25ns_25_2_1_U6.top_add_25ns_25ns_25_2_1_Adder_3_U.clk )
\add_25ns_25ns_25_2_1_U6.top_add_25ns_25ns_25_2_1_Adder_3_U.ain_s1  <= _0136_;
always @(posedge \add_25ns_25ns_25_2_1_U6.top_add_25ns_25ns_25_2_1_Adder_3_U.clk )
\add_25ns_25ns_25_2_1_U6.top_add_25ns_25ns_25_2_1_Adder_3_U.sum_s1  <= _0139_;
always @(posedge \add_25ns_25ns_25_2_1_U6.top_add_25ns_25ns_25_2_1_Adder_3_U.clk )
\add_25ns_25ns_25_2_1_U6.top_add_25ns_25ns_25_2_1_Adder_3_U.carry_s1  <= _0138_;
assign _0137_ = \add_25ns_25ns_25_2_1_U6.top_add_25ns_25ns_25_2_1_Adder_3_U.ce  ? \add_25ns_25ns_25_2_1_U6.top_add_25ns_25ns_25_2_1_Adder_3_U.b [24:12] : \add_25ns_25ns_25_2_1_U6.top_add_25ns_25ns_25_2_1_Adder_3_U.bin_s1 ;
assign _0136_ = \add_25ns_25ns_25_2_1_U6.top_add_25ns_25ns_25_2_1_Adder_3_U.ce  ? \add_25ns_25ns_25_2_1_U6.top_add_25ns_25ns_25_2_1_Adder_3_U.a [24:12] : \add_25ns_25ns_25_2_1_U6.top_add_25ns_25ns_25_2_1_Adder_3_U.ain_s1 ;
assign _0138_ = \add_25ns_25ns_25_2_1_U6.top_add_25ns_25ns_25_2_1_Adder_3_U.ce  ? \add_25ns_25ns_25_2_1_U6.top_add_25ns_25ns_25_2_1_Adder_3_U.facout_s1  : \add_25ns_25ns_25_2_1_U6.top_add_25ns_25ns_25_2_1_Adder_3_U.carry_s1 ;
assign _0139_ = \add_25ns_25ns_25_2_1_U6.top_add_25ns_25ns_25_2_1_Adder_3_U.ce  ? \add_25ns_25ns_25_2_1_U6.top_add_25ns_25ns_25_2_1_Adder_3_U.fas_s1  : \add_25ns_25ns_25_2_1_U6.top_add_25ns_25ns_25_2_1_Adder_3_U.sum_s1 ;
assign _0140_ = \add_25ns_25ns_25_2_1_U6.top_add_25ns_25ns_25_2_1_Adder_3_U.u1.a  + \add_25ns_25ns_25_2_1_U6.top_add_25ns_25ns_25_2_1_Adder_3_U.u1.b ;
assign { \add_25ns_25ns_25_2_1_U6.top_add_25ns_25ns_25_2_1_Adder_3_U.u1.cout , \add_25ns_25ns_25_2_1_U6.top_add_25ns_25ns_25_2_1_Adder_3_U.u1.s  } = _0140_ + \add_25ns_25ns_25_2_1_U6.top_add_25ns_25ns_25_2_1_Adder_3_U.u1.cin ;
assign _0141_ = \add_25ns_25ns_25_2_1_U6.top_add_25ns_25ns_25_2_1_Adder_3_U.u2.a  + \add_25ns_25ns_25_2_1_U6.top_add_25ns_25ns_25_2_1_Adder_3_U.u2.b ;
assign { \add_25ns_25ns_25_2_1_U6.top_add_25ns_25ns_25_2_1_Adder_3_U.u2.cout , \add_25ns_25ns_25_2_1_U6.top_add_25ns_25ns_25_2_1_Adder_3_U.u2.s  } = _0141_ + \add_25ns_25ns_25_2_1_U6.top_add_25ns_25ns_25_2_1_Adder_3_U.u2.cin ;
always @(posedge \add_26ns_26ns_26_2_1_U5.top_add_26ns_26ns_26_2_1_Adder_2_U.clk )
\add_26ns_26ns_26_2_1_U5.top_add_26ns_26ns_26_2_1_Adder_2_U.bin_s1  <= _0143_;
always @(posedge \add_26ns_26ns_26_2_1_U5.top_add_26ns_26ns_26_2_1_Adder_2_U.clk )
\add_26ns_26ns_26_2_1_U5.top_add_26ns_26ns_26_2_1_Adder_2_U.ain_s1  <= _0142_;
always @(posedge \add_26ns_26ns_26_2_1_U5.top_add_26ns_26ns_26_2_1_Adder_2_U.clk )
\add_26ns_26ns_26_2_1_U5.top_add_26ns_26ns_26_2_1_Adder_2_U.sum_s1  <= _0145_;
always @(posedge \add_26ns_26ns_26_2_1_U5.top_add_26ns_26ns_26_2_1_Adder_2_U.clk )
\add_26ns_26ns_26_2_1_U5.top_add_26ns_26ns_26_2_1_Adder_2_U.carry_s1  <= _0144_;
assign _0143_ = \add_26ns_26ns_26_2_1_U5.top_add_26ns_26ns_26_2_1_Adder_2_U.ce  ? \add_26ns_26ns_26_2_1_U5.top_add_26ns_26ns_26_2_1_Adder_2_U.b [25:13] : \add_26ns_26ns_26_2_1_U5.top_add_26ns_26ns_26_2_1_Adder_2_U.bin_s1 ;
assign _0142_ = \add_26ns_26ns_26_2_1_U5.top_add_26ns_26ns_26_2_1_Adder_2_U.ce  ? \add_26ns_26ns_26_2_1_U5.top_add_26ns_26ns_26_2_1_Adder_2_U.a [25:13] : \add_26ns_26ns_26_2_1_U5.top_add_26ns_26ns_26_2_1_Adder_2_U.ain_s1 ;
assign _0144_ = \add_26ns_26ns_26_2_1_U5.top_add_26ns_26ns_26_2_1_Adder_2_U.ce  ? \add_26ns_26ns_26_2_1_U5.top_add_26ns_26ns_26_2_1_Adder_2_U.facout_s1  : \add_26ns_26ns_26_2_1_U5.top_add_26ns_26ns_26_2_1_Adder_2_U.carry_s1 ;
assign _0145_ = \add_26ns_26ns_26_2_1_U5.top_add_26ns_26ns_26_2_1_Adder_2_U.ce  ? \add_26ns_26ns_26_2_1_U5.top_add_26ns_26ns_26_2_1_Adder_2_U.fas_s1  : \add_26ns_26ns_26_2_1_U5.top_add_26ns_26ns_26_2_1_Adder_2_U.sum_s1 ;
assign _0146_ = \add_26ns_26ns_26_2_1_U5.top_add_26ns_26ns_26_2_1_Adder_2_U.u1.a  + \add_26ns_26ns_26_2_1_U5.top_add_26ns_26ns_26_2_1_Adder_2_U.u1.b ;
assign { \add_26ns_26ns_26_2_1_U5.top_add_26ns_26ns_26_2_1_Adder_2_U.u1.cout , \add_26ns_26ns_26_2_1_U5.top_add_26ns_26ns_26_2_1_Adder_2_U.u1.s  } = _0146_ + \add_26ns_26ns_26_2_1_U5.top_add_26ns_26ns_26_2_1_Adder_2_U.u1.cin ;
assign _0147_ = \add_26ns_26ns_26_2_1_U5.top_add_26ns_26ns_26_2_1_Adder_2_U.u2.a  + \add_26ns_26ns_26_2_1_U5.top_add_26ns_26ns_26_2_1_Adder_2_U.u2.b ;
assign { \add_26ns_26ns_26_2_1_U5.top_add_26ns_26ns_26_2_1_Adder_2_U.u2.cout , \add_26ns_26ns_26_2_1_U5.top_add_26ns_26ns_26_2_1_Adder_2_U.u2.s  } = _0147_ + \add_26ns_26ns_26_2_1_U5.top_add_26ns_26ns_26_2_1_Adder_2_U.u2.cin ;
always @(posedge \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_1_U.clk )
\add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_1_U.bin_s1  <= _0149_;
always @(posedge \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_1_U.clk )
\add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_1_U.ain_s1  <= _0148_;
always @(posedge \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_1_U.clk )
\add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_1_U.sum_s1  <= _0151_;
always @(posedge \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_1_U.clk )
\add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_1_U.carry_s1  <= _0150_;
assign _0149_ = \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_1_U.ce  ? \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_1_U.b [1] : \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_1_U.bin_s1 ;
assign _0148_ = \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_1_U.ce  ? \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_1_U.a [1] : \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_1_U.ain_s1 ;
assign _0150_ = \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_1_U.ce  ? \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_1_U.facout_s1  : \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_1_U.carry_s1 ;
assign _0151_ = \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_1_U.ce  ? \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_1_U.fas_s1  : \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_1_U.sum_s1 ;
assign _0152_ = \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.a  + \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.b ;
assign { \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.cout , \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.s  } = _0152_ + \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.cin ;
assign _0153_ = \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.a  + \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.b ;
assign { \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.cout , \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.s  } = _0153_ + \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.cin ;
always @(posedge \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_17_U.clk )
\add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_17_U.bin_s1  <= _0155_;
always @(posedge \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_17_U.clk )
\add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_17_U.ain_s1  <= _0154_;
always @(posedge \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_17_U.clk )
\add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_17_U.sum_s1  <= _0157_;
always @(posedge \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_17_U.clk )
\add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_17_U.carry_s1  <= _0156_;
assign _0155_ = \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_17_U.ce  ? \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_17_U.b [31:16] : \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_17_U.bin_s1 ;
assign _0154_ = \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_17_U.ce  ? \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_17_U.a [31:16] : \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_17_U.ain_s1 ;
assign _0156_ = \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_17_U.ce  ? \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_17_U.facout_s1  : \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_17_U.carry_s1 ;
assign _0157_ = \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_17_U.ce  ? \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_17_U.fas_s1  : \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_17_U.sum_s1 ;
assign _0158_ = \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_17_U.u1.a  + \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_17_U.u1.b ;
assign { \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_17_U.u1.cout , \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_17_U.u1.s  } = _0158_ + \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_17_U.u1.cin ;
assign _0159_ = \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_17_U.u2.a  + \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_17_U.u2.b ;
assign { \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_17_U.u2.cout , \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_17_U.u2.s  } = _0159_ + \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_17_U.u2.cin ;
always @(posedge \add_32s_32ns_32_2_1_U24.top_add_32s_32ns_32_2_1_Adder_19_U.clk )
\add_32s_32ns_32_2_1_U24.top_add_32s_32ns_32_2_1_Adder_19_U.bin_s1  <= _0161_;
always @(posedge \add_32s_32ns_32_2_1_U24.top_add_32s_32ns_32_2_1_Adder_19_U.clk )
\add_32s_32ns_32_2_1_U24.top_add_32s_32ns_32_2_1_Adder_19_U.ain_s1  <= _0160_;
always @(posedge \add_32s_32ns_32_2_1_U24.top_add_32s_32ns_32_2_1_Adder_19_U.clk )
\add_32s_32ns_32_2_1_U24.top_add_32s_32ns_32_2_1_Adder_19_U.sum_s1  <= _0163_;
always @(posedge \add_32s_32ns_32_2_1_U24.top_add_32s_32ns_32_2_1_Adder_19_U.clk )
\add_32s_32ns_32_2_1_U24.top_add_32s_32ns_32_2_1_Adder_19_U.carry_s1  <= _0162_;
assign _0161_ = \add_32s_32ns_32_2_1_U24.top_add_32s_32ns_32_2_1_Adder_19_U.ce  ? \add_32s_32ns_32_2_1_U24.top_add_32s_32ns_32_2_1_Adder_19_U.b [31:16] : \add_32s_32ns_32_2_1_U24.top_add_32s_32ns_32_2_1_Adder_19_U.bin_s1 ;
assign _0160_ = \add_32s_32ns_32_2_1_U24.top_add_32s_32ns_32_2_1_Adder_19_U.ce  ? \add_32s_32ns_32_2_1_U24.top_add_32s_32ns_32_2_1_Adder_19_U.a [31:16] : \add_32s_32ns_32_2_1_U24.top_add_32s_32ns_32_2_1_Adder_19_U.ain_s1 ;
assign _0162_ = \add_32s_32ns_32_2_1_U24.top_add_32s_32ns_32_2_1_Adder_19_U.ce  ? \add_32s_32ns_32_2_1_U24.top_add_32s_32ns_32_2_1_Adder_19_U.facout_s1  : \add_32s_32ns_32_2_1_U24.top_add_32s_32ns_32_2_1_Adder_19_U.carry_s1 ;
assign _0163_ = \add_32s_32ns_32_2_1_U24.top_add_32s_32ns_32_2_1_Adder_19_U.ce  ? \add_32s_32ns_32_2_1_U24.top_add_32s_32ns_32_2_1_Adder_19_U.fas_s1  : \add_32s_32ns_32_2_1_U24.top_add_32s_32ns_32_2_1_Adder_19_U.sum_s1 ;
assign _0164_ = \add_32s_32ns_32_2_1_U24.top_add_32s_32ns_32_2_1_Adder_19_U.u1.a  + \add_32s_32ns_32_2_1_U24.top_add_32s_32ns_32_2_1_Adder_19_U.u1.b ;
assign { \add_32s_32ns_32_2_1_U24.top_add_32s_32ns_32_2_1_Adder_19_U.u1.cout , \add_32s_32ns_32_2_1_U24.top_add_32s_32ns_32_2_1_Adder_19_U.u1.s  } = _0164_ + \add_32s_32ns_32_2_1_U24.top_add_32s_32ns_32_2_1_Adder_19_U.u1.cin ;
assign _0165_ = \add_32s_32ns_32_2_1_U24.top_add_32s_32ns_32_2_1_Adder_19_U.u2.a  + \add_32s_32ns_32_2_1_U24.top_add_32s_32ns_32_2_1_Adder_19_U.u2.b ;
assign { \add_32s_32ns_32_2_1_U24.top_add_32s_32ns_32_2_1_Adder_19_U.u2.cout , \add_32s_32ns_32_2_1_U24.top_add_32s_32ns_32_2_1_Adder_19_U.u2.s  } = _0165_ + \add_32s_32ns_32_2_1_U24.top_add_32s_32ns_32_2_1_Adder_19_U.u2.cin ;
always @(posedge \add_33s_33s_33_2_1_U8.top_add_33s_33s_33_2_1_Adder_5_U.clk )
\add_33s_33s_33_2_1_U8.top_add_33s_33s_33_2_1_Adder_5_U.bin_s1  <= _0167_;
always @(posedge \add_33s_33s_33_2_1_U8.top_add_33s_33s_33_2_1_Adder_5_U.clk )
\add_33s_33s_33_2_1_U8.top_add_33s_33s_33_2_1_Adder_5_U.ain_s1  <= _0166_;
always @(posedge \add_33s_33s_33_2_1_U8.top_add_33s_33s_33_2_1_Adder_5_U.clk )
\add_33s_33s_33_2_1_U8.top_add_33s_33s_33_2_1_Adder_5_U.sum_s1  <= _0169_;
always @(posedge \add_33s_33s_33_2_1_U8.top_add_33s_33s_33_2_1_Adder_5_U.clk )
\add_33s_33s_33_2_1_U8.top_add_33s_33s_33_2_1_Adder_5_U.carry_s1  <= _0168_;
assign _0167_ = \add_33s_33s_33_2_1_U8.top_add_33s_33s_33_2_1_Adder_5_U.ce  ? \add_33s_33s_33_2_1_U8.top_add_33s_33s_33_2_1_Adder_5_U.b [32:16] : \add_33s_33s_33_2_1_U8.top_add_33s_33s_33_2_1_Adder_5_U.bin_s1 ;
assign _0166_ = \add_33s_33s_33_2_1_U8.top_add_33s_33s_33_2_1_Adder_5_U.ce  ? \add_33s_33s_33_2_1_U8.top_add_33s_33s_33_2_1_Adder_5_U.a [32:16] : \add_33s_33s_33_2_1_U8.top_add_33s_33s_33_2_1_Adder_5_U.ain_s1 ;
assign _0168_ = \add_33s_33s_33_2_1_U8.top_add_33s_33s_33_2_1_Adder_5_U.ce  ? \add_33s_33s_33_2_1_U8.top_add_33s_33s_33_2_1_Adder_5_U.facout_s1  : \add_33s_33s_33_2_1_U8.top_add_33s_33s_33_2_1_Adder_5_U.carry_s1 ;
assign _0169_ = \add_33s_33s_33_2_1_U8.top_add_33s_33s_33_2_1_Adder_5_U.ce  ? \add_33s_33s_33_2_1_U8.top_add_33s_33s_33_2_1_Adder_5_U.fas_s1  : \add_33s_33s_33_2_1_U8.top_add_33s_33s_33_2_1_Adder_5_U.sum_s1 ;
assign _0170_ = \add_33s_33s_33_2_1_U8.top_add_33s_33s_33_2_1_Adder_5_U.u1.a  + \add_33s_33s_33_2_1_U8.top_add_33s_33s_33_2_1_Adder_5_U.u1.b ;
assign { \add_33s_33s_33_2_1_U8.top_add_33s_33s_33_2_1_Adder_5_U.u1.cout , \add_33s_33s_33_2_1_U8.top_add_33s_33s_33_2_1_Adder_5_U.u1.s  } = _0170_ + \add_33s_33s_33_2_1_U8.top_add_33s_33s_33_2_1_Adder_5_U.u1.cin ;
assign _0171_ = \add_33s_33s_33_2_1_U8.top_add_33s_33s_33_2_1_Adder_5_U.u2.a  + \add_33s_33s_33_2_1_U8.top_add_33s_33s_33_2_1_Adder_5_U.u2.b ;
assign { \add_33s_33s_33_2_1_U8.top_add_33s_33s_33_2_1_Adder_5_U.u2.cout , \add_33s_33s_33_2_1_U8.top_add_33s_33s_33_2_1_Adder_5_U.u2.s  } = _0171_ + \add_33s_33s_33_2_1_U8.top_add_33s_33s_33_2_1_Adder_5_U.u2.cin ;
always @(posedge \add_39s_39s_39_2_1_U21.top_add_39s_39s_39_2_1_Adder_16_U.clk )
\add_39s_39s_39_2_1_U21.top_add_39s_39s_39_2_1_Adder_16_U.bin_s1  <= _0173_;
always @(posedge \add_39s_39s_39_2_1_U21.top_add_39s_39s_39_2_1_Adder_16_U.clk )
\add_39s_39s_39_2_1_U21.top_add_39s_39s_39_2_1_Adder_16_U.ain_s1  <= _0172_;
always @(posedge \add_39s_39s_39_2_1_U21.top_add_39s_39s_39_2_1_Adder_16_U.clk )
\add_39s_39s_39_2_1_U21.top_add_39s_39s_39_2_1_Adder_16_U.sum_s1  <= _0175_;
always @(posedge \add_39s_39s_39_2_1_U21.top_add_39s_39s_39_2_1_Adder_16_U.clk )
\add_39s_39s_39_2_1_U21.top_add_39s_39s_39_2_1_Adder_16_U.carry_s1  <= _0174_;
assign _0173_ = \add_39s_39s_39_2_1_U21.top_add_39s_39s_39_2_1_Adder_16_U.ce  ? \add_39s_39s_39_2_1_U21.top_add_39s_39s_39_2_1_Adder_16_U.b [38:19] : \add_39s_39s_39_2_1_U21.top_add_39s_39s_39_2_1_Adder_16_U.bin_s1 ;
assign _0172_ = \add_39s_39s_39_2_1_U21.top_add_39s_39s_39_2_1_Adder_16_U.ce  ? \add_39s_39s_39_2_1_U21.top_add_39s_39s_39_2_1_Adder_16_U.a [38:19] : \add_39s_39s_39_2_1_U21.top_add_39s_39s_39_2_1_Adder_16_U.ain_s1 ;
assign _0174_ = \add_39s_39s_39_2_1_U21.top_add_39s_39s_39_2_1_Adder_16_U.ce  ? \add_39s_39s_39_2_1_U21.top_add_39s_39s_39_2_1_Adder_16_U.facout_s1  : \add_39s_39s_39_2_1_U21.top_add_39s_39s_39_2_1_Adder_16_U.carry_s1 ;
assign _0175_ = \add_39s_39s_39_2_1_U21.top_add_39s_39s_39_2_1_Adder_16_U.ce  ? \add_39s_39s_39_2_1_U21.top_add_39s_39s_39_2_1_Adder_16_U.fas_s1  : \add_39s_39s_39_2_1_U21.top_add_39s_39s_39_2_1_Adder_16_U.sum_s1 ;
assign _0176_ = \add_39s_39s_39_2_1_U21.top_add_39s_39s_39_2_1_Adder_16_U.u1.a  + \add_39s_39s_39_2_1_U21.top_add_39s_39s_39_2_1_Adder_16_U.u1.b ;
assign { \add_39s_39s_39_2_1_U21.top_add_39s_39s_39_2_1_Adder_16_U.u1.cout , \add_39s_39s_39_2_1_U21.top_add_39s_39s_39_2_1_Adder_16_U.u1.s  } = _0176_ + \add_39s_39s_39_2_1_U21.top_add_39s_39s_39_2_1_Adder_16_U.u1.cin ;
assign _0177_ = \add_39s_39s_39_2_1_U21.top_add_39s_39s_39_2_1_Adder_16_U.u2.a  + \add_39s_39s_39_2_1_U21.top_add_39s_39s_39_2_1_Adder_16_U.u2.b ;
assign { \add_39s_39s_39_2_1_U21.top_add_39s_39s_39_2_1_Adder_16_U.u2.cout , \add_39s_39s_39_2_1_U21.top_add_39s_39s_39_2_1_Adder_16_U.u2.s  } = _0177_ + \add_39s_39s_39_2_1_U21.top_add_39s_39s_39_2_1_Adder_16_U.u2.cin ;
always @(posedge \add_3s_3ns_3_2_1_U11.top_add_3s_3ns_3_2_1_Adder_8_U.clk )
\add_3s_3ns_3_2_1_U11.top_add_3s_3ns_3_2_1_Adder_8_U.bin_s1  <= _0179_;
always @(posedge \add_3s_3ns_3_2_1_U11.top_add_3s_3ns_3_2_1_Adder_8_U.clk )
\add_3s_3ns_3_2_1_U11.top_add_3s_3ns_3_2_1_Adder_8_U.ain_s1  <= _0178_;
always @(posedge \add_3s_3ns_3_2_1_U11.top_add_3s_3ns_3_2_1_Adder_8_U.clk )
\add_3s_3ns_3_2_1_U11.top_add_3s_3ns_3_2_1_Adder_8_U.sum_s1  <= _0181_;
always @(posedge \add_3s_3ns_3_2_1_U11.top_add_3s_3ns_3_2_1_Adder_8_U.clk )
\add_3s_3ns_3_2_1_U11.top_add_3s_3ns_3_2_1_Adder_8_U.carry_s1  <= _0180_;
assign _0179_ = \add_3s_3ns_3_2_1_U11.top_add_3s_3ns_3_2_1_Adder_8_U.ce  ? \add_3s_3ns_3_2_1_U11.top_add_3s_3ns_3_2_1_Adder_8_U.b [2:1] : \add_3s_3ns_3_2_1_U11.top_add_3s_3ns_3_2_1_Adder_8_U.bin_s1 ;
assign _0178_ = \add_3s_3ns_3_2_1_U11.top_add_3s_3ns_3_2_1_Adder_8_U.ce  ? \add_3s_3ns_3_2_1_U11.top_add_3s_3ns_3_2_1_Adder_8_U.a [2:1] : \add_3s_3ns_3_2_1_U11.top_add_3s_3ns_3_2_1_Adder_8_U.ain_s1 ;
assign _0180_ = \add_3s_3ns_3_2_1_U11.top_add_3s_3ns_3_2_1_Adder_8_U.ce  ? \add_3s_3ns_3_2_1_U11.top_add_3s_3ns_3_2_1_Adder_8_U.facout_s1  : \add_3s_3ns_3_2_1_U11.top_add_3s_3ns_3_2_1_Adder_8_U.carry_s1 ;
assign _0181_ = \add_3s_3ns_3_2_1_U11.top_add_3s_3ns_3_2_1_Adder_8_U.ce  ? \add_3s_3ns_3_2_1_U11.top_add_3s_3ns_3_2_1_Adder_8_U.fas_s1  : \add_3s_3ns_3_2_1_U11.top_add_3s_3ns_3_2_1_Adder_8_U.sum_s1 ;
assign _0182_ = \add_3s_3ns_3_2_1_U11.top_add_3s_3ns_3_2_1_Adder_8_U.u1.a  + \add_3s_3ns_3_2_1_U11.top_add_3s_3ns_3_2_1_Adder_8_U.u1.b ;
assign { \add_3s_3ns_3_2_1_U11.top_add_3s_3ns_3_2_1_Adder_8_U.u1.cout , \add_3s_3ns_3_2_1_U11.top_add_3s_3ns_3_2_1_Adder_8_U.u1.s  } = _0182_ + \add_3s_3ns_3_2_1_U11.top_add_3s_3ns_3_2_1_Adder_8_U.u1.cin ;
assign _0183_ = \add_3s_3ns_3_2_1_U11.top_add_3s_3ns_3_2_1_Adder_8_U.u2.a  + \add_3s_3ns_3_2_1_U11.top_add_3s_3ns_3_2_1_Adder_8_U.u2.b ;
assign { \add_3s_3ns_3_2_1_U11.top_add_3s_3ns_3_2_1_Adder_8_U.u2.cout , \add_3s_3ns_3_2_1_U11.top_add_3s_3ns_3_2_1_Adder_8_U.u2.s  } = _0183_ + \add_3s_3ns_3_2_1_U11.top_add_3s_3ns_3_2_1_Adder_8_U.u2.cin ;
always @(posedge \add_4ns_4ns_4_2_1_U12.top_add_4ns_4ns_4_2_1_Adder_9_U.clk )
\add_4ns_4ns_4_2_1_U12.top_add_4ns_4ns_4_2_1_Adder_9_U.bin_s1  <= _0185_;
always @(posedge \add_4ns_4ns_4_2_1_U12.top_add_4ns_4ns_4_2_1_Adder_9_U.clk )
\add_4ns_4ns_4_2_1_U12.top_add_4ns_4ns_4_2_1_Adder_9_U.ain_s1  <= _0184_;
always @(posedge \add_4ns_4ns_4_2_1_U12.top_add_4ns_4ns_4_2_1_Adder_9_U.clk )
\add_4ns_4ns_4_2_1_U12.top_add_4ns_4ns_4_2_1_Adder_9_U.sum_s1  <= _0187_;
always @(posedge \add_4ns_4ns_4_2_1_U12.top_add_4ns_4ns_4_2_1_Adder_9_U.clk )
\add_4ns_4ns_4_2_1_U12.top_add_4ns_4ns_4_2_1_Adder_9_U.carry_s1  <= _0186_;
assign _0185_ = \add_4ns_4ns_4_2_1_U12.top_add_4ns_4ns_4_2_1_Adder_9_U.ce  ? \add_4ns_4ns_4_2_1_U12.top_add_4ns_4ns_4_2_1_Adder_9_U.b [3:2] : \add_4ns_4ns_4_2_1_U12.top_add_4ns_4ns_4_2_1_Adder_9_U.bin_s1 ;
assign _0184_ = \add_4ns_4ns_4_2_1_U12.top_add_4ns_4ns_4_2_1_Adder_9_U.ce  ? \add_4ns_4ns_4_2_1_U12.top_add_4ns_4ns_4_2_1_Adder_9_U.a [3:2] : \add_4ns_4ns_4_2_1_U12.top_add_4ns_4ns_4_2_1_Adder_9_U.ain_s1 ;
assign _0186_ = \add_4ns_4ns_4_2_1_U12.top_add_4ns_4ns_4_2_1_Adder_9_U.ce  ? \add_4ns_4ns_4_2_1_U12.top_add_4ns_4ns_4_2_1_Adder_9_U.facout_s1  : \add_4ns_4ns_4_2_1_U12.top_add_4ns_4ns_4_2_1_Adder_9_U.carry_s1 ;
assign _0187_ = \add_4ns_4ns_4_2_1_U12.top_add_4ns_4ns_4_2_1_Adder_9_U.ce  ? \add_4ns_4ns_4_2_1_U12.top_add_4ns_4ns_4_2_1_Adder_9_U.fas_s1  : \add_4ns_4ns_4_2_1_U12.top_add_4ns_4ns_4_2_1_Adder_9_U.sum_s1 ;
assign _0188_ = \add_4ns_4ns_4_2_1_U12.top_add_4ns_4ns_4_2_1_Adder_9_U.u1.a  + \add_4ns_4ns_4_2_1_U12.top_add_4ns_4ns_4_2_1_Adder_9_U.u1.b ;
assign { \add_4ns_4ns_4_2_1_U12.top_add_4ns_4ns_4_2_1_Adder_9_U.u1.cout , \add_4ns_4ns_4_2_1_U12.top_add_4ns_4ns_4_2_1_Adder_9_U.u1.s  } = _0188_ + \add_4ns_4ns_4_2_1_U12.top_add_4ns_4ns_4_2_1_Adder_9_U.u1.cin ;
assign _0189_ = \add_4ns_4ns_4_2_1_U12.top_add_4ns_4ns_4_2_1_Adder_9_U.u2.a  + \add_4ns_4ns_4_2_1_U12.top_add_4ns_4ns_4_2_1_Adder_9_U.u2.b ;
assign { \add_4ns_4ns_4_2_1_U12.top_add_4ns_4ns_4_2_1_Adder_9_U.u2.cout , \add_4ns_4ns_4_2_1_U12.top_add_4ns_4ns_4_2_1_Adder_9_U.u2.s  } = _0189_ + \add_4ns_4ns_4_2_1_U12.top_add_4ns_4ns_4_2_1_Adder_9_U.u2.cin ;
always @(posedge \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_9_U.clk )
\add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_9_U.bin_s1  <= _0191_;
always @(posedge \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_9_U.clk )
\add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_9_U.ain_s1  <= _0190_;
always @(posedge \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_9_U.clk )
\add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_9_U.sum_s1  <= _0193_;
always @(posedge \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_9_U.clk )
\add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_9_U.carry_s1  <= _0192_;
assign _0191_ = \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_9_U.ce  ? \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_9_U.b [3:2] : \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_9_U.bin_s1 ;
assign _0190_ = \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_9_U.ce  ? \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_9_U.a [3:2] : \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_9_U.ain_s1 ;
assign _0192_ = \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_9_U.ce  ? \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_9_U.facout_s1  : \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_9_U.carry_s1 ;
assign _0193_ = \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_9_U.ce  ? \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_9_U.fas_s1  : \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_9_U.sum_s1 ;
assign _0194_ = \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_9_U.u1.a  + \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_9_U.u1.b ;
assign { \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_9_U.u1.cout , \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_9_U.u1.s  } = _0194_ + \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_9_U.u1.cin ;
assign _0195_ = \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_9_U.u2.a  + \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_9_U.u2.b ;
assign { \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_9_U.u2.cout , \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_9_U.u2.s  } = _0195_ + \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_9_U.u2.cin ;
always @(posedge \add_4ns_4ns_4_2_1_U15.top_add_4ns_4ns_4_2_1_Adder_9_U.clk )
\add_4ns_4ns_4_2_1_U15.top_add_4ns_4ns_4_2_1_Adder_9_U.bin_s1  <= _0197_;
always @(posedge \add_4ns_4ns_4_2_1_U15.top_add_4ns_4ns_4_2_1_Adder_9_U.clk )
\add_4ns_4ns_4_2_1_U15.top_add_4ns_4ns_4_2_1_Adder_9_U.ain_s1  <= _0196_;
always @(posedge \add_4ns_4ns_4_2_1_U15.top_add_4ns_4ns_4_2_1_Adder_9_U.clk )
\add_4ns_4ns_4_2_1_U15.top_add_4ns_4ns_4_2_1_Adder_9_U.sum_s1  <= _0199_;
always @(posedge \add_4ns_4ns_4_2_1_U15.top_add_4ns_4ns_4_2_1_Adder_9_U.clk )
\add_4ns_4ns_4_2_1_U15.top_add_4ns_4ns_4_2_1_Adder_9_U.carry_s1  <= _0198_;
assign _0197_ = \add_4ns_4ns_4_2_1_U15.top_add_4ns_4ns_4_2_1_Adder_9_U.ce  ? \add_4ns_4ns_4_2_1_U15.top_add_4ns_4ns_4_2_1_Adder_9_U.b [3:2] : \add_4ns_4ns_4_2_1_U15.top_add_4ns_4ns_4_2_1_Adder_9_U.bin_s1 ;
assign _0196_ = \add_4ns_4ns_4_2_1_U15.top_add_4ns_4ns_4_2_1_Adder_9_U.ce  ? \add_4ns_4ns_4_2_1_U15.top_add_4ns_4ns_4_2_1_Adder_9_U.a [3:2] : \add_4ns_4ns_4_2_1_U15.top_add_4ns_4ns_4_2_1_Adder_9_U.ain_s1 ;
assign _0198_ = \add_4ns_4ns_4_2_1_U15.top_add_4ns_4ns_4_2_1_Adder_9_U.ce  ? \add_4ns_4ns_4_2_1_U15.top_add_4ns_4ns_4_2_1_Adder_9_U.facout_s1  : \add_4ns_4ns_4_2_1_U15.top_add_4ns_4ns_4_2_1_Adder_9_U.carry_s1 ;
assign _0199_ = \add_4ns_4ns_4_2_1_U15.top_add_4ns_4ns_4_2_1_Adder_9_U.ce  ? \add_4ns_4ns_4_2_1_U15.top_add_4ns_4ns_4_2_1_Adder_9_U.fas_s1  : \add_4ns_4ns_4_2_1_U15.top_add_4ns_4ns_4_2_1_Adder_9_U.sum_s1 ;
assign _0200_ = \add_4ns_4ns_4_2_1_U15.top_add_4ns_4ns_4_2_1_Adder_9_U.u1.a  + \add_4ns_4ns_4_2_1_U15.top_add_4ns_4ns_4_2_1_Adder_9_U.u1.b ;
assign { \add_4ns_4ns_4_2_1_U15.top_add_4ns_4ns_4_2_1_Adder_9_U.u1.cout , \add_4ns_4ns_4_2_1_U15.top_add_4ns_4ns_4_2_1_Adder_9_U.u1.s  } = _0200_ + \add_4ns_4ns_4_2_1_U15.top_add_4ns_4ns_4_2_1_Adder_9_U.u1.cin ;
assign _0201_ = \add_4ns_4ns_4_2_1_U15.top_add_4ns_4ns_4_2_1_Adder_9_U.u2.a  + \add_4ns_4ns_4_2_1_U15.top_add_4ns_4ns_4_2_1_Adder_9_U.u2.b ;
assign { \add_4ns_4ns_4_2_1_U15.top_add_4ns_4ns_4_2_1_Adder_9_U.u2.cout , \add_4ns_4ns_4_2_1_U15.top_add_4ns_4ns_4_2_1_Adder_9_U.u2.s  } = _0201_ + \add_4ns_4ns_4_2_1_U15.top_add_4ns_4ns_4_2_1_Adder_9_U.u2.cin ;
always @(posedge \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_10_U.clk )
\add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_10_U.sum_s1  <= _0205_;
always @(posedge \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_10_U.clk )
\add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_10_U.carry_s1  <= _0204_;
always @(posedge \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_10_U.clk )
\add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_10_U.bin_s1  <= _0203_;
always @(posedge \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_10_U.clk )
\add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_10_U.ain_s1  <= _0202_;
assign _0203_ = \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_10_U.ce  ? \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_10_U.b [3:2] : \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_10_U.bin_s1 ;
assign _0202_ = \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_10_U.ce  ? \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_10_U.a [3:2] : \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_10_U.ain_s1 ;
assign _0204_ = \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_10_U.ce  ? \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_10_U.facout_s1  : \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_10_U.carry_s1 ;
assign _0205_ = \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_10_U.ce  ? \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_10_U.fas_s1  : \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_10_U.sum_s1 ;
assign _0206_ = \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_10_U.u1.a  + \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_10_U.u1.b ;
assign { \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_10_U.u1.cout , \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_10_U.u1.s  } = _0206_ + \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_10_U.u1.cin ;
assign _0207_ = \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_10_U.u2.a  + \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_10_U.u2.b ;
assign { \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_10_U.u2.cout , \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_10_U.u2.s  } = _0207_ + \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_10_U.u2.cin ;
always @(posedge \add_4s_4ns_4_2_1_U16.top_add_4s_4ns_4_2_1_Adder_11_U.clk )
\add_4s_4ns_4_2_1_U16.top_add_4s_4ns_4_2_1_Adder_11_U.bin_s1  <= _0209_;
always @(posedge \add_4s_4ns_4_2_1_U16.top_add_4s_4ns_4_2_1_Adder_11_U.clk )
\add_4s_4ns_4_2_1_U16.top_add_4s_4ns_4_2_1_Adder_11_U.ain_s1  <= _0208_;
always @(posedge \add_4s_4ns_4_2_1_U16.top_add_4s_4ns_4_2_1_Adder_11_U.clk )
\add_4s_4ns_4_2_1_U16.top_add_4s_4ns_4_2_1_Adder_11_U.sum_s1  <= _0211_;
always @(posedge \add_4s_4ns_4_2_1_U16.top_add_4s_4ns_4_2_1_Adder_11_U.clk )
\add_4s_4ns_4_2_1_U16.top_add_4s_4ns_4_2_1_Adder_11_U.carry_s1  <= _0210_;
assign _0209_ = \add_4s_4ns_4_2_1_U16.top_add_4s_4ns_4_2_1_Adder_11_U.ce  ? \add_4s_4ns_4_2_1_U16.top_add_4s_4ns_4_2_1_Adder_11_U.b [3:2] : \add_4s_4ns_4_2_1_U16.top_add_4s_4ns_4_2_1_Adder_11_U.bin_s1 ;
assign _0208_ = \add_4s_4ns_4_2_1_U16.top_add_4s_4ns_4_2_1_Adder_11_U.ce  ? \add_4s_4ns_4_2_1_U16.top_add_4s_4ns_4_2_1_Adder_11_U.a [3:2] : \add_4s_4ns_4_2_1_U16.top_add_4s_4ns_4_2_1_Adder_11_U.ain_s1 ;
assign _0210_ = \add_4s_4ns_4_2_1_U16.top_add_4s_4ns_4_2_1_Adder_11_U.ce  ? \add_4s_4ns_4_2_1_U16.top_add_4s_4ns_4_2_1_Adder_11_U.facout_s1  : \add_4s_4ns_4_2_1_U16.top_add_4s_4ns_4_2_1_Adder_11_U.carry_s1 ;
assign _0211_ = \add_4s_4ns_4_2_1_U16.top_add_4s_4ns_4_2_1_Adder_11_U.ce  ? \add_4s_4ns_4_2_1_U16.top_add_4s_4ns_4_2_1_Adder_11_U.fas_s1  : \add_4s_4ns_4_2_1_U16.top_add_4s_4ns_4_2_1_Adder_11_U.sum_s1 ;
assign _0212_ = \add_4s_4ns_4_2_1_U16.top_add_4s_4ns_4_2_1_Adder_11_U.u1.a  + \add_4s_4ns_4_2_1_U16.top_add_4s_4ns_4_2_1_Adder_11_U.u1.b ;
assign { \add_4s_4ns_4_2_1_U16.top_add_4s_4ns_4_2_1_Adder_11_U.u1.cout , \add_4s_4ns_4_2_1_U16.top_add_4s_4ns_4_2_1_Adder_11_U.u1.s  } = _0212_ + \add_4s_4ns_4_2_1_U16.top_add_4s_4ns_4_2_1_Adder_11_U.u1.cin ;
assign _0213_ = \add_4s_4ns_4_2_1_U16.top_add_4s_4ns_4_2_1_Adder_11_U.u2.a  + \add_4s_4ns_4_2_1_U16.top_add_4s_4ns_4_2_1_Adder_11_U.u2.b ;
assign { \add_4s_4ns_4_2_1_U16.top_add_4s_4ns_4_2_1_Adder_11_U.u2.cout , \add_4s_4ns_4_2_1_U16.top_add_4s_4ns_4_2_1_Adder_11_U.u2.s  } = _0213_ + \add_4s_4ns_4_2_1_U16.top_add_4s_4ns_4_2_1_Adder_11_U.u2.cin ;
always @(posedge \add_5ns_5s_5_2_1_U18.top_add_5ns_5s_5_2_1_Adder_13_U.clk )
\add_5ns_5s_5_2_1_U18.top_add_5ns_5s_5_2_1_Adder_13_U.bin_s1  <= _0215_;
always @(posedge \add_5ns_5s_5_2_1_U18.top_add_5ns_5s_5_2_1_Adder_13_U.clk )
\add_5ns_5s_5_2_1_U18.top_add_5ns_5s_5_2_1_Adder_13_U.ain_s1  <= _0214_;
always @(posedge \add_5ns_5s_5_2_1_U18.top_add_5ns_5s_5_2_1_Adder_13_U.clk )
\add_5ns_5s_5_2_1_U18.top_add_5ns_5s_5_2_1_Adder_13_U.sum_s1  <= _0217_;
always @(posedge \add_5ns_5s_5_2_1_U18.top_add_5ns_5s_5_2_1_Adder_13_U.clk )
\add_5ns_5s_5_2_1_U18.top_add_5ns_5s_5_2_1_Adder_13_U.carry_s1  <= _0216_;
assign _0215_ = \add_5ns_5s_5_2_1_U18.top_add_5ns_5s_5_2_1_Adder_13_U.ce  ? \add_5ns_5s_5_2_1_U18.top_add_5ns_5s_5_2_1_Adder_13_U.b [4:2] : \add_5ns_5s_5_2_1_U18.top_add_5ns_5s_5_2_1_Adder_13_U.bin_s1 ;
assign _0214_ = \add_5ns_5s_5_2_1_U18.top_add_5ns_5s_5_2_1_Adder_13_U.ce  ? \add_5ns_5s_5_2_1_U18.top_add_5ns_5s_5_2_1_Adder_13_U.a [4:2] : \add_5ns_5s_5_2_1_U18.top_add_5ns_5s_5_2_1_Adder_13_U.ain_s1 ;
assign _0216_ = \add_5ns_5s_5_2_1_U18.top_add_5ns_5s_5_2_1_Adder_13_U.ce  ? \add_5ns_5s_5_2_1_U18.top_add_5ns_5s_5_2_1_Adder_13_U.facout_s1  : \add_5ns_5s_5_2_1_U18.top_add_5ns_5s_5_2_1_Adder_13_U.carry_s1 ;
assign _0217_ = \add_5ns_5s_5_2_1_U18.top_add_5ns_5s_5_2_1_Adder_13_U.ce  ? \add_5ns_5s_5_2_1_U18.top_add_5ns_5s_5_2_1_Adder_13_U.fas_s1  : \add_5ns_5s_5_2_1_U18.top_add_5ns_5s_5_2_1_Adder_13_U.sum_s1 ;
assign _0218_ = \add_5ns_5s_5_2_1_U18.top_add_5ns_5s_5_2_1_Adder_13_U.u1.a  + \add_5ns_5s_5_2_1_U18.top_add_5ns_5s_5_2_1_Adder_13_U.u1.b ;
assign { \add_5ns_5s_5_2_1_U18.top_add_5ns_5s_5_2_1_Adder_13_U.u1.cout , \add_5ns_5s_5_2_1_U18.top_add_5ns_5s_5_2_1_Adder_13_U.u1.s  } = _0218_ + \add_5ns_5s_5_2_1_U18.top_add_5ns_5s_5_2_1_Adder_13_U.u1.cin ;
assign _0219_ = \add_5ns_5s_5_2_1_U18.top_add_5ns_5s_5_2_1_Adder_13_U.u2.a  + \add_5ns_5s_5_2_1_U18.top_add_5ns_5s_5_2_1_Adder_13_U.u2.b ;
assign { \add_5ns_5s_5_2_1_U18.top_add_5ns_5s_5_2_1_Adder_13_U.u2.cout , \add_5ns_5s_5_2_1_U18.top_add_5ns_5s_5_2_1_Adder_13_U.u2.s  } = _0219_ + \add_5ns_5s_5_2_1_U18.top_add_5ns_5s_5_2_1_Adder_13_U.u2.cin ;
always @(posedge \add_5s_5s_5_2_1_U17.top_add_5s_5s_5_2_1_Adder_12_U.clk )
\add_5s_5s_5_2_1_U17.top_add_5s_5s_5_2_1_Adder_12_U.bin_s1  <= _0221_;
always @(posedge \add_5s_5s_5_2_1_U17.top_add_5s_5s_5_2_1_Adder_12_U.clk )
\add_5s_5s_5_2_1_U17.top_add_5s_5s_5_2_1_Adder_12_U.ain_s1  <= _0220_;
always @(posedge \add_5s_5s_5_2_1_U17.top_add_5s_5s_5_2_1_Adder_12_U.clk )
\add_5s_5s_5_2_1_U17.top_add_5s_5s_5_2_1_Adder_12_U.sum_s1  <= _0223_;
always @(posedge \add_5s_5s_5_2_1_U17.top_add_5s_5s_5_2_1_Adder_12_U.clk )
\add_5s_5s_5_2_1_U17.top_add_5s_5s_5_2_1_Adder_12_U.carry_s1  <= _0222_;
assign _0221_ = \add_5s_5s_5_2_1_U17.top_add_5s_5s_5_2_1_Adder_12_U.ce  ? \add_5s_5s_5_2_1_U17.top_add_5s_5s_5_2_1_Adder_12_U.b [4:2] : \add_5s_5s_5_2_1_U17.top_add_5s_5s_5_2_1_Adder_12_U.bin_s1 ;
assign _0220_ = \add_5s_5s_5_2_1_U17.top_add_5s_5s_5_2_1_Adder_12_U.ce  ? \add_5s_5s_5_2_1_U17.top_add_5s_5s_5_2_1_Adder_12_U.a [4:2] : \add_5s_5s_5_2_1_U17.top_add_5s_5s_5_2_1_Adder_12_U.ain_s1 ;
assign _0222_ = \add_5s_5s_5_2_1_U17.top_add_5s_5s_5_2_1_Adder_12_U.ce  ? \add_5s_5s_5_2_1_U17.top_add_5s_5s_5_2_1_Adder_12_U.facout_s1  : \add_5s_5s_5_2_1_U17.top_add_5s_5s_5_2_1_Adder_12_U.carry_s1 ;
assign _0223_ = \add_5s_5s_5_2_1_U17.top_add_5s_5s_5_2_1_Adder_12_U.ce  ? \add_5s_5s_5_2_1_U17.top_add_5s_5s_5_2_1_Adder_12_U.fas_s1  : \add_5s_5s_5_2_1_U17.top_add_5s_5s_5_2_1_Adder_12_U.sum_s1 ;
assign _0224_ = \add_5s_5s_5_2_1_U17.top_add_5s_5s_5_2_1_Adder_12_U.u1.a  + \add_5s_5s_5_2_1_U17.top_add_5s_5s_5_2_1_Adder_12_U.u1.b ;
assign { \add_5s_5s_5_2_1_U17.top_add_5s_5s_5_2_1_Adder_12_U.u1.cout , \add_5s_5s_5_2_1_U17.top_add_5s_5s_5_2_1_Adder_12_U.u1.s  } = _0224_ + \add_5s_5s_5_2_1_U17.top_add_5s_5s_5_2_1_Adder_12_U.u1.cin ;
assign _0225_ = \add_5s_5s_5_2_1_U17.top_add_5s_5s_5_2_1_Adder_12_U.u2.a  + \add_5s_5s_5_2_1_U17.top_add_5s_5s_5_2_1_Adder_12_U.u2.b ;
assign { \add_5s_5s_5_2_1_U17.top_add_5s_5s_5_2_1_Adder_12_U.u2.cout , \add_5s_5s_5_2_1_U17.top_add_5s_5s_5_2_1_Adder_12_U.u2.s  } = _0225_ + \add_5s_5s_5_2_1_U17.top_add_5s_5s_5_2_1_Adder_12_U.u2.cin ;
always @(posedge \add_6ns_6s_6_2_1_U20.top_add_6ns_6s_6_2_1_Adder_15_U.clk )
\add_6ns_6s_6_2_1_U20.top_add_6ns_6s_6_2_1_Adder_15_U.bin_s1  <= _0227_;
always @(posedge \add_6ns_6s_6_2_1_U20.top_add_6ns_6s_6_2_1_Adder_15_U.clk )
\add_6ns_6s_6_2_1_U20.top_add_6ns_6s_6_2_1_Adder_15_U.ain_s1  <= _0226_;
always @(posedge \add_6ns_6s_6_2_1_U20.top_add_6ns_6s_6_2_1_Adder_15_U.clk )
\add_6ns_6s_6_2_1_U20.top_add_6ns_6s_6_2_1_Adder_15_U.sum_s1  <= _0229_;
always @(posedge \add_6ns_6s_6_2_1_U20.top_add_6ns_6s_6_2_1_Adder_15_U.clk )
\add_6ns_6s_6_2_1_U20.top_add_6ns_6s_6_2_1_Adder_15_U.carry_s1  <= _0228_;
assign _0227_ = \add_6ns_6s_6_2_1_U20.top_add_6ns_6s_6_2_1_Adder_15_U.ce  ? \add_6ns_6s_6_2_1_U20.top_add_6ns_6s_6_2_1_Adder_15_U.b [5:3] : \add_6ns_6s_6_2_1_U20.top_add_6ns_6s_6_2_1_Adder_15_U.bin_s1 ;
assign _0226_ = \add_6ns_6s_6_2_1_U20.top_add_6ns_6s_6_2_1_Adder_15_U.ce  ? \add_6ns_6s_6_2_1_U20.top_add_6ns_6s_6_2_1_Adder_15_U.a [5:3] : \add_6ns_6s_6_2_1_U20.top_add_6ns_6s_6_2_1_Adder_15_U.ain_s1 ;
assign _0228_ = \add_6ns_6s_6_2_1_U20.top_add_6ns_6s_6_2_1_Adder_15_U.ce  ? \add_6ns_6s_6_2_1_U20.top_add_6ns_6s_6_2_1_Adder_15_U.facout_s1  : \add_6ns_6s_6_2_1_U20.top_add_6ns_6s_6_2_1_Adder_15_U.carry_s1 ;
assign _0229_ = \add_6ns_6s_6_2_1_U20.top_add_6ns_6s_6_2_1_Adder_15_U.ce  ? \add_6ns_6s_6_2_1_U20.top_add_6ns_6s_6_2_1_Adder_15_U.fas_s1  : \add_6ns_6s_6_2_1_U20.top_add_6ns_6s_6_2_1_Adder_15_U.sum_s1 ;
assign _0230_ = \add_6ns_6s_6_2_1_U20.top_add_6ns_6s_6_2_1_Adder_15_U.u1.a  + \add_6ns_6s_6_2_1_U20.top_add_6ns_6s_6_2_1_Adder_15_U.u1.b ;
assign { \add_6ns_6s_6_2_1_U20.top_add_6ns_6s_6_2_1_Adder_15_U.u1.cout , \add_6ns_6s_6_2_1_U20.top_add_6ns_6s_6_2_1_Adder_15_U.u1.s  } = _0230_ + \add_6ns_6s_6_2_1_U20.top_add_6ns_6s_6_2_1_Adder_15_U.u1.cin ;
assign _0231_ = \add_6ns_6s_6_2_1_U20.top_add_6ns_6s_6_2_1_Adder_15_U.u2.a  + \add_6ns_6s_6_2_1_U20.top_add_6ns_6s_6_2_1_Adder_15_U.u2.b ;
assign { \add_6ns_6s_6_2_1_U20.top_add_6ns_6s_6_2_1_Adder_15_U.u2.cout , \add_6ns_6s_6_2_1_U20.top_add_6ns_6s_6_2_1_Adder_15_U.u2.s  } = _0231_ + \add_6ns_6s_6_2_1_U20.top_add_6ns_6s_6_2_1_Adder_15_U.u2.cin ;
always @(posedge \add_6s_6s_6_2_1_U19.top_add_6s_6s_6_2_1_Adder_14_U.clk )
\add_6s_6s_6_2_1_U19.top_add_6s_6s_6_2_1_Adder_14_U.bin_s1  <= _0233_;
always @(posedge \add_6s_6s_6_2_1_U19.top_add_6s_6s_6_2_1_Adder_14_U.clk )
\add_6s_6s_6_2_1_U19.top_add_6s_6s_6_2_1_Adder_14_U.ain_s1  <= _0232_;
always @(posedge \add_6s_6s_6_2_1_U19.top_add_6s_6s_6_2_1_Adder_14_U.clk )
\add_6s_6s_6_2_1_U19.top_add_6s_6s_6_2_1_Adder_14_U.sum_s1  <= _0235_;
always @(posedge \add_6s_6s_6_2_1_U19.top_add_6s_6s_6_2_1_Adder_14_U.clk )
\add_6s_6s_6_2_1_U19.top_add_6s_6s_6_2_1_Adder_14_U.carry_s1  <= _0234_;
assign _0233_ = \add_6s_6s_6_2_1_U19.top_add_6s_6s_6_2_1_Adder_14_U.ce  ? \add_6s_6s_6_2_1_U19.top_add_6s_6s_6_2_1_Adder_14_U.b [5:3] : \add_6s_6s_6_2_1_U19.top_add_6s_6s_6_2_1_Adder_14_U.bin_s1 ;
assign _0232_ = \add_6s_6s_6_2_1_U19.top_add_6s_6s_6_2_1_Adder_14_U.ce  ? \add_6s_6s_6_2_1_U19.top_add_6s_6s_6_2_1_Adder_14_U.a [5:3] : \add_6s_6s_6_2_1_U19.top_add_6s_6s_6_2_1_Adder_14_U.ain_s1 ;
assign _0234_ = \add_6s_6s_6_2_1_U19.top_add_6s_6s_6_2_1_Adder_14_U.ce  ? \add_6s_6s_6_2_1_U19.top_add_6s_6s_6_2_1_Adder_14_U.facout_s1  : \add_6s_6s_6_2_1_U19.top_add_6s_6s_6_2_1_Adder_14_U.carry_s1 ;
assign _0235_ = \add_6s_6s_6_2_1_U19.top_add_6s_6s_6_2_1_Adder_14_U.ce  ? \add_6s_6s_6_2_1_U19.top_add_6s_6s_6_2_1_Adder_14_U.fas_s1  : \add_6s_6s_6_2_1_U19.top_add_6s_6s_6_2_1_Adder_14_U.sum_s1 ;
assign _0236_ = \add_6s_6s_6_2_1_U19.top_add_6s_6s_6_2_1_Adder_14_U.u1.a  + \add_6s_6s_6_2_1_U19.top_add_6s_6s_6_2_1_Adder_14_U.u1.b ;
assign { \add_6s_6s_6_2_1_U19.top_add_6s_6s_6_2_1_Adder_14_U.u1.cout , \add_6s_6s_6_2_1_U19.top_add_6s_6s_6_2_1_Adder_14_U.u1.s  } = _0236_ + \add_6s_6s_6_2_1_U19.top_add_6s_6s_6_2_1_Adder_14_U.u1.cin ;
assign _0237_ = \add_6s_6s_6_2_1_U19.top_add_6s_6s_6_2_1_Adder_14_U.u2.a  + \add_6s_6s_6_2_1_U19.top_add_6s_6s_6_2_1_Adder_14_U.u2.b ;
assign { \add_6s_6s_6_2_1_U19.top_add_6s_6s_6_2_1_Adder_14_U.u2.cout , \add_6s_6s_6_2_1_U19.top_add_6s_6s_6_2_1_Adder_14_U.u2.s  } = _0237_ + \add_6s_6s_6_2_1_U19.top_add_6s_6s_6_2_1_Adder_14_U.u2.cin ;
always @(posedge \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_4_U.clk )
\add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_4_U.bin_s1  <= _0239_;
always @(posedge \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_4_U.clk )
\add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_4_U.ain_s1  <= _0238_;
always @(posedge \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_4_U.clk )
\add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_4_U.sum_s1  <= _0241_;
always @(posedge \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_4_U.clk )
\add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_4_U.carry_s1  <= _0240_;
assign _0239_ = \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_4_U.ce  ? \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_4_U.b [7:4] : \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_4_U.bin_s1 ;
assign _0238_ = \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_4_U.ce  ? \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_4_U.a [7:4] : \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_4_U.ain_s1 ;
assign _0240_ = \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_4_U.ce  ? \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_4_U.facout_s1  : \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_4_U.carry_s1 ;
assign _0241_ = \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_4_U.ce  ? \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_4_U.fas_s1  : \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_4_U.sum_s1 ;
assign _0242_ = \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_4_U.u1.a  + \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_4_U.u1.b ;
assign { \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_4_U.u1.cout , \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_4_U.u1.s  } = _0242_ + \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_4_U.u1.cin ;
assign _0243_ = \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_4_U.u2.a  + \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_4_U.u2.b ;
assign { \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_4_U.u2.cout , \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_4_U.u2.s  } = _0243_ + \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_4_U.u2.cin ;
always @(posedge \add_9s_9ns_9_2_1_U3.top_add_9s_9ns_9_2_1_Adder_0_U.clk )
\add_9s_9ns_9_2_1_U3.top_add_9s_9ns_9_2_1_Adder_0_U.bin_s1  <= _0245_;
always @(posedge \add_9s_9ns_9_2_1_U3.top_add_9s_9ns_9_2_1_Adder_0_U.clk )
\add_9s_9ns_9_2_1_U3.top_add_9s_9ns_9_2_1_Adder_0_U.ain_s1  <= _0244_;
always @(posedge \add_9s_9ns_9_2_1_U3.top_add_9s_9ns_9_2_1_Adder_0_U.clk )
\add_9s_9ns_9_2_1_U3.top_add_9s_9ns_9_2_1_Adder_0_U.sum_s1  <= _0247_;
always @(posedge \add_9s_9ns_9_2_1_U3.top_add_9s_9ns_9_2_1_Adder_0_U.clk )
\add_9s_9ns_9_2_1_U3.top_add_9s_9ns_9_2_1_Adder_0_U.carry_s1  <= _0246_;
assign _0245_ = \add_9s_9ns_9_2_1_U3.top_add_9s_9ns_9_2_1_Adder_0_U.ce  ? \add_9s_9ns_9_2_1_U3.top_add_9s_9ns_9_2_1_Adder_0_U.b [8:4] : \add_9s_9ns_9_2_1_U3.top_add_9s_9ns_9_2_1_Adder_0_U.bin_s1 ;
assign _0244_ = \add_9s_9ns_9_2_1_U3.top_add_9s_9ns_9_2_1_Adder_0_U.ce  ? \add_9s_9ns_9_2_1_U3.top_add_9s_9ns_9_2_1_Adder_0_U.a [8:4] : \add_9s_9ns_9_2_1_U3.top_add_9s_9ns_9_2_1_Adder_0_U.ain_s1 ;
assign _0246_ = \add_9s_9ns_9_2_1_U3.top_add_9s_9ns_9_2_1_Adder_0_U.ce  ? \add_9s_9ns_9_2_1_U3.top_add_9s_9ns_9_2_1_Adder_0_U.facout_s1  : \add_9s_9ns_9_2_1_U3.top_add_9s_9ns_9_2_1_Adder_0_U.carry_s1 ;
assign _0247_ = \add_9s_9ns_9_2_1_U3.top_add_9s_9ns_9_2_1_Adder_0_U.ce  ? \add_9s_9ns_9_2_1_U3.top_add_9s_9ns_9_2_1_Adder_0_U.fas_s1  : \add_9s_9ns_9_2_1_U3.top_add_9s_9ns_9_2_1_Adder_0_U.sum_s1 ;
assign _0248_ = \add_9s_9ns_9_2_1_U3.top_add_9s_9ns_9_2_1_Adder_0_U.u1.a  + \add_9s_9ns_9_2_1_U3.top_add_9s_9ns_9_2_1_Adder_0_U.u1.b ;
assign { \add_9s_9ns_9_2_1_U3.top_add_9s_9ns_9_2_1_Adder_0_U.u1.cout , \add_9s_9ns_9_2_1_U3.top_add_9s_9ns_9_2_1_Adder_0_U.u1.s  } = _0248_ + \add_9s_9ns_9_2_1_U3.top_add_9s_9ns_9_2_1_Adder_0_U.u1.cin ;
assign _0249_ = \add_9s_9ns_9_2_1_U3.top_add_9s_9ns_9_2_1_Adder_0_U.u2.a  + \add_9s_9ns_9_2_1_U3.top_add_9s_9ns_9_2_1_Adder_0_U.u2.b ;
assign { \add_9s_9ns_9_2_1_U3.top_add_9s_9ns_9_2_1_Adder_0_U.u2.cout , \add_9s_9ns_9_2_1_U3.top_add_9s_9ns_9_2_1_Adder_0_U.u2.s  } = _0249_ + \add_9s_9ns_9_2_1_U3.top_add_9s_9ns_9_2_1_Adder_0_U.u2.cin ;
always @(posedge \add_9s_9s_9_2_1_U23.top_add_9s_9s_9_2_1_Adder_18_U.clk )
\add_9s_9s_9_2_1_U23.top_add_9s_9s_9_2_1_Adder_18_U.bin_s1  <= _0251_;
always @(posedge \add_9s_9s_9_2_1_U23.top_add_9s_9s_9_2_1_Adder_18_U.clk )
\add_9s_9s_9_2_1_U23.top_add_9s_9s_9_2_1_Adder_18_U.ain_s1  <= _0250_;
always @(posedge \add_9s_9s_9_2_1_U23.top_add_9s_9s_9_2_1_Adder_18_U.clk )
\add_9s_9s_9_2_1_U23.top_add_9s_9s_9_2_1_Adder_18_U.sum_s1  <= _0253_;
always @(posedge \add_9s_9s_9_2_1_U23.top_add_9s_9s_9_2_1_Adder_18_U.clk )
\add_9s_9s_9_2_1_U23.top_add_9s_9s_9_2_1_Adder_18_U.carry_s1  <= _0252_;
assign _0251_ = \add_9s_9s_9_2_1_U23.top_add_9s_9s_9_2_1_Adder_18_U.ce  ? \add_9s_9s_9_2_1_U23.top_add_9s_9s_9_2_1_Adder_18_U.b [8:4] : \add_9s_9s_9_2_1_U23.top_add_9s_9s_9_2_1_Adder_18_U.bin_s1 ;
assign _0250_ = \add_9s_9s_9_2_1_U23.top_add_9s_9s_9_2_1_Adder_18_U.ce  ? \add_9s_9s_9_2_1_U23.top_add_9s_9s_9_2_1_Adder_18_U.a [8:4] : \add_9s_9s_9_2_1_U23.top_add_9s_9s_9_2_1_Adder_18_U.ain_s1 ;
assign _0252_ = \add_9s_9s_9_2_1_U23.top_add_9s_9s_9_2_1_Adder_18_U.ce  ? \add_9s_9s_9_2_1_U23.top_add_9s_9s_9_2_1_Adder_18_U.facout_s1  : \add_9s_9s_9_2_1_U23.top_add_9s_9s_9_2_1_Adder_18_U.carry_s1 ;
assign _0253_ = \add_9s_9s_9_2_1_U23.top_add_9s_9s_9_2_1_Adder_18_U.ce  ? \add_9s_9s_9_2_1_U23.top_add_9s_9s_9_2_1_Adder_18_U.fas_s1  : \add_9s_9s_9_2_1_U23.top_add_9s_9s_9_2_1_Adder_18_U.sum_s1 ;
assign _0254_ = \add_9s_9s_9_2_1_U23.top_add_9s_9s_9_2_1_Adder_18_U.u1.a  + \add_9s_9s_9_2_1_U23.top_add_9s_9s_9_2_1_Adder_18_U.u1.b ;
assign { \add_9s_9s_9_2_1_U23.top_add_9s_9s_9_2_1_Adder_18_U.u1.cout , \add_9s_9s_9_2_1_U23.top_add_9s_9s_9_2_1_Adder_18_U.u1.s  } = _0254_ + \add_9s_9s_9_2_1_U23.top_add_9s_9s_9_2_1_Adder_18_U.u1.cin ;
assign _0255_ = \add_9s_9s_9_2_1_U23.top_add_9s_9s_9_2_1_Adder_18_U.u2.a  + \add_9s_9s_9_2_1_U23.top_add_9s_9s_9_2_1_Adder_18_U.u2.b ;
assign { \add_9s_9s_9_2_1_U23.top_add_9s_9s_9_2_1_Adder_18_U.u2.cout , \add_9s_9s_9_2_1_U23.top_add_9s_9s_9_2_1_Adder_18_U.u2.s  } = _0255_ + \add_9s_9s_9_2_1_U23.top_add_9s_9s_9_2_1_Adder_18_U.u2.cin ;
assign \mul_4s_4s_4_7_1_U1.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.tmp_product  = $signed(\mul_4s_4s_4_7_1_U1.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.a_reg0 ) * $signed(\mul_4s_4s_4_7_1_U1.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.b_reg0 );
always @(posedge \mul_4s_4s_4_7_1_U1.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.clk )
\mul_4s_4s_4_7_1_U1.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.a_reg0  <= _0256_;
always @(posedge \mul_4s_4s_4_7_1_U1.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.clk )
\mul_4s_4s_4_7_1_U1.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.b_reg0  <= _0257_;
always @(posedge \mul_4s_4s_4_7_1_U1.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.clk )
\mul_4s_4s_4_7_1_U1.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.buff0  <= _0258_;
always @(posedge \mul_4s_4s_4_7_1_U1.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.clk )
\mul_4s_4s_4_7_1_U1.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.buff1  <= _0259_;
always @(posedge \mul_4s_4s_4_7_1_U1.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.clk )
\mul_4s_4s_4_7_1_U1.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.buff2  <= _0260_;
always @(posedge \mul_4s_4s_4_7_1_U1.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.clk )
\mul_4s_4s_4_7_1_U1.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.buff3  <= _0261_;
always @(posedge \mul_4s_4s_4_7_1_U1.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.clk )
\mul_4s_4s_4_7_1_U1.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.buff4  <= _0262_;
assign _0262_ = \mul_4s_4s_4_7_1_U1.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.ce  ? \mul_4s_4s_4_7_1_U1.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.buff3  : \mul_4s_4s_4_7_1_U1.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.buff4 ;
assign _0261_ = \mul_4s_4s_4_7_1_U1.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.ce  ? \mul_4s_4s_4_7_1_U1.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.buff2  : \mul_4s_4s_4_7_1_U1.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.buff3 ;
assign _0260_ = \mul_4s_4s_4_7_1_U1.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.ce  ? \mul_4s_4s_4_7_1_U1.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.buff1  : \mul_4s_4s_4_7_1_U1.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.buff2 ;
assign _0259_ = \mul_4s_4s_4_7_1_U1.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.ce  ? \mul_4s_4s_4_7_1_U1.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.buff0  : \mul_4s_4s_4_7_1_U1.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.buff1 ;
assign _0258_ = \mul_4s_4s_4_7_1_U1.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.ce  ? \mul_4s_4s_4_7_1_U1.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.tmp_product  : \mul_4s_4s_4_7_1_U1.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.buff0 ;
assign _0257_ = \mul_4s_4s_4_7_1_U1.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.ce  ? \mul_4s_4s_4_7_1_U1.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.b  : \mul_4s_4s_4_7_1_U1.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.b_reg0 ;
assign _0256_ = \mul_4s_4s_4_7_1_U1.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.ce  ? \mul_4s_4s_4_7_1_U1.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.a  : \mul_4s_4s_4_7_1_U1.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.a_reg0 ;
assign \mul_4s_4s_8_7_1_U2.top_mul_4s_4s_8_7_1_Mul_DSP_1_U.tmp_product  = $signed(\mul_4s_4s_8_7_1_U2.top_mul_4s_4s_8_7_1_Mul_DSP_1_U.a_reg0 ) * $signed(\mul_4s_4s_8_7_1_U2.top_mul_4s_4s_8_7_1_Mul_DSP_1_U.b_reg0 );
always @(posedge \mul_4s_4s_8_7_1_U2.top_mul_4s_4s_8_7_1_Mul_DSP_1_U.clk )
\mul_4s_4s_8_7_1_U2.top_mul_4s_4s_8_7_1_Mul_DSP_1_U.a_reg0  <= _0263_;
always @(posedge \mul_4s_4s_8_7_1_U2.top_mul_4s_4s_8_7_1_Mul_DSP_1_U.clk )
\mul_4s_4s_8_7_1_U2.top_mul_4s_4s_8_7_1_Mul_DSP_1_U.b_reg0  <= _0264_;
always @(posedge \mul_4s_4s_8_7_1_U2.top_mul_4s_4s_8_7_1_Mul_DSP_1_U.clk )
\mul_4s_4s_8_7_1_U2.top_mul_4s_4s_8_7_1_Mul_DSP_1_U.buff0  <= _0265_;
always @(posedge \mul_4s_4s_8_7_1_U2.top_mul_4s_4s_8_7_1_Mul_DSP_1_U.clk )
\mul_4s_4s_8_7_1_U2.top_mul_4s_4s_8_7_1_Mul_DSP_1_U.buff1  <= _0266_;
always @(posedge \mul_4s_4s_8_7_1_U2.top_mul_4s_4s_8_7_1_Mul_DSP_1_U.clk )
\mul_4s_4s_8_7_1_U2.top_mul_4s_4s_8_7_1_Mul_DSP_1_U.buff2  <= _0267_;
always @(posedge \mul_4s_4s_8_7_1_U2.top_mul_4s_4s_8_7_1_Mul_DSP_1_U.clk )
\mul_4s_4s_8_7_1_U2.top_mul_4s_4s_8_7_1_Mul_DSP_1_U.buff3  <= _0268_;
always @(posedge \mul_4s_4s_8_7_1_U2.top_mul_4s_4s_8_7_1_Mul_DSP_1_U.clk )
\mul_4s_4s_8_7_1_U2.top_mul_4s_4s_8_7_1_Mul_DSP_1_U.buff4  <= _0269_;
assign _0269_ = \mul_4s_4s_8_7_1_U2.top_mul_4s_4s_8_7_1_Mul_DSP_1_U.ce  ? \mul_4s_4s_8_7_1_U2.top_mul_4s_4s_8_7_1_Mul_DSP_1_U.buff3  : \mul_4s_4s_8_7_1_U2.top_mul_4s_4s_8_7_1_Mul_DSP_1_U.buff4 ;
assign _0268_ = \mul_4s_4s_8_7_1_U2.top_mul_4s_4s_8_7_1_Mul_DSP_1_U.ce  ? \mul_4s_4s_8_7_1_U2.top_mul_4s_4s_8_7_1_Mul_DSP_1_U.buff2  : \mul_4s_4s_8_7_1_U2.top_mul_4s_4s_8_7_1_Mul_DSP_1_U.buff3 ;
assign _0267_ = \mul_4s_4s_8_7_1_U2.top_mul_4s_4s_8_7_1_Mul_DSP_1_U.ce  ? \mul_4s_4s_8_7_1_U2.top_mul_4s_4s_8_7_1_Mul_DSP_1_U.buff1  : \mul_4s_4s_8_7_1_U2.top_mul_4s_4s_8_7_1_Mul_DSP_1_U.buff2 ;
assign _0266_ = \mul_4s_4s_8_7_1_U2.top_mul_4s_4s_8_7_1_Mul_DSP_1_U.ce  ? \mul_4s_4s_8_7_1_U2.top_mul_4s_4s_8_7_1_Mul_DSP_1_U.buff0  : \mul_4s_4s_8_7_1_U2.top_mul_4s_4s_8_7_1_Mul_DSP_1_U.buff1 ;
assign _0265_ = \mul_4s_4s_8_7_1_U2.top_mul_4s_4s_8_7_1_Mul_DSP_1_U.ce  ? \mul_4s_4s_8_7_1_U2.top_mul_4s_4s_8_7_1_Mul_DSP_1_U.tmp_product  : \mul_4s_4s_8_7_1_U2.top_mul_4s_4s_8_7_1_Mul_DSP_1_U.buff0 ;
assign _0264_ = \mul_4s_4s_8_7_1_U2.top_mul_4s_4s_8_7_1_Mul_DSP_1_U.ce  ? \mul_4s_4s_8_7_1_U2.top_mul_4s_4s_8_7_1_Mul_DSP_1_U.b  : \mul_4s_4s_8_7_1_U2.top_mul_4s_4s_8_7_1_Mul_DSP_1_U.b_reg0 ;
assign _0263_ = \mul_4s_4s_8_7_1_U2.top_mul_4s_4s_8_7_1_Mul_DSP_1_U.ce  ? \mul_4s_4s_8_7_1_U2.top_mul_4s_4s_8_7_1_Mul_DSP_1_U.a  : \mul_4s_4s_8_7_1_U2.top_mul_4s_4s_8_7_1_Mul_DSP_1_U.a_reg0 ;
assign \sub_11ns_11s_11_2_1_U9.top_sub_11ns_11s_11_2_1_Adder_6_U.bin_s0  = ~ \sub_11ns_11s_11_2_1_U9.top_sub_11ns_11s_11_2_1_Adder_6_U.b ;
always @(posedge \sub_11ns_11s_11_2_1_U9.top_sub_11ns_11s_11_2_1_Adder_6_U.clk )
\sub_11ns_11s_11_2_1_U9.top_sub_11ns_11s_11_2_1_Adder_6_U.bin_s1  <= _0271_;
always @(posedge \sub_11ns_11s_11_2_1_U9.top_sub_11ns_11s_11_2_1_Adder_6_U.clk )
\sub_11ns_11s_11_2_1_U9.top_sub_11ns_11s_11_2_1_Adder_6_U.ain_s1  <= _0270_;
always @(posedge \sub_11ns_11s_11_2_1_U9.top_sub_11ns_11s_11_2_1_Adder_6_U.clk )
\sub_11ns_11s_11_2_1_U9.top_sub_11ns_11s_11_2_1_Adder_6_U.sum_s1  <= _0273_;
always @(posedge \sub_11ns_11s_11_2_1_U9.top_sub_11ns_11s_11_2_1_Adder_6_U.clk )
\sub_11ns_11s_11_2_1_U9.top_sub_11ns_11s_11_2_1_Adder_6_U.carry_s1  <= _0272_;
assign _0271_ = \sub_11ns_11s_11_2_1_U9.top_sub_11ns_11s_11_2_1_Adder_6_U.ce  ? \sub_11ns_11s_11_2_1_U9.top_sub_11ns_11s_11_2_1_Adder_6_U.bin_s0 [10:5] : \sub_11ns_11s_11_2_1_U9.top_sub_11ns_11s_11_2_1_Adder_6_U.bin_s1 ;
assign _0270_ = \sub_11ns_11s_11_2_1_U9.top_sub_11ns_11s_11_2_1_Adder_6_U.ce  ? \sub_11ns_11s_11_2_1_U9.top_sub_11ns_11s_11_2_1_Adder_6_U.a [10:5] : \sub_11ns_11s_11_2_1_U9.top_sub_11ns_11s_11_2_1_Adder_6_U.ain_s1 ;
assign _0272_ = \sub_11ns_11s_11_2_1_U9.top_sub_11ns_11s_11_2_1_Adder_6_U.ce  ? \sub_11ns_11s_11_2_1_U9.top_sub_11ns_11s_11_2_1_Adder_6_U.facout_s1  : \sub_11ns_11s_11_2_1_U9.top_sub_11ns_11s_11_2_1_Adder_6_U.carry_s1 ;
assign _0273_ = \sub_11ns_11s_11_2_1_U9.top_sub_11ns_11s_11_2_1_Adder_6_U.ce  ? \sub_11ns_11s_11_2_1_U9.top_sub_11ns_11s_11_2_1_Adder_6_U.fas_s1  : \sub_11ns_11s_11_2_1_U9.top_sub_11ns_11s_11_2_1_Adder_6_U.sum_s1 ;
assign _0274_ = \sub_11ns_11s_11_2_1_U9.top_sub_11ns_11s_11_2_1_Adder_6_U.u1.a  + \sub_11ns_11s_11_2_1_U9.top_sub_11ns_11s_11_2_1_Adder_6_U.u1.b ;
assign { \sub_11ns_11s_11_2_1_U9.top_sub_11ns_11s_11_2_1_Adder_6_U.u1.cout , \sub_11ns_11s_11_2_1_U9.top_sub_11ns_11s_11_2_1_Adder_6_U.u1.s  } = _0274_ + \sub_11ns_11s_11_2_1_U9.top_sub_11ns_11s_11_2_1_Adder_6_U.u1.cin ;
assign _0275_ = \sub_11ns_11s_11_2_1_U9.top_sub_11ns_11s_11_2_1_Adder_6_U.u2.a  + \sub_11ns_11s_11_2_1_U9.top_sub_11ns_11s_11_2_1_Adder_6_U.u2.b ;
assign { \sub_11ns_11s_11_2_1_U9.top_sub_11ns_11s_11_2_1_Adder_6_U.u2.cout , \sub_11ns_11s_11_2_1_U9.top_sub_11ns_11s_11_2_1_Adder_6_U.u2.s  } = _0275_ + \sub_11ns_11s_11_2_1_U9.top_sub_11ns_11s_11_2_1_Adder_6_U.u2.cin ;
assign \sub_9s_9s_9_2_1_U10.top_sub_9s_9s_9_2_1_Adder_7_U.bin_s0  = ~ \sub_9s_9s_9_2_1_U10.top_sub_9s_9s_9_2_1_Adder_7_U.b ;
always @(posedge \sub_9s_9s_9_2_1_U10.top_sub_9s_9s_9_2_1_Adder_7_U.clk )
\sub_9s_9s_9_2_1_U10.top_sub_9s_9s_9_2_1_Adder_7_U.bin_s1  <= _0277_;
always @(posedge \sub_9s_9s_9_2_1_U10.top_sub_9s_9s_9_2_1_Adder_7_U.clk )
\sub_9s_9s_9_2_1_U10.top_sub_9s_9s_9_2_1_Adder_7_U.ain_s1  <= _0276_;
always @(posedge \sub_9s_9s_9_2_1_U10.top_sub_9s_9s_9_2_1_Adder_7_U.clk )
\sub_9s_9s_9_2_1_U10.top_sub_9s_9s_9_2_1_Adder_7_U.sum_s1  <= _0279_;
always @(posedge \sub_9s_9s_9_2_1_U10.top_sub_9s_9s_9_2_1_Adder_7_U.clk )
\sub_9s_9s_9_2_1_U10.top_sub_9s_9s_9_2_1_Adder_7_U.carry_s1  <= _0278_;
assign _0277_ = \sub_9s_9s_9_2_1_U10.top_sub_9s_9s_9_2_1_Adder_7_U.ce  ? \sub_9s_9s_9_2_1_U10.top_sub_9s_9s_9_2_1_Adder_7_U.bin_s0 [8:4] : \sub_9s_9s_9_2_1_U10.top_sub_9s_9s_9_2_1_Adder_7_U.bin_s1 ;
assign _0276_ = \sub_9s_9s_9_2_1_U10.top_sub_9s_9s_9_2_1_Adder_7_U.ce  ? \sub_9s_9s_9_2_1_U10.top_sub_9s_9s_9_2_1_Adder_7_U.a [8:4] : \sub_9s_9s_9_2_1_U10.top_sub_9s_9s_9_2_1_Adder_7_U.ain_s1 ;
assign _0278_ = \sub_9s_9s_9_2_1_U10.top_sub_9s_9s_9_2_1_Adder_7_U.ce  ? \sub_9s_9s_9_2_1_U10.top_sub_9s_9s_9_2_1_Adder_7_U.facout_s1  : \sub_9s_9s_9_2_1_U10.top_sub_9s_9s_9_2_1_Adder_7_U.carry_s1 ;
assign _0279_ = \sub_9s_9s_9_2_1_U10.top_sub_9s_9s_9_2_1_Adder_7_U.ce  ? \sub_9s_9s_9_2_1_U10.top_sub_9s_9s_9_2_1_Adder_7_U.fas_s1  : \sub_9s_9s_9_2_1_U10.top_sub_9s_9s_9_2_1_Adder_7_U.sum_s1 ;
assign _0280_ = \sub_9s_9s_9_2_1_U10.top_sub_9s_9s_9_2_1_Adder_7_U.u1.a  + \sub_9s_9s_9_2_1_U10.top_sub_9s_9s_9_2_1_Adder_7_U.u1.b ;
assign { \sub_9s_9s_9_2_1_U10.top_sub_9s_9s_9_2_1_Adder_7_U.u1.cout , \sub_9s_9s_9_2_1_U10.top_sub_9s_9s_9_2_1_Adder_7_U.u1.s  } = _0280_ + \sub_9s_9s_9_2_1_U10.top_sub_9s_9s_9_2_1_Adder_7_U.u1.cin ;
assign _0281_ = \sub_9s_9s_9_2_1_U10.top_sub_9s_9s_9_2_1_Adder_7_U.u2.a  + \sub_9s_9s_9_2_1_U10.top_sub_9s_9s_9_2_1_Adder_7_U.u2.b ;
assign { \sub_9s_9s_9_2_1_U10.top_sub_9s_9s_9_2_1_Adder_7_U.u2.cout , \sub_9s_9s_9_2_1_U10.top_sub_9s_9s_9_2_1_Adder_7_U.u2.s  } = _0281_ + \sub_9s_9s_9_2_1_U10.top_sub_9s_9s_9_2_1_Adder_7_U.u2.cin ;
assign _0282_ = | op_6[21:0];
assign _0283_ = | p_Result_8_reg_1726;
assign _0284_ = | { tmp_reg_1832, 2'h0, p_Result_s_reg_1838 };
assign _0285_ = p_Result_s_reg_1838 != 5'h1f;
assign _0286_ = p_Result_8_reg_1726 != 8'hff;
assign _0287_ = | trunc_ln851_3_reg_2352;
assign _0288_ = | trunc_ln718_1_reg_2127;
assign _0289_ = | op_6[15:0];
assign op_4_V_fu_301_p2 = op_1[7:0] | { op_2[3], op_2[3], op_2[3], op_2[3], op_2 };
assign or_ln340_1_fu_983_p2 = or_ln340_reg_2001 | and_ln786_reg_1982;
assign or_ln340_2_fu_1008_p2 = and_ln785_2_fu_994_p2 | and_ln340_fu_1003_p2;
assign or_ln340_3_fu_1268_p2 = overflow_2_fu_1262_p2 | and_ln786_1_reg_2228;
assign or_ln340_4_fu_1344_p2 = or_ln340_3_reg_2259 | neg_src_7_fu_1339_p2;
assign or_ln340_fu_796_p2 = overflow_1_fu_791_p2 | neg_src_fu_776_p2;
assign or_ln384_1_fu_874_p2 = underflow_3_fu_869_p2 | overflow_3_reg_1995;
assign or_ln384_2_fu_1550_p2 = underflow_4_fu_1545_p2 | overflow_4_reg_2357;
assign or_ln384_fu_659_p2 = underflow_fu_654_p2 | overflow_reg_1910;
assign or_ln412_fu_682_p2 = r_reg_1806 | add_ln1192_2_reg_1932[17];
assign or_ln731_fu_317_p2 = op_2[0] | op_1[0];
assign or_ln760_fu_329_p2 = $signed(op_1[3:0]) | $signed(op_2);
assign or_ln785_1_fu_1252_p2 = xor_ln785_3_fu_1247_p2 | p_Result_37_reg_2033;
assign or_ln785_2_fu_751_p2 = p_Result_39_reg_1698 | icmp_ln768_reg_1732;
assign or_ln785_3_fu_1481_p2 = xor_ln785_6_fu_1475_p2 | p_Result_43_reg_2299;
assign or_ln785_4_fu_806_p2 = p_Result_30_reg_1755 | and_ln785_fu_802_p2;
assign or_ln785_5_fu_1377_p2 = p_Result_34_reg_2080 | and_ln785_4_fu_1373_p2;
assign or_ln785_fu_786_p2 = xor_ln785_1_fu_781_p2 | p_Result_32_reg_1893;
assign or_ln786_1_fu_1534_p2 = and_ln786_3_reg_2363 | and_ln781_2_fu_1530_p2;
assign or_ln786_fu_864_p2 = xor_ln786_fu_859_p2 | icmp_ln786_2_reg_1737;
assign or_ln788_1_fu_649_p2 = or_ln788_fu_645_p2 | icmp_ln786_reg_1916;
assign or_ln788_fu_645_p2 = icmp_ln790_reg_1879 | icmp_ln786_1_reg_1874;
assign ret_V_22_fu_1119_p2 = $signed(rhs_3_reg_2060) | $signed(op_6);
always @(posedge ap_clk)
rhs_3_reg_2060[21:0] <= 22'h000000;
always @(posedge ap_clk)
select_ln340_reg_2065 <= _0100_;
always @(posedge ap_clk)
ret_V_24_reg_2413 <= _0090_;
always @(posedge ap_clk)
ret_V_25_reg_2438 <= _0091_;
always @(posedge ap_clk)
ret_V_20_cast_reg_2443 <= _0085_;
always @(posedge ap_clk)
select_ln340_1_reg_2289 <= _0099_;
always @(posedge ap_clk)
p_Val2_13_reg_2294 <= _0073_;
always @(posedge ap_clk)
p_Result_43_reg_2299 <= _0067_;
always @(posedge ap_clk)
sext_ln850_reg_2306 <= _0102_;
always @(posedge ap_clk)
p_Result_38_reg_1720 <= _0063_;
always @(posedge ap_clk)
p_Result_8_reg_1726 <= _0070_;
always @(posedge ap_clk)
sel_tmp11_reg_2070 <= _0098_;
always @(posedge ap_clk)
p_Result_34_reg_2080 <= _0060_;
always @(posedge ap_clk)
xor_ln416_1_reg_2087 <= _0114_;
always @(posedge ap_clk)
p_Result_5_reg_2093 <= _0068_;
always @(posedge ap_clk)
p_Result_6_reg_2098 <= _0069_;
always @(posedge ap_clk)
ret_V_17_reg_2104 <= _0082_;
always @(posedge ap_clk)
p_Result_40_reg_2111 <= _0065_;
always @(posedge ap_clk)
p_Val2_12_reg_2117 <= _0072_;
always @(posedge ap_clk)
p_Result_41_reg_2122 <= _0066_;
always @(posedge ap_clk)
trunc_ln718_1_reg_2127 <= _0109_;
always @(posedge ap_clk)
p_Result_2_reg_2132 <= _0055_;
always @(posedge ap_clk)
ret_V_20_reg_2138 <= _0086_;
always @(posedge ap_clk)
ret_V_reg_2143 <= _0095_;
always @(posedge ap_clk)
trunc_ln851_1_reg_2150 <= _0111_;
always @(posedge ap_clk)
ret_V_22_reg_2155 <= _0088_;
always @(posedge ap_clk)
ret_V_7_cast_reg_2160 <= _0093_;
always @(posedge ap_clk)
trunc_ln851_2_reg_2167 <= _0112_;
always @(posedge ap_clk)
or_ln384_2_reg_2383 <= _0049_;
always @(posedge ap_clk)
or_ln340_3_reg_2259 <= _0047_;
always @(posedge ap_clk)
ret_V_18_reg_2269 <= _0083_;
always @(posedge ap_clk)
tmp_5_reg_2274 <= _0103_;
always @(posedge ap_clk)
ret_V_21_reg_2279 <= _0087_;
always @(posedge ap_clk)
ret_V_23_reg_2284 <= _0089_;
always @(posedge ap_clk)
op_3_V_reg_1816 <= _0044_;
always @(posedge ap_clk)
ret_reg_1821 <= _0096_;
always @(posedge ap_clk)
p_Result_29_reg_1826 <= _0054_;
always @(posedge ap_clk)
tmp_reg_1832 <= _0104_;
always @(posedge ap_clk)
p_Result_s_reg_1838 <= _0071_;
always @(posedge ap_clk)
trunc_ln790_reg_1844 <= _0110_;
always @(posedge ap_clk)
trunc_ln703_reg_1854 <= _0108_;
always @(posedge ap_clk)
trunc_ln1192_reg_1859 <= _0107_;
always @(posedge ap_clk)
trunc_ln1192_3_reg_1864 <= _0106_;
always @(posedge ap_clk)
op_25_V_reg_2423 <= _0043_;
always @(posedge ap_clk)
op_4_V_reg_1693 <= _0045_;
always @(posedge ap_clk)
p_Result_39_reg_1698 <= _0064_;
always @(posedge ap_clk)
op_16_V_reg_1705 <= _0040_;
always @(posedge ap_clk)
op_15_V_reg_2393 <= _0039_;
always @(posedge ap_clk)
op_23_V_reg_2398 <= _0042_;
always @(posedge ap_clk)
icmp_ln785_reg_1869 <= _0030_;
always @(posedge ap_clk)
icmp_ln786_1_reg_1874 <= _0031_;
always @(posedge ap_clk)
icmp_ln790_reg_1879 <= _0034_;
always @(posedge ap_clk)
p_Val2_3_reg_1884 <= _0075_;
always @(posedge ap_clk)
p_Result_32_reg_1893 <= _0058_;
always @(posedge ap_clk)
icmp_ln768_reg_1732 <= _0029_;
always @(posedge ap_clk)
icmp_ln786_2_reg_1737 <= _0032_;
always @(posedge ap_clk)
op_8_V_reg_1964 <= _0046_;
always @(posedge ap_clk)
deleted_zeros_reg_1970 <= _0026_;
always @(posedge ap_clk)
xor_ln785_2_reg_1976 <= _0116_;
always @(posedge ap_clk)
and_ln786_reg_1982 <= _0020_;
always @(posedge ap_clk)
overflow_3_reg_1995 <= _0051_;
always @(posedge ap_clk)
or_ln340_reg_2001 <= _0048_;
always @(posedge ap_clk)
and_ln785_1_reg_2007 <= _0017_;
always @(posedge ap_clk)
select_ln703_reg_2012 <= _0101_;
always @(posedge ap_clk)
p_Val2_8_reg_2027 <= _0077_;
always @(posedge ap_clk)
p_Result_37_reg_2033 <= _0062_;
always @(posedge ap_clk)
rhs_3_reg_2060[23:22] <= _0097_;
always @(posedge ap_clk)
and_ln414_reg_1811 <= _0016_;
always @(posedge ap_clk)
or_ln384_reg_1947 <= _0050_;
always @(posedge ap_clk)
carry_1_reg_1952 <= _0022_;
always @(posedge ap_clk)
and_ln412_reg_1959 <= _0015_;
always @(posedge ap_clk)
deleted_zeros_1_reg_2222 <= _0025_;
always @(posedge ap_clk)
and_ln786_1_reg_2228 <= _0018_;
always @(posedge ap_clk)
and_ln408_reg_2234 <= _0014_;
always @(posedge ap_clk)
ret_V_7_reg_2249 <= _0094_;
always @(posedge ap_clk)
ret_V_10_reg_2254 <= _0080_;
always @(posedge ap_clk)
overflow_4_reg_2357 <= _0052_;
always @(posedge ap_clk)
and_ln786_3_reg_2363 <= _0019_;
always @(posedge ap_clk)
ret_V_19_reg_2368 <= _0084_;
always @(posedge ap_clk)
add_ln69_reg_2373 <= _0013_;
always @(posedge ap_clk)
icmp_ln851_2_reg_2378 <= _0036_;
always @(posedge ap_clk)
ret_V_26_reg_2465 <= _0092_;
always @(posedge ap_clk)
add_ln69_3_reg_2470 <= _0012_;
always @(posedge ap_clk)
add_ln691_3_reg_2455 <= _0010_;
always @(posedge ap_clk)
overflow_reg_1910 <= _0053_;
always @(posedge ap_clk)
icmp_ln786_reg_1916 <= _0033_;
always @(posedge ap_clk)
xor_ln416_reg_1921 <= _0115_;
always @(posedge ap_clk)
add_ln1192_1_reg_1927 <= _0008_;
always @(posedge ap_clk)
add_ln1192_2_reg_1932 <= _0009_;
always @(posedge ap_clk)
p_Val2_7_reg_1937 <= _0076_;
always @(posedge ap_clk)
p_Result_36_reg_1942 <= _0061_;
always @(posedge ap_clk)
empty_reg_1750 <= _0027_;
always @(posedge ap_clk)
p_Result_30_reg_1755 <= _0056_;
always @(posedge ap_clk)
p_Val2_2_reg_1763 <= _0074_;
always @(posedge ap_clk)
p_Result_31_reg_1768 <= _0057_;
always @(posedge ap_clk)
icmp_ln414_reg_1773 <= _0028_;
always @(posedge ap_clk)
p_Result_33_reg_1778 <= _0059_;
always @(posedge ap_clk)
Range2_all_ones_reg_1784 <= _0007_;
always @(posedge ap_clk)
Range1_all_ones_reg_1789 <= _0002_;
always @(posedge ap_clk)
Range1_all_zeros_reg_1796 <= _0005_;
always @(posedge ap_clk)
trunc_ln1192_2_reg_1801 <= _0105_;
always @(posedge ap_clk)
r_reg_1806 <= _0079_;
always @(posedge ap_clk)
op_17_V_reg_2313 <= _0041_;
always @(posedge ap_clk)
carry_5_reg_2318 <= _0024_;
always @(posedge ap_clk)
Range1_all_ones_2_reg_2325 <= _0001_;
always @(posedge ap_clk)
Range1_all_zeros_2_reg_2332 <= _0004_;
always @(posedge ap_clk)
add_ln691_reg_2337 <= _0011_;
always @(posedge ap_clk)
trunc_ln851_3_reg_2352 <= _0113_;
always @(posedge ap_clk)
op_12_V_reg_2172 <= _0038_;
always @(posedge ap_clk)
ret_V_15_reg_2178 <= _0081_;
always @(posedge ap_clk)
carry_3_reg_2183 <= _0023_;
always @(posedge ap_clk)
Range2_all_ones_1_reg_2190 <= _0006_;
always @(posedge ap_clk)
Range1_all_ones_1_reg_2195 <= _0000_;
always @(posedge ap_clk)
Range1_all_zeros_1_reg_2202 <= _0003_;
always @(posedge ap_clk)
r_1_reg_2207 <= _0078_;
always @(posedge ap_clk)
icmp_ln851_reg_2212 <= _0037_;
always @(posedge ap_clk)
icmp_ln851_1_reg_2217 <= _0035_;
always @(posedge ap_clk)
ap_CS_fsm <= _0021_;
assign _0117_ = _0121_ ? 2'h2 : 2'h1;
assign _0290_ = ap_CS_fsm == 1'h1;
function [31:0] _0841_;
input [31:0] a;
input [1023:0] b;
input [31:0] s;
case (s)
32'b00000000000000000000000000000001:
_0841_ = b[31:0];
32'b00000000000000000000000000000010:
_0841_ = b[63:32];
32'b00000000000000000000000000000100:
_0841_ = b[95:64];
32'b00000000000000000000000000001000:
_0841_ = b[127:96];
32'b00000000000000000000000000010000:
_0841_ = b[159:128];
32'b00000000000000000000000000100000:
_0841_ = b[191:160];
32'b00000000000000000000000001000000:
_0841_ = b[223:192];
32'b00000000000000000000000010000000:
_0841_ = b[255:224];
32'b00000000000000000000000100000000:
_0841_ = b[287:256];
32'b00000000000000000000001000000000:
_0841_ = b[319:288];
32'b00000000000000000000010000000000:
_0841_ = b[351:320];
32'b00000000000000000000100000000000:
_0841_ = b[383:352];
32'b00000000000000000001000000000000:
_0841_ = b[415:384];
32'b00000000000000000010000000000000:
_0841_ = b[447:416];
32'b00000000000000000100000000000000:
_0841_ = b[479:448];
32'b00000000000000001000000000000000:
_0841_ = b[511:480];
32'b00000000000000010000000000000000:
_0841_ = b[543:512];
32'b00000000000000100000000000000000:
_0841_ = b[575:544];
32'b00000000000001000000000000000000:
_0841_ = b[607:576];
32'b00000000000010000000000000000000:
_0841_ = b[639:608];
32'b00000000000100000000000000000000:
_0841_ = b[671:640];
32'b00000000001000000000000000000000:
_0841_ = b[703:672];
32'b00000000010000000000000000000000:
_0841_ = b[735:704];
32'b00000000100000000000000000000000:
_0841_ = b[767:736];
32'b00000001000000000000000000000000:
_0841_ = b[799:768];
32'b00000010000000000000000000000000:
_0841_ = b[831:800];
32'b00000100000000000000000000000000:
_0841_ = b[863:832];
32'b00001000000000000000000000000000:
_0841_ = b[895:864];
32'b00010000000000000000000000000000:
_0841_ = b[927:896];
32'b00100000000000000000000000000000:
_0841_ = b[959:928];
32'b01000000000000000000000000000000:
_0841_ = b[991:960];
32'b10000000000000000000000000000000:
_0841_ = b[1023:992];
32'b00000000000000000000000000000000:
_0841_ = a;
default:
_0841_ = 32'bx;
endcase
endfunction
assign ap_NS_fsm = _0841_(32'hxxxxxxxx, { 30'h00000000, _0117_, 992'h00000004000000080000001000000020000000400000008000000100000002000000040000000800000010000000200000004000000080000001000000020000000400000008000000100000002000000040000000800000010000000200000004000000080000001000000020000000400000008000000000000001 }, { _0290_, _0321_, _0320_, _0319_, _0318_, _0317_, _0316_, _0315_, _0314_, _0313_, _0312_, _0311_, _0310_, _0309_, _0308_, _0307_, _0306_, _0305_, _0304_, _0303_, _0302_, _0301_, _0300_, _0299_, _0298_, _0297_, _0296_, _0295_, _0294_, _0293_, _0292_, _0291_ });
assign _0291_ = ap_CS_fsm == 32'd2147483648;
assign _0292_ = ap_CS_fsm == 31'h40000000;
assign _0293_ = ap_CS_fsm == 30'h20000000;
assign _0294_ = ap_CS_fsm == 29'h10000000;
assign _0295_ = ap_CS_fsm == 28'h8000000;
assign _0296_ = ap_CS_fsm == 27'h4000000;
assign _0297_ = ap_CS_fsm == 26'h2000000;
assign _0298_ = ap_CS_fsm == 25'h1000000;
assign _0299_ = ap_CS_fsm == 24'h800000;
assign _0300_ = ap_CS_fsm == 23'h400000;
assign _0301_ = ap_CS_fsm == 22'h200000;
assign _0302_ = ap_CS_fsm == 21'h100000;
assign _0303_ = ap_CS_fsm == 20'h80000;
assign _0304_ = ap_CS_fsm == 19'h40000;
assign _0305_ = ap_CS_fsm == 18'h20000;
assign _0306_ = ap_CS_fsm == 17'h10000;
assign _0307_ = ap_CS_fsm == 16'h8000;
assign _0308_ = ap_CS_fsm == 15'h4000;
assign _0309_ = ap_CS_fsm == 14'h2000;
assign _0310_ = ap_CS_fsm == 13'h1000;
assign _0311_ = ap_CS_fsm == 12'h800;
assign _0312_ = ap_CS_fsm == 11'h400;
assign _0313_ = ap_CS_fsm == 10'h200;
assign _0314_ = ap_CS_fsm == 9'h100;
assign _0315_ = ap_CS_fsm == 8'h80;
assign _0316_ = ap_CS_fsm == 7'h40;
assign _0317_ = ap_CS_fsm == 6'h20;
assign _0318_ = ap_CS_fsm == 5'h10;
assign _0319_ = ap_CS_fsm == 4'h8;
assign _0320_ = ap_CS_fsm == 3'h4;
assign _0321_ = ap_CS_fsm == 2'h2;
assign op_28_ap_vld = ap_CS_fsm[31] ? 1'h1 : 1'h0;
assign ap_idle = _0120_ ? 1'h1 : 1'h0;
assign _0100_ = _0119_ ? select_ln340_fu_987_p3 : select_ln340_reg_2065;
assign _0090_ = ap_CS_fsm[22] ? grp_fu_1582_p2 : ret_V_24_reg_2413;
assign _0085_ = ap_CS_fsm[26] ? grp_fu_1610_p2[37:6] : ret_V_20_cast_reg_2443;
assign _0091_ = ap_CS_fsm[26] ? grp_fu_1610_p2 : ret_V_25_reg_2438;
assign _0102_ = ap_CS_fsm[16] ? { tmp_5_reg_2274[2], tmp_5_reg_2274 } : sext_ln850_reg_2306;
assign _0067_ = ap_CS_fsm[16] ? grp_fu_1276_p2[3] : p_Result_43_reg_2299;
assign _0073_ = ap_CS_fsm[16] ? grp_fu_1276_p2 : p_Val2_13_reg_2294;
assign _0099_ = ap_CS_fsm[16] ? select_ln340_1_fu_1349_p3 : select_ln340_1_reg_2289;
assign _0070_ = ap_CS_fsm[2] ? grp_fu_347_p2[8:1] : p_Result_8_reg_1726;
assign _0063_ = ap_CS_fsm[2] ? grp_fu_347_p2[8] : p_Result_38_reg_1720;
assign _0112_ = ap_CS_fsm[12] ? ret_V_22_fu_1119_p2[22:0] : trunc_ln851_2_reg_2167;
assign _0093_ = ap_CS_fsm[12] ? ret_V_22_fu_1119_p2[26:23] : ret_V_7_cast_reg_2160;
assign _0088_ = ap_CS_fsm[12] ? ret_V_22_fu_1119_p2 : ret_V_22_reg_2155;
assign _0111_ = ap_CS_fsm[12] ? grp_fu_914_p2[4:0] : trunc_ln851_1_reg_2150;
assign _0095_ = ap_CS_fsm[12] ? grp_fu_914_p2[8:5] : ret_V_reg_2143;
assign _0086_ = ap_CS_fsm[12] ? grp_fu_914_p2 : ret_V_20_reg_2138;
assign _0055_ = ap_CS_fsm[12] ? grp_fu_894_p2[10:9] : p_Result_2_reg_2132;
assign _0109_ = ap_CS_fsm[12] ? grp_fu_894_p2[3:0] : trunc_ln718_1_reg_2127;
assign _0066_ = ap_CS_fsm[12] ? grp_fu_894_p2[4] : p_Result_41_reg_2122;
assign _0072_ = ap_CS_fsm[12] ? grp_fu_894_p2[8:5] : p_Val2_12_reg_2117;
assign _0065_ = ap_CS_fsm[12] ? grp_fu_894_p2[10] : p_Result_40_reg_2111;
assign _0082_ = ap_CS_fsm[12] ? grp_fu_894_p2 : ret_V_17_reg_2104;
assign _0069_ = ap_CS_fsm[12] ? grp_fu_838_p2[32:25] : p_Result_6_reg_2098;
assign _0068_ = ap_CS_fsm[12] ? grp_fu_838_p2[32:26] : p_Result_5_reg_2093;
assign _0114_ = ap_CS_fsm[12] ? xor_ln416_1_fu_1037_p2 : xor_ln416_1_reg_2087;
assign _0060_ = ap_CS_fsm[12] ? grp_fu_838_p2[32] : p_Result_34_reg_2080;
assign _0098_ = ap_CS_fsm[12] ? sel_tmp11_fu_1014_p2 : sel_tmp11_reg_2070;
assign _0049_ = ap_CS_fsm[19] ? or_ln384_2_fu_1550_p2 : or_ln384_2_reg_2383;
assign _0089_ = ap_CS_fsm[15] ? ret_V_23_fu_1322_p3 : ret_V_23_reg_2284;
assign _0087_ = ap_CS_fsm[15] ? ret_V_21_fu_1303_p3 : ret_V_21_reg_2279;
assign _0103_ = ap_CS_fsm[15] ? grp_fu_1241_p2[3:1] : tmp_5_reg_2274;
assign _0083_ = ap_CS_fsm[15] ? grp_fu_1241_p2 : ret_V_18_reg_2269;
assign _0047_ = ap_CS_fsm[15] ? or_ln340_3_fu_1268_p2 : or_ln340_3_reg_2259;
assign _0106_ = ap_CS_fsm[6] ? grp_fu_279_p2[2:0] : trunc_ln1192_3_reg_1864;
assign _0107_ = ap_CS_fsm[6] ? grp_fu_279_p2[1:0] : trunc_ln1192_reg_1859;
assign _0108_ = ap_CS_fsm[6] ? grp_fu_279_p2[0] : trunc_ln703_reg_1854;
assign _0110_ = ap_CS_fsm[6] ? grp_fu_307_p2[1:0] : trunc_ln790_reg_1844;
assign _0071_ = ap_CS_fsm[6] ? grp_fu_307_p2[7:3] : p_Result_s_reg_1838;
assign _0104_ = ap_CS_fsm[6] ? grp_fu_307_p2[2] : tmp_reg_1832;
assign _0054_ = ap_CS_fsm[6] ? grp_fu_307_p2[7] : p_Result_29_reg_1826;
assign _0096_ = ap_CS_fsm[6] ? grp_fu_307_p2 : ret_reg_1821;
assign _0044_ = ap_CS_fsm[6] ? grp_fu_279_p2 : op_3_V_reg_1816;
assign _0043_ = ap_CS_fsm[24] ? grp_fu_1591_p2 : op_25_V_reg_2423;
assign _0040_ = ap_CS_fsm[0] ? op_16_V_fu_335_p2 : op_16_V_reg_1705;
assign _0064_ = ap_CS_fsm[0] ? p_Result_39_fu_323_p2 : p_Result_39_reg_1698;
assign _0045_ = ap_CS_fsm[0] ? op_4_V_fu_301_p2 : op_4_V_reg_1693;
assign _0042_ = ap_CS_fsm[20] ? grp_fu_1558_p2 : op_23_V_reg_2398;
assign _0039_ = ap_CS_fsm[20] ? op_15_V_fu_1570_p3 : op_15_V_reg_2393;
assign _0058_ = ap_CS_fsm[7] ? grp_fu_518_p2[1] : p_Result_32_reg_1893;
assign _0075_ = ap_CS_fsm[7] ? grp_fu_518_p2 : p_Val2_3_reg_1884;
assign _0034_ = ap_CS_fsm[7] ? icmp_ln790_fu_561_p2 : icmp_ln790_reg_1879;
assign _0031_ = ap_CS_fsm[7] ? icmp_ln786_1_fu_549_p2 : icmp_ln786_1_reg_1874;
assign _0030_ = ap_CS_fsm[7] ? icmp_ln785_fu_543_p2 : icmp_ln785_reg_1869;
assign _0032_ = ap_CS_fsm[3] ? icmp_ln786_2_fu_376_p2 : icmp_ln786_2_reg_1737;
assign _0029_ = ap_CS_fsm[3] ? icmp_ln768_fu_371_p2 : icmp_ln768_reg_1732;
assign _0051_ = ap_CS_fsm[10] ? overflow_3_fu_760_p2 : overflow_3_reg_1995;
assign _0020_ = ap_CS_fsm[10] ? and_ln786_fu_738_p2 : and_ln786_reg_1982;
assign _0116_ = ap_CS_fsm[10] ? xor_ln785_2_fu_733_p2 : xor_ln785_2_reg_1976;
assign _0026_ = ap_CS_fsm[10] ? deleted_zeros_fu_712_p3 : deleted_zeros_reg_1970;
assign _0046_ = ap_CS_fsm[10] ? op_8_V_fu_705_p3 : op_8_V_reg_1964;
assign _0097_ = ap_CS_fsm[11] ? select_ln384_5_fu_927_p3 : rhs_3_reg_2060[23:22];
assign _0062_ = ap_CS_fsm[11] ? grp_fu_746_p2[7] : p_Result_37_reg_2033;
assign _0077_ = ap_CS_fsm[11] ? grp_fu_746_p2 : p_Val2_8_reg_2027;
assign _0101_ = ap_CS_fsm[11] ? select_ln703_fu_816_p3 : select_ln703_reg_2012;
assign _0017_ = ap_CS_fsm[11] ? and_ln785_1_fu_811_p2 : and_ln785_1_reg_2007;
assign _0048_ = ap_CS_fsm[11] ? or_ln340_fu_796_p2 : or_ln340_reg_2001;
assign _0016_ = ap_CS_fsm[5] ? and_ln414_fu_481_p2 : and_ln414_reg_1811;
assign _0015_ = ap_CS_fsm[9] ? and_ln412_fu_687_p2 : and_ln412_reg_1959;
assign _0022_ = ap_CS_fsm[9] ? carry_1_fu_664_p2 : carry_1_reg_1952;
assign _0050_ = ap_CS_fsm[9] ? or_ln384_fu_659_p2 : or_ln384_reg_1947;
assign _0080_ = ap_CS_fsm[14] ? grp_fu_1188_p2 : ret_V_10_reg_2254;
assign _0094_ = ap_CS_fsm[14] ? grp_fu_1178_p2 : ret_V_7_reg_2249;
assign _0014_ = ap_CS_fsm[14] ? and_ln408_fu_1227_p2 : and_ln408_reg_2234;
assign _0018_ = ap_CS_fsm[14] ? and_ln786_1_fu_1222_p2 : and_ln786_1_reg_2228;
assign _0025_ = ap_CS_fsm[14] ? deleted_zeros_1_fu_1193_p3 : deleted_zeros_1_reg_2222;
assign _0036_ = ap_CS_fsm[18] ? icmp_ln851_2_fu_1525_p2 : icmp_ln851_2_reg_2378;
assign _0013_ = ap_CS_fsm[18] ? grp_fu_1428_p2 : add_ln69_reg_2373;
assign _0084_ = ap_CS_fsm[18] ? ret_V_19_fu_1518_p3 : ret_V_19_reg_2368;
assign _0019_ = ap_CS_fsm[18] ? and_ln786_3_fu_1497_p2 : and_ln786_3_reg_2363;
assign _0052_ = ap_CS_fsm[18] ? overflow_4_fu_1491_p2 : overflow_4_reg_2357;
assign _0012_ = ap_CS_fsm[29] ? grp_fu_1638_p2 : add_ln69_3_reg_2470;
assign _0092_ = ap_CS_fsm[29] ? ret_V_26_fu_1656_p3 : ret_V_26_reg_2465;
assign _0010_ = _0118_ ? grp_fu_1626_p2 : add_ln691_3_reg_2455;
assign _0061_ = ap_CS_fsm[8] ? grp_fu_594_p2[24] : p_Result_36_reg_1942;
assign _0076_ = ap_CS_fsm[8] ? grp_fu_594_p2[24:17] : p_Val2_7_reg_1937;
assign _0009_ = ap_CS_fsm[8] ? grp_fu_594_p2 : add_ln1192_2_reg_1932;
assign _0008_ = ap_CS_fsm[8] ? grp_fu_589_p2 : add_ln1192_1_reg_1927;
assign _0115_ = ap_CS_fsm[8] ? xor_ln416_fu_622_p2 : xor_ln416_reg_1921;
assign _0033_ = ap_CS_fsm[8] ? icmp_ln786_fu_616_p2 : icmp_ln786_reg_1916;
assign _0053_ = ap_CS_fsm[8] ? overflow_fu_611_p2 : overflow_reg_1910;
assign _0079_ = ap_CS_fsm[4] ? r_fu_475_p2 : r_reg_1806;
assign _0105_ = ap_CS_fsm[4] ? op_6[25:0] : trunc_ln1192_2_reg_1801;
assign _0005_ = ap_CS_fsm[4] ? Range1_all_zeros_fu_461_p2 : Range1_all_zeros_reg_1796;
assign _0002_ = ap_CS_fsm[4] ? Range1_all_ones_fu_455_p2 : Range1_all_ones_reg_1789;
assign _0007_ = ap_CS_fsm[4] ? Range2_all_ones_fu_439_p2 : Range2_all_ones_reg_1784;
assign _0059_ = ap_CS_fsm[4] ? op_6[24] : p_Result_33_reg_1778;
assign _0028_ = ap_CS_fsm[4] ? icmp_ln414_fu_415_p2 : icmp_ln414_reg_1773;
assign _0057_ = ap_CS_fsm[4] ? op_6[23] : p_Result_31_reg_1768;
assign _0074_ = ap_CS_fsm[4] ? op_6[23:22] : p_Val2_2_reg_1763;
assign _0056_ = ap_CS_fsm[4] ? op_6[31] : p_Result_30_reg_1755;
assign _0027_ = ap_CS_fsm[4] ? op_6[24:0] : empty_reg_1750;
assign _0113_ = ap_CS_fsm[17] ? op_17_V_fu_1387_p3[5:0] : trunc_ln851_3_reg_2352;
assign _0011_ = ap_CS_fsm[17] ? grp_fu_1367_p2 : add_ln691_reg_2337;
assign _0004_ = ap_CS_fsm[17] ? Range1_all_zeros_2_fu_1416_p2 : Range1_all_zeros_2_reg_2332;
assign _0001_ = ap_CS_fsm[17] ? Range1_all_ones_2_fu_1411_p2 : Range1_all_ones_2_reg_2325;
assign _0024_ = ap_CS_fsm[17] ? carry_5_fu_1405_p2 : carry_5_reg_2318;
assign _0041_ = ap_CS_fsm[17] ? op_17_V_fu_1387_p3 : op_17_V_reg_2313;
assign _0035_ = ap_CS_fsm[13] ? icmp_ln851_1_fu_1183_p2 : icmp_ln851_1_reg_2217;
assign _0037_ = ap_CS_fsm[13] ? icmp_ln851_fu_1173_p2 : icmp_ln851_reg_2212;
assign _0078_ = ap_CS_fsm[13] ? r_1_fu_1168_p2 : r_1_reg_2207;
assign _0003_ = ap_CS_fsm[13] ? Range1_all_zeros_1_fu_1163_p2 : Range1_all_zeros_1_reg_2202;
assign _0000_ = ap_CS_fsm[13] ? Range1_all_ones_1_fu_1158_p2 : Range1_all_ones_1_reg_2195;
assign _0006_ = ap_CS_fsm[13] ? Range2_all_ones_1_fu_1153_p2 : Range2_all_ones_1_reg_2190;
assign _0023_ = ap_CS_fsm[13] ? carry_3_fu_1149_p2 : carry_3_reg_2183;
assign _0081_ = ap_CS_fsm[13] ? grp_fu_1024_p2 : ret_V_15_reg_2178;
assign _0038_ = ap_CS_fsm[13] ? op_12_V_fu_1143_p3 : op_12_V_reg_2172;
assign _0021_ = ap_rst ? 32'd1 : ap_NS_fsm;
assign Range1_all_ones_1_fu_1158_p2 = _0124_ ? 1'h1 : 1'h0;
assign Range1_all_ones_2_fu_1411_p2 = _0125_ ? 1'h1 : 1'h0;
assign Range1_all_ones_fu_455_p2 = _0126_ ? 1'h1 : 1'h0;
assign Range1_all_zeros_1_fu_1163_p2 = _0127_ ? 1'h1 : 1'h0;
assign Range1_all_zeros_2_fu_1416_p2 = _0128_ ? 1'h1 : 1'h0;
assign Range1_all_zeros_fu_461_p2 = _0129_ ? 1'h1 : 1'h0;
assign Range2_all_ones_1_fu_1153_p2 = _0130_ ? 1'h1 : 1'h0;
assign Range2_all_ones_fu_439_p2 = _0131_ ? 1'h1 : 1'h0;
assign deleted_ones_1_fu_1216_p3 = carry_3_reg_2183 ? and_ln780_1_fu_1211_p2 : Range1_all_ones_1_reg_2195;
assign deleted_ones_2_fu_1469_p3 = carry_5_reg_2318 ? and_ln780_2_fu_1463_p2 : Range1_all_ones_2_reg_2325;
assign deleted_ones_fu_727_p3 = carry_1_reg_1952 ? and_ln780_fu_722_p2 : Range1_all_ones_reg_1789;
assign deleted_zeros_1_fu_1193_p3 = carry_3_reg_2183 ? Range1_all_ones_1_reg_2195 : Range1_all_zeros_1_reg_2202;
assign deleted_zeros_2_fu_1445_p3 = carry_5_reg_2318 ? Range1_all_ones_2_reg_2325 : Range1_all_zeros_2_reg_2332;
assign deleted_zeros_fu_712_p3 = carry_1_reg_1952 ? Range1_all_ones_reg_1789 : Range1_all_zeros_reg_1796;
assign icmp_ln414_fu_415_p2 = _0282_ ? 1'h1 : 1'h0;
assign icmp_ln768_fu_371_p2 = _0283_ ? 1'h1 : 1'h0;
assign icmp_ln785_fu_543_p2 = _0284_ ? 1'h1 : 1'h0;
assign icmp_ln786_1_fu_549_p2 = _0285_ ? 1'h1 : 1'h0;
assign icmp_ln786_2_fu_376_p2 = _0286_ ? 1'h1 : 1'h0;
assign icmp_ln786_fu_616_p2 = _0132_ ? 1'h1 : 1'h0;
assign icmp_ln790_fu_561_p2 = _0133_ ? 1'h1 : 1'h0;
assign icmp_ln851_1_fu_1183_p2 = _0134_ ? 1'h1 : 1'h0;
assign icmp_ln851_2_fu_1525_p2 = _0287_ ? 1'h1 : 1'h0;
assign icmp_ln851_fu_1173_p2 = _0135_ ? 1'h1 : 1'h0;
assign op_12_V_fu_1143_p3 = sel_tmp11_reg_2070 ? p_Val2_3_reg_1884 : select_ln785_fu_1138_p3;
assign op_15_V_fu_1570_p3 = or_ln384_2_reg_2383 ? select_ln384_2_fu_1563_p3 : p_Val2_13_reg_2294;
assign op_17_V_fu_1387_p3 = and_ln785_5_fu_1382_p2 ? p_Val2_8_reg_2027 : select_ln340_1_reg_2289;
assign op_8_V_fu_705_p3 = or_ln384_reg_1947 ? select_ln384_fu_698_p3 : { ret_reg_1821[2:0], 5'h00 };
assign r_1_fu_1168_p2 = _0288_ ? 1'h1 : 1'h0;
assign r_fu_475_p2 = _0289_ ? 1'h1 : 1'h0;
assign ret_V_19_fu_1518_p3 = ret_V_18_reg_2269[3] ? select_ln850_fu_1512_p3 : sext_ln850_reg_2306;
assign ret_V_21_fu_1303_p3 = ret_V_20_reg_2138[8] ? select_ln850_1_fu_1298_p3 : ret_V_reg_2143;
assign ret_V_23_fu_1322_p3 = ret_V_22_reg_2155[31] ? select_ln850_2_fu_1317_p3 : ret_V_7_cast_reg_2160;
assign ret_V_26_fu_1656_p3 = ret_V_25_reg_2438[38] ? select_ln850_3_fu_1651_p3 : ret_V_20_cast_reg_2443;
assign select_ln340_1_fu_1349_p3 = or_ln340_4_fu_1344_p2 ? 8'h00 : p_Val2_8_reg_2027;
assign select_ln340_fu_987_p3 = or_ln340_1_fu_983_p2 ? { p_Result_33_reg_1778, p_Val2_4_fu_969_p2 } : p_Val2_3_reg_1884;
assign select_ln384_2_fu_1563_p3 = overflow_4_reg_2357 ? 4'h7 : 4'h8;
assign select_ln384_4_fu_920_p3 = overflow_3_reg_1995 ? 2'h1 : 2'h2;
assign select_ln384_5_fu_927_p3 = or_ln384_1_fu_874_p2 ? select_ln384_4_fu_920_p3 : { p_Result_39_reg_1698, 1'h0 };
assign select_ln384_fu_698_p3 = overflow_reg_1910 ? 8'h7f : 8'h81;
assign select_ln703_fu_816_p3 = op_0 ? 3'h7 : 3'h0;
assign select_ln785_fu_1138_p3 = and_ln785_1_reg_2007 ? p_Val2_3_reg_1884 : select_ln340_reg_2065;
assign select_ln850_1_fu_1298_p3 = icmp_ln851_reg_2212 ? ret_V_reg_2143 : ret_V_7_reg_2249;
assign select_ln850_2_fu_1317_p3 = icmp_ln851_1_reg_2217 ? ret_V_7_cast_reg_2160 : ret_V_10_reg_2254;
assign select_ln850_3_fu_1651_p3 = icmp_ln851_2_reg_2378 ? add_ln691_3_reg_2455 : ret_V_20_cast_reg_2443;
assign select_ln850_fu_1512_p3 = op_12_V_reg_2172[0] ? add_ln691_reg_2337 : sext_ln850_reg_2306;
assign p_Result_39_fu_323_p2 = op_5[0] ^ or_ln731_fu_317_p2;
assign xor_ln365_fu_957_p2 = p_Val2_3_reg_1884[1] ^ op_6[24];
assign Range2_all_ones_2_fu_1438_p3 = ret_V_17_reg_2104[10];
assign and_ln_fu_599_p3 = { tmp_reg_1832, 7'h00 };
assign ap_CS_fsm_state1 = ap_CS_fsm[0];
assign ap_CS_fsm_state10 = ap_CS_fsm[9];
assign ap_CS_fsm_state11 = ap_CS_fsm[10];
assign ap_CS_fsm_state12 = ap_CS_fsm[11];
assign ap_CS_fsm_state13 = ap_CS_fsm[12];
assign ap_CS_fsm_state14 = ap_CS_fsm[13];
assign ap_CS_fsm_state15 = ap_CS_fsm[14];
assign ap_CS_fsm_state16 = ap_CS_fsm[15];
assign ap_CS_fsm_state17 = ap_CS_fsm[16];
assign ap_CS_fsm_state18 = ap_CS_fsm[17];
assign ap_CS_fsm_state19 = ap_CS_fsm[18];
assign ap_CS_fsm_state2 = ap_CS_fsm[1];
assign ap_CS_fsm_state20 = ap_CS_fsm[19];
assign ap_CS_fsm_state21 = ap_CS_fsm[20];
assign ap_CS_fsm_state22 = ap_CS_fsm[21];
assign ap_CS_fsm_state23 = ap_CS_fsm[22];
assign ap_CS_fsm_state24 = ap_CS_fsm[23];
assign ap_CS_fsm_state25 = ap_CS_fsm[24];
assign ap_CS_fsm_state26 = ap_CS_fsm[25];
assign ap_CS_fsm_state27 = ap_CS_fsm[26];
assign ap_CS_fsm_state28 = ap_CS_fsm[27];
assign ap_CS_fsm_state29 = ap_CS_fsm[28];
assign ap_CS_fsm_state3 = ap_CS_fsm[2];
assign ap_CS_fsm_state30 = ap_CS_fsm[29];
assign ap_CS_fsm_state31 = ap_CS_fsm[30];
assign ap_CS_fsm_state32 = ap_CS_fsm[31];
assign ap_CS_fsm_state4 = ap_CS_fsm[3];
assign ap_CS_fsm_state5 = ap_CS_fsm[4];
assign ap_CS_fsm_state6 = ap_CS_fsm[5];
assign ap_CS_fsm_state7 = ap_CS_fsm[6];
assign ap_CS_fsm_state8 = ap_CS_fsm[7];
assign ap_CS_fsm_state9 = ap_CS_fsm[8];
assign ap_done = op_28_ap_vld;
assign ap_ready = op_28_ap_vld;
assign empty_fu_381_p0 = op_6;
assign empty_fu_381_p1 = op_6[24:0];
assign grp_fu_1024_p0 = { op_9[1], op_9 };
assign grp_fu_1241_p0 = { ret_V_15_reg_2178, 1'h0 };
assign grp_fu_1241_p1 = { op_12_V_reg_2172[1], op_12_V_reg_2172[1], op_12_V_reg_2172 };
assign grp_fu_1276_p1 = { 3'h0, and_ln408_reg_2234 };
assign grp_fu_1367_p0 = { tmp_5_reg_2274[2], tmp_5_reg_2274 };
assign grp_fu_1428_p0 = { ret_V_23_reg_2284[3], ret_V_23_reg_2284 };
assign grp_fu_1428_p1 = { op_13[1], op_13[1], op_13[1], op_13 };
assign grp_fu_1558_p1 = { ret_V_19_reg_2368[3], ret_V_19_reg_2368 };
assign grp_fu_1582_p0 = { op_23_V_reg_2398[4], op_23_V_reg_2398 };
assign grp_fu_1582_p1 = { op_15_V_reg_2393[3], op_15_V_reg_2393[3], op_15_V_reg_2393 };
assign grp_fu_1591_p1 = { op_16_V_reg_1705[3], op_16_V_reg_1705[3], op_16_V_reg_1705 };
assign grp_fu_1610_p0 = { op_25_V_reg_2423[5], op_25_V_reg_2423[5], op_25_V_reg_2423[5], op_25_V_reg_2423[5], op_25_V_reg_2423[5], op_25_V_reg_2423[5], op_25_V_reg_2423[5], op_25_V_reg_2423[5], op_25_V_reg_2423[5], op_25_V_reg_2423[5], op_25_V_reg_2423[5], op_25_V_reg_2423[5], op_25_V_reg_2423[5], op_25_V_reg_2423[5], op_25_V_reg_2423[5], op_25_V_reg_2423[5], op_25_V_reg_2423[5], op_25_V_reg_2423[5], op_25_V_reg_2423[5], op_25_V_reg_2423[5], op_25_V_reg_2423[5], op_25_V_reg_2423[5], op_25_V_reg_2423[5], op_25_V_reg_2423[5], op_25_V_reg_2423[5], op_25_V_reg_2423[5], op_25_V_reg_2423[5], op_25_V_reg_2423, 6'h00 };
assign grp_fu_1610_p1 = { op_17_V_reg_2313[7], op_17_V_reg_2313[7], op_17_V_reg_2313[7], op_17_V_reg_2313[7], op_17_V_reg_2313[7], op_17_V_reg_2313[7], op_17_V_reg_2313[7], op_17_V_reg_2313[7], op_17_V_reg_2313[7], op_17_V_reg_2313[7], op_17_V_reg_2313[7], op_17_V_reg_2313[7], op_17_V_reg_2313[7], op_17_V_reg_2313[7], op_17_V_reg_2313[7], op_17_V_reg_2313[7], op_17_V_reg_2313[7], op_17_V_reg_2313[7], op_17_V_reg_2313[7], op_17_V_reg_2313[7], op_17_V_reg_2313[7], op_17_V_reg_2313[7], op_17_V_reg_2313[7], op_17_V_reg_2313[7], op_17_V_reg_2313[7], op_17_V_reg_2313[7], op_17_V_reg_2313[7], op_17_V_reg_2313[7], op_17_V_reg_2313[7], op_17_V_reg_2313[7], op_17_V_reg_2313[7], op_17_V_reg_2313 };
assign grp_fu_1638_p0 = { op_19[7], op_19 };
assign grp_fu_1638_p1 = { ret_V_21_reg_2279[3], ret_V_21_reg_2279[3], ret_V_21_reg_2279[3], ret_V_21_reg_2279[3], ret_V_21_reg_2279[3], ret_V_21_reg_2279 };
assign grp_fu_1666_p0 = { add_ln69_3_reg_2470[8], add_ln69_3_reg_2470[8], add_ln69_3_reg_2470[8], add_ln69_3_reg_2470[8], add_ln69_3_reg_2470[8], add_ln69_3_reg_2470[8], add_ln69_3_reg_2470[8], add_ln69_3_reg_2470[8], add_ln69_3_reg_2470[8], add_ln69_3_reg_2470[8], add_ln69_3_reg_2470[8], add_ln69_3_reg_2470[8], add_ln69_3_reg_2470[8], add_ln69_3_reg_2470[8], add_ln69_3_reg_2470[8], add_ln69_3_reg_2470[8], add_ln69_3_reg_2470[8], add_ln69_3_reg_2470[8], add_ln69_3_reg_2470[8], add_ln69_3_reg_2470[8], add_ln69_3_reg_2470[8], add_ln69_3_reg_2470[8], add_ln69_3_reg_2470[8], add_ln69_3_reg_2470 };
assign grp_fu_307_p0 = op_2;
assign grp_fu_307_p1 = op_2;
assign grp_fu_347_p0 = { op_4_V_reg_1693[7], op_4_V_reg_1693 };
assign grp_fu_347_p1 = { 7'h00, op_5 };
assign grp_fu_518_p1 = { 1'h0, and_ln414_reg_1811 };
assign grp_fu_589_p0 = { trunc_ln1192_3_reg_1864, 23'h000000 };
assign grp_fu_594_p0 = { trunc_ln1192_reg_1859, 23'h000000 };
assign grp_fu_746_p1 = { 7'h00, and_ln412_reg_1959 };
assign grp_fu_838_p0 = { op_3_V_reg_1816[3], op_3_V_reg_1816[3], op_3_V_reg_1816[3], op_3_V_reg_1816[3], op_3_V_reg_1816[3], op_3_V_reg_1816[3], op_3_V_reg_1816, 23'h000000 };
assign grp_fu_838_p1 = { op_6[31], op_6 };
assign grp_fu_894_p0 = { 2'h0, op_7, 5'h00 };
assign grp_fu_894_p1 = { op_8_V_reg_1964[7], op_8_V_reg_1964[7], op_8_V_reg_1964[7], op_8_V_reg_1964 };
assign grp_fu_914_p0 = { op_8_V_reg_1964[7], op_8_V_reg_1964 };
assign grp_fu_914_p1 = { trunc_ln703_reg_1854, trunc_ln703_reg_1854, trunc_ln703_reg_1854, 6'h00 };
assign lhs_V_1_fu_824_p3 = { op_3_V_reg_1816, 23'h000000 };
assign lhs_V_3_fu_879_p3 = { op_7, 5'h00 };
assign op_28 = grp_fu_1666_p2;
assign or_ln760_fu_329_p1 = op_2;
assign or_ln_fu_535_p4 = { tmp_reg_1832, 2'h0, p_Result_s_reg_1838 };
assign p_Result_12_fu_974_p4 = { p_Result_33_reg_1778, p_Val2_4_fu_969_p2 };
assign p_Result_17_fu_668_p3 = add_ln1192_2_reg_1932[17];
assign p_Result_1_fu_429_p1 = op_6;
assign p_Result_1_fu_429_p4 = op_6[31:25];
assign p_Result_25_fu_1502_p3 = ret_V_18_reg_2269[3];
assign p_Result_26_fu_1291_p3 = ret_V_20_reg_2138[8];
assign p_Result_27_fu_1310_p3 = ret_V_22_reg_2155[31];
assign p_Result_28_fu_1644_p3 = ret_V_25_reg_2438[38];
assign p_Result_30_fu_385_p1 = op_6;
assign p_Result_31_fu_403_p1 = op_6;
assign p_Result_33_fu_421_p1 = op_6;
assign p_Result_35_fu_675_p1 = op_6;
assign p_Result_35_fu_675_p3 = op_6[16];
assign p_Result_3_fu_445_p1 = op_6;
assign p_Result_3_fu_445_p4 = op_6[31:24];
assign p_Result_42_fu_1393_p3 = ret_V_17_reg_2104[8];
assign p_Result_s_20_fu_554_p3 = { trunc_ln790_reg_1844, 5'h00 };
assign p_Val2_10_fu_852_p3 = { p_Result_39_reg_1698, 1'h0 };
assign p_Val2_1_fu_693_p2 = { ret_reg_1821[2:0], 5'h00 };
assign p_Val2_2_fu_393_p1 = op_6;
assign ret_V_22_fu_1119_p1 = op_6;
assign rhs_3_fu_935_p3 = { select_ln384_5_fu_927_p3, 22'h000000 };
assign rhs_fu_903_p3 = { trunc_ln703_reg_1854, 6'h00 };
assign sext_ln1195_fu_1116_p1 = { rhs_3_reg_2060[23], rhs_3_reg_2060[23], rhs_3_reg_2060[23], rhs_3_reg_2060[23], rhs_3_reg_2060[23], rhs_3_reg_2060[23], rhs_3_reg_2060[23], rhs_3_reg_2060[23], rhs_3_reg_2060 };
assign sext_ln69_fu_289_p0 = op_2;
assign sext_ln69_fu_289_p1 = { op_2[3], op_2[3], op_2[3], op_2[3], op_2 };
assign sext_ln703_1_fu_835_p0 = op_6;
assign sext_ln850_fu_1364_p1 = { tmp_5_reg_2274[2], tmp_5_reg_2274 };
assign tmp_14_fu_1198_p3 = add_ln1192_1_reg_1927[25];
assign tmp_21_fu_1450_p3 = ret_V_17_reg_2104[9];
assign tmp_25_fu_1599_p3 = { op_25_V_reg_2423, 6'h00 };
assign tmp_6_fu_943_p1 = op_6;
assign tmp_6_fu_943_p3 = op_6[24];
assign tmp_7_fu_950_p3 = p_Val2_3_reg_1884[1];
assign trunc_ln1192_2_fu_467_p0 = op_6;
assign trunc_ln1192_2_fu_467_p1 = op_6[25:0];
assign trunc_ln1192_3_fu_531_p1 = grp_fu_279_p2[2:0];
assign trunc_ln1192_fu_527_p1 = grp_fu_279_p2[1:0];
assign trunc_ln414_fu_411_p0 = op_6;
assign trunc_ln414_fu_411_p1 = op_6[21:0];
assign trunc_ln69_1_fu_285_p1 = op_1[7:0];
assign trunc_ln69_2_fu_293_p1 = op_1[0];
assign trunc_ln69_3_fu_297_p0 = op_2;
assign trunc_ln69_3_fu_297_p1 = op_2[0];
assign trunc_ln69_fu_275_p1 = op_1[3:0];
assign trunc_ln703_fu_523_p1 = grp_fu_279_p2[0];
assign trunc_ln718_1_fu_1088_p1 = grp_fu_894_p2[3:0];
assign trunc_ln718_fu_471_p0 = op_6;
assign trunc_ln718_fu_471_p1 = op_6[15:0];
assign trunc_ln731_fu_313_p1 = op_5[0];
assign trunc_ln790_fu_511_p1 = grp_fu_307_p2[1:0];
assign trunc_ln851_1_fu_1112_p1 = grp_fu_914_p2[4:0];
assign trunc_ln851_2_fu_1134_p1 = ret_V_22_fu_1119_p2[22:0];
assign trunc_ln851_3_fu_1434_p1 = op_17_V_fu_1387_p3[5:0];
assign trunc_ln851_fu_1509_p1 = op_12_V_reg_2172[0];
assign \sub_9s_9s_9_2_1_U10.top_sub_9s_9s_9_2_1_Adder_7_U.ain_s0  = \sub_9s_9s_9_2_1_U10.top_sub_9s_9s_9_2_1_Adder_7_U.a ;
assign \sub_9s_9s_9_2_1_U10.top_sub_9s_9s_9_2_1_Adder_7_U.s  = { \sub_9s_9s_9_2_1_U10.top_sub_9s_9s_9_2_1_Adder_7_U.fas_s2 , \sub_9s_9s_9_2_1_U10.top_sub_9s_9s_9_2_1_Adder_7_U.sum_s1  };
assign \sub_9s_9s_9_2_1_U10.top_sub_9s_9s_9_2_1_Adder_7_U.u2.a  = \sub_9s_9s_9_2_1_U10.top_sub_9s_9s_9_2_1_Adder_7_U.ain_s1 ;
assign \sub_9s_9s_9_2_1_U10.top_sub_9s_9s_9_2_1_Adder_7_U.u2.b  = \sub_9s_9s_9_2_1_U10.top_sub_9s_9s_9_2_1_Adder_7_U.bin_s1 ;
assign \sub_9s_9s_9_2_1_U10.top_sub_9s_9s_9_2_1_Adder_7_U.u2.cin  = \sub_9s_9s_9_2_1_U10.top_sub_9s_9s_9_2_1_Adder_7_U.carry_s1 ;
assign \sub_9s_9s_9_2_1_U10.top_sub_9s_9s_9_2_1_Adder_7_U.facout_s2  = \sub_9s_9s_9_2_1_U10.top_sub_9s_9s_9_2_1_Adder_7_U.u2.cout ;
assign \sub_9s_9s_9_2_1_U10.top_sub_9s_9s_9_2_1_Adder_7_U.fas_s2  = \sub_9s_9s_9_2_1_U10.top_sub_9s_9s_9_2_1_Adder_7_U.u2.s ;
assign \sub_9s_9s_9_2_1_U10.top_sub_9s_9s_9_2_1_Adder_7_U.u1.a  = \sub_9s_9s_9_2_1_U10.top_sub_9s_9s_9_2_1_Adder_7_U.a [3:0];
assign \sub_9s_9s_9_2_1_U10.top_sub_9s_9s_9_2_1_Adder_7_U.u1.b  = \sub_9s_9s_9_2_1_U10.top_sub_9s_9s_9_2_1_Adder_7_U.bin_s0 [3:0];
assign \sub_9s_9s_9_2_1_U10.top_sub_9s_9s_9_2_1_Adder_7_U.u1.cin  = 1'h1;
assign \sub_9s_9s_9_2_1_U10.top_sub_9s_9s_9_2_1_Adder_7_U.facout_s1  = \sub_9s_9s_9_2_1_U10.top_sub_9s_9s_9_2_1_Adder_7_U.u1.cout ;
assign \sub_9s_9s_9_2_1_U10.top_sub_9s_9s_9_2_1_Adder_7_U.fas_s1  = \sub_9s_9s_9_2_1_U10.top_sub_9s_9s_9_2_1_Adder_7_U.u1.s ;
assign \sub_9s_9s_9_2_1_U10.top_sub_9s_9s_9_2_1_Adder_7_U.a  = \sub_9s_9s_9_2_1_U10.din0 ;
assign \sub_9s_9s_9_2_1_U10.top_sub_9s_9s_9_2_1_Adder_7_U.b  = \sub_9s_9s_9_2_1_U10.din1 ;
assign \sub_9s_9s_9_2_1_U10.top_sub_9s_9s_9_2_1_Adder_7_U.ce  = \sub_9s_9s_9_2_1_U10.ce ;
assign \sub_9s_9s_9_2_1_U10.top_sub_9s_9s_9_2_1_Adder_7_U.clk  = \sub_9s_9s_9_2_1_U10.clk ;
assign \sub_9s_9s_9_2_1_U10.top_sub_9s_9s_9_2_1_Adder_7_U.reset  = \sub_9s_9s_9_2_1_U10.reset ;
assign \sub_9s_9s_9_2_1_U10.dout  = \sub_9s_9s_9_2_1_U10.top_sub_9s_9s_9_2_1_Adder_7_U.s ;
assign \sub_9s_9s_9_2_1_U10.ce  = 1'h1;
assign \sub_9s_9s_9_2_1_U10.clk  = ap_clk;
assign \sub_9s_9s_9_2_1_U10.din0  = { op_8_V_reg_1964[7], op_8_V_reg_1964 };
assign \sub_9s_9s_9_2_1_U10.din1  = { trunc_ln703_reg_1854, trunc_ln703_reg_1854, trunc_ln703_reg_1854, 6'h00 };
assign grp_fu_914_p2 = \sub_9s_9s_9_2_1_U10.dout ;
assign \sub_9s_9s_9_2_1_U10.reset  = ap_rst;
assign \sub_11ns_11s_11_2_1_U9.top_sub_11ns_11s_11_2_1_Adder_6_U.ain_s0  = \sub_11ns_11s_11_2_1_U9.top_sub_11ns_11s_11_2_1_Adder_6_U.a ;
assign \sub_11ns_11s_11_2_1_U9.top_sub_11ns_11s_11_2_1_Adder_6_U.s  = { \sub_11ns_11s_11_2_1_U9.top_sub_11ns_11s_11_2_1_Adder_6_U.fas_s2 , \sub_11ns_11s_11_2_1_U9.top_sub_11ns_11s_11_2_1_Adder_6_U.sum_s1  };
assign \sub_11ns_11s_11_2_1_U9.top_sub_11ns_11s_11_2_1_Adder_6_U.u2.a  = \sub_11ns_11s_11_2_1_U9.top_sub_11ns_11s_11_2_1_Adder_6_U.ain_s1 ;
assign \sub_11ns_11s_11_2_1_U9.top_sub_11ns_11s_11_2_1_Adder_6_U.u2.b  = \sub_11ns_11s_11_2_1_U9.top_sub_11ns_11s_11_2_1_Adder_6_U.bin_s1 ;
assign \sub_11ns_11s_11_2_1_U9.top_sub_11ns_11s_11_2_1_Adder_6_U.u2.cin  = \sub_11ns_11s_11_2_1_U9.top_sub_11ns_11s_11_2_1_Adder_6_U.carry_s1 ;
assign \sub_11ns_11s_11_2_1_U9.top_sub_11ns_11s_11_2_1_Adder_6_U.facout_s2  = \sub_11ns_11s_11_2_1_U9.top_sub_11ns_11s_11_2_1_Adder_6_U.u2.cout ;
assign \sub_11ns_11s_11_2_1_U9.top_sub_11ns_11s_11_2_1_Adder_6_U.fas_s2  = \sub_11ns_11s_11_2_1_U9.top_sub_11ns_11s_11_2_1_Adder_6_U.u2.s ;
assign \sub_11ns_11s_11_2_1_U9.top_sub_11ns_11s_11_2_1_Adder_6_U.u1.a  = \sub_11ns_11s_11_2_1_U9.top_sub_11ns_11s_11_2_1_Adder_6_U.a [4:0];
assign \sub_11ns_11s_11_2_1_U9.top_sub_11ns_11s_11_2_1_Adder_6_U.u1.b  = \sub_11ns_11s_11_2_1_U9.top_sub_11ns_11s_11_2_1_Adder_6_U.bin_s0 [4:0];
assign \sub_11ns_11s_11_2_1_U9.top_sub_11ns_11s_11_2_1_Adder_6_U.u1.cin  = 1'h1;
assign \sub_11ns_11s_11_2_1_U9.top_sub_11ns_11s_11_2_1_Adder_6_U.facout_s1  = \sub_11ns_11s_11_2_1_U9.top_sub_11ns_11s_11_2_1_Adder_6_U.u1.cout ;
assign \sub_11ns_11s_11_2_1_U9.top_sub_11ns_11s_11_2_1_Adder_6_U.fas_s1  = \sub_11ns_11s_11_2_1_U9.top_sub_11ns_11s_11_2_1_Adder_6_U.u1.s ;
assign \sub_11ns_11s_11_2_1_U9.top_sub_11ns_11s_11_2_1_Adder_6_U.a  = \sub_11ns_11s_11_2_1_U9.din0 ;
assign \sub_11ns_11s_11_2_1_U9.top_sub_11ns_11s_11_2_1_Adder_6_U.b  = \sub_11ns_11s_11_2_1_U9.din1 ;
assign \sub_11ns_11s_11_2_1_U9.top_sub_11ns_11s_11_2_1_Adder_6_U.ce  = \sub_11ns_11s_11_2_1_U9.ce ;
assign \sub_11ns_11s_11_2_1_U9.top_sub_11ns_11s_11_2_1_Adder_6_U.clk  = \sub_11ns_11s_11_2_1_U9.clk ;
assign \sub_11ns_11s_11_2_1_U9.top_sub_11ns_11s_11_2_1_Adder_6_U.reset  = \sub_11ns_11s_11_2_1_U9.reset ;
assign \sub_11ns_11s_11_2_1_U9.dout  = \sub_11ns_11s_11_2_1_U9.top_sub_11ns_11s_11_2_1_Adder_6_U.s ;
assign \sub_11ns_11s_11_2_1_U9.ce  = 1'h1;
assign \sub_11ns_11s_11_2_1_U9.clk  = ap_clk;
assign \sub_11ns_11s_11_2_1_U9.din0  = { 2'h0, op_7, 5'h00 };
assign \sub_11ns_11s_11_2_1_U9.din1  = { op_8_V_reg_1964[7], op_8_V_reg_1964[7], op_8_V_reg_1964[7], op_8_V_reg_1964 };
assign grp_fu_894_p2 = \sub_11ns_11s_11_2_1_U9.dout ;
assign \sub_11ns_11s_11_2_1_U9.reset  = ap_rst;
assign \mul_4s_4s_8_7_1_U2.top_mul_4s_4s_8_7_1_Mul_DSP_1_U.p  = \mul_4s_4s_8_7_1_U2.top_mul_4s_4s_8_7_1_Mul_DSP_1_U.buff4 ;
assign \mul_4s_4s_8_7_1_U2.top_mul_4s_4s_8_7_1_Mul_DSP_1_U.a  = \mul_4s_4s_8_7_1_U2.din0 ;
assign \mul_4s_4s_8_7_1_U2.top_mul_4s_4s_8_7_1_Mul_DSP_1_U.b  = \mul_4s_4s_8_7_1_U2.din1 ;
assign \mul_4s_4s_8_7_1_U2.top_mul_4s_4s_8_7_1_Mul_DSP_1_U.ce  = \mul_4s_4s_8_7_1_U2.ce ;
assign \mul_4s_4s_8_7_1_U2.top_mul_4s_4s_8_7_1_Mul_DSP_1_U.clk  = \mul_4s_4s_8_7_1_U2.clk ;
assign \mul_4s_4s_8_7_1_U2.dout  = \mul_4s_4s_8_7_1_U2.top_mul_4s_4s_8_7_1_Mul_DSP_1_U.p ;
assign \mul_4s_4s_8_7_1_U2.ce  = 1'h1;
assign \mul_4s_4s_8_7_1_U2.clk  = ap_clk;
assign \mul_4s_4s_8_7_1_U2.din0  = op_2;
assign \mul_4s_4s_8_7_1_U2.din1  = op_2;
assign grp_fu_307_p2 = \mul_4s_4s_8_7_1_U2.dout ;
assign \mul_4s_4s_8_7_1_U2.reset  = ap_rst;
assign \mul_4s_4s_4_7_1_U1.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.p  = \mul_4s_4s_4_7_1_U1.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.buff4 ;
assign \mul_4s_4s_4_7_1_U1.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.a  = \mul_4s_4s_4_7_1_U1.din0 ;
assign \mul_4s_4s_4_7_1_U1.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.b  = \mul_4s_4s_4_7_1_U1.din1 ;
assign \mul_4s_4s_4_7_1_U1.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.ce  = \mul_4s_4s_4_7_1_U1.ce ;
assign \mul_4s_4s_4_7_1_U1.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.clk  = \mul_4s_4s_4_7_1_U1.clk ;
assign \mul_4s_4s_4_7_1_U1.dout  = \mul_4s_4s_4_7_1_U1.top_mul_4s_4s_4_7_1_Mul_DSP_0_U.p ;
assign \mul_4s_4s_4_7_1_U1.ce  = 1'h1;
assign \mul_4s_4s_4_7_1_U1.clk  = ap_clk;
assign \mul_4s_4s_4_7_1_U1.din0  = op_1[3:0];
assign \mul_4s_4s_4_7_1_U1.din1  = op_2;
assign grp_fu_279_p2 = \mul_4s_4s_4_7_1_U1.dout ;
assign \mul_4s_4s_4_7_1_U1.reset  = ap_rst;
assign \add_9s_9s_9_2_1_U23.top_add_9s_9s_9_2_1_Adder_18_U.ain_s0  = \add_9s_9s_9_2_1_U23.top_add_9s_9s_9_2_1_Adder_18_U.a ;
assign \add_9s_9s_9_2_1_U23.top_add_9s_9s_9_2_1_Adder_18_U.bin_s0  = \add_9s_9s_9_2_1_U23.top_add_9s_9s_9_2_1_Adder_18_U.b ;
assign \add_9s_9s_9_2_1_U23.top_add_9s_9s_9_2_1_Adder_18_U.s  = { \add_9s_9s_9_2_1_U23.top_add_9s_9s_9_2_1_Adder_18_U.fas_s2 , \add_9s_9s_9_2_1_U23.top_add_9s_9s_9_2_1_Adder_18_U.sum_s1  };
assign \add_9s_9s_9_2_1_U23.top_add_9s_9s_9_2_1_Adder_18_U.u2.a  = \add_9s_9s_9_2_1_U23.top_add_9s_9s_9_2_1_Adder_18_U.ain_s1 ;
assign \add_9s_9s_9_2_1_U23.top_add_9s_9s_9_2_1_Adder_18_U.u2.b  = \add_9s_9s_9_2_1_U23.top_add_9s_9s_9_2_1_Adder_18_U.bin_s1 ;
assign \add_9s_9s_9_2_1_U23.top_add_9s_9s_9_2_1_Adder_18_U.u2.cin  = \add_9s_9s_9_2_1_U23.top_add_9s_9s_9_2_1_Adder_18_U.carry_s1 ;
assign \add_9s_9s_9_2_1_U23.top_add_9s_9s_9_2_1_Adder_18_U.facout_s2  = \add_9s_9s_9_2_1_U23.top_add_9s_9s_9_2_1_Adder_18_U.u2.cout ;
assign \add_9s_9s_9_2_1_U23.top_add_9s_9s_9_2_1_Adder_18_U.fas_s2  = \add_9s_9s_9_2_1_U23.top_add_9s_9s_9_2_1_Adder_18_U.u2.s ;
assign \add_9s_9s_9_2_1_U23.top_add_9s_9s_9_2_1_Adder_18_U.u1.a  = \add_9s_9s_9_2_1_U23.top_add_9s_9s_9_2_1_Adder_18_U.a [3:0];
assign \add_9s_9s_9_2_1_U23.top_add_9s_9s_9_2_1_Adder_18_U.u1.b  = \add_9s_9s_9_2_1_U23.top_add_9s_9s_9_2_1_Adder_18_U.b [3:0];
assign \add_9s_9s_9_2_1_U23.top_add_9s_9s_9_2_1_Adder_18_U.u1.cin  = 1'h0;
assign \add_9s_9s_9_2_1_U23.top_add_9s_9s_9_2_1_Adder_18_U.facout_s1  = \add_9s_9s_9_2_1_U23.top_add_9s_9s_9_2_1_Adder_18_U.u1.cout ;
assign \add_9s_9s_9_2_1_U23.top_add_9s_9s_9_2_1_Adder_18_U.fas_s1  = \add_9s_9s_9_2_1_U23.top_add_9s_9s_9_2_1_Adder_18_U.u1.s ;
assign \add_9s_9s_9_2_1_U23.top_add_9s_9s_9_2_1_Adder_18_U.a  = \add_9s_9s_9_2_1_U23.din0 ;
assign \add_9s_9s_9_2_1_U23.top_add_9s_9s_9_2_1_Adder_18_U.b  = \add_9s_9s_9_2_1_U23.din1 ;
assign \add_9s_9s_9_2_1_U23.top_add_9s_9s_9_2_1_Adder_18_U.ce  = \add_9s_9s_9_2_1_U23.ce ;
assign \add_9s_9s_9_2_1_U23.top_add_9s_9s_9_2_1_Adder_18_U.clk  = \add_9s_9s_9_2_1_U23.clk ;
assign \add_9s_9s_9_2_1_U23.top_add_9s_9s_9_2_1_Adder_18_U.reset  = \add_9s_9s_9_2_1_U23.reset ;
assign \add_9s_9s_9_2_1_U23.dout  = \add_9s_9s_9_2_1_U23.top_add_9s_9s_9_2_1_Adder_18_U.s ;
assign \add_9s_9s_9_2_1_U23.ce  = 1'h1;
assign \add_9s_9s_9_2_1_U23.clk  = ap_clk;
assign \add_9s_9s_9_2_1_U23.din0  = { op_19[7], op_19 };
assign \add_9s_9s_9_2_1_U23.din1  = { ret_V_21_reg_2279[3], ret_V_21_reg_2279[3], ret_V_21_reg_2279[3], ret_V_21_reg_2279[3], ret_V_21_reg_2279[3], ret_V_21_reg_2279 };
assign grp_fu_1638_p2 = \add_9s_9s_9_2_1_U23.dout ;
assign \add_9s_9s_9_2_1_U23.reset  = ap_rst;
assign \add_9s_9ns_9_2_1_U3.top_add_9s_9ns_9_2_1_Adder_0_U.ain_s0  = \add_9s_9ns_9_2_1_U3.top_add_9s_9ns_9_2_1_Adder_0_U.a ;
assign \add_9s_9ns_9_2_1_U3.top_add_9s_9ns_9_2_1_Adder_0_U.bin_s0  = \add_9s_9ns_9_2_1_U3.top_add_9s_9ns_9_2_1_Adder_0_U.b ;
assign \add_9s_9ns_9_2_1_U3.top_add_9s_9ns_9_2_1_Adder_0_U.s  = { \add_9s_9ns_9_2_1_U3.top_add_9s_9ns_9_2_1_Adder_0_U.fas_s2 , \add_9s_9ns_9_2_1_U3.top_add_9s_9ns_9_2_1_Adder_0_U.sum_s1  };
assign \add_9s_9ns_9_2_1_U3.top_add_9s_9ns_9_2_1_Adder_0_U.u2.a  = \add_9s_9ns_9_2_1_U3.top_add_9s_9ns_9_2_1_Adder_0_U.ain_s1 ;
assign \add_9s_9ns_9_2_1_U3.top_add_9s_9ns_9_2_1_Adder_0_U.u2.b  = \add_9s_9ns_9_2_1_U3.top_add_9s_9ns_9_2_1_Adder_0_U.bin_s1 ;
assign \add_9s_9ns_9_2_1_U3.top_add_9s_9ns_9_2_1_Adder_0_U.u2.cin  = \add_9s_9ns_9_2_1_U3.top_add_9s_9ns_9_2_1_Adder_0_U.carry_s1 ;
assign \add_9s_9ns_9_2_1_U3.top_add_9s_9ns_9_2_1_Adder_0_U.facout_s2  = \add_9s_9ns_9_2_1_U3.top_add_9s_9ns_9_2_1_Adder_0_U.u2.cout ;
assign \add_9s_9ns_9_2_1_U3.top_add_9s_9ns_9_2_1_Adder_0_U.fas_s2  = \add_9s_9ns_9_2_1_U3.top_add_9s_9ns_9_2_1_Adder_0_U.u2.s ;
assign \add_9s_9ns_9_2_1_U3.top_add_9s_9ns_9_2_1_Adder_0_U.u1.a  = \add_9s_9ns_9_2_1_U3.top_add_9s_9ns_9_2_1_Adder_0_U.a [3:0];
assign \add_9s_9ns_9_2_1_U3.top_add_9s_9ns_9_2_1_Adder_0_U.u1.b  = \add_9s_9ns_9_2_1_U3.top_add_9s_9ns_9_2_1_Adder_0_U.b [3:0];
assign \add_9s_9ns_9_2_1_U3.top_add_9s_9ns_9_2_1_Adder_0_U.u1.cin  = 1'h0;
assign \add_9s_9ns_9_2_1_U3.top_add_9s_9ns_9_2_1_Adder_0_U.facout_s1  = \add_9s_9ns_9_2_1_U3.top_add_9s_9ns_9_2_1_Adder_0_U.u1.cout ;
assign \add_9s_9ns_9_2_1_U3.top_add_9s_9ns_9_2_1_Adder_0_U.fas_s1  = \add_9s_9ns_9_2_1_U3.top_add_9s_9ns_9_2_1_Adder_0_U.u1.s ;
assign \add_9s_9ns_9_2_1_U3.top_add_9s_9ns_9_2_1_Adder_0_U.a  = \add_9s_9ns_9_2_1_U3.din0 ;
assign \add_9s_9ns_9_2_1_U3.top_add_9s_9ns_9_2_1_Adder_0_U.b  = \add_9s_9ns_9_2_1_U3.din1 ;
assign \add_9s_9ns_9_2_1_U3.top_add_9s_9ns_9_2_1_Adder_0_U.ce  = \add_9s_9ns_9_2_1_U3.ce ;
assign \add_9s_9ns_9_2_1_U3.top_add_9s_9ns_9_2_1_Adder_0_U.clk  = \add_9s_9ns_9_2_1_U3.clk ;
assign \add_9s_9ns_9_2_1_U3.top_add_9s_9ns_9_2_1_Adder_0_U.reset  = \add_9s_9ns_9_2_1_U3.reset ;
assign \add_9s_9ns_9_2_1_U3.dout  = \add_9s_9ns_9_2_1_U3.top_add_9s_9ns_9_2_1_Adder_0_U.s ;
assign \add_9s_9ns_9_2_1_U3.ce  = 1'h1;
assign \add_9s_9ns_9_2_1_U3.clk  = ap_clk;
assign \add_9s_9ns_9_2_1_U3.din0  = { op_4_V_reg_1693[7], op_4_V_reg_1693 };
assign \add_9s_9ns_9_2_1_U3.din1  = { 7'h00, op_5 };
assign grp_fu_347_p2 = \add_9s_9ns_9_2_1_U3.dout ;
assign \add_9s_9ns_9_2_1_U3.reset  = ap_rst;
assign \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_4_U.ain_s0  = \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_4_U.a ;
assign \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_4_U.bin_s0  = \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_4_U.b ;
assign \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_4_U.s  = { \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_4_U.fas_s2 , \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_4_U.sum_s1  };
assign \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_4_U.u2.a  = \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_4_U.ain_s1 ;
assign \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_4_U.u2.b  = \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_4_U.bin_s1 ;
assign \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_4_U.u2.cin  = \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_4_U.carry_s1 ;
assign \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_4_U.facout_s2  = \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_4_U.u2.cout ;
assign \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_4_U.fas_s2  = \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_4_U.u2.s ;
assign \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_4_U.u1.a  = \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_4_U.a [3:0];
assign \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_4_U.u1.b  = \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_4_U.b [3:0];
assign \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_4_U.u1.cin  = 1'h0;
assign \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_4_U.facout_s1  = \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_4_U.u1.cout ;
assign \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_4_U.fas_s1  = \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_4_U.u1.s ;
assign \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_4_U.a  = \add_8ns_8ns_8_2_1_U7.din0 ;
assign \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_4_U.b  = \add_8ns_8ns_8_2_1_U7.din1 ;
assign \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_4_U.ce  = \add_8ns_8ns_8_2_1_U7.ce ;
assign \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_4_U.clk  = \add_8ns_8ns_8_2_1_U7.clk ;
assign \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_4_U.reset  = \add_8ns_8ns_8_2_1_U7.reset ;
assign \add_8ns_8ns_8_2_1_U7.dout  = \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_4_U.s ;
assign \add_8ns_8ns_8_2_1_U7.ce  = 1'h1;
assign \add_8ns_8ns_8_2_1_U7.clk  = ap_clk;
assign \add_8ns_8ns_8_2_1_U7.din0  = p_Val2_7_reg_1937;
assign \add_8ns_8ns_8_2_1_U7.din1  = { 7'h00, and_ln412_reg_1959 };
assign grp_fu_746_p2 = \add_8ns_8ns_8_2_1_U7.dout ;
assign \add_8ns_8ns_8_2_1_U7.reset  = ap_rst;
assign \add_6s_6s_6_2_1_U19.top_add_6s_6s_6_2_1_Adder_14_U.ain_s0  = \add_6s_6s_6_2_1_U19.top_add_6s_6s_6_2_1_Adder_14_U.a ;
assign \add_6s_6s_6_2_1_U19.top_add_6s_6s_6_2_1_Adder_14_U.bin_s0  = \add_6s_6s_6_2_1_U19.top_add_6s_6s_6_2_1_Adder_14_U.b ;
assign \add_6s_6s_6_2_1_U19.top_add_6s_6s_6_2_1_Adder_14_U.s  = { \add_6s_6s_6_2_1_U19.top_add_6s_6s_6_2_1_Adder_14_U.fas_s2 , \add_6s_6s_6_2_1_U19.top_add_6s_6s_6_2_1_Adder_14_U.sum_s1  };
assign \add_6s_6s_6_2_1_U19.top_add_6s_6s_6_2_1_Adder_14_U.u2.a  = \add_6s_6s_6_2_1_U19.top_add_6s_6s_6_2_1_Adder_14_U.ain_s1 ;
assign \add_6s_6s_6_2_1_U19.top_add_6s_6s_6_2_1_Adder_14_U.u2.b  = \add_6s_6s_6_2_1_U19.top_add_6s_6s_6_2_1_Adder_14_U.bin_s1 ;
assign \add_6s_6s_6_2_1_U19.top_add_6s_6s_6_2_1_Adder_14_U.u2.cin  = \add_6s_6s_6_2_1_U19.top_add_6s_6s_6_2_1_Adder_14_U.carry_s1 ;
assign \add_6s_6s_6_2_1_U19.top_add_6s_6s_6_2_1_Adder_14_U.facout_s2  = \add_6s_6s_6_2_1_U19.top_add_6s_6s_6_2_1_Adder_14_U.u2.cout ;
assign \add_6s_6s_6_2_1_U19.top_add_6s_6s_6_2_1_Adder_14_U.fas_s2  = \add_6s_6s_6_2_1_U19.top_add_6s_6s_6_2_1_Adder_14_U.u2.s ;
assign \add_6s_6s_6_2_1_U19.top_add_6s_6s_6_2_1_Adder_14_U.u1.a  = \add_6s_6s_6_2_1_U19.top_add_6s_6s_6_2_1_Adder_14_U.a [2:0];
assign \add_6s_6s_6_2_1_U19.top_add_6s_6s_6_2_1_Adder_14_U.u1.b  = \add_6s_6s_6_2_1_U19.top_add_6s_6s_6_2_1_Adder_14_U.b [2:0];
assign \add_6s_6s_6_2_1_U19.top_add_6s_6s_6_2_1_Adder_14_U.u1.cin  = 1'h0;
assign \add_6s_6s_6_2_1_U19.top_add_6s_6s_6_2_1_Adder_14_U.facout_s1  = \add_6s_6s_6_2_1_U19.top_add_6s_6s_6_2_1_Adder_14_U.u1.cout ;
assign \add_6s_6s_6_2_1_U19.top_add_6s_6s_6_2_1_Adder_14_U.fas_s1  = \add_6s_6s_6_2_1_U19.top_add_6s_6s_6_2_1_Adder_14_U.u1.s ;
assign \add_6s_6s_6_2_1_U19.top_add_6s_6s_6_2_1_Adder_14_U.a  = \add_6s_6s_6_2_1_U19.din0 ;
assign \add_6s_6s_6_2_1_U19.top_add_6s_6s_6_2_1_Adder_14_U.b  = \add_6s_6s_6_2_1_U19.din1 ;
assign \add_6s_6s_6_2_1_U19.top_add_6s_6s_6_2_1_Adder_14_U.ce  = \add_6s_6s_6_2_1_U19.ce ;
assign \add_6s_6s_6_2_1_U19.top_add_6s_6s_6_2_1_Adder_14_U.clk  = \add_6s_6s_6_2_1_U19.clk ;
assign \add_6s_6s_6_2_1_U19.top_add_6s_6s_6_2_1_Adder_14_U.reset  = \add_6s_6s_6_2_1_U19.reset ;
assign \add_6s_6s_6_2_1_U19.dout  = \add_6s_6s_6_2_1_U19.top_add_6s_6s_6_2_1_Adder_14_U.s ;
assign \add_6s_6s_6_2_1_U19.ce  = 1'h1;
assign \add_6s_6s_6_2_1_U19.clk  = ap_clk;
assign \add_6s_6s_6_2_1_U19.din0  = { op_23_V_reg_2398[4], op_23_V_reg_2398 };
assign \add_6s_6s_6_2_1_U19.din1  = { op_15_V_reg_2393[3], op_15_V_reg_2393[3], op_15_V_reg_2393 };
assign grp_fu_1582_p2 = \add_6s_6s_6_2_1_U19.dout ;
assign \add_6s_6s_6_2_1_U19.reset  = ap_rst;
assign \add_6ns_6s_6_2_1_U20.top_add_6ns_6s_6_2_1_Adder_15_U.ain_s0  = \add_6ns_6s_6_2_1_U20.top_add_6ns_6s_6_2_1_Adder_15_U.a ;
assign \add_6ns_6s_6_2_1_U20.top_add_6ns_6s_6_2_1_Adder_15_U.bin_s0  = \add_6ns_6s_6_2_1_U20.top_add_6ns_6s_6_2_1_Adder_15_U.b ;
assign \add_6ns_6s_6_2_1_U20.top_add_6ns_6s_6_2_1_Adder_15_U.s  = { \add_6ns_6s_6_2_1_U20.top_add_6ns_6s_6_2_1_Adder_15_U.fas_s2 , \add_6ns_6s_6_2_1_U20.top_add_6ns_6s_6_2_1_Adder_15_U.sum_s1  };
assign \add_6ns_6s_6_2_1_U20.top_add_6ns_6s_6_2_1_Adder_15_U.u2.a  = \add_6ns_6s_6_2_1_U20.top_add_6ns_6s_6_2_1_Adder_15_U.ain_s1 ;
assign \add_6ns_6s_6_2_1_U20.top_add_6ns_6s_6_2_1_Adder_15_U.u2.b  = \add_6ns_6s_6_2_1_U20.top_add_6ns_6s_6_2_1_Adder_15_U.bin_s1 ;
assign \add_6ns_6s_6_2_1_U20.top_add_6ns_6s_6_2_1_Adder_15_U.u2.cin  = \add_6ns_6s_6_2_1_U20.top_add_6ns_6s_6_2_1_Adder_15_U.carry_s1 ;
assign \add_6ns_6s_6_2_1_U20.top_add_6ns_6s_6_2_1_Adder_15_U.facout_s2  = \add_6ns_6s_6_2_1_U20.top_add_6ns_6s_6_2_1_Adder_15_U.u2.cout ;
assign \add_6ns_6s_6_2_1_U20.top_add_6ns_6s_6_2_1_Adder_15_U.fas_s2  = \add_6ns_6s_6_2_1_U20.top_add_6ns_6s_6_2_1_Adder_15_U.u2.s ;
assign \add_6ns_6s_6_2_1_U20.top_add_6ns_6s_6_2_1_Adder_15_U.u1.a  = \add_6ns_6s_6_2_1_U20.top_add_6ns_6s_6_2_1_Adder_15_U.a [2:0];
assign \add_6ns_6s_6_2_1_U20.top_add_6ns_6s_6_2_1_Adder_15_U.u1.b  = \add_6ns_6s_6_2_1_U20.top_add_6ns_6s_6_2_1_Adder_15_U.b [2:0];
assign \add_6ns_6s_6_2_1_U20.top_add_6ns_6s_6_2_1_Adder_15_U.u1.cin  = 1'h0;
assign \add_6ns_6s_6_2_1_U20.top_add_6ns_6s_6_2_1_Adder_15_U.facout_s1  = \add_6ns_6s_6_2_1_U20.top_add_6ns_6s_6_2_1_Adder_15_U.u1.cout ;
assign \add_6ns_6s_6_2_1_U20.top_add_6ns_6s_6_2_1_Adder_15_U.fas_s1  = \add_6ns_6s_6_2_1_U20.top_add_6ns_6s_6_2_1_Adder_15_U.u1.s ;
assign \add_6ns_6s_6_2_1_U20.top_add_6ns_6s_6_2_1_Adder_15_U.a  = \add_6ns_6s_6_2_1_U20.din0 ;
assign \add_6ns_6s_6_2_1_U20.top_add_6ns_6s_6_2_1_Adder_15_U.b  = \add_6ns_6s_6_2_1_U20.din1 ;
assign \add_6ns_6s_6_2_1_U20.top_add_6ns_6s_6_2_1_Adder_15_U.ce  = \add_6ns_6s_6_2_1_U20.ce ;
assign \add_6ns_6s_6_2_1_U20.top_add_6ns_6s_6_2_1_Adder_15_U.clk  = \add_6ns_6s_6_2_1_U20.clk ;
assign \add_6ns_6s_6_2_1_U20.top_add_6ns_6s_6_2_1_Adder_15_U.reset  = \add_6ns_6s_6_2_1_U20.reset ;
assign \add_6ns_6s_6_2_1_U20.dout  = \add_6ns_6s_6_2_1_U20.top_add_6ns_6s_6_2_1_Adder_15_U.s ;
assign \add_6ns_6s_6_2_1_U20.ce  = 1'h1;
assign \add_6ns_6s_6_2_1_U20.clk  = ap_clk;
assign \add_6ns_6s_6_2_1_U20.din0  = ret_V_24_reg_2413;
assign \add_6ns_6s_6_2_1_U20.din1  = { op_16_V_reg_1705[3], op_16_V_reg_1705[3], op_16_V_reg_1705 };
assign grp_fu_1591_p2 = \add_6ns_6s_6_2_1_U20.dout ;
assign \add_6ns_6s_6_2_1_U20.reset  = ap_rst;
assign \add_5s_5s_5_2_1_U17.top_add_5s_5s_5_2_1_Adder_12_U.ain_s0  = \add_5s_5s_5_2_1_U17.top_add_5s_5s_5_2_1_Adder_12_U.a ;
assign \add_5s_5s_5_2_1_U17.top_add_5s_5s_5_2_1_Adder_12_U.bin_s0  = \add_5s_5s_5_2_1_U17.top_add_5s_5s_5_2_1_Adder_12_U.b ;
assign \add_5s_5s_5_2_1_U17.top_add_5s_5s_5_2_1_Adder_12_U.s  = { \add_5s_5s_5_2_1_U17.top_add_5s_5s_5_2_1_Adder_12_U.fas_s2 , \add_5s_5s_5_2_1_U17.top_add_5s_5s_5_2_1_Adder_12_U.sum_s1  };
assign \add_5s_5s_5_2_1_U17.top_add_5s_5s_5_2_1_Adder_12_U.u2.a  = \add_5s_5s_5_2_1_U17.top_add_5s_5s_5_2_1_Adder_12_U.ain_s1 ;
assign \add_5s_5s_5_2_1_U17.top_add_5s_5s_5_2_1_Adder_12_U.u2.b  = \add_5s_5s_5_2_1_U17.top_add_5s_5s_5_2_1_Adder_12_U.bin_s1 ;
assign \add_5s_5s_5_2_1_U17.top_add_5s_5s_5_2_1_Adder_12_U.u2.cin  = \add_5s_5s_5_2_1_U17.top_add_5s_5s_5_2_1_Adder_12_U.carry_s1 ;
assign \add_5s_5s_5_2_1_U17.top_add_5s_5s_5_2_1_Adder_12_U.facout_s2  = \add_5s_5s_5_2_1_U17.top_add_5s_5s_5_2_1_Adder_12_U.u2.cout ;
assign \add_5s_5s_5_2_1_U17.top_add_5s_5s_5_2_1_Adder_12_U.fas_s2  = \add_5s_5s_5_2_1_U17.top_add_5s_5s_5_2_1_Adder_12_U.u2.s ;
assign \add_5s_5s_5_2_1_U17.top_add_5s_5s_5_2_1_Adder_12_U.u1.a  = \add_5s_5s_5_2_1_U17.top_add_5s_5s_5_2_1_Adder_12_U.a [1:0];
assign \add_5s_5s_5_2_1_U17.top_add_5s_5s_5_2_1_Adder_12_U.u1.b  = \add_5s_5s_5_2_1_U17.top_add_5s_5s_5_2_1_Adder_12_U.b [1:0];
assign \add_5s_5s_5_2_1_U17.top_add_5s_5s_5_2_1_Adder_12_U.u1.cin  = 1'h0;
assign \add_5s_5s_5_2_1_U17.top_add_5s_5s_5_2_1_Adder_12_U.facout_s1  = \add_5s_5s_5_2_1_U17.top_add_5s_5s_5_2_1_Adder_12_U.u1.cout ;
assign \add_5s_5s_5_2_1_U17.top_add_5s_5s_5_2_1_Adder_12_U.fas_s1  = \add_5s_5s_5_2_1_U17.top_add_5s_5s_5_2_1_Adder_12_U.u1.s ;
assign \add_5s_5s_5_2_1_U17.top_add_5s_5s_5_2_1_Adder_12_U.a  = \add_5s_5s_5_2_1_U17.din0 ;
assign \add_5s_5s_5_2_1_U17.top_add_5s_5s_5_2_1_Adder_12_U.b  = \add_5s_5s_5_2_1_U17.din1 ;
assign \add_5s_5s_5_2_1_U17.top_add_5s_5s_5_2_1_Adder_12_U.ce  = \add_5s_5s_5_2_1_U17.ce ;
assign \add_5s_5s_5_2_1_U17.top_add_5s_5s_5_2_1_Adder_12_U.clk  = \add_5s_5s_5_2_1_U17.clk ;
assign \add_5s_5s_5_2_1_U17.top_add_5s_5s_5_2_1_Adder_12_U.reset  = \add_5s_5s_5_2_1_U17.reset ;
assign \add_5s_5s_5_2_1_U17.dout  = \add_5s_5s_5_2_1_U17.top_add_5s_5s_5_2_1_Adder_12_U.s ;
assign \add_5s_5s_5_2_1_U17.ce  = 1'h1;
assign \add_5s_5s_5_2_1_U17.clk  = ap_clk;
assign \add_5s_5s_5_2_1_U17.din0  = { ret_V_23_reg_2284[3], ret_V_23_reg_2284 };
assign \add_5s_5s_5_2_1_U17.din1  = { op_13[1], op_13[1], op_13[1], op_13 };
assign grp_fu_1428_p2 = \add_5s_5s_5_2_1_U17.dout ;
assign \add_5s_5s_5_2_1_U17.reset  = ap_rst;
assign \add_5ns_5s_5_2_1_U18.top_add_5ns_5s_5_2_1_Adder_13_U.ain_s0  = \add_5ns_5s_5_2_1_U18.top_add_5ns_5s_5_2_1_Adder_13_U.a ;
assign \add_5ns_5s_5_2_1_U18.top_add_5ns_5s_5_2_1_Adder_13_U.bin_s0  = \add_5ns_5s_5_2_1_U18.top_add_5ns_5s_5_2_1_Adder_13_U.b ;
assign \add_5ns_5s_5_2_1_U18.top_add_5ns_5s_5_2_1_Adder_13_U.s  = { \add_5ns_5s_5_2_1_U18.top_add_5ns_5s_5_2_1_Adder_13_U.fas_s2 , \add_5ns_5s_5_2_1_U18.top_add_5ns_5s_5_2_1_Adder_13_U.sum_s1  };
assign \add_5ns_5s_5_2_1_U18.top_add_5ns_5s_5_2_1_Adder_13_U.u2.a  = \add_5ns_5s_5_2_1_U18.top_add_5ns_5s_5_2_1_Adder_13_U.ain_s1 ;
assign \add_5ns_5s_5_2_1_U18.top_add_5ns_5s_5_2_1_Adder_13_U.u2.b  = \add_5ns_5s_5_2_1_U18.top_add_5ns_5s_5_2_1_Adder_13_U.bin_s1 ;
assign \add_5ns_5s_5_2_1_U18.top_add_5ns_5s_5_2_1_Adder_13_U.u2.cin  = \add_5ns_5s_5_2_1_U18.top_add_5ns_5s_5_2_1_Adder_13_U.carry_s1 ;
assign \add_5ns_5s_5_2_1_U18.top_add_5ns_5s_5_2_1_Adder_13_U.facout_s2  = \add_5ns_5s_5_2_1_U18.top_add_5ns_5s_5_2_1_Adder_13_U.u2.cout ;
assign \add_5ns_5s_5_2_1_U18.top_add_5ns_5s_5_2_1_Adder_13_U.fas_s2  = \add_5ns_5s_5_2_1_U18.top_add_5ns_5s_5_2_1_Adder_13_U.u2.s ;
assign \add_5ns_5s_5_2_1_U18.top_add_5ns_5s_5_2_1_Adder_13_U.u1.a  = \add_5ns_5s_5_2_1_U18.top_add_5ns_5s_5_2_1_Adder_13_U.a [1:0];
assign \add_5ns_5s_5_2_1_U18.top_add_5ns_5s_5_2_1_Adder_13_U.u1.b  = \add_5ns_5s_5_2_1_U18.top_add_5ns_5s_5_2_1_Adder_13_U.b [1:0];
assign \add_5ns_5s_5_2_1_U18.top_add_5ns_5s_5_2_1_Adder_13_U.u1.cin  = 1'h0;
assign \add_5ns_5s_5_2_1_U18.top_add_5ns_5s_5_2_1_Adder_13_U.facout_s1  = \add_5ns_5s_5_2_1_U18.top_add_5ns_5s_5_2_1_Adder_13_U.u1.cout ;
assign \add_5ns_5s_5_2_1_U18.top_add_5ns_5s_5_2_1_Adder_13_U.fas_s1  = \add_5ns_5s_5_2_1_U18.top_add_5ns_5s_5_2_1_Adder_13_U.u1.s ;
assign \add_5ns_5s_5_2_1_U18.top_add_5ns_5s_5_2_1_Adder_13_U.a  = \add_5ns_5s_5_2_1_U18.din0 ;
assign \add_5ns_5s_5_2_1_U18.top_add_5ns_5s_5_2_1_Adder_13_U.b  = \add_5ns_5s_5_2_1_U18.din1 ;
assign \add_5ns_5s_5_2_1_U18.top_add_5ns_5s_5_2_1_Adder_13_U.ce  = \add_5ns_5s_5_2_1_U18.ce ;
assign \add_5ns_5s_5_2_1_U18.top_add_5ns_5s_5_2_1_Adder_13_U.clk  = \add_5ns_5s_5_2_1_U18.clk ;
assign \add_5ns_5s_5_2_1_U18.top_add_5ns_5s_5_2_1_Adder_13_U.reset  = \add_5ns_5s_5_2_1_U18.reset ;
assign \add_5ns_5s_5_2_1_U18.dout  = \add_5ns_5s_5_2_1_U18.top_add_5ns_5s_5_2_1_Adder_13_U.s ;
assign \add_5ns_5s_5_2_1_U18.ce  = 1'h1;
assign \add_5ns_5s_5_2_1_U18.clk  = ap_clk;
assign \add_5ns_5s_5_2_1_U18.din0  = add_ln69_reg_2373;
assign \add_5ns_5s_5_2_1_U18.din1  = { ret_V_19_reg_2368[3], ret_V_19_reg_2368 };
assign grp_fu_1558_p2 = \add_5ns_5s_5_2_1_U18.dout ;
assign \add_5ns_5s_5_2_1_U18.reset  = ap_rst;
assign \add_4s_4ns_4_2_1_U16.top_add_4s_4ns_4_2_1_Adder_11_U.ain_s0  = \add_4s_4ns_4_2_1_U16.top_add_4s_4ns_4_2_1_Adder_11_U.a ;
assign \add_4s_4ns_4_2_1_U16.top_add_4s_4ns_4_2_1_Adder_11_U.bin_s0  = \add_4s_4ns_4_2_1_U16.top_add_4s_4ns_4_2_1_Adder_11_U.b ;
assign \add_4s_4ns_4_2_1_U16.top_add_4s_4ns_4_2_1_Adder_11_U.s  = { \add_4s_4ns_4_2_1_U16.top_add_4s_4ns_4_2_1_Adder_11_U.fas_s2 , \add_4s_4ns_4_2_1_U16.top_add_4s_4ns_4_2_1_Adder_11_U.sum_s1  };
assign \add_4s_4ns_4_2_1_U16.top_add_4s_4ns_4_2_1_Adder_11_U.u2.a  = \add_4s_4ns_4_2_1_U16.top_add_4s_4ns_4_2_1_Adder_11_U.ain_s1 ;
assign \add_4s_4ns_4_2_1_U16.top_add_4s_4ns_4_2_1_Adder_11_U.u2.b  = \add_4s_4ns_4_2_1_U16.top_add_4s_4ns_4_2_1_Adder_11_U.bin_s1 ;
assign \add_4s_4ns_4_2_1_U16.top_add_4s_4ns_4_2_1_Adder_11_U.u2.cin  = \add_4s_4ns_4_2_1_U16.top_add_4s_4ns_4_2_1_Adder_11_U.carry_s1 ;
assign \add_4s_4ns_4_2_1_U16.top_add_4s_4ns_4_2_1_Adder_11_U.facout_s2  = \add_4s_4ns_4_2_1_U16.top_add_4s_4ns_4_2_1_Adder_11_U.u2.cout ;
assign \add_4s_4ns_4_2_1_U16.top_add_4s_4ns_4_2_1_Adder_11_U.fas_s2  = \add_4s_4ns_4_2_1_U16.top_add_4s_4ns_4_2_1_Adder_11_U.u2.s ;
assign \add_4s_4ns_4_2_1_U16.top_add_4s_4ns_4_2_1_Adder_11_U.u1.a  = \add_4s_4ns_4_2_1_U16.top_add_4s_4ns_4_2_1_Adder_11_U.a [1:0];
assign \add_4s_4ns_4_2_1_U16.top_add_4s_4ns_4_2_1_Adder_11_U.u1.b  = \add_4s_4ns_4_2_1_U16.top_add_4s_4ns_4_2_1_Adder_11_U.b [1:0];
assign \add_4s_4ns_4_2_1_U16.top_add_4s_4ns_4_2_1_Adder_11_U.u1.cin  = 1'h0;
assign \add_4s_4ns_4_2_1_U16.top_add_4s_4ns_4_2_1_Adder_11_U.facout_s1  = \add_4s_4ns_4_2_1_U16.top_add_4s_4ns_4_2_1_Adder_11_U.u1.cout ;
assign \add_4s_4ns_4_2_1_U16.top_add_4s_4ns_4_2_1_Adder_11_U.fas_s1  = \add_4s_4ns_4_2_1_U16.top_add_4s_4ns_4_2_1_Adder_11_U.u1.s ;
assign \add_4s_4ns_4_2_1_U16.top_add_4s_4ns_4_2_1_Adder_11_U.a  = \add_4s_4ns_4_2_1_U16.din0 ;
assign \add_4s_4ns_4_2_1_U16.top_add_4s_4ns_4_2_1_Adder_11_U.b  = \add_4s_4ns_4_2_1_U16.din1 ;
assign \add_4s_4ns_4_2_1_U16.top_add_4s_4ns_4_2_1_Adder_11_U.ce  = \add_4s_4ns_4_2_1_U16.ce ;
assign \add_4s_4ns_4_2_1_U16.top_add_4s_4ns_4_2_1_Adder_11_U.clk  = \add_4s_4ns_4_2_1_U16.clk ;
assign \add_4s_4ns_4_2_1_U16.top_add_4s_4ns_4_2_1_Adder_11_U.reset  = \add_4s_4ns_4_2_1_U16.reset ;
assign \add_4s_4ns_4_2_1_U16.dout  = \add_4s_4ns_4_2_1_U16.top_add_4s_4ns_4_2_1_Adder_11_U.s ;
assign \add_4s_4ns_4_2_1_U16.ce  = 1'h1;
assign \add_4s_4ns_4_2_1_U16.clk  = ap_clk;
assign \add_4s_4ns_4_2_1_U16.din0  = { tmp_5_reg_2274[2], tmp_5_reg_2274 };
assign \add_4s_4ns_4_2_1_U16.din1  = 4'h1;
assign grp_fu_1367_p2 = \add_4s_4ns_4_2_1_U16.dout ;
assign \add_4s_4ns_4_2_1_U16.reset  = ap_rst;
assign \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_10_U.ain_s0  = \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_10_U.a ;
assign \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_10_U.bin_s0  = \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_10_U.b ;
assign \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_10_U.s  = { \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_10_U.fas_s2 , \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_10_U.sum_s1  };
assign \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_10_U.u2.a  = \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_10_U.ain_s1 ;
assign \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_10_U.u2.b  = \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_10_U.bin_s1 ;
assign \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_10_U.u2.cin  = \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_10_U.carry_s1 ;
assign \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_10_U.facout_s2  = \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_10_U.u2.cout ;
assign \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_10_U.fas_s2  = \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_10_U.u2.s ;
assign \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_10_U.u1.a  = \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_10_U.a [1:0];
assign \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_10_U.u1.b  = \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_10_U.b [1:0];
assign \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_10_U.u1.cin  = 1'h0;
assign \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_10_U.facout_s1  = \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_10_U.u1.cout ;
assign \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_10_U.fas_s1  = \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_10_U.u1.s ;
assign \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_10_U.a  = \add_4ns_4s_4_2_1_U14.din0 ;
assign \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_10_U.b  = \add_4ns_4s_4_2_1_U14.din1 ;
assign \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_10_U.ce  = \add_4ns_4s_4_2_1_U14.ce ;
assign \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_10_U.clk  = \add_4ns_4s_4_2_1_U14.clk ;
assign \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_10_U.reset  = \add_4ns_4s_4_2_1_U14.reset ;
assign \add_4ns_4s_4_2_1_U14.dout  = \add_4ns_4s_4_2_1_U14.top_add_4ns_4s_4_2_1_Adder_10_U.s ;
assign \add_4ns_4s_4_2_1_U14.ce  = 1'h1;
assign \add_4ns_4s_4_2_1_U14.clk  = ap_clk;
assign \add_4ns_4s_4_2_1_U14.din0  = { ret_V_15_reg_2178, 1'h0 };
assign \add_4ns_4s_4_2_1_U14.din1  = { op_12_V_reg_2172[1], op_12_V_reg_2172[1], op_12_V_reg_2172 };
assign grp_fu_1241_p2 = \add_4ns_4s_4_2_1_U14.dout ;
assign \add_4ns_4s_4_2_1_U14.reset  = ap_rst;
assign \add_4ns_4ns_4_2_1_U15.top_add_4ns_4ns_4_2_1_Adder_9_U.ain_s0  = \add_4ns_4ns_4_2_1_U15.top_add_4ns_4ns_4_2_1_Adder_9_U.a ;
assign \add_4ns_4ns_4_2_1_U15.top_add_4ns_4ns_4_2_1_Adder_9_U.bin_s0  = \add_4ns_4ns_4_2_1_U15.top_add_4ns_4ns_4_2_1_Adder_9_U.b ;
assign \add_4ns_4ns_4_2_1_U15.top_add_4ns_4ns_4_2_1_Adder_9_U.s  = { \add_4ns_4ns_4_2_1_U15.top_add_4ns_4ns_4_2_1_Adder_9_U.fas_s2 , \add_4ns_4ns_4_2_1_U15.top_add_4ns_4ns_4_2_1_Adder_9_U.sum_s1  };
assign \add_4ns_4ns_4_2_1_U15.top_add_4ns_4ns_4_2_1_Adder_9_U.u2.a  = \add_4ns_4ns_4_2_1_U15.top_add_4ns_4ns_4_2_1_Adder_9_U.ain_s1 ;
assign \add_4ns_4ns_4_2_1_U15.top_add_4ns_4ns_4_2_1_Adder_9_U.u2.b  = \add_4ns_4ns_4_2_1_U15.top_add_4ns_4ns_4_2_1_Adder_9_U.bin_s1 ;
assign \add_4ns_4ns_4_2_1_U15.top_add_4ns_4ns_4_2_1_Adder_9_U.u2.cin  = \add_4ns_4ns_4_2_1_U15.top_add_4ns_4ns_4_2_1_Adder_9_U.carry_s1 ;
assign \add_4ns_4ns_4_2_1_U15.top_add_4ns_4ns_4_2_1_Adder_9_U.facout_s2  = \add_4ns_4ns_4_2_1_U15.top_add_4ns_4ns_4_2_1_Adder_9_U.u2.cout ;
assign \add_4ns_4ns_4_2_1_U15.top_add_4ns_4ns_4_2_1_Adder_9_U.fas_s2  = \add_4ns_4ns_4_2_1_U15.top_add_4ns_4ns_4_2_1_Adder_9_U.u2.s ;
assign \add_4ns_4ns_4_2_1_U15.top_add_4ns_4ns_4_2_1_Adder_9_U.u1.a  = \add_4ns_4ns_4_2_1_U15.top_add_4ns_4ns_4_2_1_Adder_9_U.a [1:0];
assign \add_4ns_4ns_4_2_1_U15.top_add_4ns_4ns_4_2_1_Adder_9_U.u1.b  = \add_4ns_4ns_4_2_1_U15.top_add_4ns_4ns_4_2_1_Adder_9_U.b [1:0];
assign \add_4ns_4ns_4_2_1_U15.top_add_4ns_4ns_4_2_1_Adder_9_U.u1.cin  = 1'h0;
assign \add_4ns_4ns_4_2_1_U15.top_add_4ns_4ns_4_2_1_Adder_9_U.facout_s1  = \add_4ns_4ns_4_2_1_U15.top_add_4ns_4ns_4_2_1_Adder_9_U.u1.cout ;
assign \add_4ns_4ns_4_2_1_U15.top_add_4ns_4ns_4_2_1_Adder_9_U.fas_s1  = \add_4ns_4ns_4_2_1_U15.top_add_4ns_4ns_4_2_1_Adder_9_U.u1.s ;
assign \add_4ns_4ns_4_2_1_U15.top_add_4ns_4ns_4_2_1_Adder_9_U.a  = \add_4ns_4ns_4_2_1_U15.din0 ;
assign \add_4ns_4ns_4_2_1_U15.top_add_4ns_4ns_4_2_1_Adder_9_U.b  = \add_4ns_4ns_4_2_1_U15.din1 ;
assign \add_4ns_4ns_4_2_1_U15.top_add_4ns_4ns_4_2_1_Adder_9_U.ce  = \add_4ns_4ns_4_2_1_U15.ce ;
assign \add_4ns_4ns_4_2_1_U15.top_add_4ns_4ns_4_2_1_Adder_9_U.clk  = \add_4ns_4ns_4_2_1_U15.clk ;
assign \add_4ns_4ns_4_2_1_U15.top_add_4ns_4ns_4_2_1_Adder_9_U.reset  = \add_4ns_4ns_4_2_1_U15.reset ;
assign \add_4ns_4ns_4_2_1_U15.dout  = \add_4ns_4ns_4_2_1_U15.top_add_4ns_4ns_4_2_1_Adder_9_U.s ;
assign \add_4ns_4ns_4_2_1_U15.ce  = 1'h1;
assign \add_4ns_4ns_4_2_1_U15.clk  = ap_clk;
assign \add_4ns_4ns_4_2_1_U15.din0  = p_Val2_12_reg_2117;
assign \add_4ns_4ns_4_2_1_U15.din1  = { 3'h0, and_ln408_reg_2234 };
assign grp_fu_1276_p2 = \add_4ns_4ns_4_2_1_U15.dout ;
assign \add_4ns_4ns_4_2_1_U15.reset  = ap_rst;
assign \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_9_U.ain_s0  = \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_9_U.a ;
assign \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_9_U.bin_s0  = \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_9_U.b ;
assign \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_9_U.s  = { \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_9_U.fas_s2 , \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_9_U.sum_s1  };
assign \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_9_U.u2.a  = \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_9_U.ain_s1 ;
assign \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_9_U.u2.b  = \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_9_U.bin_s1 ;
assign \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_9_U.u2.cin  = \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_9_U.carry_s1 ;
assign \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_9_U.facout_s2  = \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_9_U.u2.cout ;
assign \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_9_U.fas_s2  = \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_9_U.u2.s ;
assign \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_9_U.u1.a  = \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_9_U.a [1:0];
assign \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_9_U.u1.b  = \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_9_U.b [1:0];
assign \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_9_U.u1.cin  = 1'h0;
assign \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_9_U.facout_s1  = \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_9_U.u1.cout ;
assign \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_9_U.fas_s1  = \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_9_U.u1.s ;
assign \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_9_U.a  = \add_4ns_4ns_4_2_1_U13.din0 ;
assign \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_9_U.b  = \add_4ns_4ns_4_2_1_U13.din1 ;
assign \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_9_U.ce  = \add_4ns_4ns_4_2_1_U13.ce ;
assign \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_9_U.clk  = \add_4ns_4ns_4_2_1_U13.clk ;
assign \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_9_U.reset  = \add_4ns_4ns_4_2_1_U13.reset ;
assign \add_4ns_4ns_4_2_1_U13.dout  = \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_9_U.s ;
assign \add_4ns_4ns_4_2_1_U13.ce  = 1'h1;
assign \add_4ns_4ns_4_2_1_U13.clk  = ap_clk;
assign \add_4ns_4ns_4_2_1_U13.din0  = ret_V_7_cast_reg_2160;
assign \add_4ns_4ns_4_2_1_U13.din1  = 4'h1;
assign grp_fu_1188_p2 = \add_4ns_4ns_4_2_1_U13.dout ;
assign \add_4ns_4ns_4_2_1_U13.reset  = ap_rst;
assign \add_4ns_4ns_4_2_1_U12.top_add_4ns_4ns_4_2_1_Adder_9_U.ain_s0  = \add_4ns_4ns_4_2_1_U12.top_add_4ns_4ns_4_2_1_Adder_9_U.a ;
assign \add_4ns_4ns_4_2_1_U12.top_add_4ns_4ns_4_2_1_Adder_9_U.bin_s0  = \add_4ns_4ns_4_2_1_U12.top_add_4ns_4ns_4_2_1_Adder_9_U.b ;
assign \add_4ns_4ns_4_2_1_U12.top_add_4ns_4ns_4_2_1_Adder_9_U.s  = { \add_4ns_4ns_4_2_1_U12.top_add_4ns_4ns_4_2_1_Adder_9_U.fas_s2 , \add_4ns_4ns_4_2_1_U12.top_add_4ns_4ns_4_2_1_Adder_9_U.sum_s1  };
assign \add_4ns_4ns_4_2_1_U12.top_add_4ns_4ns_4_2_1_Adder_9_U.u2.a  = \add_4ns_4ns_4_2_1_U12.top_add_4ns_4ns_4_2_1_Adder_9_U.ain_s1 ;
assign \add_4ns_4ns_4_2_1_U12.top_add_4ns_4ns_4_2_1_Adder_9_U.u2.b  = \add_4ns_4ns_4_2_1_U12.top_add_4ns_4ns_4_2_1_Adder_9_U.bin_s1 ;
assign \add_4ns_4ns_4_2_1_U12.top_add_4ns_4ns_4_2_1_Adder_9_U.u2.cin  = \add_4ns_4ns_4_2_1_U12.top_add_4ns_4ns_4_2_1_Adder_9_U.carry_s1 ;
assign \add_4ns_4ns_4_2_1_U12.top_add_4ns_4ns_4_2_1_Adder_9_U.facout_s2  = \add_4ns_4ns_4_2_1_U12.top_add_4ns_4ns_4_2_1_Adder_9_U.u2.cout ;
assign \add_4ns_4ns_4_2_1_U12.top_add_4ns_4ns_4_2_1_Adder_9_U.fas_s2  = \add_4ns_4ns_4_2_1_U12.top_add_4ns_4ns_4_2_1_Adder_9_U.u2.s ;
assign \add_4ns_4ns_4_2_1_U12.top_add_4ns_4ns_4_2_1_Adder_9_U.u1.a  = \add_4ns_4ns_4_2_1_U12.top_add_4ns_4ns_4_2_1_Adder_9_U.a [1:0];
assign \add_4ns_4ns_4_2_1_U12.top_add_4ns_4ns_4_2_1_Adder_9_U.u1.b  = \add_4ns_4ns_4_2_1_U12.top_add_4ns_4ns_4_2_1_Adder_9_U.b [1:0];
assign \add_4ns_4ns_4_2_1_U12.top_add_4ns_4ns_4_2_1_Adder_9_U.u1.cin  = 1'h0;
assign \add_4ns_4ns_4_2_1_U12.top_add_4ns_4ns_4_2_1_Adder_9_U.facout_s1  = \add_4ns_4ns_4_2_1_U12.top_add_4ns_4ns_4_2_1_Adder_9_U.u1.cout ;
assign \add_4ns_4ns_4_2_1_U12.top_add_4ns_4ns_4_2_1_Adder_9_U.fas_s1  = \add_4ns_4ns_4_2_1_U12.top_add_4ns_4ns_4_2_1_Adder_9_U.u1.s ;
assign \add_4ns_4ns_4_2_1_U12.top_add_4ns_4ns_4_2_1_Adder_9_U.a  = \add_4ns_4ns_4_2_1_U12.din0 ;
assign \add_4ns_4ns_4_2_1_U12.top_add_4ns_4ns_4_2_1_Adder_9_U.b  = \add_4ns_4ns_4_2_1_U12.din1 ;
assign \add_4ns_4ns_4_2_1_U12.top_add_4ns_4ns_4_2_1_Adder_9_U.ce  = \add_4ns_4ns_4_2_1_U12.ce ;
assign \add_4ns_4ns_4_2_1_U12.top_add_4ns_4ns_4_2_1_Adder_9_U.clk  = \add_4ns_4ns_4_2_1_U12.clk ;
assign \add_4ns_4ns_4_2_1_U12.top_add_4ns_4ns_4_2_1_Adder_9_U.reset  = \add_4ns_4ns_4_2_1_U12.reset ;
assign \add_4ns_4ns_4_2_1_U12.dout  = \add_4ns_4ns_4_2_1_U12.top_add_4ns_4ns_4_2_1_Adder_9_U.s ;
assign \add_4ns_4ns_4_2_1_U12.ce  = 1'h1;
assign \add_4ns_4ns_4_2_1_U12.clk  = ap_clk;
assign \add_4ns_4ns_4_2_1_U12.din0  = ret_V_reg_2143;
assign \add_4ns_4ns_4_2_1_U12.din1  = 4'h1;
assign grp_fu_1178_p2 = \add_4ns_4ns_4_2_1_U12.dout ;
assign \add_4ns_4ns_4_2_1_U12.reset  = ap_rst;
assign \add_3s_3ns_3_2_1_U11.top_add_3s_3ns_3_2_1_Adder_8_U.ain_s0  = \add_3s_3ns_3_2_1_U11.top_add_3s_3ns_3_2_1_Adder_8_U.a ;
assign \add_3s_3ns_3_2_1_U11.top_add_3s_3ns_3_2_1_Adder_8_U.bin_s0  = \add_3s_3ns_3_2_1_U11.top_add_3s_3ns_3_2_1_Adder_8_U.b ;
assign \add_3s_3ns_3_2_1_U11.top_add_3s_3ns_3_2_1_Adder_8_U.s  = { \add_3s_3ns_3_2_1_U11.top_add_3s_3ns_3_2_1_Adder_8_U.fas_s2 , \add_3s_3ns_3_2_1_U11.top_add_3s_3ns_3_2_1_Adder_8_U.sum_s1  };
assign \add_3s_3ns_3_2_1_U11.top_add_3s_3ns_3_2_1_Adder_8_U.u2.a  = \add_3s_3ns_3_2_1_U11.top_add_3s_3ns_3_2_1_Adder_8_U.ain_s1 ;
assign \add_3s_3ns_3_2_1_U11.top_add_3s_3ns_3_2_1_Adder_8_U.u2.b  = \add_3s_3ns_3_2_1_U11.top_add_3s_3ns_3_2_1_Adder_8_U.bin_s1 ;
assign \add_3s_3ns_3_2_1_U11.top_add_3s_3ns_3_2_1_Adder_8_U.u2.cin  = \add_3s_3ns_3_2_1_U11.top_add_3s_3ns_3_2_1_Adder_8_U.carry_s1 ;
assign \add_3s_3ns_3_2_1_U11.top_add_3s_3ns_3_2_1_Adder_8_U.facout_s2  = \add_3s_3ns_3_2_1_U11.top_add_3s_3ns_3_2_1_Adder_8_U.u2.cout ;
assign \add_3s_3ns_3_2_1_U11.top_add_3s_3ns_3_2_1_Adder_8_U.fas_s2  = \add_3s_3ns_3_2_1_U11.top_add_3s_3ns_3_2_1_Adder_8_U.u2.s ;
assign \add_3s_3ns_3_2_1_U11.top_add_3s_3ns_3_2_1_Adder_8_U.u1.a  = \add_3s_3ns_3_2_1_U11.top_add_3s_3ns_3_2_1_Adder_8_U.a [0];
assign \add_3s_3ns_3_2_1_U11.top_add_3s_3ns_3_2_1_Adder_8_U.u1.b  = \add_3s_3ns_3_2_1_U11.top_add_3s_3ns_3_2_1_Adder_8_U.b [0];
assign \add_3s_3ns_3_2_1_U11.top_add_3s_3ns_3_2_1_Adder_8_U.u1.cin  = 1'h0;
assign \add_3s_3ns_3_2_1_U11.top_add_3s_3ns_3_2_1_Adder_8_U.facout_s1  = \add_3s_3ns_3_2_1_U11.top_add_3s_3ns_3_2_1_Adder_8_U.u1.cout ;
assign \add_3s_3ns_3_2_1_U11.top_add_3s_3ns_3_2_1_Adder_8_U.fas_s1  = \add_3s_3ns_3_2_1_U11.top_add_3s_3ns_3_2_1_Adder_8_U.u1.s ;
assign \add_3s_3ns_3_2_1_U11.top_add_3s_3ns_3_2_1_Adder_8_U.a  = \add_3s_3ns_3_2_1_U11.din0 ;
assign \add_3s_3ns_3_2_1_U11.top_add_3s_3ns_3_2_1_Adder_8_U.b  = \add_3s_3ns_3_2_1_U11.din1 ;
assign \add_3s_3ns_3_2_1_U11.top_add_3s_3ns_3_2_1_Adder_8_U.ce  = \add_3s_3ns_3_2_1_U11.ce ;
assign \add_3s_3ns_3_2_1_U11.top_add_3s_3ns_3_2_1_Adder_8_U.clk  = \add_3s_3ns_3_2_1_U11.clk ;
assign \add_3s_3ns_3_2_1_U11.top_add_3s_3ns_3_2_1_Adder_8_U.reset  = \add_3s_3ns_3_2_1_U11.reset ;
assign \add_3s_3ns_3_2_1_U11.dout  = \add_3s_3ns_3_2_1_U11.top_add_3s_3ns_3_2_1_Adder_8_U.s ;
assign \add_3s_3ns_3_2_1_U11.ce  = 1'h1;
assign \add_3s_3ns_3_2_1_U11.clk  = ap_clk;
assign \add_3s_3ns_3_2_1_U11.din0  = { op_9[1], op_9 };
assign \add_3s_3ns_3_2_1_U11.din1  = select_ln703_reg_2012;
assign grp_fu_1024_p2 = \add_3s_3ns_3_2_1_U11.dout ;
assign \add_3s_3ns_3_2_1_U11.reset  = ap_rst;
assign \add_39s_39s_39_2_1_U21.top_add_39s_39s_39_2_1_Adder_16_U.ain_s0  = \add_39s_39s_39_2_1_U21.top_add_39s_39s_39_2_1_Adder_16_U.a ;
assign \add_39s_39s_39_2_1_U21.top_add_39s_39s_39_2_1_Adder_16_U.bin_s0  = \add_39s_39s_39_2_1_U21.top_add_39s_39s_39_2_1_Adder_16_U.b ;
assign \add_39s_39s_39_2_1_U21.top_add_39s_39s_39_2_1_Adder_16_U.s  = { \add_39s_39s_39_2_1_U21.top_add_39s_39s_39_2_1_Adder_16_U.fas_s2 , \add_39s_39s_39_2_1_U21.top_add_39s_39s_39_2_1_Adder_16_U.sum_s1  };
assign \add_39s_39s_39_2_1_U21.top_add_39s_39s_39_2_1_Adder_16_U.u2.a  = \add_39s_39s_39_2_1_U21.top_add_39s_39s_39_2_1_Adder_16_U.ain_s1 ;
assign \add_39s_39s_39_2_1_U21.top_add_39s_39s_39_2_1_Adder_16_U.u2.b  = \add_39s_39s_39_2_1_U21.top_add_39s_39s_39_2_1_Adder_16_U.bin_s1 ;
assign \add_39s_39s_39_2_1_U21.top_add_39s_39s_39_2_1_Adder_16_U.u2.cin  = \add_39s_39s_39_2_1_U21.top_add_39s_39s_39_2_1_Adder_16_U.carry_s1 ;
assign \add_39s_39s_39_2_1_U21.top_add_39s_39s_39_2_1_Adder_16_U.facout_s2  = \add_39s_39s_39_2_1_U21.top_add_39s_39s_39_2_1_Adder_16_U.u2.cout ;
assign \add_39s_39s_39_2_1_U21.top_add_39s_39s_39_2_1_Adder_16_U.fas_s2  = \add_39s_39s_39_2_1_U21.top_add_39s_39s_39_2_1_Adder_16_U.u2.s ;
assign \add_39s_39s_39_2_1_U21.top_add_39s_39s_39_2_1_Adder_16_U.u1.a  = \add_39s_39s_39_2_1_U21.top_add_39s_39s_39_2_1_Adder_16_U.a [18:0];
assign \add_39s_39s_39_2_1_U21.top_add_39s_39s_39_2_1_Adder_16_U.u1.b  = \add_39s_39s_39_2_1_U21.top_add_39s_39s_39_2_1_Adder_16_U.b [18:0];
assign \add_39s_39s_39_2_1_U21.top_add_39s_39s_39_2_1_Adder_16_U.u1.cin  = 1'h0;
assign \add_39s_39s_39_2_1_U21.top_add_39s_39s_39_2_1_Adder_16_U.facout_s1  = \add_39s_39s_39_2_1_U21.top_add_39s_39s_39_2_1_Adder_16_U.u1.cout ;
assign \add_39s_39s_39_2_1_U21.top_add_39s_39s_39_2_1_Adder_16_U.fas_s1  = \add_39s_39s_39_2_1_U21.top_add_39s_39s_39_2_1_Adder_16_U.u1.s ;
assign \add_39s_39s_39_2_1_U21.top_add_39s_39s_39_2_1_Adder_16_U.a  = \add_39s_39s_39_2_1_U21.din0 ;
assign \add_39s_39s_39_2_1_U21.top_add_39s_39s_39_2_1_Adder_16_U.b  = \add_39s_39s_39_2_1_U21.din1 ;
assign \add_39s_39s_39_2_1_U21.top_add_39s_39s_39_2_1_Adder_16_U.ce  = \add_39s_39s_39_2_1_U21.ce ;
assign \add_39s_39s_39_2_1_U21.top_add_39s_39s_39_2_1_Adder_16_U.clk  = \add_39s_39s_39_2_1_U21.clk ;
assign \add_39s_39s_39_2_1_U21.top_add_39s_39s_39_2_1_Adder_16_U.reset  = \add_39s_39s_39_2_1_U21.reset ;
assign \add_39s_39s_39_2_1_U21.dout  = \add_39s_39s_39_2_1_U21.top_add_39s_39s_39_2_1_Adder_16_U.s ;
assign \add_39s_39s_39_2_1_U21.ce  = 1'h1;
assign \add_39s_39s_39_2_1_U21.clk  = ap_clk;
assign \add_39s_39s_39_2_1_U21.din0  = { op_25_V_reg_2423[5], op_25_V_reg_2423[5], op_25_V_reg_2423[5], op_25_V_reg_2423[5], op_25_V_reg_2423[5], op_25_V_reg_2423[5], op_25_V_reg_2423[5], op_25_V_reg_2423[5], op_25_V_reg_2423[5], op_25_V_reg_2423[5], op_25_V_reg_2423[5], op_25_V_reg_2423[5], op_25_V_reg_2423[5], op_25_V_reg_2423[5], op_25_V_reg_2423[5], op_25_V_reg_2423[5], op_25_V_reg_2423[5], op_25_V_reg_2423[5], op_25_V_reg_2423[5], op_25_V_reg_2423[5], op_25_V_reg_2423[5], op_25_V_reg_2423[5], op_25_V_reg_2423[5], op_25_V_reg_2423[5], op_25_V_reg_2423[5], op_25_V_reg_2423[5], op_25_V_reg_2423[5], op_25_V_reg_2423, 6'h00 };
assign \add_39s_39s_39_2_1_U21.din1  = { op_17_V_reg_2313[7], op_17_V_reg_2313[7], op_17_V_reg_2313[7], op_17_V_reg_2313[7], op_17_V_reg_2313[7], op_17_V_reg_2313[7], op_17_V_reg_2313[7], op_17_V_reg_2313[7], op_17_V_reg_2313[7], op_17_V_reg_2313[7], op_17_V_reg_2313[7], op_17_V_reg_2313[7], op_17_V_reg_2313[7], op_17_V_reg_2313[7], op_17_V_reg_2313[7], op_17_V_reg_2313[7], op_17_V_reg_2313[7], op_17_V_reg_2313[7], op_17_V_reg_2313[7], op_17_V_reg_2313[7], op_17_V_reg_2313[7], op_17_V_reg_2313[7], op_17_V_reg_2313[7], op_17_V_reg_2313[7], op_17_V_reg_2313[7], op_17_V_reg_2313[7], op_17_V_reg_2313[7], op_17_V_reg_2313[7], op_17_V_reg_2313[7], op_17_V_reg_2313[7], op_17_V_reg_2313[7], op_17_V_reg_2313 };
assign grp_fu_1610_p2 = \add_39s_39s_39_2_1_U21.dout ;
assign \add_39s_39s_39_2_1_U21.reset  = ap_rst;
assign \add_33s_33s_33_2_1_U8.top_add_33s_33s_33_2_1_Adder_5_U.ain_s0  = \add_33s_33s_33_2_1_U8.top_add_33s_33s_33_2_1_Adder_5_U.a ;
assign \add_33s_33s_33_2_1_U8.top_add_33s_33s_33_2_1_Adder_5_U.bin_s0  = \add_33s_33s_33_2_1_U8.top_add_33s_33s_33_2_1_Adder_5_U.b ;
assign \add_33s_33s_33_2_1_U8.top_add_33s_33s_33_2_1_Adder_5_U.s  = { \add_33s_33s_33_2_1_U8.top_add_33s_33s_33_2_1_Adder_5_U.fas_s2 , \add_33s_33s_33_2_1_U8.top_add_33s_33s_33_2_1_Adder_5_U.sum_s1  };
assign \add_33s_33s_33_2_1_U8.top_add_33s_33s_33_2_1_Adder_5_U.u2.a  = \add_33s_33s_33_2_1_U8.top_add_33s_33s_33_2_1_Adder_5_U.ain_s1 ;
assign \add_33s_33s_33_2_1_U8.top_add_33s_33s_33_2_1_Adder_5_U.u2.b  = \add_33s_33s_33_2_1_U8.top_add_33s_33s_33_2_1_Adder_5_U.bin_s1 ;
assign \add_33s_33s_33_2_1_U8.top_add_33s_33s_33_2_1_Adder_5_U.u2.cin  = \add_33s_33s_33_2_1_U8.top_add_33s_33s_33_2_1_Adder_5_U.carry_s1 ;
assign \add_33s_33s_33_2_1_U8.top_add_33s_33s_33_2_1_Adder_5_U.facout_s2  = \add_33s_33s_33_2_1_U8.top_add_33s_33s_33_2_1_Adder_5_U.u2.cout ;
assign \add_33s_33s_33_2_1_U8.top_add_33s_33s_33_2_1_Adder_5_U.fas_s2  = \add_33s_33s_33_2_1_U8.top_add_33s_33s_33_2_1_Adder_5_U.u2.s ;
assign \add_33s_33s_33_2_1_U8.top_add_33s_33s_33_2_1_Adder_5_U.u1.a  = \add_33s_33s_33_2_1_U8.top_add_33s_33s_33_2_1_Adder_5_U.a [15:0];
assign \add_33s_33s_33_2_1_U8.top_add_33s_33s_33_2_1_Adder_5_U.u1.b  = \add_33s_33s_33_2_1_U8.top_add_33s_33s_33_2_1_Adder_5_U.b [15:0];
assign \add_33s_33s_33_2_1_U8.top_add_33s_33s_33_2_1_Adder_5_U.u1.cin  = 1'h0;
assign \add_33s_33s_33_2_1_U8.top_add_33s_33s_33_2_1_Adder_5_U.facout_s1  = \add_33s_33s_33_2_1_U8.top_add_33s_33s_33_2_1_Adder_5_U.u1.cout ;
assign \add_33s_33s_33_2_1_U8.top_add_33s_33s_33_2_1_Adder_5_U.fas_s1  = \add_33s_33s_33_2_1_U8.top_add_33s_33s_33_2_1_Adder_5_U.u1.s ;
assign \add_33s_33s_33_2_1_U8.top_add_33s_33s_33_2_1_Adder_5_U.a  = \add_33s_33s_33_2_1_U8.din0 ;
assign \add_33s_33s_33_2_1_U8.top_add_33s_33s_33_2_1_Adder_5_U.b  = \add_33s_33s_33_2_1_U8.din1 ;
assign \add_33s_33s_33_2_1_U8.top_add_33s_33s_33_2_1_Adder_5_U.ce  = \add_33s_33s_33_2_1_U8.ce ;
assign \add_33s_33s_33_2_1_U8.top_add_33s_33s_33_2_1_Adder_5_U.clk  = \add_33s_33s_33_2_1_U8.clk ;
assign \add_33s_33s_33_2_1_U8.top_add_33s_33s_33_2_1_Adder_5_U.reset  = \add_33s_33s_33_2_1_U8.reset ;
assign \add_33s_33s_33_2_1_U8.dout  = \add_33s_33s_33_2_1_U8.top_add_33s_33s_33_2_1_Adder_5_U.s ;
assign \add_33s_33s_33_2_1_U8.ce  = 1'h1;
assign \add_33s_33s_33_2_1_U8.clk  = ap_clk;
assign \add_33s_33s_33_2_1_U8.din0  = { op_3_V_reg_1816[3], op_3_V_reg_1816[3], op_3_V_reg_1816[3], op_3_V_reg_1816[3], op_3_V_reg_1816[3], op_3_V_reg_1816[3], op_3_V_reg_1816, 23'h000000 };
assign \add_33s_33s_33_2_1_U8.din1  = { op_6[31], op_6 };
assign grp_fu_838_p2 = \add_33s_33s_33_2_1_U8.dout ;
assign \add_33s_33s_33_2_1_U8.reset  = ap_rst;
assign \add_32s_32ns_32_2_1_U24.top_add_32s_32ns_32_2_1_Adder_19_U.ain_s0  = \add_32s_32ns_32_2_1_U24.top_add_32s_32ns_32_2_1_Adder_19_U.a ;
assign \add_32s_32ns_32_2_1_U24.top_add_32s_32ns_32_2_1_Adder_19_U.bin_s0  = \add_32s_32ns_32_2_1_U24.top_add_32s_32ns_32_2_1_Adder_19_U.b ;
assign \add_32s_32ns_32_2_1_U24.top_add_32s_32ns_32_2_1_Adder_19_U.s  = { \add_32s_32ns_32_2_1_U24.top_add_32s_32ns_32_2_1_Adder_19_U.fas_s2 , \add_32s_32ns_32_2_1_U24.top_add_32s_32ns_32_2_1_Adder_19_U.sum_s1  };
assign \add_32s_32ns_32_2_1_U24.top_add_32s_32ns_32_2_1_Adder_19_U.u2.a  = \add_32s_32ns_32_2_1_U24.top_add_32s_32ns_32_2_1_Adder_19_U.ain_s1 ;
assign \add_32s_32ns_32_2_1_U24.top_add_32s_32ns_32_2_1_Adder_19_U.u2.b  = \add_32s_32ns_32_2_1_U24.top_add_32s_32ns_32_2_1_Adder_19_U.bin_s1 ;
assign \add_32s_32ns_32_2_1_U24.top_add_32s_32ns_32_2_1_Adder_19_U.u2.cin  = \add_32s_32ns_32_2_1_U24.top_add_32s_32ns_32_2_1_Adder_19_U.carry_s1 ;
assign \add_32s_32ns_32_2_1_U24.top_add_32s_32ns_32_2_1_Adder_19_U.facout_s2  = \add_32s_32ns_32_2_1_U24.top_add_32s_32ns_32_2_1_Adder_19_U.u2.cout ;
assign \add_32s_32ns_32_2_1_U24.top_add_32s_32ns_32_2_1_Adder_19_U.fas_s2  = \add_32s_32ns_32_2_1_U24.top_add_32s_32ns_32_2_1_Adder_19_U.u2.s ;
assign \add_32s_32ns_32_2_1_U24.top_add_32s_32ns_32_2_1_Adder_19_U.u1.a  = \add_32s_32ns_32_2_1_U24.top_add_32s_32ns_32_2_1_Adder_19_U.a [15:0];
assign \add_32s_32ns_32_2_1_U24.top_add_32s_32ns_32_2_1_Adder_19_U.u1.b  = \add_32s_32ns_32_2_1_U24.top_add_32s_32ns_32_2_1_Adder_19_U.b [15:0];
assign \add_32s_32ns_32_2_1_U24.top_add_32s_32ns_32_2_1_Adder_19_U.u1.cin  = 1'h0;
assign \add_32s_32ns_32_2_1_U24.top_add_32s_32ns_32_2_1_Adder_19_U.facout_s1  = \add_32s_32ns_32_2_1_U24.top_add_32s_32ns_32_2_1_Adder_19_U.u1.cout ;
assign \add_32s_32ns_32_2_1_U24.top_add_32s_32ns_32_2_1_Adder_19_U.fas_s1  = \add_32s_32ns_32_2_1_U24.top_add_32s_32ns_32_2_1_Adder_19_U.u1.s ;
assign \add_32s_32ns_32_2_1_U24.top_add_32s_32ns_32_2_1_Adder_19_U.a  = \add_32s_32ns_32_2_1_U24.din0 ;
assign \add_32s_32ns_32_2_1_U24.top_add_32s_32ns_32_2_1_Adder_19_U.b  = \add_32s_32ns_32_2_1_U24.din1 ;
assign \add_32s_32ns_32_2_1_U24.top_add_32s_32ns_32_2_1_Adder_19_U.ce  = \add_32s_32ns_32_2_1_U24.ce ;
assign \add_32s_32ns_32_2_1_U24.top_add_32s_32ns_32_2_1_Adder_19_U.clk  = \add_32s_32ns_32_2_1_U24.clk ;
assign \add_32s_32ns_32_2_1_U24.top_add_32s_32ns_32_2_1_Adder_19_U.reset  = \add_32s_32ns_32_2_1_U24.reset ;
assign \add_32s_32ns_32_2_1_U24.dout  = \add_32s_32ns_32_2_1_U24.top_add_32s_32ns_32_2_1_Adder_19_U.s ;
assign \add_32s_32ns_32_2_1_U24.ce  = 1'h1;
assign \add_32s_32ns_32_2_1_U24.clk  = ap_clk;
assign \add_32s_32ns_32_2_1_U24.din0  = { add_ln69_3_reg_2470[8], add_ln69_3_reg_2470[8], add_ln69_3_reg_2470[8], add_ln69_3_reg_2470[8], add_ln69_3_reg_2470[8], add_ln69_3_reg_2470[8], add_ln69_3_reg_2470[8], add_ln69_3_reg_2470[8], add_ln69_3_reg_2470[8], add_ln69_3_reg_2470[8], add_ln69_3_reg_2470[8], add_ln69_3_reg_2470[8], add_ln69_3_reg_2470[8], add_ln69_3_reg_2470[8], add_ln69_3_reg_2470[8], add_ln69_3_reg_2470[8], add_ln69_3_reg_2470[8], add_ln69_3_reg_2470[8], add_ln69_3_reg_2470[8], add_ln69_3_reg_2470[8], add_ln69_3_reg_2470[8], add_ln69_3_reg_2470[8], add_ln69_3_reg_2470[8], add_ln69_3_reg_2470 };
assign \add_32s_32ns_32_2_1_U24.din1  = ret_V_26_reg_2465;
assign grp_fu_1666_p2 = \add_32s_32ns_32_2_1_U24.dout ;
assign \add_32s_32ns_32_2_1_U24.reset  = ap_rst;
assign \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_17_U.ain_s0  = \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_17_U.a ;
assign \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_17_U.bin_s0  = \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_17_U.b ;
assign \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_17_U.s  = { \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_17_U.fas_s2 , \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_17_U.sum_s1  };
assign \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_17_U.u2.a  = \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_17_U.ain_s1 ;
assign \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_17_U.u2.b  = \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_17_U.bin_s1 ;
assign \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_17_U.u2.cin  = \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_17_U.carry_s1 ;
assign \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_17_U.facout_s2  = \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_17_U.u2.cout ;
assign \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_17_U.fas_s2  = \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_17_U.u2.s ;
assign \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_17_U.u1.a  = \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_17_U.a [15:0];
assign \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_17_U.u1.b  = \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_17_U.b [15:0];
assign \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_17_U.u1.cin  = 1'h0;
assign \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_17_U.facout_s1  = \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_17_U.u1.cout ;
assign \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_17_U.fas_s1  = \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_17_U.u1.s ;
assign \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_17_U.a  = \add_32ns_32ns_32_2_1_U22.din0 ;
assign \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_17_U.b  = \add_32ns_32ns_32_2_1_U22.din1 ;
assign \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_17_U.ce  = \add_32ns_32ns_32_2_1_U22.ce ;
assign \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_17_U.clk  = \add_32ns_32ns_32_2_1_U22.clk ;
assign \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_17_U.reset  = \add_32ns_32ns_32_2_1_U22.reset ;
assign \add_32ns_32ns_32_2_1_U22.dout  = \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_17_U.s ;
assign \add_32ns_32ns_32_2_1_U22.ce  = 1'h1;
assign \add_32ns_32ns_32_2_1_U22.clk  = ap_clk;
assign \add_32ns_32ns_32_2_1_U22.din0  = ret_V_20_cast_reg_2443;
assign \add_32ns_32ns_32_2_1_U22.din1  = 32'd1;
assign grp_fu_1626_p2 = \add_32ns_32ns_32_2_1_U22.dout ;
assign \add_32ns_32ns_32_2_1_U22.reset  = ap_rst;
assign \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_1_U.ain_s0  = \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_1_U.a ;
assign \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_1_U.bin_s0  = \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_1_U.b ;
assign \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_1_U.s  = { \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_1_U.fas_s2 , \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_1_U.sum_s1  };
assign \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.a  = \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_1_U.ain_s1 ;
assign \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.b  = \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_1_U.bin_s1 ;
assign \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.cin  = \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_1_U.carry_s1 ;
assign \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_1_U.facout_s2  = \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.cout ;
assign \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_1_U.fas_s2  = \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.s ;
assign \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.a  = \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_1_U.a [0];
assign \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.b  = \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_1_U.b [0];
assign \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.cin  = 1'h0;
assign \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_1_U.facout_s1  = \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.cout ;
assign \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_1_U.fas_s1  = \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.s ;
assign \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_1_U.a  = \add_2ns_2ns_2_2_1_U4.din0 ;
assign \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_1_U.b  = \add_2ns_2ns_2_2_1_U4.din1 ;
assign \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_1_U.ce  = \add_2ns_2ns_2_2_1_U4.ce ;
assign \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_1_U.clk  = \add_2ns_2ns_2_2_1_U4.clk ;
assign \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_1_U.reset  = \add_2ns_2ns_2_2_1_U4.reset ;
assign \add_2ns_2ns_2_2_1_U4.dout  = \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_1_U.s ;
assign \add_2ns_2ns_2_2_1_U4.ce  = 1'h1;
assign \add_2ns_2ns_2_2_1_U4.clk  = ap_clk;
assign \add_2ns_2ns_2_2_1_U4.din0  = p_Val2_2_reg_1763;
assign \add_2ns_2ns_2_2_1_U4.din1  = { 1'h0, and_ln414_reg_1811 };
assign grp_fu_518_p2 = \add_2ns_2ns_2_2_1_U4.dout ;
assign \add_2ns_2ns_2_2_1_U4.reset  = ap_rst;
assign \add_26ns_26ns_26_2_1_U5.top_add_26ns_26ns_26_2_1_Adder_2_U.ain_s0  = \add_26ns_26ns_26_2_1_U5.top_add_26ns_26ns_26_2_1_Adder_2_U.a ;
assign \add_26ns_26ns_26_2_1_U5.top_add_26ns_26ns_26_2_1_Adder_2_U.bin_s0  = \add_26ns_26ns_26_2_1_U5.top_add_26ns_26ns_26_2_1_Adder_2_U.b ;
assign \add_26ns_26ns_26_2_1_U5.top_add_26ns_26ns_26_2_1_Adder_2_U.s  = { \add_26ns_26ns_26_2_1_U5.top_add_26ns_26ns_26_2_1_Adder_2_U.fas_s2 , \add_26ns_26ns_26_2_1_U5.top_add_26ns_26ns_26_2_1_Adder_2_U.sum_s1  };
assign \add_26ns_26ns_26_2_1_U5.top_add_26ns_26ns_26_2_1_Adder_2_U.u2.a  = \add_26ns_26ns_26_2_1_U5.top_add_26ns_26ns_26_2_1_Adder_2_U.ain_s1 ;
assign \add_26ns_26ns_26_2_1_U5.top_add_26ns_26ns_26_2_1_Adder_2_U.u2.b  = \add_26ns_26ns_26_2_1_U5.top_add_26ns_26ns_26_2_1_Adder_2_U.bin_s1 ;
assign \add_26ns_26ns_26_2_1_U5.top_add_26ns_26ns_26_2_1_Adder_2_U.u2.cin  = \add_26ns_26ns_26_2_1_U5.top_add_26ns_26ns_26_2_1_Adder_2_U.carry_s1 ;
assign \add_26ns_26ns_26_2_1_U5.top_add_26ns_26ns_26_2_1_Adder_2_U.facout_s2  = \add_26ns_26ns_26_2_1_U5.top_add_26ns_26ns_26_2_1_Adder_2_U.u2.cout ;
assign \add_26ns_26ns_26_2_1_U5.top_add_26ns_26ns_26_2_1_Adder_2_U.fas_s2  = \add_26ns_26ns_26_2_1_U5.top_add_26ns_26ns_26_2_1_Adder_2_U.u2.s ;
assign \add_26ns_26ns_26_2_1_U5.top_add_26ns_26ns_26_2_1_Adder_2_U.u1.a  = \add_26ns_26ns_26_2_1_U5.top_add_26ns_26ns_26_2_1_Adder_2_U.a [12:0];
assign \add_26ns_26ns_26_2_1_U5.top_add_26ns_26ns_26_2_1_Adder_2_U.u1.b  = \add_26ns_26ns_26_2_1_U5.top_add_26ns_26ns_26_2_1_Adder_2_U.b [12:0];
assign \add_26ns_26ns_26_2_1_U5.top_add_26ns_26ns_26_2_1_Adder_2_U.u1.cin  = 1'h0;
assign \add_26ns_26ns_26_2_1_U5.top_add_26ns_26ns_26_2_1_Adder_2_U.facout_s1  = \add_26ns_26ns_26_2_1_U5.top_add_26ns_26ns_26_2_1_Adder_2_U.u1.cout ;
assign \add_26ns_26ns_26_2_1_U5.top_add_26ns_26ns_26_2_1_Adder_2_U.fas_s1  = \add_26ns_26ns_26_2_1_U5.top_add_26ns_26ns_26_2_1_Adder_2_U.u1.s ;
assign \add_26ns_26ns_26_2_1_U5.top_add_26ns_26ns_26_2_1_Adder_2_U.a  = \add_26ns_26ns_26_2_1_U5.din0 ;
assign \add_26ns_26ns_26_2_1_U5.top_add_26ns_26ns_26_2_1_Adder_2_U.b  = \add_26ns_26ns_26_2_1_U5.din1 ;
assign \add_26ns_26ns_26_2_1_U5.top_add_26ns_26ns_26_2_1_Adder_2_U.ce  = \add_26ns_26ns_26_2_1_U5.ce ;
assign \add_26ns_26ns_26_2_1_U5.top_add_26ns_26ns_26_2_1_Adder_2_U.clk  = \add_26ns_26ns_26_2_1_U5.clk ;
assign \add_26ns_26ns_26_2_1_U5.top_add_26ns_26ns_26_2_1_Adder_2_U.reset  = \add_26ns_26ns_26_2_1_U5.reset ;
assign \add_26ns_26ns_26_2_1_U5.dout  = \add_26ns_26ns_26_2_1_U5.top_add_26ns_26ns_26_2_1_Adder_2_U.s ;
assign \add_26ns_26ns_26_2_1_U5.ce  = 1'h1;
assign \add_26ns_26ns_26_2_1_U5.clk  = ap_clk;
assign \add_26ns_26ns_26_2_1_U5.din0  = { trunc_ln1192_3_reg_1864, 23'h000000 };
assign \add_26ns_26ns_26_2_1_U5.din1  = trunc_ln1192_2_reg_1801;
assign grp_fu_589_p2 = \add_26ns_26ns_26_2_1_U5.dout ;
assign \add_26ns_26ns_26_2_1_U5.reset  = ap_rst;
assign \add_25ns_25ns_25_2_1_U6.top_add_25ns_25ns_25_2_1_Adder_3_U.ain_s0  = \add_25ns_25ns_25_2_1_U6.top_add_25ns_25ns_25_2_1_Adder_3_U.a ;
assign \add_25ns_25ns_25_2_1_U6.top_add_25ns_25ns_25_2_1_Adder_3_U.bin_s0  = \add_25ns_25ns_25_2_1_U6.top_add_25ns_25ns_25_2_1_Adder_3_U.b ;
assign \add_25ns_25ns_25_2_1_U6.top_add_25ns_25ns_25_2_1_Adder_3_U.s  = { \add_25ns_25ns_25_2_1_U6.top_add_25ns_25ns_25_2_1_Adder_3_U.fas_s2 , \add_25ns_25ns_25_2_1_U6.top_add_25ns_25ns_25_2_1_Adder_3_U.sum_s1  };
assign \add_25ns_25ns_25_2_1_U6.top_add_25ns_25ns_25_2_1_Adder_3_U.u2.a  = \add_25ns_25ns_25_2_1_U6.top_add_25ns_25ns_25_2_1_Adder_3_U.ain_s1 ;
assign \add_25ns_25ns_25_2_1_U6.top_add_25ns_25ns_25_2_1_Adder_3_U.u2.b  = \add_25ns_25ns_25_2_1_U6.top_add_25ns_25ns_25_2_1_Adder_3_U.bin_s1 ;
assign \add_25ns_25ns_25_2_1_U6.top_add_25ns_25ns_25_2_1_Adder_3_U.u2.cin  = \add_25ns_25ns_25_2_1_U6.top_add_25ns_25ns_25_2_1_Adder_3_U.carry_s1 ;
assign \add_25ns_25ns_25_2_1_U6.top_add_25ns_25ns_25_2_1_Adder_3_U.facout_s2  = \add_25ns_25ns_25_2_1_U6.top_add_25ns_25ns_25_2_1_Adder_3_U.u2.cout ;
assign \add_25ns_25ns_25_2_1_U6.top_add_25ns_25ns_25_2_1_Adder_3_U.fas_s2  = \add_25ns_25ns_25_2_1_U6.top_add_25ns_25ns_25_2_1_Adder_3_U.u2.s ;
assign \add_25ns_25ns_25_2_1_U6.top_add_25ns_25ns_25_2_1_Adder_3_U.u1.a  = \add_25ns_25ns_25_2_1_U6.top_add_25ns_25ns_25_2_1_Adder_3_U.a [11:0];
assign \add_25ns_25ns_25_2_1_U6.top_add_25ns_25ns_25_2_1_Adder_3_U.u1.b  = \add_25ns_25ns_25_2_1_U6.top_add_25ns_25ns_25_2_1_Adder_3_U.b [11:0];
assign \add_25ns_25ns_25_2_1_U6.top_add_25ns_25ns_25_2_1_Adder_3_U.u1.cin  = 1'h0;
assign \add_25ns_25ns_25_2_1_U6.top_add_25ns_25ns_25_2_1_Adder_3_U.facout_s1  = \add_25ns_25ns_25_2_1_U6.top_add_25ns_25ns_25_2_1_Adder_3_U.u1.cout ;
assign \add_25ns_25ns_25_2_1_U6.top_add_25ns_25ns_25_2_1_Adder_3_U.fas_s1  = \add_25ns_25ns_25_2_1_U6.top_add_25ns_25ns_25_2_1_Adder_3_U.u1.s ;
assign \add_25ns_25ns_25_2_1_U6.top_add_25ns_25ns_25_2_1_Adder_3_U.a  = \add_25ns_25ns_25_2_1_U6.din0 ;
assign \add_25ns_25ns_25_2_1_U6.top_add_25ns_25ns_25_2_1_Adder_3_U.b  = \add_25ns_25ns_25_2_1_U6.din1 ;
assign \add_25ns_25ns_25_2_1_U6.top_add_25ns_25ns_25_2_1_Adder_3_U.ce  = \add_25ns_25ns_25_2_1_U6.ce ;
assign \add_25ns_25ns_25_2_1_U6.top_add_25ns_25ns_25_2_1_Adder_3_U.clk  = \add_25ns_25ns_25_2_1_U6.clk ;
assign \add_25ns_25ns_25_2_1_U6.top_add_25ns_25ns_25_2_1_Adder_3_U.reset  = \add_25ns_25ns_25_2_1_U6.reset ;
assign \add_25ns_25ns_25_2_1_U6.dout  = \add_25ns_25ns_25_2_1_U6.top_add_25ns_25ns_25_2_1_Adder_3_U.s ;
assign \add_25ns_25ns_25_2_1_U6.ce  = 1'h1;
assign \add_25ns_25ns_25_2_1_U6.clk  = ap_clk;
assign \add_25ns_25ns_25_2_1_U6.din0  = { trunc_ln1192_reg_1859, 23'h000000 };
assign \add_25ns_25ns_25_2_1_U6.din1  = empty_reg_1750;
assign grp_fu_594_p2 = \add_25ns_25ns_25_2_1_U6.dout ;
assign \add_25ns_25ns_25_2_1_U6.reset  = ap_rst;
endmodule


// Machine B:
// Processed by function `add_clk_enable_signal` in `verilog_tricks.py`.
// Processed by function `remove_reset_signal` in `verilog_tricks.py`.
module top_B (
  ap_clk,
  ap_start,
  ap_done,
  ap_idle,
  ap_ready,
  op_0,
  op_1,
  op_2,
  op_5,
  op_6,
  op_7,
  op_9,
  op_13,
  op_19,
  op_28,
  op_28_ap_vld,
clk_enable
);
input clk_enable;


input ap_clk;
wire ap_rst;
assign ap_rst = op_28_ap_vld;
input ap_start;
input op_0;
input [31:0] op_1;
input [1:0] op_13;
input [7:0] op_19;
input [3:0] op_2;
input [1:0] op_5;
input [31:0] op_6;
input [3:0] op_7;
input [1:0] op_9;
output ap_done;
output ap_idle;
output ap_ready;
output [31:0] op_28;
output op_28_ap_vld;


reg Range1_all_ones_1_reg_1972;
reg Range1_all_ones_reg_1898;
reg Range1_all_zeros_reg_1905;
reg Range2_all_ones_reg_1893;
reg [8:0] add_ln69_3_reg_2079;
reg and_ln786_1_reg_1983;
reg [6:0] ap_CS_fsm = 7'h01;
reg carry_3_reg_1967;
reg deleted_zeros_1_reg_1977;
reg icmp_ln768_reg_1801;
reg icmp_ln785_reg_1839;
reg icmp_ln786_1_reg_1844;
reg icmp_ln786_2_reg_1806;
reg icmp_ln790_reg_1849;
reg icmp_ln851_2_reg_2035;
reg icmp_ln851_reg_2057;
reg [1:0] op_12_V_reg_1944;
reg [3:0] op_15_V_reg_2040;
reg [3:0] op_16_V_reg_1811;
reg [7:0] op_17_V_reg_1994;
reg [4:0] op_23_V_reg_2062;
reg [3:0] op_3_V_reg_1762;
reg [7:0] op_8_V_reg_1938;
reg p_Result_29_reg_1828;
reg [1:0] p_Result_2_reg_2024;
reg p_Result_30_reg_1854;
reg p_Result_31_reg_1861;
reg p_Result_32_reg_1875;
reg p_Result_33_reg_1887;
reg p_Result_34_reg_1955;
reg p_Result_36_reg_1915;
reg p_Result_37_reg_1926;
reg p_Result_38_reg_1788;
reg p_Result_39_reg_1794;
reg p_Result_40_reg_2006;
reg p_Result_43_reg_2017;
reg [3:0] p_Val2_13_reg_2012;
reg [1:0] p_Val2_3_reg_1866;
reg [7:0] p_Val2_8_reg_1920;
reg [2:0] ret_V_15_reg_1950;
reg [10:0] ret_V_17_reg_1999;
reg [3:0] ret_V_19_reg_2030;
reg [31:0] ret_V_20_cast_reg_2072;
reg [8:0] ret_V_20_reg_2045;
reg [3:0] ret_V_23_reg_1989;
reg [38:0] ret_V_25_reg_2067;
reg [3:0] ret_V_reg_2050;
reg [7:0] ret_reg_1823;
reg [23:0] rhs_3_reg_1933;
reg [7:0] sext_ln69_reg_1767;
reg tmp_reg_1834;
reg [25:0] trunc_ln1192_2_reg_1910;
reg [2:0] trunc_ln1192_3_reg_1783;
reg [1:0] trunc_ln1192_reg_1778;
reg trunc_ln703_reg_1773;
reg xor_ln416_1_reg_1962;
reg xor_ln416_reg_1881;
wire _000_;
wire _001_;
wire _002_;
wire _003_;
wire [8:0] _004_;
wire _005_;
wire [6:0] _006_;
wire _007_;
wire _008_;
wire _009_;
wire _010_;
wire _011_;
wire _012_;
wire _013_;
wire _014_;
wire _015_;
wire [1:0] _016_;
wire [3:0] _017_;
wire [3:0] _018_;
wire [7:0] _019_;
wire [4:0] _020_;
wire [3:0] _021_;
wire [7:0] _022_;
wire _023_;
wire [1:0] _024_;
wire _025_;
wire _026_;
wire _027_;
wire _028_;
wire _029_;
wire _030_;
wire _031_;
wire _032_;
wire _033_;
wire _034_;
wire _035_;
wire [3:0] _036_;
wire [1:0] _037_;
wire [7:0] _038_;
wire [2:0] _039_;
wire [10:0] _040_;
wire [3:0] _041_;
wire [31:0] _042_;
wire [8:0] _043_;
wire [3:0] _044_;
wire [38:0] _045_;
wire [3:0] _046_;
wire [7:0] _047_;
wire [1:0] _048_;
wire [7:0] _049_;
wire _050_;
wire [25:0] _051_;
wire [2:0] _052_;
wire [1:0] _053_;
wire _054_;
wire _055_;
wire _056_;
wire [1:0] _057_;
wire _058_;
wire _059_;
wire _060_;
wire _061_;
wire _062_;
wire _063_;
wire _064_;
wire _065_;
wire _066_;
wire _067_;
wire _068_;
wire _069_;
wire _070_;
wire _071_;
wire _072_;
wire _073_;
wire _074_;
wire _075_;
wire _076_;
wire _077_;
wire _078_;
wire _079_;
wire _080_;
wire _081_;
wire _082_;
wire _083_;
wire _084_;
wire _085_;
wire _086_;
wire _087_;
wire Range1_all_ones_1_fu_1083_p2;
wire Range1_all_ones_2_fu_1458_p2;
wire Range1_all_ones_fu_565_p2;
wire Range1_all_zeros_1_fu_1089_p2;
wire Range1_all_zeros_2_fu_1463_p2;
wire Range1_all_zeros_fu_571_p2;
wire Range2_all_ones_1_fu_1067_p2;
wire Range2_all_ones_2_fu_1451_p3;
wire Range2_all_ones_fu_549_p2;
wire [25:0] add_ln1192_1_fu_1034_p2;
wire [24:0] add_ln1192_2_fu_588_p2;
wire [31:0] add_ln691_3_fu_1734_p2;
wire [3:0] add_ln691_fu_1401_p2;
wire [8:0] add_ln69_3_fu_1721_p2;
wire [4:0] add_ln69_fu_1624_p2;
wire and_ln340_fu_964_p2;
wire and_ln408_fu_1326_p2;
wire and_ln412_fu_644_p2;
wire and_ln414_fu_501_p2;
wire and_ln780_1_fu_1117_p2;
wire and_ln780_2_fu_1489_p2;
wire and_ln780_fu_815_p2;
wire and_ln781_1_fu_1194_p2;
wire and_ln781_2_fu_1503_p2;
wire and_ln781_fu_827_p2;
wire and_ln785_1_fu_939_p2;
wire and_ln785_2_fu_952_p2;
wire and_ln785_4_fu_1248_p2;
wire and_ln785_5_fu_1257_p2;
wire and_ln785_fu_929_p2;
wire and_ln786_1_fu_1131_p2;
wire and_ln786_3_fu_1531_p2;
wire and_ln786_fu_865_p2;
wire [7:0] and_ln_fu_740_p3;
wire ap_CS_fsm_state1;
wire ap_CS_fsm_state2;
wire ap_CS_fsm_state3;
wire ap_CS_fsm_state4;
wire ap_CS_fsm_state5;
wire ap_CS_fsm_state6;
wire ap_CS_fsm_state7;
wire [6:0] ap_NS_fsm;
wire ap_clk;
wire ap_done;
wire ap_idle;
wire ap_ready;
wire ap_rst;
wire ap_start;
wire carry_1_fu_800_p2;
wire carry_3_fu_1052_p2;
wire carry_5_fu_1445_p2;
wire deleted_ones_1_fu_1123_p3;
wire deleted_ones_2_fu_1495_p3;
wire deleted_ones_fu_820_p3;
wire deleted_zeros_1_fu_1095_p3;
wire deleted_zeros_2_fu_1468_p3;
wire deleted_zeros_fu_804_p3;
wire [31:0] empty_fu_391_p0;
wire [24:0] empty_fu_391_p1;
wire icmp_ln414_fu_495_p2;
wire icmp_ln768_fu_367_p2;
wire icmp_ln785_fu_435_p2;
wire icmp_ln786_1_fu_441_p2;
wire icmp_ln786_2_fu_373_p2;
wire icmp_ln786_fu_757_p2;
wire icmp_ln790_fu_459_p2;
wire icmp_ln851_1_fu_1166_p2;
wire icmp_ln851_2_fu_1427_p2;
wire icmp_ln851_fu_1611_p2;
wire [26:0] lhs_V_1_fu_1007_p3;
wire [8:0] lhs_V_3_fu_1269_p3;
wire [3:0] \mul_4s_4s_4_1_1_U1.din0 ;
wire [3:0] \mul_4s_4s_4_1_1_U1.din1 ;
wire [3:0] \mul_4s_4s_4_1_1_U1.dout ;
wire [3:0] \mul_4s_4s_4_1_1_U1.top_mul_4s_4s_4_1_1_Multiplier_0_U.a ;
wire [3:0] \mul_4s_4s_4_1_1_U1.top_mul_4s_4s_4_1_1_Multiplier_0_U.b ;
wire [3:0] \mul_4s_4s_4_1_1_U1.top_mul_4s_4s_4_1_1_Multiplier_0_U.p ;
wire [3:0] \mul_4s_4s_8_1_1_U2.din0 ;
wire [3:0] \mul_4s_4s_8_1_1_U2.din1 ;
wire [7:0] \mul_4s_4s_8_1_1_U2.dout ;
wire [3:0] \mul_4s_4s_8_1_1_U2.top_mul_4s_4s_8_1_1_Multiplier_1_U.a ;
wire [3:0] \mul_4s_4s_8_1_1_U2.top_mul_4s_4s_8_1_1_Multiplier_1_U.b ;
wire [7:0] \mul_4s_4s_8_1_1_U2.top_mul_4s_4s_8_1_1_Multiplier_1_U.p ;
wire neg_src_7_fu_1204_p2;
wire neg_src_fu_838_p2;
wire op_0;
wire [31:0] op_1;
wire [1:0] op_12_V_fu_982_p3;
wire [1:0] op_13;
wire [3:0] op_15_V_fu_1567_p3;
wire [3:0] op_16_V_fu_385_p2;
wire [7:0] op_17_V_fu_1262_p3;
wire [7:0] op_19;
wire [3:0] op_2;
wire [4:0] op_23_V_fu_1630_p2;
wire [5:0] op_25_V_fu_1680_p2;
wire [31:0] op_28;
wire op_28_ap_vld;
wire [3:0] op_3_V_fu_279_p2;
wire [7:0] op_4_V_fu_301_p2;
wire [1:0] op_5;
wire [31:0] op_6;
wire [3:0] op_7;
wire [7:0] op_8_V_fu_792_p3;
wire [1:0] op_9;
wire or_ln340_1_fu_916_p2;
wire or_ln340_2_fu_970_p2;
wire or_ln340_3_fu_1230_p2;
wire or_ln340_4_fu_1235_p2;
wire or_ln340_fu_870_p2;
wire or_ln384_1_fu_705_p2;
wire or_ln384_2_fu_1561_p2;
wire or_ln384_fu_786_p2;
wire or_ln412_fu_638_p2;
wire or_ln731_fu_345_p2;
wire [3:0] or_ln760_fu_379_p1;
wire [3:0] or_ln760_fu_379_p2;
wire or_ln785_1_fu_1214_p2;
wire or_ln785_2_fu_675_p2;
wire or_ln785_3_fu_1515_p2;
wire or_ln785_4_fu_934_p2;
wire or_ln785_5_fu_1252_p2;
wire or_ln785_fu_849_p2;
wire or_ln786_1_fu_1536_p2;
wire or_ln786_fu_695_p2;
wire or_ln788_1_fu_767_p2;
wire or_ln788_fu_763_p2;
wire [7:0] or_ln_fu_425_p4;
wire overflow_1_fu_859_p2;
wire overflow_2_fu_1224_p2;
wire overflow_3_fu_684_p2;
wire overflow_4_fu_1525_p2;
wire overflow_fu_752_p2;
wire [1:0] p_Result_12_fu_907_p4;
wire p_Result_17_fu_604_p3;
wire [31:0] p_Result_1_fu_539_p1;
wire [6:0] p_Result_1_fu_539_p4;
wire p_Result_25_fu_1390_p3;
wire p_Result_26_fu_1636_p3;
wire p_Result_27_fu_1154_p3;
wire p_Result_28_fu_1727_p3;
wire [31:0] p_Result_30_fu_465_p1;
wire p_Result_30_fu_465_p3;
wire [31:0] p_Result_31_fu_483_p1;
wire p_Result_32_fu_517_p3;
wire [31:0] p_Result_33_fu_531_p1;
wire [31:0] p_Result_35_fu_612_p1;
wire p_Result_35_fu_612_p3;
wire p_Result_39_fu_351_p2;
wire [31:0] p_Result_3_fu_555_p1;
wire [7:0] p_Result_3_fu_555_p4;
wire p_Result_41_fu_1308_p3;
wire p_Result_42_fu_1433_p3;
wire [6:0] p_Result_5_fu_1057_p4;
wire [7:0] p_Result_6_fu_1073_p4;
wire [7:0] p_Result_8_fu_357_p4;
wire [6:0] p_Result_s_20_fu_451_p3;
wire [4:0] p_Result_s_fu_415_p4;
wire [1:0] p_Val2_10_fu_668_p3;
wire [3:0] p_Val2_12_fu_1298_p4;
wire [3:0] p_Val2_13_fu_1336_p2;
wire [7:0] p_Val2_1_fu_735_p2;
wire [31:0] p_Val2_2_fu_473_p1;
wire [1:0] p_Val2_2_fu_473_p4;
wire [1:0] p_Val2_3_fu_511_p2;
wire p_Val2_4_fu_902_p2;
wire [7:0] p_Val2_7_fu_594_p4;
wire [7:0] p_Val2_8_fu_654_p2;
wire r_1_fu_1320_p2;
wire r_fu_624_p2;
wire [8:0] ret_2_fu_327_p2;
wire [3:0] ret_V_10_fu_1172_p2;
wire [2:0] ret_V_15_fu_1001_p2;
wire [32:0] ret_V_16_fu_1028_p2;
wire [10:0] ret_V_17_fu_1284_p2;
wire [3:0] ret_V_18_fu_1370_p2;
wire [3:0] ret_V_19_fu_1415_p3;
wire [8:0] ret_V_20_fu_1591_p2;
wire [3:0] ret_V_21_fu_1654_p3;
wire [31:0] ret_V_22_fu_1139_p1;
wire [31:0] ret_V_22_fu_1139_p2;
wire [3:0] ret_V_23_fu_1186_p3;
wire [5:0] ret_V_24_fu_1671_p2;
wire [38:0] ret_V_25_fu_1701_p2;
wire [31:0] ret_V_26_fu_1745_p3;
wire [3:0] ret_V_7_cast_fu_1144_p4;
wire [3:0] ret_V_7_fu_1643_p2;
wire [3:0] ret_fu_395_p0;
wire [3:0] ret_fu_395_p1;
wire [7:0] ret_fu_395_p2;
wire [3:0] rhs_2_fu_1363_p3;
wire [23:0] rhs_3_fu_727_p3;
wire [6:0] rhs_fu_1580_p3;
wire sel_tmp11_fu_976_p2;
wire [7:0] select_ln340_1_fu_1241_p3;
wire [1:0] select_ln340_fu_922_p3;
wire [3:0] select_ln384_2_fu_1553_p3;
wire [1:0] select_ln384_4_fu_711_p3;
wire [1:0] select_ln384_5_fu_719_p3;
wire [7:0] select_ln384_fu_778_p3;
wire [2:0] select_ln703_fu_989_p3;
wire [1:0] select_ln785_fu_945_p3;
wire [3:0] select_ln850_1_fu_1648_p3;
wire [3:0] select_ln850_2_fu_1178_p3;
wire [31:0] select_ln850_3_fu_1739_p3;
wire [3:0] select_ln850_fu_1407_p3;
wire [3:0] sext_ln1192_1_fu_1360_p1;
wire [5:0] sext_ln1192_2_fu_1668_p1;
wire [38:0] sext_ln1192_3_fu_1697_p1;
wire [32:0] sext_ln1192_fu_1014_p1;
wire [8:0] sext_ln1193_fu_1587_p1;
wire [31:0] sext_ln1195_fu_1136_p1;
wire [8:0] sext_ln19_fu_1661_p1;
wire [8:0] sext_ln215_fu_319_p1;
wire [5:0] sext_ln23_fu_1665_p1;
wire [4:0] sext_ln69_1_fu_1617_p1;
wire [4:0] sext_ln69_2_fu_1621_p1;
wire [5:0] sext_ln69_3_fu_1677_p1;
wire [8:0] sext_ln69_4_fu_1717_p1;
wire [31:0] sext_ln69_5_fu_1752_p1;
wire [3:0] sext_ln69_fu_289_p0;
wire [7:0] sext_ln69_fu_289_p1;
wire [31:0] sext_ln703_1_fu_1018_p0;
wire [32:0] sext_ln703_1_fu_1018_p1;
wire [10:0] sext_ln703_2_fu_1281_p1;
wire [8:0] sext_ln703_3_fu_1577_p1;
wire [38:0] sext_ln703_4_fu_1686_p1;
wire [2:0] sext_ln703_fu_997_p1;
wire [4:0] sext_ln831_fu_1574_p1;
wire [3:0] sext_ln850_fu_1386_p1;
wire tmp_14_fu_1103_p3;
wire tmp_21_fu_1476_p3;
wire [11:0] tmp_25_fu_1689_p3;
wire [2:0] tmp_5_fu_1376_p4;
wire [31:0] tmp_6_fu_876_p1;
wire tmp_6_fu_876_p3;
wire tmp_7_fu_883_p3;
wire tmp_fu_407_p3;
wire [24:0] trunc_ln1192_1_fu_577_p3;
wire [31:0] trunc_ln1192_2_fu_584_p0;
wire [25:0] trunc_ln1192_2_fu_584_p1;
wire [2:0] trunc_ln1192_3_fu_315_p1;
wire [25:0] trunc_ln1192_4_fu_1021_p3;
wire [1:0] trunc_ln1192_fu_311_p1;
wire [31:0] trunc_ln414_fu_491_p0;
wire [21:0] trunc_ln414_fu_491_p1;
wire [7:0] trunc_ln69_1_fu_285_p1;
wire trunc_ln69_2_fu_293_p1;
wire [3:0] trunc_ln69_3_fu_297_p0;
wire trunc_ln69_3_fu_297_p1;
wire [3:0] trunc_ln69_fu_275_p1;
wire trunc_ln703_fu_307_p1;
wire [3:0] trunc_ln718_1_fu_1316_p1;
wire [31:0] trunc_ln718_fu_620_p0;
wire [15:0] trunc_ln718_fu_620_p1;
wire trunc_ln731_fu_341_p1;
wire [1:0] trunc_ln790_fu_447_p1;
wire [4:0] trunc_ln851_1_fu_1607_p1;
wire [22:0] trunc_ln851_2_fu_1162_p1;
wire [5:0] trunc_ln851_3_fu_1423_p1;
wire trunc_ln851_fu_1398_p1;
wire underflow_3_fu_700_p2;
wire underflow_4_fu_1548_p2;
wire underflow_fu_773_p2;
wire xor_ln365_1_fu_896_p2;
wire xor_ln365_fu_890_p2;
wire xor_ln416_1_fu_1047_p2;
wire xor_ln416_2_fu_1440_p2;
wire xor_ln416_fu_525_p2;
wire xor_ln780_1_fu_1111_p2;
wire xor_ln780_2_fu_1483_p2;
wire xor_ln780_fu_810_p2;
wire xor_ln781_1_fu_1198_p2;
wire xor_ln781_fu_832_p2;
wire xor_ln785_1_fu_843_p2;
wire xor_ln785_2_fu_854_p2;
wire xor_ln785_3_fu_1209_p2;
wire xor_ln785_4_fu_1219_p2;
wire xor_ln785_5_fu_679_p2;
wire xor_ln785_6_fu_1509_p2;
wire xor_ln785_7_fu_1520_p2;
wire xor_ln785_fu_747_p2;
wire xor_ln786_1_fu_958_p2;
wire xor_ln786_2_fu_1542_p2;
wire xor_ln786_fu_690_p2;
wire [10:0] zext_ln1193_fu_1277_p1;
wire [8:0] zext_ln215_fu_323_p1;
wire [7:0] zext_ln415_1_fu_650_p1;
wire [3:0] zext_ln415_2_fu_1332_p1;
wire [1:0] zext_ln415_fu_507_p1;


assign add_ln1192_1_fu_1034_p2 = { trunc_ln1192_3_reg_1783, 23'h000000 } + trunc_ln1192_2_reg_1910;
assign add_ln1192_2_fu_588_p2 = { trunc_ln1192_reg_1778, 23'h000000 } + op_6[24:0];
assign add_ln691_3_fu_1734_p2 = ret_V_20_cast_reg_2072 + 1'h1;
assign add_ln691_fu_1401_p2 = $signed(ret_V_18_fu_1370_p2[3:1]) + $signed(2'h1);
assign add_ln69_3_fu_1721_p2 = $signed(op_19) + $signed(ret_V_21_fu_1654_p3);
assign add_ln69_fu_1624_p2 = $signed(ret_V_23_reg_1989) + $signed(op_13);
assign op_23_V_fu_1630_p2 = $signed(add_ln69_fu_1624_p2) + $signed(ret_V_19_reg_2030);
assign op_25_V_fu_1680_p2 = $signed(ret_V_24_fu_1671_p2) + $signed(op_16_V_reg_1811);
assign op_28 = $signed(add_ln69_3_reg_2079) + $signed(ret_V_26_fu_1745_p3);
assign p_Val2_13_fu_1336_p2 = ret_V_17_fu_1284_p2[8:5] + and_ln408_fu_1326_p2;
assign p_Val2_3_fu_511_p2 = op_6[23:22] + and_ln414_fu_501_p2;
assign p_Val2_8_fu_654_p2 = add_ln1192_2_fu_588_p2[24:17] + and_ln412_fu_644_p2;
assign ret_2_fu_327_p2 = $signed(op_4_V_fu_301_p2) + $signed({ 1'h0, op_5 });
assign ret_V_10_fu_1172_p2 = ret_V_22_fu_1139_p2[26:23] + 1'h1;
assign ret_V_15_fu_1001_p2 = $signed(op_9) + $signed(select_ln703_fu_989_p3);
assign ret_V_16_fu_1028_p2 = $signed({ op_3_V_reg_1762, 23'h000000 }) + $signed(op_6);
assign ret_V_18_fu_1370_p2 = $signed({ ret_V_15_reg_1950, 1'h0 }) + $signed(op_12_V_reg_1944);
assign ret_V_24_fu_1671_p2 = $signed(op_23_V_reg_2062) + $signed(op_15_V_reg_2040);
assign { ret_V_25_fu_1701_p2[38], ret_V_25_fu_1701_p2[11:0] } = $signed({ op_25_V_fu_1680_p2, 6'h00 }) + $signed(op_17_V_reg_1994);
assign ret_V_7_fu_1643_p2 = ret_V_reg_2050 + 1'h1;
assign underflow_3_fu_700_p2 = p_Result_38_reg_1788 & or_ln786_fu_695_p2;
assign underflow_4_fu_1548_p2 = xor_ln786_2_fu_1542_p2 & p_Result_40_reg_2006;
assign underflow_fu_773_p2 = p_Result_29_reg_1828 & or_ln788_1_fu_767_p2;
assign _058_ = ap_CS_fsm[0] & _060_;
assign _059_ = ap_CS_fsm[0] & ap_start;
assign and_ln340_fu_964_p2 = xor_ln786_1_fu_958_p2 & or_ln340_fu_870_p2;
assign and_ln408_fu_1326_p2 = r_1_fu_1320_p2 & ret_V_17_fu_1284_p2[4];
assign and_ln412_fu_644_p2 = op_6[16] & or_ln412_fu_638_p2;
assign and_ln414_fu_501_p2 = op_6[31] & icmp_ln414_fu_495_p2;
assign and_ln780_1_fu_1117_p2 = xor_ln780_1_fu_1111_p2 & Range2_all_ones_1_fu_1067_p2;
assign and_ln780_2_fu_1489_p2 = xor_ln780_2_fu_1483_p2 & ret_V_17_reg_1999[10];
assign and_ln780_fu_815_p2 = xor_ln780_fu_810_p2 & Range2_all_ones_reg_1893;
assign and_ln781_1_fu_1194_p2 = carry_3_reg_1967 & Range1_all_ones_1_reg_1972;
assign and_ln781_2_fu_1503_p2 = carry_5_fu_1445_p2 & Range1_all_ones_2_fu_1458_p2;
assign and_ln781_fu_827_p2 = carry_1_fu_800_p2 & Range1_all_ones_reg_1898;
assign and_ln785_1_fu_939_p2 = or_ln785_4_fu_934_p2 & and_ln786_fu_865_p2;
assign and_ln785_2_fu_952_p2 = xor_ln785_2_fu_854_p2 & and_ln786_fu_865_p2;
assign and_ln785_4_fu_1248_p2 = xor_ln416_1_reg_1962 & deleted_zeros_1_reg_1977;
assign and_ln785_5_fu_1257_p2 = or_ln785_5_fu_1252_p2 & and_ln786_1_reg_1983;
assign and_ln785_fu_929_p2 = xor_ln416_reg_1881 & deleted_zeros_fu_804_p3;
assign and_ln786_1_fu_1131_p2 = p_Result_37_reg_1926 & deleted_ones_1_fu_1123_p3;
assign and_ln786_3_fu_1531_p2 = p_Result_43_reg_2017 & deleted_ones_2_fu_1495_p3;
assign and_ln786_fu_865_p2 = p_Result_32_reg_1875 & deleted_ones_fu_820_p3;
assign carry_1_fu_800_p2 = xor_ln416_reg_1881 & p_Result_31_reg_1861;
assign carry_3_fu_1052_p2 = xor_ln416_1_fu_1047_p2 & p_Result_36_reg_1915;
assign carry_5_fu_1445_p2 = xor_ln416_2_fu_1440_p2 & ret_V_17_reg_1999[8];
assign neg_src_7_fu_1204_p2 = xor_ln781_1_fu_1198_p2 & p_Result_34_reg_1955;
assign neg_src_fu_838_p2 = xor_ln781_fu_832_p2 & p_Result_30_reg_1854;
assign overflow_1_fu_859_p2 = xor_ln785_2_fu_854_p2 & or_ln785_fu_849_p2;
assign overflow_2_fu_1224_p2 = xor_ln785_4_fu_1219_p2 & or_ln785_1_fu_1214_p2;
assign overflow_3_fu_684_p2 = xor_ln785_5_fu_679_p2 & or_ln785_2_fu_675_p2;
assign overflow_4_fu_1525_p2 = xor_ln785_7_fu_1520_p2 & or_ln785_3_fu_1515_p2;
assign overflow_fu_752_p2 = xor_ln785_fu_747_p2 & icmp_ln785_reg_1839;
assign sel_tmp11_fu_976_p2 = xor_ln365_1_fu_896_p2 & or_ln340_2_fu_970_p2;
assign xor_ln781_fu_832_p2 = ~ and_ln781_fu_827_p2;
assign xor_ln785_1_fu_843_p2 = ~ deleted_zeros_fu_804_p3;
assign xor_ln785_2_fu_854_p2 = ~ p_Result_30_reg_1854;
assign xor_ln780_fu_810_p2 = ~ p_Result_33_reg_1887;
assign xor_ln786_1_fu_958_p2 = ~ and_ln786_fu_865_p2;
assign xor_ln780_1_fu_1111_p2 = ~ add_ln1192_1_fu_1034_p2[25];
assign xor_ln780_2_fu_1483_p2 = ~ ret_V_17_reg_1999[9];
assign xor_ln416_2_fu_1440_p2 = ~ p_Result_43_reg_2017;
assign xor_ln416_1_fu_1047_p2 = ~ p_Result_37_reg_1926;
assign xor_ln781_1_fu_1198_p2 = ~ and_ln781_1_fu_1194_p2;
assign xor_ln785_3_fu_1209_p2 = ~ deleted_zeros_1_reg_1977;
assign xor_ln785_4_fu_1219_p2 = ~ p_Result_34_reg_1955;
assign xor_ln365_1_fu_896_p2 = ~ xor_ln365_fu_890_p2;
assign xor_ln785_6_fu_1509_p2 = ~ deleted_zeros_2_fu_1468_p3;
assign xor_ln785_7_fu_1520_p2 = ~ p_Result_40_reg_2006;
assign xor_ln786_2_fu_1542_p2 = ~ or_ln786_1_fu_1536_p2;
assign xor_ln785_fu_747_p2 = ~ p_Result_29_reg_1828;
assign xor_ln785_5_fu_679_p2 = ~ p_Result_38_reg_1788;
assign xor_ln786_fu_690_p2 = ~ p_Result_39_reg_1794;
assign xor_ln416_fu_525_p2 = ~ p_Val2_3_fu_511_p2[1];
assign p_Val2_4_fu_902_p2 = ~ p_Val2_3_reg_1866[0];
assign op_16_V_fu_385_p2 = ~ or_ln760_fu_379_p2;
assign _060_ = ~ ap_start;
assign _061_ = ret_V_16_fu_1028_p2[32:25] == 8'hff;
assign _062_ = p_Result_2_reg_2024 == 2'h3;
assign _063_ = op_6[31:24] == 8'hff;
assign _064_ = ! ret_V_16_fu_1028_p2[32:25];
assign _065_ = ! p_Result_2_reg_2024;
assign _066_ = ! op_6[31:24];
assign _067_ = ret_V_16_fu_1028_p2[32:26] == 7'h7f;
assign _068_ = op_6[31:25] == 7'h7f;
assign _069_ = ! { tmp_reg_1834, 7'h00 };
assign _070_ = ! { ret_fu_395_p2[1:0], 5'h00 };
assign _071_ = ! ret_V_22_fu_1139_p2[22:0];
assign _072_ = ! ret_V_20_fu_1591_p2[4:0];
assign \mul_4s_4s_4_1_1_U1.top_mul_4s_4s_4_1_1_Multiplier_0_U.p  = $signed(\mul_4s_4s_4_1_1_U1.top_mul_4s_4s_4_1_1_Multiplier_0_U.a ) * $signed(\mul_4s_4s_4_1_1_U1.top_mul_4s_4s_4_1_1_Multiplier_0_U.b );
assign \mul_4s_4s_8_1_1_U2.top_mul_4s_4s_8_1_1_Multiplier_1_U.p  = $signed(\mul_4s_4s_8_1_1_U2.top_mul_4s_4s_8_1_1_Multiplier_1_U.a ) * $signed(\mul_4s_4s_8_1_1_U2.top_mul_4s_4s_8_1_1_Multiplier_1_U.b );
assign _073_ = | op_6[21:0];
assign _074_ = | ret_2_fu_327_p2[8:1];
assign _075_ = | { ret_fu_395_p2[2], 2'h0, ret_fu_395_p2[7:3] };
assign _076_ = ret_fu_395_p2[7:3] != 5'h1f;
assign _077_ = ret_2_fu_327_p2[8:1] != 8'hff;
assign _078_ = | op_17_V_fu_1262_p3[5:0];
assign _079_ = | ret_V_17_fu_1284_p2[3:0];
assign _080_ = | op_6[15:0];
assign op_4_V_fu_301_p2 = op_1[7:0] | { op_2[3], op_2[3], op_2[3], op_2[3], op_2 };
assign or_ln340_1_fu_916_p2 = or_ln340_fu_870_p2 | and_ln786_fu_865_p2;
assign or_ln340_2_fu_970_p2 = and_ln785_2_fu_952_p2 | and_ln340_fu_964_p2;
assign or_ln340_3_fu_1230_p2 = overflow_2_fu_1224_p2 | and_ln786_1_reg_1983;
assign or_ln340_4_fu_1235_p2 = or_ln340_3_fu_1230_p2 | neg_src_7_fu_1204_p2;
assign or_ln340_fu_870_p2 = overflow_1_fu_859_p2 | neg_src_fu_838_p2;
assign or_ln384_1_fu_705_p2 = underflow_3_fu_700_p2 | overflow_3_fu_684_p2;
assign or_ln384_2_fu_1561_p2 = underflow_4_fu_1548_p2 | overflow_4_fu_1525_p2;
assign or_ln384_fu_786_p2 = underflow_fu_773_p2 | overflow_fu_752_p2;
assign or_ln412_fu_638_p2 = r_fu_624_p2 | add_ln1192_2_fu_588_p2[17];
assign or_ln731_fu_345_p2 = op_2[0] | op_1[0];
assign or_ln760_fu_379_p2 = $signed(op_1[3:0]) | $signed(op_2);
assign or_ln785_1_fu_1214_p2 = xor_ln785_3_fu_1209_p2 | p_Result_37_reg_1926;
assign or_ln785_2_fu_675_p2 = p_Result_39_reg_1794 | icmp_ln768_reg_1801;
assign or_ln785_3_fu_1515_p2 = xor_ln785_6_fu_1509_p2 | p_Result_43_reg_2017;
assign or_ln785_4_fu_934_p2 = p_Result_30_reg_1854 | and_ln785_fu_929_p2;
assign or_ln785_5_fu_1252_p2 = p_Result_34_reg_1955 | and_ln785_4_fu_1248_p2;
assign or_ln785_fu_849_p2 = xor_ln785_1_fu_843_p2 | p_Result_32_reg_1875;
assign or_ln786_1_fu_1536_p2 = and_ln786_3_fu_1531_p2 | and_ln781_2_fu_1503_p2;
assign or_ln786_fu_695_p2 = xor_ln786_fu_690_p2 | icmp_ln786_2_reg_1806;
assign or_ln788_1_fu_767_p2 = or_ln788_fu_763_p2 | icmp_ln786_fu_757_p2;
assign or_ln788_fu_763_p2 = icmp_ln790_reg_1849 | icmp_ln786_1_reg_1844;
assign ret_V_22_fu_1139_p2 = $signed(rhs_3_reg_1933) | $signed(op_6);
always @(posedge ap_clk)
rhs_3_reg_1933[21:0] <= 22'h000000;
always @(posedge ap_clk)
op_15_V_reg_2040 <= _017_;
always @(posedge ap_clk)
ret_V_20_reg_2045 <= _043_;
always @(posedge ap_clk)
ret_V_reg_2050 <= _046_;
always @(posedge ap_clk)
icmp_ln851_reg_2057 <= _015_;
always @(posedge ap_clk)
op_23_V_reg_2062 <= _020_;
always @(posedge ap_clk)
op_17_V_reg_1994 <= _019_;
always @(posedge ap_clk)
ret_V_17_reg_1999 <= _040_;
always @(posedge ap_clk)
p_Result_40_reg_2006 <= _034_;
always @(posedge ap_clk)
p_Val2_13_reg_2012 <= _036_;
always @(posedge ap_clk)
p_Result_43_reg_2017 <= _035_;
always @(posedge ap_clk)
p_Result_2_reg_2024 <= _024_;
always @(posedge ap_clk)
ret_V_19_reg_2030 <= _041_;
always @(posedge ap_clk)
icmp_ln851_2_reg_2035 <= _014_;
always @(posedge ap_clk)
op_3_V_reg_1762 <= _021_;
always @(posedge ap_clk)
sext_ln69_reg_1767 <= _049_;
always @(posedge ap_clk)
trunc_ln703_reg_1773 <= _054_;
always @(posedge ap_clk)
trunc_ln1192_reg_1778 <= _053_;
always @(posedge ap_clk)
trunc_ln1192_3_reg_1783 <= _052_;
always @(posedge ap_clk)
p_Result_38_reg_1788 <= _032_;
always @(posedge ap_clk)
p_Result_39_reg_1794 <= _033_;
always @(posedge ap_clk)
icmp_ln768_reg_1801 <= _009_;
always @(posedge ap_clk)
icmp_ln786_2_reg_1806 <= _012_;
always @(posedge ap_clk)
op_16_V_reg_1811 <= _018_;
always @(posedge ap_clk)
ret_V_25_reg_2067 <= _045_;
always @(posedge ap_clk)
ret_V_20_cast_reg_2072 <= _042_;
always @(posedge ap_clk)
add_ln69_3_reg_2079 <= _004_;
always @(posedge ap_clk)
ret_reg_1823 <= _047_;
always @(posedge ap_clk)
p_Result_29_reg_1828 <= _023_;
always @(posedge ap_clk)
tmp_reg_1834 <= _050_;
always @(posedge ap_clk)
icmp_ln785_reg_1839 <= _010_;
always @(posedge ap_clk)
icmp_ln786_1_reg_1844 <= _011_;
always @(posedge ap_clk)
icmp_ln790_reg_1849 <= _013_;
always @(posedge ap_clk)
p_Result_30_reg_1854 <= _025_;
always @(posedge ap_clk)
p_Result_31_reg_1861 <= _026_;
always @(posedge ap_clk)
p_Val2_3_reg_1866 <= _037_;
always @(posedge ap_clk)
p_Result_32_reg_1875 <= _027_;
always @(posedge ap_clk)
xor_ln416_reg_1881 <= _056_;
always @(posedge ap_clk)
p_Result_33_reg_1887 <= _028_;
always @(posedge ap_clk)
Range2_all_ones_reg_1893 <= _003_;
always @(posedge ap_clk)
Range1_all_ones_reg_1898 <= _001_;
always @(posedge ap_clk)
Range1_all_zeros_reg_1905 <= _002_;
always @(posedge ap_clk)
trunc_ln1192_2_reg_1910 <= _051_;
always @(posedge ap_clk)
p_Result_36_reg_1915 <= _030_;
always @(posedge ap_clk)
p_Val2_8_reg_1920 <= _038_;
always @(posedge ap_clk)
p_Result_37_reg_1926 <= _031_;
always @(posedge ap_clk)
rhs_3_reg_1933[23:22] <= _048_;
always @(posedge ap_clk)
op_8_V_reg_1938 <= _022_;
always @(posedge ap_clk)
op_12_V_reg_1944 <= _016_;
always @(posedge ap_clk)
ret_V_15_reg_1950 <= _039_;
always @(posedge ap_clk)
p_Result_34_reg_1955 <= _029_;
always @(posedge ap_clk)
xor_ln416_1_reg_1962 <= _055_;
always @(posedge ap_clk)
carry_3_reg_1967 <= _007_;
always @(posedge ap_clk)
Range1_all_ones_1_reg_1972 <= _000_;
always @(posedge ap_clk)
deleted_zeros_1_reg_1977 <= _008_;
always @(posedge ap_clk)
and_ln786_1_reg_1983 <= _005_;
always @(posedge ap_clk)
ret_V_23_reg_1989 <= _044_;
always @(posedge ap_clk)
ap_CS_fsm <= _006_;
assign _057_ = _059_ ? 2'h2 : 2'h1;
assign _081_ = ap_CS_fsm == 1'h1;
function [6:0] _270_;
input [6:0] a;
input [48:0] b;
input [6:0] s;
case (s)
7'b0000001:
_270_ = b[6:0];
7'b0000010:
_270_ = b[13:7];
7'b0000100:
_270_ = b[20:14];
7'b0001000:
_270_ = b[27:21];
7'b0010000:
_270_ = b[34:28];
7'b0100000:
_270_ = b[41:35];
7'b1000000:
_270_ = b[48:42];
7'b0000000:
_270_ = a;
default:
_270_ = 7'bx;
endcase
endfunction
assign ap_NS_fsm = _270_(7'hxx, { 5'h00, _057_, 42'h02082082001 }, { _081_, _087_, _086_, _085_, _084_, _083_, _082_ });
assign _082_ = ap_CS_fsm == 7'h40;
assign _083_ = ap_CS_fsm == 6'h20;
assign _084_ = ap_CS_fsm == 5'h10;
assign _085_ = ap_CS_fsm == 4'h8;
assign _086_ = ap_CS_fsm == 3'h4;
assign _087_ = ap_CS_fsm == 2'h2;
assign op_28_ap_vld = ap_CS_fsm[6] ? 1'h1 : 1'h0;
assign ap_idle = _058_ ? 1'h1 : 1'h0;
assign _020_ = ap_CS_fsm[4] ? op_23_V_fu_1630_p2 : op_23_V_reg_2062;
assign _015_ = ap_CS_fsm[4] ? icmp_ln851_fu_1611_p2 : icmp_ln851_reg_2057;
assign _046_ = ap_CS_fsm[4] ? ret_V_20_fu_1591_p2[8:5] : ret_V_reg_2050;
assign _043_ = ap_CS_fsm[4] ? ret_V_20_fu_1591_p2 : ret_V_20_reg_2045;
assign _017_ = ap_CS_fsm[4] ? op_15_V_fu_1567_p3 : op_15_V_reg_2040;
assign _014_ = ap_CS_fsm[3] ? icmp_ln851_2_fu_1427_p2 : icmp_ln851_2_reg_2035;
assign _041_ = ap_CS_fsm[3] ? ret_V_19_fu_1415_p3 : ret_V_19_reg_2030;
assign _024_ = ap_CS_fsm[3] ? ret_V_17_fu_1284_p2[10:9] : p_Result_2_reg_2024;
assign _035_ = ap_CS_fsm[3] ? p_Val2_13_fu_1336_p2[3] : p_Result_43_reg_2017;
assign _036_ = ap_CS_fsm[3] ? p_Val2_13_fu_1336_p2 : p_Val2_13_reg_2012;
assign _034_ = ap_CS_fsm[3] ? ret_V_17_fu_1284_p2[10] : p_Result_40_reg_2006;
assign _040_ = ap_CS_fsm[3] ? ret_V_17_fu_1284_p2 : ret_V_17_reg_1999;
assign _019_ = ap_CS_fsm[3] ? op_17_V_fu_1262_p3 : op_17_V_reg_1994;
assign _018_ = ap_CS_fsm[0] ? op_16_V_fu_385_p2 : op_16_V_reg_1811;
assign _012_ = ap_CS_fsm[0] ? icmp_ln786_2_fu_373_p2 : icmp_ln786_2_reg_1806;
assign _009_ = ap_CS_fsm[0] ? icmp_ln768_fu_367_p2 : icmp_ln768_reg_1801;
assign _033_ = ap_CS_fsm[0] ? p_Result_39_fu_351_p2 : p_Result_39_reg_1794;
assign _032_ = ap_CS_fsm[0] ? ret_2_fu_327_p2[8] : p_Result_38_reg_1788;
assign _052_ = ap_CS_fsm[0] ? op_3_V_fu_279_p2[2:0] : trunc_ln1192_3_reg_1783;
assign _053_ = ap_CS_fsm[0] ? op_3_V_fu_279_p2[1:0] : trunc_ln1192_reg_1778;
assign _054_ = ap_CS_fsm[0] ? op_3_V_fu_279_p2[0] : trunc_ln703_reg_1773;
assign _049_ = ap_CS_fsm[0] ? { op_2[3], op_2[3], op_2[3], op_2[3], op_2 } : sext_ln69_reg_1767;
assign _021_ = ap_CS_fsm[0] ? op_3_V_fu_279_p2 : op_3_V_reg_1762;
assign _004_ = ap_CS_fsm[5] ? add_ln69_3_fu_1721_p2 : add_ln69_3_reg_2079;
assign _042_ = ap_CS_fsm[5] ? { ret_V_25_fu_1701_p2[38], ret_V_25_fu_1701_p2[38], ret_V_25_fu_1701_p2[38], ret_V_25_fu_1701_p2[38], ret_V_25_fu_1701_p2[38], ret_V_25_fu_1701_p2[38], ret_V_25_fu_1701_p2[38], ret_V_25_fu_1701_p2[38], ret_V_25_fu_1701_p2[38], ret_V_25_fu_1701_p2[38], ret_V_25_fu_1701_p2[38], ret_V_25_fu_1701_p2[38], ret_V_25_fu_1701_p2[38], ret_V_25_fu_1701_p2[38], ret_V_25_fu_1701_p2[38], ret_V_25_fu_1701_p2[38], ret_V_25_fu_1701_p2[38], ret_V_25_fu_1701_p2[38], ret_V_25_fu_1701_p2[38], ret_V_25_fu_1701_p2[38], ret_V_25_fu_1701_p2[38], ret_V_25_fu_1701_p2[38], ret_V_25_fu_1701_p2[38], ret_V_25_fu_1701_p2[38], ret_V_25_fu_1701_p2[38], ret_V_25_fu_1701_p2[38], ret_V_25_fu_1701_p2[11:6] } : ret_V_20_cast_reg_2072;
assign _045_ = ap_CS_fsm[5] ? { ret_V_25_fu_1701_p2[38], ret_V_25_fu_1701_p2[38], ret_V_25_fu_1701_p2[38], ret_V_25_fu_1701_p2[38], ret_V_25_fu_1701_p2[38], ret_V_25_fu_1701_p2[38], ret_V_25_fu_1701_p2[38], ret_V_25_fu_1701_p2[38], ret_V_25_fu_1701_p2[38], ret_V_25_fu_1701_p2[38], ret_V_25_fu_1701_p2[38], ret_V_25_fu_1701_p2[38], ret_V_25_fu_1701_p2[38], ret_V_25_fu_1701_p2[38], ret_V_25_fu_1701_p2[38], ret_V_25_fu_1701_p2[38], ret_V_25_fu_1701_p2[38], ret_V_25_fu_1701_p2[38], ret_V_25_fu_1701_p2[38], ret_V_25_fu_1701_p2[38], ret_V_25_fu_1701_p2[38], ret_V_25_fu_1701_p2[38], ret_V_25_fu_1701_p2[38], ret_V_25_fu_1701_p2[38], ret_V_25_fu_1701_p2[38], ret_V_25_fu_1701_p2[38], ret_V_25_fu_1701_p2[38], ret_V_25_fu_1701_p2[11:0] } : ret_V_25_reg_2067;
assign _048_ = ap_CS_fsm[1] ? select_ln384_5_fu_719_p3 : rhs_3_reg_1933[23:22];
assign _031_ = ap_CS_fsm[1] ? p_Val2_8_fu_654_p2[7] : p_Result_37_reg_1926;
assign _038_ = ap_CS_fsm[1] ? p_Val2_8_fu_654_p2 : p_Val2_8_reg_1920;
assign _030_ = ap_CS_fsm[1] ? add_ln1192_2_fu_588_p2[24] : p_Result_36_reg_1915;
assign _051_ = ap_CS_fsm[1] ? op_6[25:0] : trunc_ln1192_2_reg_1910;
assign _002_ = ap_CS_fsm[1] ? Range1_all_zeros_fu_571_p2 : Range1_all_zeros_reg_1905;
assign _001_ = ap_CS_fsm[1] ? Range1_all_ones_fu_565_p2 : Range1_all_ones_reg_1898;
assign _003_ = ap_CS_fsm[1] ? Range2_all_ones_fu_549_p2 : Range2_all_ones_reg_1893;
assign _028_ = ap_CS_fsm[1] ? op_6[24] : p_Result_33_reg_1887;
assign _056_ = ap_CS_fsm[1] ? xor_ln416_fu_525_p2 : xor_ln416_reg_1881;
assign _027_ = ap_CS_fsm[1] ? p_Val2_3_fu_511_p2[1] : p_Result_32_reg_1875;
assign _037_ = ap_CS_fsm[1] ? p_Val2_3_fu_511_p2 : p_Val2_3_reg_1866;
assign _026_ = ap_CS_fsm[1] ? op_6[23] : p_Result_31_reg_1861;
assign _025_ = ap_CS_fsm[1] ? op_6[31] : p_Result_30_reg_1854;
assign _013_ = ap_CS_fsm[1] ? icmp_ln790_fu_459_p2 : icmp_ln790_reg_1849;
assign _011_ = ap_CS_fsm[1] ? icmp_ln786_1_fu_441_p2 : icmp_ln786_1_reg_1844;
assign _010_ = ap_CS_fsm[1] ? icmp_ln785_fu_435_p2 : icmp_ln785_reg_1839;
assign _050_ = ap_CS_fsm[1] ? ret_fu_395_p2[2] : tmp_reg_1834;
assign _023_ = ap_CS_fsm[1] ? ret_fu_395_p2[7] : p_Result_29_reg_1828;
assign _047_ = ap_CS_fsm[1] ? ret_fu_395_p2 : ret_reg_1823;
assign _044_ = ap_CS_fsm[2] ? ret_V_23_fu_1186_p3 : ret_V_23_reg_1989;
assign _005_ = ap_CS_fsm[2] ? and_ln786_1_fu_1131_p2 : and_ln786_1_reg_1983;
assign _008_ = ap_CS_fsm[2] ? deleted_zeros_1_fu_1095_p3 : deleted_zeros_1_reg_1977;
assign _000_ = ap_CS_fsm[2] ? Range1_all_ones_1_fu_1083_p2 : Range1_all_ones_1_reg_1972;
assign _007_ = ap_CS_fsm[2] ? carry_3_fu_1052_p2 : carry_3_reg_1967;
assign _055_ = ap_CS_fsm[2] ? xor_ln416_1_fu_1047_p2 : xor_ln416_1_reg_1962;
assign _029_ = ap_CS_fsm[2] ? ret_V_16_fu_1028_p2[32] : p_Result_34_reg_1955;
assign _039_ = ap_CS_fsm[2] ? ret_V_15_fu_1001_p2 : ret_V_15_reg_1950;
assign _016_ = ap_CS_fsm[2] ? op_12_V_fu_982_p3 : op_12_V_reg_1944;
assign _022_ = ap_CS_fsm[2] ? op_8_V_fu_792_p3 : op_8_V_reg_1938;
assign _006_ = ap_rst ? 7'h01 : ap_NS_fsm;
assign ret_V_17_fu_1284_p2 = $signed({ 1'h0, op_7, 5'h00 }) - $signed(op_8_V_reg_1938);
assign ret_V_20_fu_1591_p2 = $signed(op_8_V_reg_1938) - $signed({ trunc_ln703_reg_1773, 6'h00 });
assign Range1_all_ones_1_fu_1083_p2 = _061_ ? 1'h1 : 1'h0;
assign Range1_all_ones_2_fu_1458_p2 = _062_ ? 1'h1 : 1'h0;
assign Range1_all_ones_fu_565_p2 = _063_ ? 1'h1 : 1'h0;
assign Range1_all_zeros_1_fu_1089_p2 = _064_ ? 1'h1 : 1'h0;
assign Range1_all_zeros_2_fu_1463_p2 = _065_ ? 1'h1 : 1'h0;
assign Range1_all_zeros_fu_571_p2 = _066_ ? 1'h1 : 1'h0;
assign Range2_all_ones_1_fu_1067_p2 = _067_ ? 1'h1 : 1'h0;
assign Range2_all_ones_fu_549_p2 = _068_ ? 1'h1 : 1'h0;
assign deleted_ones_1_fu_1123_p3 = carry_3_fu_1052_p2 ? and_ln780_1_fu_1117_p2 : Range1_all_ones_1_fu_1083_p2;
assign deleted_ones_2_fu_1495_p3 = carry_5_fu_1445_p2 ? and_ln780_2_fu_1489_p2 : Range1_all_ones_2_fu_1458_p2;
assign deleted_ones_fu_820_p3 = carry_1_fu_800_p2 ? and_ln780_fu_815_p2 : Range1_all_ones_reg_1898;
assign deleted_zeros_1_fu_1095_p3 = carry_3_fu_1052_p2 ? Range1_all_ones_1_fu_1083_p2 : Range1_all_zeros_1_fu_1089_p2;
assign deleted_zeros_2_fu_1468_p3 = carry_5_fu_1445_p2 ? Range1_all_ones_2_fu_1458_p2 : Range1_all_zeros_2_fu_1463_p2;
assign deleted_zeros_fu_804_p3 = carry_1_fu_800_p2 ? Range1_all_ones_reg_1898 : Range1_all_zeros_reg_1905;
assign icmp_ln414_fu_495_p2 = _073_ ? 1'h1 : 1'h0;
assign icmp_ln768_fu_367_p2 = _074_ ? 1'h1 : 1'h0;
assign icmp_ln785_fu_435_p2 = _075_ ? 1'h1 : 1'h0;
assign icmp_ln786_1_fu_441_p2 = _076_ ? 1'h1 : 1'h0;
assign icmp_ln786_2_fu_373_p2 = _077_ ? 1'h1 : 1'h0;
assign icmp_ln786_fu_757_p2 = _069_ ? 1'h1 : 1'h0;
assign icmp_ln790_fu_459_p2 = _070_ ? 1'h1 : 1'h0;
assign icmp_ln851_1_fu_1166_p2 = _071_ ? 1'h1 : 1'h0;
assign icmp_ln851_2_fu_1427_p2 = _078_ ? 1'h1 : 1'h0;
assign icmp_ln851_fu_1611_p2 = _072_ ? 1'h1 : 1'h0;
assign op_12_V_fu_982_p3 = sel_tmp11_fu_976_p2 ? p_Val2_3_reg_1866 : select_ln785_fu_945_p3;
assign op_15_V_fu_1567_p3 = or_ln384_2_fu_1561_p2 ? select_ln384_2_fu_1553_p3 : p_Val2_13_reg_2012;
assign op_17_V_fu_1262_p3 = and_ln785_5_fu_1257_p2 ? p_Val2_8_reg_1920 : select_ln340_1_fu_1241_p3;
assign op_8_V_fu_792_p3 = or_ln384_fu_786_p2 ? select_ln384_fu_778_p3 : { ret_reg_1823[2:0], 5'h00 };
assign r_1_fu_1320_p2 = _079_ ? 1'h1 : 1'h0;
assign r_fu_624_p2 = _080_ ? 1'h1 : 1'h0;
assign ret_V_19_fu_1415_p3 = ret_V_18_fu_1370_p2[3] ? select_ln850_fu_1407_p3 : { 2'h0, ret_V_18_fu_1370_p2[2:1] };
assign ret_V_21_fu_1654_p3 = ret_V_20_reg_2045[8] ? select_ln850_1_fu_1648_p3 : ret_V_reg_2050;
assign ret_V_23_fu_1186_p3 = ret_V_22_fu_1139_p2[31] ? select_ln850_2_fu_1178_p3 : ret_V_22_fu_1139_p2[26:23];
assign ret_V_26_fu_1745_p3 = ret_V_25_reg_2067[38] ? select_ln850_3_fu_1739_p3 : ret_V_20_cast_reg_2072;
assign select_ln340_1_fu_1241_p3 = or_ln340_4_fu_1235_p2 ? 8'h00 : p_Val2_8_reg_1920;
assign select_ln340_fu_922_p3 = or_ln340_1_fu_916_p2 ? { p_Result_33_reg_1887, p_Val2_4_fu_902_p2 } : p_Val2_3_reg_1866;
assign select_ln384_2_fu_1553_p3 = overflow_4_fu_1525_p2 ? 4'h7 : 4'h8;
assign select_ln384_4_fu_711_p3 = overflow_3_fu_684_p2 ? 2'h1 : 2'h2;
assign select_ln384_5_fu_719_p3 = or_ln384_1_fu_705_p2 ? select_ln384_4_fu_711_p3 : { p_Result_39_reg_1794, 1'h0 };
assign select_ln384_fu_778_p3 = overflow_fu_752_p2 ? 8'h7f : 8'h81;
assign select_ln703_fu_989_p3 = op_0 ? 3'h7 : 3'h0;
assign select_ln785_fu_945_p3 = and_ln785_1_fu_939_p2 ? p_Val2_3_reg_1866 : select_ln340_fu_922_p3;
assign select_ln850_1_fu_1648_p3 = icmp_ln851_reg_2057 ? ret_V_reg_2050 : ret_V_7_fu_1643_p2;
assign select_ln850_2_fu_1178_p3 = icmp_ln851_1_fu_1166_p2 ? ret_V_22_fu_1139_p2[26:23] : ret_V_10_fu_1172_p2;
assign select_ln850_3_fu_1739_p3 = icmp_ln851_2_reg_2035 ? add_ln691_3_fu_1734_p2 : ret_V_20_cast_reg_2072;
assign select_ln850_fu_1407_p3 = op_12_V_reg_1944[0] ? add_ln691_fu_1401_p2 : { 2'h3, ret_V_18_fu_1370_p2[2:1] };
assign xor_ln365_fu_890_p2 = p_Val2_3_reg_1866[1] ^ op_6[24];
assign p_Result_39_fu_351_p2 = op_5[0] ^ or_ln731_fu_345_p2;
assign Range2_all_ones_2_fu_1451_p3 = ret_V_17_reg_1999[10];
assign and_ln_fu_740_p3 = { tmp_reg_1834, 7'h00 };
assign ap_CS_fsm_state1 = ap_CS_fsm[0];
assign ap_CS_fsm_state2 = ap_CS_fsm[1];
assign ap_CS_fsm_state3 = ap_CS_fsm[2];
assign ap_CS_fsm_state4 = ap_CS_fsm[3];
assign ap_CS_fsm_state5 = ap_CS_fsm[4];
assign ap_CS_fsm_state6 = ap_CS_fsm[5];
assign ap_CS_fsm_state7 = ap_CS_fsm[6];
assign ap_done = op_28_ap_vld;
assign ap_ready = op_28_ap_vld;
assign empty_fu_391_p0 = op_6;
assign empty_fu_391_p1 = op_6[24:0];
assign lhs_V_1_fu_1007_p3 = { op_3_V_reg_1762, 23'h000000 };
assign lhs_V_3_fu_1269_p3 = { op_7, 5'h00 };
assign or_ln760_fu_379_p1 = op_2;
assign or_ln_fu_425_p4 = { ret_fu_395_p2[2], 2'h0, ret_fu_395_p2[7:3] };
assign p_Result_12_fu_907_p4 = { p_Result_33_reg_1887, p_Val2_4_fu_902_p2 };
assign p_Result_17_fu_604_p3 = add_ln1192_2_fu_588_p2[17];
assign p_Result_1_fu_539_p1 = op_6;
assign p_Result_1_fu_539_p4 = op_6[31:25];
assign p_Result_25_fu_1390_p3 = ret_V_18_fu_1370_p2[3];
assign p_Result_26_fu_1636_p3 = ret_V_20_reg_2045[8];
assign p_Result_27_fu_1154_p3 = ret_V_22_fu_1139_p2[31];
assign p_Result_28_fu_1727_p3 = ret_V_25_reg_2067[38];
assign p_Result_30_fu_465_p1 = op_6;
assign p_Result_30_fu_465_p3 = op_6[31];
assign p_Result_31_fu_483_p1 = op_6;
assign p_Result_32_fu_517_p3 = p_Val2_3_fu_511_p2[1];
assign p_Result_33_fu_531_p1 = op_6;
assign p_Result_35_fu_612_p1 = op_6;
assign p_Result_35_fu_612_p3 = op_6[16];
assign p_Result_3_fu_555_p1 = op_6;
assign p_Result_3_fu_555_p4 = op_6[31:24];
assign p_Result_41_fu_1308_p3 = ret_V_17_fu_1284_p2[4];
assign p_Result_42_fu_1433_p3 = ret_V_17_reg_1999[8];
assign p_Result_5_fu_1057_p4 = ret_V_16_fu_1028_p2[32:26];
assign p_Result_6_fu_1073_p4 = ret_V_16_fu_1028_p2[32:25];
assign p_Result_8_fu_357_p4 = ret_2_fu_327_p2[8:1];
assign p_Result_s_20_fu_451_p3 = { ret_fu_395_p2[1:0], 5'h00 };
assign p_Result_s_fu_415_p4 = ret_fu_395_p2[7:3];
assign p_Val2_10_fu_668_p3 = { p_Result_39_reg_1794, 1'h0 };
assign p_Val2_12_fu_1298_p4 = ret_V_17_fu_1284_p2[8:5];
assign p_Val2_1_fu_735_p2 = { ret_reg_1823[2:0], 5'h00 };
assign p_Val2_2_fu_473_p1 = op_6;
assign p_Val2_2_fu_473_p4 = op_6[23:22];
assign p_Val2_7_fu_594_p4 = add_ln1192_2_fu_588_p2[24:17];
assign ret_V_22_fu_1139_p1 = op_6;
assign ret_V_25_fu_1701_p2[37:12] = { ret_V_25_fu_1701_p2[38], ret_V_25_fu_1701_p2[38], ret_V_25_fu_1701_p2[38], ret_V_25_fu_1701_p2[38], ret_V_25_fu_1701_p2[38], ret_V_25_fu_1701_p2[38], ret_V_25_fu_1701_p2[38], ret_V_25_fu_1701_p2[38], ret_V_25_fu_1701_p2[38], ret_V_25_fu_1701_p2[38], ret_V_25_fu_1701_p2[38], ret_V_25_fu_1701_p2[38], ret_V_25_fu_1701_p2[38], ret_V_25_fu_1701_p2[38], ret_V_25_fu_1701_p2[38], ret_V_25_fu_1701_p2[38], ret_V_25_fu_1701_p2[38], ret_V_25_fu_1701_p2[38], ret_V_25_fu_1701_p2[38], ret_V_25_fu_1701_p2[38], ret_V_25_fu_1701_p2[38], ret_V_25_fu_1701_p2[38], ret_V_25_fu_1701_p2[38], ret_V_25_fu_1701_p2[38], ret_V_25_fu_1701_p2[38], ret_V_25_fu_1701_p2[38] };
assign ret_V_7_cast_fu_1144_p4 = ret_V_22_fu_1139_p2[26:23];
assign ret_fu_395_p0 = sext_ln69_reg_1767[3:0];
assign ret_fu_395_p1 = sext_ln69_reg_1767[3:0];
assign rhs_2_fu_1363_p3 = { ret_V_15_reg_1950, 1'h0 };
assign rhs_3_fu_727_p3 = { select_ln384_5_fu_719_p3, 22'h000000 };
assign rhs_fu_1580_p3 = { trunc_ln703_reg_1773, 6'h00 };
assign sext_ln1192_1_fu_1360_p1 = { op_12_V_reg_1944[1], op_12_V_reg_1944[1], op_12_V_reg_1944 };
assign sext_ln1192_2_fu_1668_p1 = { op_15_V_reg_2040[3], op_15_V_reg_2040[3], op_15_V_reg_2040 };
assign sext_ln1192_3_fu_1697_p1 = { op_25_V_fu_1680_p2[5], op_25_V_fu_1680_p2[5], op_25_V_fu_1680_p2[5], op_25_V_fu_1680_p2[5], op_25_V_fu_1680_p2[5], op_25_V_fu_1680_p2[5], op_25_V_fu_1680_p2[5], op_25_V_fu_1680_p2[5], op_25_V_fu_1680_p2[5], op_25_V_fu_1680_p2[5], op_25_V_fu_1680_p2[5], op_25_V_fu_1680_p2[5], op_25_V_fu_1680_p2[5], op_25_V_fu_1680_p2[5], op_25_V_fu_1680_p2[5], op_25_V_fu_1680_p2[5], op_25_V_fu_1680_p2[5], op_25_V_fu_1680_p2[5], op_25_V_fu_1680_p2[5], op_25_V_fu_1680_p2[5], op_25_V_fu_1680_p2[5], op_25_V_fu_1680_p2[5], op_25_V_fu_1680_p2[5], op_25_V_fu_1680_p2[5], op_25_V_fu_1680_p2[5], op_25_V_fu_1680_p2[5], op_25_V_fu_1680_p2[5], op_25_V_fu_1680_p2, 6'h00 };
assign sext_ln1192_fu_1014_p1 = { op_3_V_reg_1762[3], op_3_V_reg_1762[3], op_3_V_reg_1762[3], op_3_V_reg_1762[3], op_3_V_reg_1762[3], op_3_V_reg_1762[3], op_3_V_reg_1762, 23'h000000 };
assign sext_ln1193_fu_1587_p1 = { trunc_ln703_reg_1773, trunc_ln703_reg_1773, trunc_ln703_reg_1773, 6'h00 };
assign sext_ln1195_fu_1136_p1 = { rhs_3_reg_1933[23], rhs_3_reg_1933[23], rhs_3_reg_1933[23], rhs_3_reg_1933[23], rhs_3_reg_1933[23], rhs_3_reg_1933[23], rhs_3_reg_1933[23], rhs_3_reg_1933[23], rhs_3_reg_1933 };
assign sext_ln19_fu_1661_p1 = { ret_V_21_fu_1654_p3[3], ret_V_21_fu_1654_p3[3], ret_V_21_fu_1654_p3[3], ret_V_21_fu_1654_p3[3], ret_V_21_fu_1654_p3[3], ret_V_21_fu_1654_p3 };
assign sext_ln215_fu_319_p1 = { op_4_V_fu_301_p2[7], op_4_V_fu_301_p2 };
assign sext_ln23_fu_1665_p1 = { op_23_V_reg_2062[4], op_23_V_reg_2062 };
assign sext_ln69_1_fu_1617_p1 = { op_13[1], op_13[1], op_13[1], op_13 };
assign sext_ln69_2_fu_1621_p1 = { ret_V_23_reg_1989[3], ret_V_23_reg_1989 };
assign sext_ln69_3_fu_1677_p1 = { op_16_V_reg_1811[3], op_16_V_reg_1811[3], op_16_V_reg_1811 };
assign sext_ln69_4_fu_1717_p1 = { op_19[7], op_19 };
assign sext_ln69_5_fu_1752_p1 = { add_ln69_3_reg_2079[8], add_ln69_3_reg_2079[8], add_ln69_3_reg_2079[8], add_ln69_3_reg_2079[8], add_ln69_3_reg_2079[8], add_ln69_3_reg_2079[8], add_ln69_3_reg_2079[8], add_ln69_3_reg_2079[8], add_ln69_3_reg_2079[8], add_ln69_3_reg_2079[8], add_ln69_3_reg_2079[8], add_ln69_3_reg_2079[8], add_ln69_3_reg_2079[8], add_ln69_3_reg_2079[8], add_ln69_3_reg_2079[8], add_ln69_3_reg_2079[8], add_ln69_3_reg_2079[8], add_ln69_3_reg_2079[8], add_ln69_3_reg_2079[8], add_ln69_3_reg_2079[8], add_ln69_3_reg_2079[8], add_ln69_3_reg_2079[8], add_ln69_3_reg_2079[8], add_ln69_3_reg_2079 };
assign sext_ln69_fu_289_p0 = op_2;
assign sext_ln69_fu_289_p1 = { op_2[3], op_2[3], op_2[3], op_2[3], op_2 };
assign sext_ln703_1_fu_1018_p0 = op_6;
assign sext_ln703_1_fu_1018_p1 = { op_6[31], op_6 };
assign sext_ln703_2_fu_1281_p1 = { op_8_V_reg_1938[7], op_8_V_reg_1938[7], op_8_V_reg_1938[7], op_8_V_reg_1938 };
assign sext_ln703_3_fu_1577_p1 = { op_8_V_reg_1938[7], op_8_V_reg_1938 };
assign sext_ln703_4_fu_1686_p1 = { op_17_V_reg_1994[7], op_17_V_reg_1994[7], op_17_V_reg_1994[7], op_17_V_reg_1994[7], op_17_V_reg_1994[7], op_17_V_reg_1994[7], op_17_V_reg_1994[7], op_17_V_reg_1994[7], op_17_V_reg_1994[7], op_17_V_reg_1994[7], op_17_V_reg_1994[7], op_17_V_reg_1994[7], op_17_V_reg_1994[7], op_17_V_reg_1994[7], op_17_V_reg_1994[7], op_17_V_reg_1994[7], op_17_V_reg_1994[7], op_17_V_reg_1994[7], op_17_V_reg_1994[7], op_17_V_reg_1994[7], op_17_V_reg_1994[7], op_17_V_reg_1994[7], op_17_V_reg_1994[7], op_17_V_reg_1994[7], op_17_V_reg_1994[7], op_17_V_reg_1994[7], op_17_V_reg_1994[7], op_17_V_reg_1994[7], op_17_V_reg_1994[7], op_17_V_reg_1994[7], op_17_V_reg_1994[7], op_17_V_reg_1994 };
assign sext_ln703_fu_997_p1 = { op_9[1], op_9 };
assign sext_ln831_fu_1574_p1 = { ret_V_19_reg_2030[3], ret_V_19_reg_2030 };
assign sext_ln850_fu_1386_p1 = { ret_V_18_fu_1370_p2[3], ret_V_18_fu_1370_p2[3:1] };
assign tmp_14_fu_1103_p3 = add_ln1192_1_fu_1034_p2[25];
assign tmp_21_fu_1476_p3 = ret_V_17_reg_1999[9];
assign tmp_25_fu_1689_p3 = { op_25_V_fu_1680_p2, 6'h00 };
assign tmp_5_fu_1376_p4 = ret_V_18_fu_1370_p2[3:1];
assign tmp_6_fu_876_p1 = op_6;
assign tmp_6_fu_876_p3 = op_6[24];
assign tmp_7_fu_883_p3 = p_Val2_3_reg_1866[1];
assign tmp_fu_407_p3 = ret_fu_395_p2[2];
assign trunc_ln1192_1_fu_577_p3 = { trunc_ln1192_reg_1778, 23'h000000 };
assign trunc_ln1192_2_fu_584_p0 = op_6;
assign trunc_ln1192_2_fu_584_p1 = op_6[25:0];
assign trunc_ln1192_3_fu_315_p1 = op_3_V_fu_279_p2[2:0];
assign trunc_ln1192_4_fu_1021_p3 = { trunc_ln1192_3_reg_1783, 23'h000000 };
assign trunc_ln1192_fu_311_p1 = op_3_V_fu_279_p2[1:0];
assign trunc_ln414_fu_491_p0 = op_6;
assign trunc_ln414_fu_491_p1 = op_6[21:0];
assign trunc_ln69_1_fu_285_p1 = op_1[7:0];
assign trunc_ln69_2_fu_293_p1 = op_1[0];
assign trunc_ln69_3_fu_297_p0 = op_2;
assign trunc_ln69_3_fu_297_p1 = op_2[0];
assign trunc_ln69_fu_275_p1 = op_1[3:0];
assign trunc_ln703_fu_307_p1 = op_3_V_fu_279_p2[0];
assign trunc_ln718_1_fu_1316_p1 = ret_V_17_fu_1284_p2[3:0];
assign trunc_ln718_fu_620_p0 = op_6;
assign trunc_ln718_fu_620_p1 = op_6[15:0];
assign trunc_ln731_fu_341_p1 = op_5[0];
assign trunc_ln790_fu_447_p1 = ret_fu_395_p2[1:0];
assign trunc_ln851_1_fu_1607_p1 = ret_V_20_fu_1591_p2[4:0];
assign trunc_ln851_2_fu_1162_p1 = ret_V_22_fu_1139_p2[22:0];
assign trunc_ln851_3_fu_1423_p1 = op_17_V_fu_1262_p3[5:0];
assign trunc_ln851_fu_1398_p1 = op_12_V_reg_1944[0];
assign zext_ln1193_fu_1277_p1 = { 2'h0, op_7, 5'h00 };
assign zext_ln215_fu_323_p1 = { 7'h00, op_5 };
assign zext_ln415_1_fu_650_p1 = { 7'h00, and_ln412_fu_644_p2 };
assign zext_ln415_2_fu_1332_p1 = { 3'h0, and_ln408_fu_1326_p2 };
assign zext_ln415_fu_507_p1 = { 1'h0, and_ln414_fu_501_p2 };
assign \mul_4s_4s_8_1_1_U2.top_mul_4s_4s_8_1_1_Multiplier_1_U.a  = \mul_4s_4s_8_1_1_U2.din0 ;
assign \mul_4s_4s_8_1_1_U2.top_mul_4s_4s_8_1_1_Multiplier_1_U.b  = \mul_4s_4s_8_1_1_U2.din1 ;
assign \mul_4s_4s_8_1_1_U2.dout  = \mul_4s_4s_8_1_1_U2.top_mul_4s_4s_8_1_1_Multiplier_1_U.p ;
assign \mul_4s_4s_8_1_1_U2.din0  = sext_ln69_reg_1767[3:0];
assign \mul_4s_4s_8_1_1_U2.din1  = sext_ln69_reg_1767[3:0];
assign ret_fu_395_p2 = \mul_4s_4s_8_1_1_U2.dout ;
assign \mul_4s_4s_4_1_1_U1.top_mul_4s_4s_4_1_1_Multiplier_0_U.a  = \mul_4s_4s_4_1_1_U1.din0 ;
assign \mul_4s_4s_4_1_1_U1.top_mul_4s_4s_4_1_1_Multiplier_0_U.b  = \mul_4s_4s_4_1_1_U1.din1 ;
assign \mul_4s_4s_4_1_1_U1.dout  = \mul_4s_4s_4_1_1_U1.top_mul_4s_4s_4_1_1_Multiplier_0_U.p ;
assign \mul_4s_4s_4_1_1_U1.din0  = op_1[3:0];
assign \mul_4s_4s_4_1_1_U1.din1  = op_2;
assign op_3_V_fu_279_p2 = \mul_4s_4s_4_1_1_U1.dout ;
endmodule


// Product machine:
module top_A_times_top_B (ap_start, op_0, op_1, op_13, op_19, op_2, op_5, op_6, op_7, op_9, ap_clk, unsafe_signal);
input ap_start;
input op_0;
input [31:0] op_1;
input [1:0] op_13;
input [7:0] op_19;
input [3:0] op_2;
input [1:0] op_5;
input [31:0] op_6;
input [3:0] op_7;
input [1:0] op_9;
input ap_clk;
output unsafe_signal;
reg _setup;
initial _setup = 1'b0;
always @ (posedge ap_clk) _setup <= 1'b1;
reg ap_start_internal;
always @ (posedge ap_clk) if (!_setup) ap_start_internal <= ap_start;
reg op_0_internal;
always @ (posedge ap_clk) if (!_setup) op_0_internal <= op_0;
reg [31:0] op_1_internal;
always @ (posedge ap_clk) if (!_setup) op_1_internal <= op_1;
reg [1:0] op_13_internal;
always @ (posedge ap_clk) if (!_setup) op_13_internal <= op_13;
reg [7:0] op_19_internal;
always @ (posedge ap_clk) if (!_setup) op_19_internal <= op_19;
reg [3:0] op_2_internal;
always @ (posedge ap_clk) if (!_setup) op_2_internal <= op_2;
reg [1:0] op_5_internal;
always @ (posedge ap_clk) if (!_setup) op_5_internal <= op_5;
reg [31:0] op_6_internal;
always @ (posedge ap_clk) if (!_setup) op_6_internal <= op_6;
reg [3:0] op_7_internal;
always @ (posedge ap_clk) if (!_setup) op_7_internal <= op_7;
reg [1:0] op_9_internal;
always @ (posedge ap_clk) if (!_setup) op_9_internal <= op_9;
wire ap_done_A;
wire ap_done_B;
wire ap_done_eq;
assign ap_done_eq = ap_done_A == ap_done_B;
wire ap_idle_A;
wire ap_idle_B;
wire ap_idle_eq;
assign ap_idle_eq = ap_idle_A == ap_idle_B;
wire ap_ready_A;
wire ap_ready_B;
wire ap_ready_eq;
assign ap_ready_eq = ap_ready_A == ap_ready_B;
wire [31:0] op_28_A;
wire [31:0] op_28_B;
wire op_28_eq;
assign op_28_eq = op_28_A == op_28_B;
wire op_28_ap_vld_A;
wire op_28_ap_vld_B;
wire clk_enable_A;
wire clk_enable_B;
assign clk_enable_A = _setup & (~op_28_ap_vld_A | op_28_ap_vld_B);
assign clk_enable_B = _setup;
wire divergent;
assign divergent = ~(ap_done_eq & ap_idle_eq & ap_ready_eq & op_28_eq);
assign unsafe_signal = op_28_ap_vld_A & op_28_ap_vld_B & divergent;
top_A instance_A (
    .ap_clk(ap_clk),
    .clk_enable(clk_enable_A),
    .ap_start(ap_start_internal),
    .op_0(op_0_internal),
    .op_1(op_1_internal),
    .op_13(op_13_internal),
    .op_19(op_19_internal),
    .op_2(op_2_internal),
    .op_5(op_5_internal),
    .op_6(op_6_internal),
    .op_7(op_7_internal),
    .op_9(op_9_internal),
    .ap_done(ap_done_A),
    .ap_idle(ap_idle_A),
    .ap_ready(ap_ready_A),
    .op_28(op_28_A),
    .op_28_ap_vld(op_28_ap_vld_A)
);
top_B instance_B (
    .ap_clk(ap_clk),
    .clk_enable(clk_enable_B),
    .ap_start(ap_start_internal),
    .op_0(op_0_internal),
    .op_1(op_1_internal),
    .op_13(op_13_internal),
    .op_19(op_19_internal),
    .op_2(op_2_internal),
    .op_5(op_5_internal),
    .op_6(op_6_internal),
    .op_7(op_7_internal),
    .op_9(op_9_internal),
    .ap_done(ap_done_B),
    .ap_idle(ap_idle_B),
    .ap_ready(ap_ready_B),
    .op_28(op_28_B),
    .op_28_ap_vld(op_28_ap_vld_B)
);
endmodule
