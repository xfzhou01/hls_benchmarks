// Processed by function `construct_kairos` in `verilog_tricks.py`.
// Machine A:
// Processed by function `add_clk_enable_signal` in `verilog_tricks.py`.
// Processed by function `remove_reset_signal` in `verilog_tricks.py`.
module top_A (
  ap_clk,
  ap_start,
  ap_done,
  ap_idle,
  ap_ready,
  op_0,
  op_1,
  op_2,
  op_5,
  op_7,
  op_8,
  op_9,
  op_10,
  op_13,
  op_15,
  op_28,
  op_28_ap_vld,
clk_enable
);
input clk_enable;


input ap_clk;
wire ap_rst;
assign ap_rst = op_28_ap_vld;
input ap_start;
input [7:0] op_0;
input [15:0] op_1;
input [1:0] op_10;
input [1:0] op_13;
input [1:0] op_15;
input [7:0] op_2;
input [3:0] op_5;
input [3:0] op_7;
input [15:0] op_8;
input [3:0] op_9;
output ap_done;
output ap_idle;
output ap_ready;
output [31:0] op_28;
output op_28_ap_vld;


reg [7:0] \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.ain_s1 ;
reg [7:0] \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.bin_s1 ;
reg \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.carry_s1 ;
reg [7:0] \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.sum_s1 ;
reg [8:0] \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.ain_s1 ;
reg [8:0] \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.bin_s1 ;
reg \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.carry_s1 ;
reg [7:0] \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.sum_s1 ;
reg [8:0] \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.ain_s1 ;
reg [8:0] \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.bin_s1 ;
reg \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.carry_s1 ;
reg [8:0] \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.sum_s1 ;
reg [8:0] \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.ain_s1 ;
reg [8:0] \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.bin_s1 ;
reg \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.carry_s1 ;
reg [8:0] \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.sum_s1 ;
reg [8:0] \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.ain_s1 ;
reg [8:0] \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.bin_s1 ;
reg \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.carry_s1 ;
reg [8:0] \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.sum_s1 ;
reg [9:0] \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.ain_s1 ;
reg [9:0] \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.bin_s1 ;
reg \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.carry_s1 ;
reg [9:0] \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.sum_s1 ;
reg [9:0] \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.ain_s1 ;
reg [9:0] \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.bin_s1 ;
reg \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.carry_s1 ;
reg [9:0] \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.sum_s1 ;
reg [9:0] \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.ain_s1 ;
reg [9:0] \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.bin_s1 ;
reg \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.carry_s1 ;
reg [9:0] \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.sum_s1 ;
reg [9:0] \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.ain_s1 ;
reg [9:0] \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.bin_s1 ;
reg \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.carry_s1 ;
reg [9:0] \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.sum_s1 ;
reg [9:0] \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.ain_s1 ;
reg [9:0] \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.bin_s1 ;
reg \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.carry_s1 ;
reg [9:0] \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.sum_s1 ;
reg \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.ain_s1 ;
reg \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.bin_s1 ;
reg \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.carry_s1 ;
reg \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.sum_s1 ;
reg \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.ain_s1 ;
reg \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.bin_s1 ;
reg \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.carry_s1 ;
reg \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.sum_s1 ;
reg [1:0] \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.ain_s1 ;
reg [1:0] \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.bin_s1 ;
reg \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.carry_s1 ;
reg [1:0] \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.sum_s1 ;
reg [19:0] add_ln691_reg_980;
reg [3:0] add_ln69_1_reg_933;
reg [19:0] add_ln69_3_reg_995;
reg [16:0] add_ln69_4_reg_809;
reg [17:0] add_ln69_reg_928;
reg [24:0] ap_CS_fsm = 25'h0000001;
reg [3:0] \ashr_9ns_4ns_9_7_1_U7.din1_cast_array[0] ;
reg [3:0] \ashr_9ns_4ns_9_7_1_U7.din1_cast_array[1] ;
reg [3:0] \ashr_9ns_4ns_9_7_1_U7.din1_cast_array[2] ;
reg [3:0] \ashr_9ns_4ns_9_7_1_U7.din1_cast_array[3] ;
reg [3:0] \ashr_9ns_4ns_9_7_1_U7.din1_cast_array[4] ;
reg [3:0] \ashr_9ns_4ns_9_7_1_U7.din1_cast_array[5] ;
reg [8:0] \ashr_9ns_4ns_9_7_1_U7.dout_array[0] ;
reg [8:0] \ashr_9ns_4ns_9_7_1_U7.dout_array[1] ;
reg [8:0] \ashr_9ns_4ns_9_7_1_U7.dout_array[2] ;
reg [8:0] \ashr_9ns_4ns_9_7_1_U7.dout_array[3] ;
reg [8:0] \ashr_9ns_4ns_9_7_1_U7.dout_array[4] ;
reg [8:0] \ashr_9ns_4ns_9_7_1_U7.dout_array[5] ;
reg [8:0] ashr_ln1333_reg_871;
reg icmp_ln851_1_reg_876;
reg icmp_ln851_2_reg_834;
reg icmp_ln851_3_reg_784;
reg icmp_ln851_reg_726;
reg isNeg_reg_693;
reg [15:0] \mul_16s_4ns_16_7_1_U1.top_mul_16s_4ns_16_7_1_Mul_DSP_0_U.a_reg0 ;
reg [3:0] \mul_16s_4ns_16_7_1_U1.top_mul_16s_4ns_16_7_1_Mul_DSP_0_U.b_reg0 ;
reg [15:0] \mul_16s_4ns_16_7_1_U1.top_mul_16s_4ns_16_7_1_Mul_DSP_0_U.buff0 ;
reg [15:0] \mul_16s_4ns_16_7_1_U1.top_mul_16s_4ns_16_7_1_Mul_DSP_0_U.buff1 ;
reg [15:0] \mul_16s_4ns_16_7_1_U1.top_mul_16s_4ns_16_7_1_Mul_DSP_0_U.buff2 ;
reg [15:0] \mul_16s_4ns_16_7_1_U1.top_mul_16s_4ns_16_7_1_Mul_DSP_0_U.buff3 ;
reg [15:0] \mul_16s_4ns_16_7_1_U1.top_mul_16s_4ns_16_7_1_Mul_DSP_0_U.buff4 ;
reg [5:0] \mul_6s_6s_6_7_1_U3.top_mul_6s_6s_6_7_1_Mul_DSP_1_U.a_reg0 ;
reg [5:0] \mul_6s_6s_6_7_1_U3.top_mul_6s_6s_6_7_1_Mul_DSP_1_U.b_reg0 ;
reg [5:0] \mul_6s_6s_6_7_1_U3.top_mul_6s_6s_6_7_1_Mul_DSP_1_U.buff0 ;
reg [5:0] \mul_6s_6s_6_7_1_U3.top_mul_6s_6s_6_7_1_Mul_DSP_1_U.buff1 ;
reg [5:0] \mul_6s_6s_6_7_1_U3.top_mul_6s_6s_6_7_1_Mul_DSP_1_U.buff2 ;
reg [5:0] \mul_6s_6s_6_7_1_U3.top_mul_6s_6s_6_7_1_Mul_DSP_1_U.buff3 ;
reg [5:0] \mul_6s_6s_6_7_1_U3.top_mul_6s_6s_6_7_1_Mul_DSP_1_U.buff4 ;
reg [15:0] mul_ln728_reg_814;
reg [5:0] mul_ln731_reg_819;
reg [17:0] op_23_V_reg_943;
reg op_25_V_reg_898;
reg [3:0] r_reg_774;
reg [1:0] ret_V_12_reg_789;
reg [15:0] ret_V_17_reg_779;
reg [1:0] ret_V_19_reg_903;
reg [19:0] ret_V_20_reg_856;
reg [1:0] ret_V_21_cast_reg_756;
reg [17:0] ret_V_21_reg_908;
reg [16:0] ret_V_22_reg_751;
reg [1:0] ret_V_23_reg_804;
reg [19:0] ret_V_24_reg_963;
reg [19:0] ret_V_25_reg_985;
reg [15:0] ret_V_2_reg_746;
reg [1:0] ret_V_4_cast_reg_844;
reg [1:0] ret_V_5_reg_888;
reg [16:0] ret_V_8_reg_861;
reg [17:0] ret_V_9_reg_893;
reg [15:0] ret_V_reg_699;
reg [17:0] sext_ln835_reg_881;
reg [19:0] sext_ln850_reg_973;
reg [3:0] \shl_9ns_4ns_9_7_1_U6.din1_cast_array[0] ;
reg [3:0] \shl_9ns_4ns_9_7_1_U6.din1_cast_array[1] ;
reg [3:0] \shl_9ns_4ns_9_7_1_U6.din1_cast_array[2] ;
reg [3:0] \shl_9ns_4ns_9_7_1_U6.din1_cast_array[3] ;
reg [3:0] \shl_9ns_4ns_9_7_1_U6.din1_cast_array[4] ;
reg [3:0] \shl_9ns_4ns_9_7_1_U6.din1_cast_array[5] ;
reg [8:0] \shl_9ns_4ns_9_7_1_U6.dout_array[0] ;
reg [8:0] \shl_9ns_4ns_9_7_1_U6.dout_array[1] ;
reg [8:0] \shl_9ns_4ns_9_7_1_U6.dout_array[2] ;
reg [8:0] \shl_9ns_4ns_9_7_1_U6.dout_array[3] ;
reg [8:0] \shl_9ns_4ns_9_7_1_U6.dout_array[4] ;
reg [8:0] \shl_9ns_4ns_9_7_1_U6.dout_array[5] ;
reg [8:0] shl_ln1299_reg_866;
reg [8:0] \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.ain_s1 ;
reg [8:0] \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.bin_s1 ;
reg \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.carry_s1 ;
reg [7:0] \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.sum_s1 ;
reg [1:0] \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.ain_s1 ;
reg [1:0] \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.bin_s1 ;
reg \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.carry_s1 ;
reg [1:0] \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.sum_s1 ;
reg [3:0] sub_ln1367_reg_721;
reg [18:0] tmp_3_reg_968;
reg [8:0] trunc_ln1118_reg_682;
reg [1:0] trunc_ln851_1_reg_851;
reg [7:0] trunc_ln851_3_reg_763;
reg [24:0] trunc_ln851_reg_706;
reg [3:0] ush_reg_741;
reg [7:0] _561_;
wire [19:0] _000_;
wire [3:0] _001_;
wire [19:0] _002_;
wire [16:0] _003_;
wire [17:0] _004_;
wire [24:0] _005_;
wire [8:0] _006_;
wire _007_;
wire _008_;
wire _009_;
wire _010_;
wire _011_;
wire [15:0] _012_;
wire [5:0] _013_;
wire [17:0] _014_;
wire _015_;
wire [3:0] _016_;
wire [1:0] _017_;
wire [15:0] _018_;
wire [7:0] _019_;
wire [1:0] _020_;
wire [19:0] _021_;
wire [1:0] _022_;
wire [17:0] _023_;
wire [16:0] _024_;
wire [1:0] _025_;
wire [19:0] _026_;
wire [19:0] _027_;
wire [15:0] _028_;
wire [1:0] _029_;
wire [1:0] _030_;
wire [16:0] _031_;
wire [17:0] _032_;
wire [15:0] _033_;
wire [17:0] _034_;
wire [19:0] _035_;
wire [8:0] _036_;
wire [3:0] _037_;
wire [18:0] _038_;
wire [8:0] _039_;
wire [7:0] _040_;
wire [24:0] _041_;
wire [3:0] _042_;
wire [1:0] _043_;
wire _044_;
wire _045_;
wire _046_;
wire _047_;
wire _048_;
wire _049_;
wire _050_;
wire _051_;
wire _052_;
wire _053_;
wire _054_;
wire _055_;
wire [7:0] _056_;
wire [7:0] _057_;
wire _058_;
wire [7:0] _059_;
wire [8:0] _060_;
wire [8:0] _061_;
wire [8:0] _062_;
wire [8:0] _063_;
wire _064_;
wire [7:0] _065_;
wire [8:0] _066_;
wire [9:0] _067_;
wire [8:0] _068_;
wire [8:0] _069_;
wire _070_;
wire [8:0] _071_;
wire [9:0] _072_;
wire [9:0] _073_;
wire [8:0] _074_;
wire [8:0] _075_;
wire _076_;
wire [8:0] _077_;
wire [9:0] _078_;
wire [9:0] _079_;
wire [8:0] _080_;
wire [8:0] _081_;
wire _082_;
wire [8:0] _083_;
wire [9:0] _084_;
wire [9:0] _085_;
wire [9:0] _086_;
wire [9:0] _087_;
wire _088_;
wire [9:0] _089_;
wire [10:0] _090_;
wire [10:0] _091_;
wire [9:0] _092_;
wire [9:0] _093_;
wire _094_;
wire [9:0] _095_;
wire [10:0] _096_;
wire [10:0] _097_;
wire [9:0] _098_;
wire [9:0] _099_;
wire _100_;
wire [9:0] _101_;
wire [10:0] _102_;
wire [10:0] _103_;
wire [9:0] _104_;
wire [9:0] _105_;
wire _106_;
wire [9:0] _107_;
wire [10:0] _108_;
wire [10:0] _109_;
wire [9:0] _110_;
wire [9:0] _111_;
wire _112_;
wire [9:0] _113_;
wire [10:0] _114_;
wire [10:0] _115_;
wire _116_;
wire _117_;
wire _118_;
wire _119_;
wire [1:0] _120_;
wire [1:0] _121_;
wire _122_;
wire _123_;
wire _124_;
wire _125_;
wire [1:0] _126_;
wire [1:0] _127_;
wire [1:0] _128_;
wire [1:0] _129_;
wire _130_;
wire [1:0] _131_;
wire [2:0] _132_;
wire [2:0] _133_;
wire [3:0] _134_;
wire [3:0] _135_;
wire [3:0] _136_;
wire [3:0] _137_;
wire [3:0] _138_;
wire [3:0] _139_;
wire [8:0] _140_;
wire [8:0] _141_;
wire [8:0] _142_;
wire [8:0] _143_;
wire [8:0] _144_;
wire [8:0] _145_;
wire [3:0] _146_;
wire [8:0] _147_;
wire [3:0] _148_;
wire [8:0] _149_;
wire [3:0] _150_;
wire [8:0] _151_;
wire [3:0] _152_;
wire [8:0] _153_;
wire [3:0] _154_;
wire [8:0] _155_;
wire [3:0] _156_;
wire [8:0] _157_;
wire [8:0] _158_;
wire [8:0] _159_;
wire [8:0] _160_;
wire [15:0] _161_;
wire [3:0] _162_;
wire [15:0] _163_;
wire [15:0] _164_;
wire [15:0] _165_;
wire [15:0] _166_;
wire [15:0] _167_;
wire [5:0] _168_;
wire [5:0] _169_;
wire [5:0] _170_;
wire [5:0] _171_;
wire [5:0] _172_;
wire [5:0] _173_;
wire [5:0] _174_;
wire [3:0] _175_;
wire [3:0] _176_;
wire [3:0] _177_;
wire [3:0] _178_;
wire [3:0] _179_;
wire [3:0] _180_;
wire [8:0] _181_;
wire [8:0] _182_;
wire [8:0] _183_;
wire [8:0] _184_;
wire [8:0] _185_;
wire [8:0] _186_;
wire [3:0] _187_;
wire [8:0] _188_;
wire [3:0] _189_;
wire [8:0] _190_;
wire [3:0] _191_;
wire [8:0] _192_;
wire [3:0] _193_;
wire [8:0] _194_;
wire [3:0] _195_;
wire [8:0] _196_;
wire [3:0] _197_;
wire [8:0] _198_;
wire [8:0] _199_;
wire [8:0] _200_;
wire [8:0] _201_;
wire [8:0] _202_;
wire [8:0] _203_;
wire _204_;
wire [7:0] _205_;
wire [8:0] _206_;
wire [9:0] _207_;
wire [1:0] _208_;
wire [1:0] _209_;
wire _210_;
wire [1:0] _211_;
wire [2:0] _212_;
wire [2:0] _213_;
wire _214_;
wire _215_;
wire _216_;
wire _217_;
wire _218_;
wire _219_;
wire _220_;
wire _221_;
wire _222_;
wire _223_;
wire _224_;
wire _225_;
wire _226_;
wire _227_;
wire _228_;
wire _229_;
wire _230_;
wire _231_;
wire _232_;
wire _233_;
wire _234_;
wire _235_;
wire _236_;
wire _237_;
wire _238_;
wire \add_16ns_16ns_16_2_1_U4.ce ;
wire \add_16ns_16ns_16_2_1_U4.clk ;
wire [15:0] \add_16ns_16ns_16_2_1_U4.din0 ;
wire [15:0] \add_16ns_16ns_16_2_1_U4.din1 ;
wire [15:0] \add_16ns_16ns_16_2_1_U4.dout ;
wire \add_16ns_16ns_16_2_1_U4.reset ;
wire [15:0] \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.a ;
wire [15:0] \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.ain_s0 ;
wire [15:0] \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.b ;
wire [15:0] \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.bin_s0 ;
wire \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.ce ;
wire \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.clk ;
wire \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.facout_s1 ;
wire \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.facout_s2 ;
wire [7:0] \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.fas_s1 ;
wire [7:0] \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.fas_s2 ;
wire \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.reset ;
wire [15:0] \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.s ;
wire [7:0] \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.u1.a ;
wire [7:0] \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.u1.b ;
wire \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.u1.cin ;
wire \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.u1.cout ;
wire [7:0] \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.u1.s ;
wire [7:0] \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.u2.a ;
wire [7:0] \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.u2.b ;
wire \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.u2.cin ;
wire \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.u2.cout ;
wire [7:0] \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.u2.s ;
wire \add_17s_17s_17_2_1_U9.ce ;
wire \add_17s_17s_17_2_1_U9.clk ;
wire [16:0] \add_17s_17s_17_2_1_U9.din0 ;
wire [16:0] \add_17s_17s_17_2_1_U9.din1 ;
wire [16:0] \add_17s_17s_17_2_1_U9.dout ;
wire \add_17s_17s_17_2_1_U9.reset ;
wire [16:0] \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.a ;
wire [16:0] \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.ain_s0 ;
wire [16:0] \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.b ;
wire [16:0] \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.bin_s0 ;
wire \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.ce ;
wire \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.clk ;
wire \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.facout_s1 ;
wire \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.facout_s2 ;
wire [7:0] \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.fas_s1 ;
wire [8:0] \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.fas_s2 ;
wire \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.reset ;
wire [16:0] \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.s ;
wire [7:0] \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.u1.a ;
wire [7:0] \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.u1.b ;
wire \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.u1.cin ;
wire \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.u1.cout ;
wire [7:0] \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.u1.s ;
wire [8:0] \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.u2.a ;
wire [8:0] \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.u2.b ;
wire \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.u2.cin ;
wire \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.u2.cout ;
wire [8:0] \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.u2.s ;
wire \add_18ns_18ns_18_2_1_U13.ce ;
wire \add_18ns_18ns_18_2_1_U13.clk ;
wire [17:0] \add_18ns_18ns_18_2_1_U13.din0 ;
wire [17:0] \add_18ns_18ns_18_2_1_U13.din1 ;
wire [17:0] \add_18ns_18ns_18_2_1_U13.dout ;
wire \add_18ns_18ns_18_2_1_U13.reset ;
wire [17:0] \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.a ;
wire [17:0] \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.ain_s0 ;
wire [17:0] \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.b ;
wire [17:0] \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.bin_s0 ;
wire \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.ce ;
wire \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.clk ;
wire \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.facout_s1 ;
wire \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.facout_s2 ;
wire [8:0] \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.fas_s1 ;
wire [8:0] \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.fas_s2 ;
wire \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.reset ;
wire [17:0] \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.s ;
wire [8:0] \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.u1.a ;
wire [8:0] \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.u1.b ;
wire \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.u1.cin ;
wire \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.u1.cout ;
wire [8:0] \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.u1.s ;
wire [8:0] \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.u2.a ;
wire [8:0] \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.u2.b ;
wire \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.u2.cin ;
wire \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.u2.cout ;
wire [8:0] \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.u2.s ;
wire \add_18s_18ns_18_2_1_U12.ce ;
wire \add_18s_18ns_18_2_1_U12.clk ;
wire [17:0] \add_18s_18ns_18_2_1_U12.din0 ;
wire [17:0] \add_18s_18ns_18_2_1_U12.din1 ;
wire [17:0] \add_18s_18ns_18_2_1_U12.dout ;
wire \add_18s_18ns_18_2_1_U12.reset ;
wire [17:0] \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.a ;
wire [17:0] \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.ain_s0 ;
wire [17:0] \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.b ;
wire [17:0] \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.bin_s0 ;
wire \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.ce ;
wire \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.clk ;
wire \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.facout_s1 ;
wire \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.facout_s2 ;
wire [8:0] \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.fas_s1 ;
wire [8:0] \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.fas_s2 ;
wire \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.reset ;
wire [17:0] \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.s ;
wire [8:0] \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.u1.a ;
wire [8:0] \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.u1.b ;
wire \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.u1.cin ;
wire \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.u1.cout ;
wire [8:0] \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.u1.s ;
wire [8:0] \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.u2.a ;
wire [8:0] \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.u2.b ;
wire \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.u2.cin ;
wire \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.u2.cout ;
wire [8:0] \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.u2.s ;
wire \add_18s_18ns_18_2_1_U15.ce ;
wire \add_18s_18ns_18_2_1_U15.clk ;
wire [17:0] \add_18s_18ns_18_2_1_U15.din0 ;
wire [17:0] \add_18s_18ns_18_2_1_U15.din1 ;
wire [17:0] \add_18s_18ns_18_2_1_U15.dout ;
wire \add_18s_18ns_18_2_1_U15.reset ;
wire [17:0] \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.a ;
wire [17:0] \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.ain_s0 ;
wire [17:0] \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.b ;
wire [17:0] \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.bin_s0 ;
wire \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.ce ;
wire \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.clk ;
wire \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.facout_s1 ;
wire \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.facout_s2 ;
wire [8:0] \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.fas_s1 ;
wire [8:0] \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.fas_s2 ;
wire \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.reset ;
wire [17:0] \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.s ;
wire [8:0] \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.u1.a ;
wire [8:0] \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.u1.b ;
wire \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.u1.cin ;
wire \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.u1.cout ;
wire [8:0] \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.u1.s ;
wire [8:0] \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.u2.a ;
wire [8:0] \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.u2.b ;
wire \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.u2.cin ;
wire \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.u2.cout ;
wire [8:0] \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.u2.s ;
wire \add_20ns_20ns_20_2_1_U18.ce ;
wire \add_20ns_20ns_20_2_1_U18.clk ;
wire [19:0] \add_20ns_20ns_20_2_1_U18.din0 ;
wire [19:0] \add_20ns_20ns_20_2_1_U18.din1 ;
wire [19:0] \add_20ns_20ns_20_2_1_U18.dout ;
wire \add_20ns_20ns_20_2_1_U18.reset ;
wire [19:0] \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.a ;
wire [19:0] \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.ain_s0 ;
wire [19:0] \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.b ;
wire [19:0] \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.bin_s0 ;
wire \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.ce ;
wire \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.clk ;
wire \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.facout_s1 ;
wire \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.facout_s2 ;
wire [9:0] \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.fas_s1 ;
wire [9:0] \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.fas_s2 ;
wire \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.reset ;
wire [19:0] \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.s ;
wire [9:0] \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.u1.a ;
wire [9:0] \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.u1.b ;
wire \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.u1.cin ;
wire \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.u1.cout ;
wire [9:0] \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.u1.s ;
wire [9:0] \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.u2.a ;
wire [9:0] \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.u2.b ;
wire \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.u2.cin ;
wire \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.u2.cout ;
wire [9:0] \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.u2.s ;
wire \add_20ns_20s_20_2_1_U10.ce ;
wire \add_20ns_20s_20_2_1_U10.clk ;
wire [19:0] \add_20ns_20s_20_2_1_U10.din0 ;
wire [19:0] \add_20ns_20s_20_2_1_U10.din1 ;
wire [19:0] \add_20ns_20s_20_2_1_U10.dout ;
wire \add_20ns_20s_20_2_1_U10.reset ;
wire [19:0] \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.a ;
wire [19:0] \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.ain_s0 ;
wire [19:0] \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.b ;
wire [19:0] \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.bin_s0 ;
wire \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.ce ;
wire \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.clk ;
wire \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.facout_s1 ;
wire \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.facout_s2 ;
wire [9:0] \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.fas_s1 ;
wire [9:0] \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.fas_s2 ;
wire \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.reset ;
wire [19:0] \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.s ;
wire [9:0] \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.u1.a ;
wire [9:0] \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.u1.b ;
wire \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.u1.cin ;
wire \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.u1.cout ;
wire [9:0] \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.u1.s ;
wire [9:0] \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.u2.a ;
wire [9:0] \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.u2.b ;
wire \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.u2.cin ;
wire \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.u2.cout ;
wire [9:0] \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.u2.s ;
wire \add_20s_20ns_20_2_1_U17.ce ;
wire \add_20s_20ns_20_2_1_U17.clk ;
wire [19:0] \add_20s_20ns_20_2_1_U17.din0 ;
wire [19:0] \add_20s_20ns_20_2_1_U17.din1 ;
wire [19:0] \add_20s_20ns_20_2_1_U17.dout ;
wire \add_20s_20ns_20_2_1_U17.reset ;
wire [19:0] \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.a ;
wire [19:0] \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.ain_s0 ;
wire [19:0] \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.b ;
wire [19:0] \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.bin_s0 ;
wire \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.ce ;
wire \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.clk ;
wire \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.facout_s1 ;
wire \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.facout_s2 ;
wire [9:0] \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.fas_s1 ;
wire [9:0] \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.fas_s2 ;
wire \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.reset ;
wire [19:0] \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.s ;
wire [9:0] \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.u1.a ;
wire [9:0] \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.u1.b ;
wire \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.u1.cin ;
wire \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.u1.cout ;
wire [9:0] \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.u1.s ;
wire [9:0] \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.u2.a ;
wire [9:0] \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.u2.b ;
wire \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.u2.cin ;
wire \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.u2.cout ;
wire [9:0] \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.u2.s ;
wire \add_20s_20ns_20_2_1_U19.ce ;
wire \add_20s_20ns_20_2_1_U19.clk ;
wire [19:0] \add_20s_20ns_20_2_1_U19.din0 ;
wire [19:0] \add_20s_20ns_20_2_1_U19.din1 ;
wire [19:0] \add_20s_20ns_20_2_1_U19.dout ;
wire \add_20s_20ns_20_2_1_U19.reset ;
wire [19:0] \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.a ;
wire [19:0] \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.ain_s0 ;
wire [19:0] \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.b ;
wire [19:0] \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.bin_s0 ;
wire \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.ce ;
wire \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.clk ;
wire \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.facout_s1 ;
wire \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.facout_s2 ;
wire [9:0] \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.fas_s1 ;
wire [9:0] \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.fas_s2 ;
wire \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.reset ;
wire [19:0] \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.s ;
wire [9:0] \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.u1.a ;
wire [9:0] \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.u1.b ;
wire \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.u1.cin ;
wire \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.u1.cout ;
wire [9:0] \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.u1.s ;
wire [9:0] \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.u2.a ;
wire [9:0] \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.u2.b ;
wire \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.u2.cin ;
wire \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.u2.cout ;
wire [9:0] \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.u2.s ;
wire \add_20s_20s_20_2_1_U16.ce ;
wire \add_20s_20s_20_2_1_U16.clk ;
wire [19:0] \add_20s_20s_20_2_1_U16.din0 ;
wire [19:0] \add_20s_20s_20_2_1_U16.din1 ;
wire [19:0] \add_20s_20s_20_2_1_U16.dout ;
wire \add_20s_20s_20_2_1_U16.reset ;
wire [19:0] \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.a ;
wire [19:0] \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.ain_s0 ;
wire [19:0] \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.b ;
wire [19:0] \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.bin_s0 ;
wire \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.ce ;
wire \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.clk ;
wire \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.facout_s1 ;
wire \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.facout_s2 ;
wire [9:0] \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.fas_s1 ;
wire [9:0] \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.fas_s2 ;
wire \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.reset ;
wire [19:0] \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.s ;
wire [9:0] \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.u1.a ;
wire [9:0] \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.u1.b ;
wire \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.u1.cin ;
wire \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.u1.cout ;
wire [9:0] \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.u1.s ;
wire [9:0] \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.u2.a ;
wire [9:0] \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.u2.b ;
wire \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.u2.cin ;
wire \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.u2.cout ;
wire [9:0] \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.u2.s ;
wire \add_2ns_2ns_2_2_1_U11.ce ;
wire \add_2ns_2ns_2_2_1_U11.clk ;
wire [1:0] \add_2ns_2ns_2_2_1_U11.din0 ;
wire [1:0] \add_2ns_2ns_2_2_1_U11.din1 ;
wire [1:0] \add_2ns_2ns_2_2_1_U11.dout ;
wire \add_2ns_2ns_2_2_1_U11.reset ;
wire [1:0] \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.a ;
wire [1:0] \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.ain_s0 ;
wire [1:0] \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.b ;
wire [1:0] \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.bin_s0 ;
wire \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.ce ;
wire \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.clk ;
wire \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.facout_s1 ;
wire \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.facout_s2 ;
wire \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.fas_s1 ;
wire \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.fas_s2 ;
wire \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.reset ;
wire [1:0] \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.s ;
wire \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.u1.a ;
wire \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.u1.b ;
wire \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.u1.cin ;
wire \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.u1.cout ;
wire \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.u1.s ;
wire \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.u2.a ;
wire \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.u2.b ;
wire \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.u2.cin ;
wire \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.u2.cout ;
wire \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.u2.s ;
wire \add_2ns_2ns_2_2_1_U8.ce ;
wire \add_2ns_2ns_2_2_1_U8.clk ;
wire [1:0] \add_2ns_2ns_2_2_1_U8.din0 ;
wire [1:0] \add_2ns_2ns_2_2_1_U8.din1 ;
wire [1:0] \add_2ns_2ns_2_2_1_U8.dout ;
wire \add_2ns_2ns_2_2_1_U8.reset ;
wire [1:0] \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.a ;
wire [1:0] \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.ain_s0 ;
wire [1:0] \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.b ;
wire [1:0] \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.bin_s0 ;
wire \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.ce ;
wire \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.clk ;
wire \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.facout_s1 ;
wire \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.facout_s2 ;
wire \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.fas_s1 ;
wire \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.fas_s2 ;
wire \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.reset ;
wire [1:0] \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.s ;
wire \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.u1.a ;
wire \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.u1.b ;
wire \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.u1.cin ;
wire \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.u1.cout ;
wire \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.u1.s ;
wire \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.u2.a ;
wire \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.u2.b ;
wire \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.u2.cin ;
wire \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.u2.cout ;
wire \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.u2.s ;
wire \add_4s_4ns_4_2_1_U14.ce ;
wire \add_4s_4ns_4_2_1_U14.clk ;
wire [3:0] \add_4s_4ns_4_2_1_U14.din0 ;
wire [3:0] \add_4s_4ns_4_2_1_U14.din1 ;
wire [3:0] \add_4s_4ns_4_2_1_U14.dout ;
wire \add_4s_4ns_4_2_1_U14.reset ;
wire [3:0] \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.a ;
wire [3:0] \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.ain_s0 ;
wire [3:0] \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.b ;
wire [3:0] \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.bin_s0 ;
wire \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.ce ;
wire \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.clk ;
wire \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.facout_s1 ;
wire \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.facout_s2 ;
wire [1:0] \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.fas_s1 ;
wire [1:0] \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.fas_s2 ;
wire \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.reset ;
wire [3:0] \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.s ;
wire [1:0] \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.u1.a ;
wire [1:0] \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.u1.b ;
wire \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.u1.cin ;
wire \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.u1.cout ;
wire [1:0] \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.u1.s ;
wire [1:0] \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.u2.a ;
wire [1:0] \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.u2.b ;
wire \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.u2.cin ;
wire \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.u2.cout ;
wire [1:0] \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.u2.s ;
wire ap_CS_fsm_state1;
wire ap_CS_fsm_state10;
wire ap_CS_fsm_state11;
wire ap_CS_fsm_state12;
wire ap_CS_fsm_state13;
wire ap_CS_fsm_state14;
wire ap_CS_fsm_state15;
wire ap_CS_fsm_state16;
wire ap_CS_fsm_state17;
wire ap_CS_fsm_state18;
wire ap_CS_fsm_state19;
wire ap_CS_fsm_state2;
wire ap_CS_fsm_state20;
wire ap_CS_fsm_state21;
wire ap_CS_fsm_state22;
wire ap_CS_fsm_state23;
wire ap_CS_fsm_state24;
wire ap_CS_fsm_state25;
wire ap_CS_fsm_state3;
wire ap_CS_fsm_state4;
wire ap_CS_fsm_state5;
wire ap_CS_fsm_state6;
wire ap_CS_fsm_state7;
wire ap_CS_fsm_state8;
wire ap_CS_fsm_state9;
wire [24:0] ap_NS_fsm;
wire ap_clk;
wire ap_done;
wire ap_idle;
wire ap_ready;
wire ap_rst;
wire ap_start;
wire \ashr_9ns_4ns_9_7_1_U7.ce ;
wire \ashr_9ns_4ns_9_7_1_U7.clk ;
wire [8:0] \ashr_9ns_4ns_9_7_1_U7.din0 ;
wire [8:0] \ashr_9ns_4ns_9_7_1_U7.din1 ;
wire [3:0] \ashr_9ns_4ns_9_7_1_U7.din1_cast ;
wire [3:0] \ashr_9ns_4ns_9_7_1_U7.din1_mask ;
wire [8:0] \ashr_9ns_4ns_9_7_1_U7.dout ;
wire \ashr_9ns_4ns_9_7_1_U7.reset ;
wire [3:0] grp_fu_201_p1;
wire [15:0] grp_fu_201_p10;
wire [15:0] grp_fu_201_p2;
wire [3:0] grp_fu_215_p2;
wire [5:0] grp_fu_257_p0;
wire [5:0] grp_fu_257_p1;
wire [5:0] grp_fu_257_p2;
wire [15:0] grp_fu_276_p2;
wire [16:0] grp_fu_297_p0;
wire [16:0] grp_fu_297_p1;
wire [16:0] grp_fu_297_p2;
wire [8:0] grp_fu_325_p2;
wire [8:0] grp_fu_330_p2;
wire [1:0] grp_fu_364_p2;
wire [16:0] grp_fu_375_p0;
wire [16:0] grp_fu_375_p1;
wire [16:0] grp_fu_375_p2;
wire [19:0] grp_fu_415_p0;
wire [19:0] grp_fu_415_p1;
wire [19:0] grp_fu_415_p2;
wire [1:0] grp_fu_485_p2;
wire [17:0] grp_fu_493_p0;
wire [17:0] grp_fu_493_p2;
wire [17:0] grp_fu_566_p1;
wire [17:0] grp_fu_566_p2;
wire [3:0] grp_fu_571_p0;
wire [3:0] grp_fu_571_p1;
wire [3:0] grp_fu_571_p2;
wire [17:0] grp_fu_580_p0;
wire [17:0] grp_fu_580_p2;
wire [19:0] grp_fu_600_p0;
wire [19:0] grp_fu_600_p1;
wire [19:0] grp_fu_600_p2;
wire [19:0] grp_fu_619_p0;
wire [19:0] grp_fu_619_p2;
wire [19:0] grp_fu_651_p0;
wire [19:0] grp_fu_651_p2;
wire [19:0] grp_fu_659_p0;
wire [19:0] grp_fu_659_p2;
wire icmp_ln851_1_fu_480_p2;
wire icmp_ln851_2_fu_425_p2;
wire icmp_ln851_3_fu_359_p2;
wire icmp_ln851_fu_271_p2;
wire [9:0] lhs_V_fu_438_p3;
wire \mul_16s_4ns_16_7_1_U1.ce ;
wire \mul_16s_4ns_16_7_1_U1.clk ;
wire [15:0] \mul_16s_4ns_16_7_1_U1.din0 ;
wire [3:0] \mul_16s_4ns_16_7_1_U1.din1 ;
wire [15:0] \mul_16s_4ns_16_7_1_U1.dout ;
wire \mul_16s_4ns_16_7_1_U1.reset ;
wire [15:0] \mul_16s_4ns_16_7_1_U1.top_mul_16s_4ns_16_7_1_Mul_DSP_0_U.a ;
wire [3:0] \mul_16s_4ns_16_7_1_U1.top_mul_16s_4ns_16_7_1_Mul_DSP_0_U.b ;
wire \mul_16s_4ns_16_7_1_U1.top_mul_16s_4ns_16_7_1_Mul_DSP_0_U.ce ;
wire \mul_16s_4ns_16_7_1_U1.top_mul_16s_4ns_16_7_1_Mul_DSP_0_U.clk ;
wire [15:0] \mul_16s_4ns_16_7_1_U1.top_mul_16s_4ns_16_7_1_Mul_DSP_0_U.p ;
wire [15:0] \mul_16s_4ns_16_7_1_U1.top_mul_16s_4ns_16_7_1_Mul_DSP_0_U.tmp_product ;
wire \mul_6s_6s_6_7_1_U3.ce ;
wire \mul_6s_6s_6_7_1_U3.clk ;
wire [5:0] \mul_6s_6s_6_7_1_U3.din0 ;
wire [5:0] \mul_6s_6s_6_7_1_U3.din1 ;
wire [5:0] \mul_6s_6s_6_7_1_U3.dout ;
wire \mul_6s_6s_6_7_1_U3.reset ;
wire [5:0] \mul_6s_6s_6_7_1_U3.top_mul_6s_6s_6_7_1_Mul_DSP_1_U.a ;
wire [5:0] \mul_6s_6s_6_7_1_U3.top_mul_6s_6s_6_7_1_Mul_DSP_1_U.b ;
wire \mul_6s_6s_6_7_1_U3.top_mul_6s_6s_6_7_1_Mul_DSP_1_U.ce ;
wire \mul_6s_6s_6_7_1_U3.top_mul_6s_6s_6_7_1_Mul_DSP_1_U.clk ;
wire [5:0] \mul_6s_6s_6_7_1_U3.top_mul_6s_6s_6_7_1_Mul_DSP_1_U.p ;
wire [5:0] \mul_6s_6s_6_7_1_U3.top_mul_6s_6s_6_7_1_Mul_DSP_1_U.tmp_product ;
wire [7:0] op_0;
wire [15:0] op_1;
wire [1:0] op_10;
wire [1:0] op_13;
wire [1:0] op_15;
wire op_16_V_fu_505_p3;
wire [7:0] op_2;
wire op_25_V_fu_512_p2;
wire [31:0] op_28;
wire op_28_ap_vld;
wire [7:0] op_4_V_fu_431_p3;
wire [3:0] op_5;
wire [15:0] op_6_V_fu_263_p3;
wire [3:0] op_7;
wire [15:0] op_8;
wire [3:0] op_9;
wire p_Result_1_fu_518_p3;
wire p_Result_2_fu_537_p3;
wire p_Result_3_fu_381_p3;
wire p_Result_4_fu_625_p3;
wire [15:0] p_Result_s_fu_340_p1;
wire p_Result_s_fu_340_p3;
wire [3:0] r_fu_335_p2;
wire [40:0] ret_V_16_fu_229_p2;
wire [15:0] ret_V_17_fu_352_p3;
wire [9:0] ret_V_18_fu_450_p2;
wire [9:0] ret_V_18_reg_839;
wire [1:0] ret_V_19_fu_530_p3;
wire [17:0] ret_V_21_fu_549_p3;
wire [1:0] ret_V_23_fu_393_p3;
wire [19:0] ret_V_25_fu_641_p3;
wire [18:0] rhs_2_fu_404_p3;
wire [9:0] rhs_3_fu_285_p3;
wire [15:0] rhs_fu_221_p1;
wire [40:0] rhs_fu_221_p3;
wire [1:0] select_ln850_1_fu_525_p3;
wire [17:0] select_ln850_2_fu_544_p3;
wire [1:0] select_ln850_3_fu_388_p3;
wire [19:0] select_ln850_4_fu_635_p3;
wire [15:0] select_ln850_fu_347_p3;
wire [1:0] sext_ln1192_1_fu_585_p0;
wire [3:0] sext_ln1192_fu_400_p0;
wire [9:0] sext_ln703_fu_446_p1;
wire [17:0] sext_ln835_fu_490_p1;
wire [19:0] sext_ln850_fu_616_p1;
wire \shl_9ns_4ns_9_7_1_U6.ce ;
wire \shl_9ns_4ns_9_7_1_U6.clk ;
wire [8:0] \shl_9ns_4ns_9_7_1_U6.din0 ;
wire [8:0] \shl_9ns_4ns_9_7_1_U6.din1 ;
wire [3:0] \shl_9ns_4ns_9_7_1_U6.din1_cast ;
wire [3:0] \shl_9ns_4ns_9_7_1_U6.din1_mask ;
wire [8:0] \shl_9ns_4ns_9_7_1_U6.dout ;
wire \shl_9ns_4ns_9_7_1_U6.reset ;
wire \sub_17ns_17ns_17_2_1_U5.ce ;
wire \sub_17ns_17ns_17_2_1_U5.clk ;
wire [16:0] \sub_17ns_17ns_17_2_1_U5.din0 ;
wire [16:0] \sub_17ns_17ns_17_2_1_U5.din1 ;
wire [16:0] \sub_17ns_17ns_17_2_1_U5.dout ;
wire \sub_17ns_17ns_17_2_1_U5.reset ;
wire [16:0] \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.a ;
wire [16:0] \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.ain_s0 ;
wire [16:0] \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.b ;
wire [16:0] \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.bin_s0 ;
wire \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.ce ;
wire \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.clk ;
wire \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.facout_s1 ;
wire \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.facout_s2 ;
wire [7:0] \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.fas_s1 ;
wire [8:0] \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.fas_s2 ;
wire \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.reset ;
wire [16:0] \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.s ;
wire [7:0] \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.u1.a ;
wire [7:0] \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.u1.b ;
wire \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.u1.cin ;
wire \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.u1.cout ;
wire [7:0] \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.u1.s ;
wire [8:0] \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.u2.a ;
wire [8:0] \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.u2.b ;
wire \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.u2.cin ;
wire \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.u2.cout ;
wire [8:0] \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.u2.s ;
wire \sub_4ns_4ns_4_2_1_U2.ce ;
wire \sub_4ns_4ns_4_2_1_U2.clk ;
wire [3:0] \sub_4ns_4ns_4_2_1_U2.din0 ;
wire [3:0] \sub_4ns_4ns_4_2_1_U2.din1 ;
wire [3:0] \sub_4ns_4ns_4_2_1_U2.dout ;
wire \sub_4ns_4ns_4_2_1_U2.reset ;
wire [3:0] \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.a ;
wire [3:0] \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.ain_s0 ;
wire [3:0] \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.b ;
wire [3:0] \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.bin_s0 ;
wire \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.ce ;
wire \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.clk ;
wire \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.facout_s1 ;
wire \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.facout_s2 ;
wire [1:0] \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.fas_s1 ;
wire [1:0] \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.fas_s2 ;
wire \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.reset ;
wire [3:0] \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.s ;
wire [1:0] \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.u1.a ;
wire [1:0] \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.u1.b ;
wire \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.u1.cin ;
wire \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.u1.cout ;
wire [1:0] \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.u1.s ;
wire [1:0] \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.u2.a ;
wire [1:0] \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.u2.b ;
wire \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.u2.cin ;
wire \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.u2.cout ;
wire [1:0] \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.u2.s ;
wire [18:0] tmp_fu_589_p3;
wire [15:0] trunc_ln1118_fu_193_p0;
wire [8:0] trunc_ln1118_fu_193_p1;
wire trunc_ln1368_1_fu_502_p1;
wire trunc_ln1368_fu_499_p1;
wire [1:0] trunc_ln851_1_fu_466_p1;
wire [3:0] trunc_ln851_2_fu_421_p0;
wire [2:0] trunc_ln851_2_fu_421_p1;
wire [7:0] trunc_ln851_3_fu_318_p1;
wire [1:0] trunc_ln851_4_fu_632_p0;
wire trunc_ln851_4_fu_632_p1;
wire [24:0] trunc_ln851_fu_245_p1;
wire [3:0] ush_fu_303_p3;
wire [8:0] zext_ln1367_fu_322_p1;


assign _044_ = _049_ & ap_CS_fsm[9];
assign _045_ = ap_CS_fsm[10] & _050_;
assign _046_ = isNeg_reg_693 & ap_CS_fsm[9];
assign _047_ = _051_ & ap_CS_fsm[0];
assign _048_ = ap_start & ap_CS_fsm[0];
assign op_25_V_fu_512_p2 = ~ op_16_V_fu_505_p3;
assign r_fu_335_p2 = ~ op_9;
assign ret_V_16_fu_229_p2[25] = ~ op_8[0];
assign _049_ = ~ isNeg_reg_693;
assign _050_ = ~ icmp_ln851_2_reg_834;
assign _051_ = ~ ap_start;
assign _052_ = ! trunc_ln851_1_reg_851;
assign _053_ = ! op_7[2:0];
assign _054_ = ! trunc_ln851_3_reg_763;
assign _055_ = ! trunc_ln851_reg_706;
always @(posedge \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.clk )
\add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.bin_s1  <= _057_;
always @(posedge \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.clk )
\add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.ain_s1  <= _056_;
always @(posedge \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.clk )
\add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.sum_s1  <= _059_;
always @(posedge \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.clk )
\add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.carry_s1  <= _058_;
assign _057_ = \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.ce  ? \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.b [15:8] : \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.bin_s1 ;
assign _056_ = \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.ce  ? \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.a [15:8] : \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.ain_s1 ;
assign _058_ = \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.ce  ? \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.facout_s1  : \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.carry_s1 ;
assign _059_ = \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.ce  ? \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.fas_s1  : \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.sum_s1 ;
assign _060_ = \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.u1.a  + \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.u1.b ;
assign { \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.u1.cout , \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.u1.s  } = _060_ + \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.u1.cin ;
assign _061_ = \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.u2.a  + \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.u2.b ;
assign { \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.u2.cout , \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.u2.s  } = _061_ + \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.u2.cin ;
always @(posedge \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.clk )
\add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.bin_s1  <= _063_;
always @(posedge \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.clk )
\add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.ain_s1  <= _062_;
always @(posedge \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.clk )
\add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.sum_s1  <= _065_;
always @(posedge \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.clk )
\add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.carry_s1  <= _064_;
assign _063_ = \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.ce  ? \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.b [16:8] : \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.bin_s1 ;
assign _062_ = \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.ce  ? \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.a [16:8] : \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.ain_s1 ;
assign _064_ = \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.ce  ? \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.facout_s1  : \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.carry_s1 ;
assign _065_ = \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.ce  ? \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.fas_s1  : \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.sum_s1 ;
assign _066_ = \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.u1.a  + \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.u1.b ;
assign { \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.u1.cout , \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.u1.s  } = _066_ + \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.u1.cin ;
assign _067_ = \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.u2.a  + \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.u2.b ;
assign { \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.u2.cout , \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.u2.s  } = _067_ + \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.u2.cin ;
always @(posedge \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.clk )
\add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.bin_s1  <= _069_;
always @(posedge \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.clk )
\add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.ain_s1  <= _068_;
always @(posedge \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.clk )
\add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.sum_s1  <= _071_;
always @(posedge \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.clk )
\add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.carry_s1  <= _070_;
assign _069_ = \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.ce  ? \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.b [17:9] : \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.bin_s1 ;
assign _068_ = \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.ce  ? \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.a [17:9] : \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.ain_s1 ;
assign _070_ = \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.ce  ? \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.facout_s1  : \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.carry_s1 ;
assign _071_ = \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.ce  ? \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.fas_s1  : \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.sum_s1 ;
assign _072_ = \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.u1.a  + \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.u1.b ;
assign { \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.u1.cout , \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.u1.s  } = _072_ + \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.u1.cin ;
assign _073_ = \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.u2.a  + \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.u2.b ;
assign { \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.u2.cout , \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.u2.s  } = _073_ + \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.u2.cin ;
always @(posedge \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.clk )
\add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.bin_s1  <= _075_;
always @(posedge \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.clk )
\add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.ain_s1  <= _074_;
always @(posedge \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.clk )
\add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.sum_s1  <= _077_;
always @(posedge \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.clk )
\add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.carry_s1  <= _076_;
assign _075_ = \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.ce  ? \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.b [17:9] : \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.bin_s1 ;
assign _074_ = \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.ce  ? \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.a [17:9] : \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.ain_s1 ;
assign _076_ = \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.ce  ? \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.facout_s1  : \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.carry_s1 ;
assign _077_ = \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.ce  ? \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.fas_s1  : \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.sum_s1 ;
assign _078_ = \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.u1.a  + \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.u1.b ;
assign { \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.u1.cout , \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.u1.s  } = _078_ + \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.u1.cin ;
assign _079_ = \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.u2.a  + \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.u2.b ;
assign { \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.u2.cout , \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.u2.s  } = _079_ + \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.u2.cin ;
always @(posedge \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.clk )
\add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.bin_s1  <= _081_;
always @(posedge \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.clk )
\add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.ain_s1  <= _080_;
always @(posedge \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.clk )
\add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.sum_s1  <= _083_;
always @(posedge \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.clk )
\add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.carry_s1  <= _082_;
assign _081_ = \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.ce  ? \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.b [17:9] : \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.bin_s1 ;
assign _080_ = \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.ce  ? \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.a [17:9] : \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.ain_s1 ;
assign _082_ = \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.ce  ? \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.facout_s1  : \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.carry_s1 ;
assign _083_ = \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.ce  ? \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.fas_s1  : \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.sum_s1 ;
assign _084_ = \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.u1.a  + \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.u1.b ;
assign { \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.u1.cout , \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.u1.s  } = _084_ + \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.u1.cin ;
assign _085_ = \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.u2.a  + \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.u2.b ;
assign { \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.u2.cout , \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.u2.s  } = _085_ + \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.u2.cin ;
always @(posedge \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.clk )
\add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.bin_s1  <= _087_;
always @(posedge \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.clk )
\add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.ain_s1  <= _086_;
always @(posedge \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.clk )
\add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.sum_s1  <= _089_;
always @(posedge \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.clk )
\add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.carry_s1  <= _088_;
assign _087_ = \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.ce  ? \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.b [19:10] : \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.bin_s1 ;
assign _086_ = \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.ce  ? \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.a [19:10] : \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.ain_s1 ;
assign _088_ = \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.ce  ? \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.facout_s1  : \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.carry_s1 ;
assign _089_ = \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.ce  ? \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.fas_s1  : \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.sum_s1 ;
assign _090_ = \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.u1.a  + \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.u1.b ;
assign { \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.u1.cout , \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.u1.s  } = _090_ + \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.u1.cin ;
assign _091_ = \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.u2.a  + \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.u2.b ;
assign { \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.u2.cout , \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.u2.s  } = _091_ + \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.u2.cin ;
always @(posedge \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.clk )
\add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.bin_s1  <= _093_;
always @(posedge \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.clk )
\add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.ain_s1  <= _092_;
always @(posedge \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.clk )
\add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.sum_s1  <= _095_;
always @(posedge \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.clk )
\add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.carry_s1  <= _094_;
assign _093_ = \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.ce  ? \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.b [19:10] : \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.bin_s1 ;
assign _092_ = \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.ce  ? \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.a [19:10] : \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.ain_s1 ;
assign _094_ = \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.ce  ? \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.facout_s1  : \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.carry_s1 ;
assign _095_ = \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.ce  ? \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.fas_s1  : \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.sum_s1 ;
assign _096_ = \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.u1.a  + \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.u1.b ;
assign { \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.u1.cout , \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.u1.s  } = _096_ + \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.u1.cin ;
assign _097_ = \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.u2.a  + \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.u2.b ;
assign { \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.u2.cout , \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.u2.s  } = _097_ + \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.u2.cin ;
always @(posedge \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.clk )
\add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.bin_s1  <= _099_;
always @(posedge \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.clk )
\add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.ain_s1  <= _098_;
always @(posedge \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.clk )
\add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.sum_s1  <= _101_;
always @(posedge \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.clk )
\add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.carry_s1  <= _100_;
assign _099_ = \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.ce  ? \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.b [19:10] : \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.bin_s1 ;
assign _098_ = \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.ce  ? \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.a [19:10] : \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.ain_s1 ;
assign _100_ = \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.ce  ? \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.facout_s1  : \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.carry_s1 ;
assign _101_ = \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.ce  ? \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.fas_s1  : \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.sum_s1 ;
assign _102_ = \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.u1.a  + \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.u1.b ;
assign { \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.u1.cout , \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.u1.s  } = _102_ + \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.u1.cin ;
assign _103_ = \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.u2.a  + \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.u2.b ;
assign { \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.u2.cout , \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.u2.s  } = _103_ + \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.u2.cin ;
always @(posedge \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.clk )
\add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.bin_s1  <= _105_;
always @(posedge \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.clk )
\add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.ain_s1  <= _104_;
always @(posedge \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.clk )
\add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.sum_s1  <= _107_;
always @(posedge \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.clk )
\add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.carry_s1  <= _106_;
assign _105_ = \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.ce  ? \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.b [19:10] : \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.bin_s1 ;
assign _104_ = \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.ce  ? \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.a [19:10] : \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.ain_s1 ;
assign _106_ = \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.ce  ? \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.facout_s1  : \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.carry_s1 ;
assign _107_ = \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.ce  ? \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.fas_s1  : \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.sum_s1 ;
assign _108_ = \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.u1.a  + \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.u1.b ;
assign { \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.u1.cout , \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.u1.s  } = _108_ + \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.u1.cin ;
assign _109_ = \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.u2.a  + \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.u2.b ;
assign { \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.u2.cout , \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.u2.s  } = _109_ + \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.u2.cin ;
always @(posedge \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.clk )
\add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.bin_s1  <= _111_;
always @(posedge \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.clk )
\add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.ain_s1  <= _110_;
always @(posedge \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.clk )
\add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.sum_s1  <= _113_;
always @(posedge \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.clk )
\add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.carry_s1  <= _112_;
assign _111_ = \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.ce  ? \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.b [19:10] : \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.bin_s1 ;
assign _110_ = \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.ce  ? \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.a [19:10] : \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.ain_s1 ;
assign _112_ = \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.ce  ? \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.facout_s1  : \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.carry_s1 ;
assign _113_ = \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.ce  ? \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.fas_s1  : \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.sum_s1 ;
assign _114_ = \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.u1.a  + \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.u1.b ;
assign { \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.u1.cout , \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.u1.s  } = _114_ + \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.u1.cin ;
assign _115_ = \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.u2.a  + \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.u2.b ;
assign { \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.u2.cout , \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.u2.s  } = _115_ + \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.u2.cin ;
always @(posedge \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.clk )
\add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.bin_s1  <= _117_;
always @(posedge \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.clk )
\add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.ain_s1  <= _116_;
always @(posedge \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.clk )
\add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.sum_s1  <= _119_;
always @(posedge \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.clk )
\add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.carry_s1  <= _118_;
assign _117_ = \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.ce  ? \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.b [1] : \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.bin_s1 ;
assign _116_ = \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.ce  ? \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.a [1] : \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.ain_s1 ;
assign _118_ = \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.ce  ? \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.facout_s1  : \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.carry_s1 ;
assign _119_ = \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.ce  ? \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.fas_s1  : \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.sum_s1 ;
assign _120_ = \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.u1.a  + \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.u1.b ;
assign { \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.u1.cout , \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.u1.s  } = _120_ + \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.u1.cin ;
assign _121_ = \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.u2.a  + \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.u2.b ;
assign { \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.u2.cout , \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.u2.s  } = _121_ + \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.u2.cin ;
always @(posedge \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.clk )
\add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.bin_s1  <= _123_;
always @(posedge \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.clk )
\add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.ain_s1  <= _122_;
always @(posedge \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.clk )
\add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.sum_s1  <= _125_;
always @(posedge \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.clk )
\add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.carry_s1  <= _124_;
assign _123_ = \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.ce  ? \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.b [1] : \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.bin_s1 ;
assign _122_ = \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.ce  ? \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.a [1] : \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.ain_s1 ;
assign _124_ = \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.ce  ? \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.facout_s1  : \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.carry_s1 ;
assign _125_ = \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.ce  ? \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.fas_s1  : \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.sum_s1 ;
assign _126_ = \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.u1.a  + \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.u1.b ;
assign { \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.u1.cout , \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.u1.s  } = _126_ + \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.u1.cin ;
assign _127_ = \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.u2.a  + \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.u2.b ;
assign { \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.u2.cout , \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.u2.s  } = _127_ + \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.u2.cin ;
always @(posedge \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.clk )
\add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.bin_s1  <= _129_;
always @(posedge \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.clk )
\add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.ain_s1  <= _128_;
always @(posedge \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.clk )
\add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.sum_s1  <= _131_;
always @(posedge \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.clk )
\add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.carry_s1  <= _130_;
assign _129_ = \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.ce  ? \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.b [3:2] : \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.bin_s1 ;
assign _128_ = \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.ce  ? \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.a [3:2] : \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.ain_s1 ;
assign _130_ = \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.ce  ? \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.facout_s1  : \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.carry_s1 ;
assign _131_ = \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.ce  ? \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.fas_s1  : \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.sum_s1 ;
assign _132_ = \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.u1.a  + \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.u1.b ;
assign { \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.u1.cout , \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.u1.s  } = _132_ + \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.u1.cin ;
assign _133_ = \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.u2.a  + \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.u2.b ;
assign { \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.u2.cout , \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.u2.s  } = _133_ + \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.u2.cin ;
always @(posedge \ashr_9ns_4ns_9_7_1_U7.clk )
\ashr_9ns_4ns_9_7_1_U7.dout_array[5]  <= _145_;
always @(posedge \ashr_9ns_4ns_9_7_1_U7.clk )
\ashr_9ns_4ns_9_7_1_U7.din1_cast_array[5]  <= _139_;
always @(posedge \ashr_9ns_4ns_9_7_1_U7.clk )
\ashr_9ns_4ns_9_7_1_U7.dout_array[4]  <= _144_;
always @(posedge \ashr_9ns_4ns_9_7_1_U7.clk )
\ashr_9ns_4ns_9_7_1_U7.din1_cast_array[4]  <= _138_;
always @(posedge \ashr_9ns_4ns_9_7_1_U7.clk )
\ashr_9ns_4ns_9_7_1_U7.dout_array[3]  <= _143_;
always @(posedge \ashr_9ns_4ns_9_7_1_U7.clk )
\ashr_9ns_4ns_9_7_1_U7.din1_cast_array[3]  <= _137_;
always @(posedge \ashr_9ns_4ns_9_7_1_U7.clk )
\ashr_9ns_4ns_9_7_1_U7.dout_array[2]  <= _142_;
always @(posedge \ashr_9ns_4ns_9_7_1_U7.clk )
\ashr_9ns_4ns_9_7_1_U7.din1_cast_array[2]  <= _136_;
always @(posedge \ashr_9ns_4ns_9_7_1_U7.clk )
\ashr_9ns_4ns_9_7_1_U7.dout_array[1]  <= _141_;
always @(posedge \ashr_9ns_4ns_9_7_1_U7.clk )
\ashr_9ns_4ns_9_7_1_U7.din1_cast_array[1]  <= _135_;
always @(posedge \ashr_9ns_4ns_9_7_1_U7.clk )
\ashr_9ns_4ns_9_7_1_U7.dout_array[0]  <= _140_;
always @(posedge \ashr_9ns_4ns_9_7_1_U7.clk )
\ashr_9ns_4ns_9_7_1_U7.din1_cast_array[0]  <= _134_;
assign _146_ = \ashr_9ns_4ns_9_7_1_U7.ce  ? \ashr_9ns_4ns_9_7_1_U7.din1_cast_array[4]  : \ashr_9ns_4ns_9_7_1_U7.din1_cast_array[5] ;
assign _139_ = \ashr_9ns_4ns_9_7_1_U7.reset  ? 4'h0 : _146_;
assign _147_ = \ashr_9ns_4ns_9_7_1_U7.ce  ? _160_ : \ashr_9ns_4ns_9_7_1_U7.dout_array[5] ;
assign _145_ = \ashr_9ns_4ns_9_7_1_U7.reset  ? 9'h000 : _147_;
assign _148_ = \ashr_9ns_4ns_9_7_1_U7.ce  ? \ashr_9ns_4ns_9_7_1_U7.din1_cast_array[3]  : \ashr_9ns_4ns_9_7_1_U7.din1_cast_array[4] ;
assign _138_ = \ashr_9ns_4ns_9_7_1_U7.reset  ? 4'h0 : _148_;
assign _149_ = \ashr_9ns_4ns_9_7_1_U7.ce  ? _159_ : \ashr_9ns_4ns_9_7_1_U7.dout_array[4] ;
assign _144_ = \ashr_9ns_4ns_9_7_1_U7.reset  ? 9'h000 : _149_;
assign _150_ = \ashr_9ns_4ns_9_7_1_U7.ce  ? \ashr_9ns_4ns_9_7_1_U7.din1_cast_array[2]  : \ashr_9ns_4ns_9_7_1_U7.din1_cast_array[3] ;
assign _137_ = \ashr_9ns_4ns_9_7_1_U7.reset  ? 4'h0 : _150_;
assign _151_ = \ashr_9ns_4ns_9_7_1_U7.ce  ? _158_ : \ashr_9ns_4ns_9_7_1_U7.dout_array[3] ;
assign _143_ = \ashr_9ns_4ns_9_7_1_U7.reset  ? 9'h000 : _151_;
assign _152_ = \ashr_9ns_4ns_9_7_1_U7.ce  ? \ashr_9ns_4ns_9_7_1_U7.din1_cast_array[1]  : \ashr_9ns_4ns_9_7_1_U7.din1_cast_array[2] ;
assign _136_ = \ashr_9ns_4ns_9_7_1_U7.reset  ? 4'h0 : _152_;
assign _153_ = \ashr_9ns_4ns_9_7_1_U7.ce  ? \ashr_9ns_4ns_9_7_1_U7.dout_array[1]  : \ashr_9ns_4ns_9_7_1_U7.dout_array[2] ;
assign _142_ = \ashr_9ns_4ns_9_7_1_U7.reset  ? 9'h000 : _153_;
assign _154_ = \ashr_9ns_4ns_9_7_1_U7.ce  ? \ashr_9ns_4ns_9_7_1_U7.din1_cast_array[0]  : \ashr_9ns_4ns_9_7_1_U7.din1_cast_array[1] ;
assign _135_ = \ashr_9ns_4ns_9_7_1_U7.reset  ? 4'h0 : _154_;
assign _155_ = \ashr_9ns_4ns_9_7_1_U7.ce  ? \ashr_9ns_4ns_9_7_1_U7.dout_array[0]  : \ashr_9ns_4ns_9_7_1_U7.dout_array[1] ;
assign _141_ = \ashr_9ns_4ns_9_7_1_U7.reset  ? 9'h000 : _155_;
assign _156_ = \ashr_9ns_4ns_9_7_1_U7.ce  ? \ashr_9ns_4ns_9_7_1_U7.din1 [3:0] : \ashr_9ns_4ns_9_7_1_U7.din1_cast_array[0] ;
assign _134_ = \ashr_9ns_4ns_9_7_1_U7.reset  ? 4'h0 : _156_;
assign _157_ = \ashr_9ns_4ns_9_7_1_U7.ce  ? \ashr_9ns_4ns_9_7_1_U7.din0  : \ashr_9ns_4ns_9_7_1_U7.dout_array[0] ;
assign _140_ = \ashr_9ns_4ns_9_7_1_U7.reset  ? 9'h000 : _157_;
assign _158_ = $signed(\ashr_9ns_4ns_9_7_1_U7.dout_array[2] ) >>> { \ashr_9ns_4ns_9_7_1_U7.din1_cast_array[2] [3], 3'h0 };
assign _159_ = $signed(\ashr_9ns_4ns_9_7_1_U7.dout_array[3] ) >>> { \ashr_9ns_4ns_9_7_1_U7.din1_cast_array[3] [2], 2'h0 };
assign _160_ = $signed(\ashr_9ns_4ns_9_7_1_U7.dout_array[4] ) >>> { \ashr_9ns_4ns_9_7_1_U7.din1_cast_array[4] [1], 1'h0 };
assign \ashr_9ns_4ns_9_7_1_U7.dout  = $signed(\ashr_9ns_4ns_9_7_1_U7.dout_array[5] ) >>> \ashr_9ns_4ns_9_7_1_U7.din1_cast_array[5] [0];
assign \mul_16s_4ns_16_7_1_U1.top_mul_16s_4ns_16_7_1_Mul_DSP_0_U.tmp_product  = $signed(\mul_16s_4ns_16_7_1_U1.top_mul_16s_4ns_16_7_1_Mul_DSP_0_U.a_reg0 ) * $signed({ 1'h0, \mul_16s_4ns_16_7_1_U1.top_mul_16s_4ns_16_7_1_Mul_DSP_0_U.b_reg0  });
always @(posedge \mul_16s_4ns_16_7_1_U1.top_mul_16s_4ns_16_7_1_Mul_DSP_0_U.clk )
\mul_16s_4ns_16_7_1_U1.top_mul_16s_4ns_16_7_1_Mul_DSP_0_U.a_reg0  <= _161_;
always @(posedge \mul_16s_4ns_16_7_1_U1.top_mul_16s_4ns_16_7_1_Mul_DSP_0_U.clk )
\mul_16s_4ns_16_7_1_U1.top_mul_16s_4ns_16_7_1_Mul_DSP_0_U.b_reg0  <= _162_;
always @(posedge \mul_16s_4ns_16_7_1_U1.top_mul_16s_4ns_16_7_1_Mul_DSP_0_U.clk )
\mul_16s_4ns_16_7_1_U1.top_mul_16s_4ns_16_7_1_Mul_DSP_0_U.buff0  <= _163_;
always @(posedge \mul_16s_4ns_16_7_1_U1.top_mul_16s_4ns_16_7_1_Mul_DSP_0_U.clk )
\mul_16s_4ns_16_7_1_U1.top_mul_16s_4ns_16_7_1_Mul_DSP_0_U.buff1  <= _164_;
always @(posedge \mul_16s_4ns_16_7_1_U1.top_mul_16s_4ns_16_7_1_Mul_DSP_0_U.clk )
\mul_16s_4ns_16_7_1_U1.top_mul_16s_4ns_16_7_1_Mul_DSP_0_U.buff2  <= _165_;
always @(posedge \mul_16s_4ns_16_7_1_U1.top_mul_16s_4ns_16_7_1_Mul_DSP_0_U.clk )
\mul_16s_4ns_16_7_1_U1.top_mul_16s_4ns_16_7_1_Mul_DSP_0_U.buff3  <= _166_;
always @(posedge \mul_16s_4ns_16_7_1_U1.top_mul_16s_4ns_16_7_1_Mul_DSP_0_U.clk )
\mul_16s_4ns_16_7_1_U1.top_mul_16s_4ns_16_7_1_Mul_DSP_0_U.buff4  <= _167_;
assign _167_ = \mul_16s_4ns_16_7_1_U1.top_mul_16s_4ns_16_7_1_Mul_DSP_0_U.ce  ? \mul_16s_4ns_16_7_1_U1.top_mul_16s_4ns_16_7_1_Mul_DSP_0_U.buff3  : \mul_16s_4ns_16_7_1_U1.top_mul_16s_4ns_16_7_1_Mul_DSP_0_U.buff4 ;
assign _166_ = \mul_16s_4ns_16_7_1_U1.top_mul_16s_4ns_16_7_1_Mul_DSP_0_U.ce  ? \mul_16s_4ns_16_7_1_U1.top_mul_16s_4ns_16_7_1_Mul_DSP_0_U.buff2  : \mul_16s_4ns_16_7_1_U1.top_mul_16s_4ns_16_7_1_Mul_DSP_0_U.buff3 ;
assign _165_ = \mul_16s_4ns_16_7_1_U1.top_mul_16s_4ns_16_7_1_Mul_DSP_0_U.ce  ? \mul_16s_4ns_16_7_1_U1.top_mul_16s_4ns_16_7_1_Mul_DSP_0_U.buff1  : \mul_16s_4ns_16_7_1_U1.top_mul_16s_4ns_16_7_1_Mul_DSP_0_U.buff2 ;
assign _164_ = \mul_16s_4ns_16_7_1_U1.top_mul_16s_4ns_16_7_1_Mul_DSP_0_U.ce  ? \mul_16s_4ns_16_7_1_U1.top_mul_16s_4ns_16_7_1_Mul_DSP_0_U.buff0  : \mul_16s_4ns_16_7_1_U1.top_mul_16s_4ns_16_7_1_Mul_DSP_0_U.buff1 ;
assign _163_ = \mul_16s_4ns_16_7_1_U1.top_mul_16s_4ns_16_7_1_Mul_DSP_0_U.ce  ? \mul_16s_4ns_16_7_1_U1.top_mul_16s_4ns_16_7_1_Mul_DSP_0_U.tmp_product  : \mul_16s_4ns_16_7_1_U1.top_mul_16s_4ns_16_7_1_Mul_DSP_0_U.buff0 ;
assign _162_ = \mul_16s_4ns_16_7_1_U1.top_mul_16s_4ns_16_7_1_Mul_DSP_0_U.ce  ? \mul_16s_4ns_16_7_1_U1.top_mul_16s_4ns_16_7_1_Mul_DSP_0_U.b  : \mul_16s_4ns_16_7_1_U1.top_mul_16s_4ns_16_7_1_Mul_DSP_0_U.b_reg0 ;
assign _161_ = \mul_16s_4ns_16_7_1_U1.top_mul_16s_4ns_16_7_1_Mul_DSP_0_U.ce  ? \mul_16s_4ns_16_7_1_U1.top_mul_16s_4ns_16_7_1_Mul_DSP_0_U.a  : \mul_16s_4ns_16_7_1_U1.top_mul_16s_4ns_16_7_1_Mul_DSP_0_U.a_reg0 ;
assign \mul_6s_6s_6_7_1_U3.top_mul_6s_6s_6_7_1_Mul_DSP_1_U.tmp_product  = $signed(\mul_6s_6s_6_7_1_U3.top_mul_6s_6s_6_7_1_Mul_DSP_1_U.a_reg0 ) * $signed(\mul_6s_6s_6_7_1_U3.top_mul_6s_6s_6_7_1_Mul_DSP_1_U.b_reg0 );
always @(posedge \mul_6s_6s_6_7_1_U3.top_mul_6s_6s_6_7_1_Mul_DSP_1_U.clk )
\mul_6s_6s_6_7_1_U3.top_mul_6s_6s_6_7_1_Mul_DSP_1_U.a_reg0  <= _168_;
always @(posedge \mul_6s_6s_6_7_1_U3.top_mul_6s_6s_6_7_1_Mul_DSP_1_U.clk )
\mul_6s_6s_6_7_1_U3.top_mul_6s_6s_6_7_1_Mul_DSP_1_U.b_reg0  <= _169_;
always @(posedge \mul_6s_6s_6_7_1_U3.top_mul_6s_6s_6_7_1_Mul_DSP_1_U.clk )
\mul_6s_6s_6_7_1_U3.top_mul_6s_6s_6_7_1_Mul_DSP_1_U.buff0  <= _170_;
always @(posedge \mul_6s_6s_6_7_1_U3.top_mul_6s_6s_6_7_1_Mul_DSP_1_U.clk )
\mul_6s_6s_6_7_1_U3.top_mul_6s_6s_6_7_1_Mul_DSP_1_U.buff1  <= _171_;
always @(posedge \mul_6s_6s_6_7_1_U3.top_mul_6s_6s_6_7_1_Mul_DSP_1_U.clk )
\mul_6s_6s_6_7_1_U3.top_mul_6s_6s_6_7_1_Mul_DSP_1_U.buff2  <= _172_;
always @(posedge \mul_6s_6s_6_7_1_U3.top_mul_6s_6s_6_7_1_Mul_DSP_1_U.clk )
\mul_6s_6s_6_7_1_U3.top_mul_6s_6s_6_7_1_Mul_DSP_1_U.buff3  <= _173_;
always @(posedge \mul_6s_6s_6_7_1_U3.top_mul_6s_6s_6_7_1_Mul_DSP_1_U.clk )
\mul_6s_6s_6_7_1_U3.top_mul_6s_6s_6_7_1_Mul_DSP_1_U.buff4  <= _174_;
assign _174_ = \mul_6s_6s_6_7_1_U3.top_mul_6s_6s_6_7_1_Mul_DSP_1_U.ce  ? \mul_6s_6s_6_7_1_U3.top_mul_6s_6s_6_7_1_Mul_DSP_1_U.buff3  : \mul_6s_6s_6_7_1_U3.top_mul_6s_6s_6_7_1_Mul_DSP_1_U.buff4 ;
assign _173_ = \mul_6s_6s_6_7_1_U3.top_mul_6s_6s_6_7_1_Mul_DSP_1_U.ce  ? \mul_6s_6s_6_7_1_U3.top_mul_6s_6s_6_7_1_Mul_DSP_1_U.buff2  : \mul_6s_6s_6_7_1_U3.top_mul_6s_6s_6_7_1_Mul_DSP_1_U.buff3 ;
assign _172_ = \mul_6s_6s_6_7_1_U3.top_mul_6s_6s_6_7_1_Mul_DSP_1_U.ce  ? \mul_6s_6s_6_7_1_U3.top_mul_6s_6s_6_7_1_Mul_DSP_1_U.buff1  : \mul_6s_6s_6_7_1_U3.top_mul_6s_6s_6_7_1_Mul_DSP_1_U.buff2 ;
assign _171_ = \mul_6s_6s_6_7_1_U3.top_mul_6s_6s_6_7_1_Mul_DSP_1_U.ce  ? \mul_6s_6s_6_7_1_U3.top_mul_6s_6s_6_7_1_Mul_DSP_1_U.buff0  : \mul_6s_6s_6_7_1_U3.top_mul_6s_6s_6_7_1_Mul_DSP_1_U.buff1 ;
assign _170_ = \mul_6s_6s_6_7_1_U3.top_mul_6s_6s_6_7_1_Mul_DSP_1_U.ce  ? \mul_6s_6s_6_7_1_U3.top_mul_6s_6s_6_7_1_Mul_DSP_1_U.tmp_product  : \mul_6s_6s_6_7_1_U3.top_mul_6s_6s_6_7_1_Mul_DSP_1_U.buff0 ;
assign _169_ = \mul_6s_6s_6_7_1_U3.top_mul_6s_6s_6_7_1_Mul_DSP_1_U.ce  ? \mul_6s_6s_6_7_1_U3.top_mul_6s_6s_6_7_1_Mul_DSP_1_U.b  : \mul_6s_6s_6_7_1_U3.top_mul_6s_6s_6_7_1_Mul_DSP_1_U.b_reg0 ;
assign _168_ = \mul_6s_6s_6_7_1_U3.top_mul_6s_6s_6_7_1_Mul_DSP_1_U.ce  ? \mul_6s_6s_6_7_1_U3.top_mul_6s_6s_6_7_1_Mul_DSP_1_U.a  : \mul_6s_6s_6_7_1_U3.top_mul_6s_6s_6_7_1_Mul_DSP_1_U.a_reg0 ;
always @(posedge \shl_9ns_4ns_9_7_1_U6.clk )
\shl_9ns_4ns_9_7_1_U6.dout_array[5]  <= _186_;
always @(posedge \shl_9ns_4ns_9_7_1_U6.clk )
\shl_9ns_4ns_9_7_1_U6.din1_cast_array[5]  <= _180_;
always @(posedge \shl_9ns_4ns_9_7_1_U6.clk )
\shl_9ns_4ns_9_7_1_U6.dout_array[4]  <= _185_;
always @(posedge \shl_9ns_4ns_9_7_1_U6.clk )
\shl_9ns_4ns_9_7_1_U6.din1_cast_array[4]  <= _179_;
always @(posedge \shl_9ns_4ns_9_7_1_U6.clk )
\shl_9ns_4ns_9_7_1_U6.dout_array[3]  <= _184_;
always @(posedge \shl_9ns_4ns_9_7_1_U6.clk )
\shl_9ns_4ns_9_7_1_U6.din1_cast_array[3]  <= _178_;
always @(posedge \shl_9ns_4ns_9_7_1_U6.clk )
\shl_9ns_4ns_9_7_1_U6.dout_array[2]  <= _183_;
always @(posedge \shl_9ns_4ns_9_7_1_U6.clk )
\shl_9ns_4ns_9_7_1_U6.din1_cast_array[2]  <= _177_;
always @(posedge \shl_9ns_4ns_9_7_1_U6.clk )
\shl_9ns_4ns_9_7_1_U6.dout_array[1]  <= _182_;
always @(posedge \shl_9ns_4ns_9_7_1_U6.clk )
\shl_9ns_4ns_9_7_1_U6.din1_cast_array[1]  <= _176_;
always @(posedge \shl_9ns_4ns_9_7_1_U6.clk )
\shl_9ns_4ns_9_7_1_U6.dout_array[0]  <= _181_;
always @(posedge \shl_9ns_4ns_9_7_1_U6.clk )
\shl_9ns_4ns_9_7_1_U6.din1_cast_array[0]  <= _175_;
assign _187_ = \shl_9ns_4ns_9_7_1_U6.ce  ? \shl_9ns_4ns_9_7_1_U6.din1_cast_array[4]  : \shl_9ns_4ns_9_7_1_U6.din1_cast_array[5] ;
assign _180_ = \shl_9ns_4ns_9_7_1_U6.reset  ? 4'h0 : _187_;
assign _188_ = \shl_9ns_4ns_9_7_1_U6.ce  ? _201_ : \shl_9ns_4ns_9_7_1_U6.dout_array[5] ;
assign _186_ = \shl_9ns_4ns_9_7_1_U6.reset  ? 9'h000 : _188_;
assign _189_ = \shl_9ns_4ns_9_7_1_U6.ce  ? \shl_9ns_4ns_9_7_1_U6.din1_cast_array[3]  : \shl_9ns_4ns_9_7_1_U6.din1_cast_array[4] ;
assign _179_ = \shl_9ns_4ns_9_7_1_U6.reset  ? 4'h0 : _189_;
assign _190_ = \shl_9ns_4ns_9_7_1_U6.ce  ? _200_ : \shl_9ns_4ns_9_7_1_U6.dout_array[4] ;
assign _185_ = \shl_9ns_4ns_9_7_1_U6.reset  ? 9'h000 : _190_;
assign _191_ = \shl_9ns_4ns_9_7_1_U6.ce  ? \shl_9ns_4ns_9_7_1_U6.din1_cast_array[2]  : \shl_9ns_4ns_9_7_1_U6.din1_cast_array[3] ;
assign _178_ = \shl_9ns_4ns_9_7_1_U6.reset  ? 4'h0 : _191_;
assign _192_ = \shl_9ns_4ns_9_7_1_U6.ce  ? _199_ : \shl_9ns_4ns_9_7_1_U6.dout_array[3] ;
assign _184_ = \shl_9ns_4ns_9_7_1_U6.reset  ? 9'h000 : _192_;
assign _193_ = \shl_9ns_4ns_9_7_1_U6.ce  ? \shl_9ns_4ns_9_7_1_U6.din1_cast_array[1]  : \shl_9ns_4ns_9_7_1_U6.din1_cast_array[2] ;
assign _177_ = \shl_9ns_4ns_9_7_1_U6.reset  ? 4'h0 : _193_;
assign _194_ = \shl_9ns_4ns_9_7_1_U6.ce  ? \shl_9ns_4ns_9_7_1_U6.dout_array[1]  : \shl_9ns_4ns_9_7_1_U6.dout_array[2] ;
assign _183_ = \shl_9ns_4ns_9_7_1_U6.reset  ? 9'h000 : _194_;
assign _195_ = \shl_9ns_4ns_9_7_1_U6.ce  ? \shl_9ns_4ns_9_7_1_U6.din1_cast_array[0]  : \shl_9ns_4ns_9_7_1_U6.din1_cast_array[1] ;
assign _176_ = \shl_9ns_4ns_9_7_1_U6.reset  ? 4'h0 : _195_;
assign _196_ = \shl_9ns_4ns_9_7_1_U6.ce  ? \shl_9ns_4ns_9_7_1_U6.dout_array[0]  : \shl_9ns_4ns_9_7_1_U6.dout_array[1] ;
assign _182_ = \shl_9ns_4ns_9_7_1_U6.reset  ? 9'h000 : _196_;
assign _197_ = \shl_9ns_4ns_9_7_1_U6.ce  ? \shl_9ns_4ns_9_7_1_U6.din1 [3:0] : \shl_9ns_4ns_9_7_1_U6.din1_cast_array[0] ;
assign _175_ = \shl_9ns_4ns_9_7_1_U6.reset  ? 4'h0 : _197_;
assign _198_ = \shl_9ns_4ns_9_7_1_U6.ce  ? \shl_9ns_4ns_9_7_1_U6.din0  : \shl_9ns_4ns_9_7_1_U6.dout_array[0] ;
assign _181_ = \shl_9ns_4ns_9_7_1_U6.reset  ? 9'h000 : _198_;
assign _199_ = \shl_9ns_4ns_9_7_1_U6.dout_array[2]  << { \shl_9ns_4ns_9_7_1_U6.din1_cast_array[2] [3], 3'h0 };
assign _200_ = \shl_9ns_4ns_9_7_1_U6.dout_array[3]  << { \shl_9ns_4ns_9_7_1_U6.din1_cast_array[3] [2], 2'h0 };
assign _201_ = \shl_9ns_4ns_9_7_1_U6.dout_array[4]  << { \shl_9ns_4ns_9_7_1_U6.din1_cast_array[4] [1], 1'h0 };
assign \shl_9ns_4ns_9_7_1_U6.dout  = \shl_9ns_4ns_9_7_1_U6.dout_array[5]  << \shl_9ns_4ns_9_7_1_U6.din1_cast_array[5] [0];
assign \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.bin_s0  = ~ \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.b ;
always @(posedge \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.clk )
\sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.bin_s1  <= _203_;
always @(posedge \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.clk )
\sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.ain_s1  <= _202_;
always @(posedge \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.clk )
\sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.sum_s1  <= _205_;
always @(posedge \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.clk )
\sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.carry_s1  <= _204_;
assign _203_ = \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.ce  ? \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.bin_s0 [16:8] : \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.bin_s1 ;
assign _202_ = \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.ce  ? \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.a [16:8] : \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.ain_s1 ;
assign _204_ = \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.ce  ? \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.facout_s1  : \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.carry_s1 ;
assign _205_ = \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.ce  ? \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.fas_s1  : \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.sum_s1 ;
assign _206_ = \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.u1.a  + \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.u1.b ;
assign { \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.u1.cout , \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.u1.s  } = _206_ + \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.u1.cin ;
assign _207_ = \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.u2.a  + \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.u2.b ;
assign { \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.u2.cout , \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.u2.s  } = _207_ + \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.u2.cin ;
assign \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.bin_s0  = ~ \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.b ;
always @(posedge \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.clk )
\sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.bin_s1  <= _209_;
always @(posedge \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.clk )
\sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.ain_s1  <= _208_;
always @(posedge \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.clk )
\sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.sum_s1  <= _211_;
always @(posedge \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.clk )
\sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.carry_s1  <= _210_;
assign _209_ = \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.ce  ? \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.bin_s0 [3:2] : \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.bin_s1 ;
assign _208_ = \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.ce  ? \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.a [3:2] : \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.ain_s1 ;
assign _210_ = \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.ce  ? \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.facout_s1  : \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.carry_s1 ;
assign _211_ = \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.ce  ? \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.fas_s1  : \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.sum_s1 ;
assign _212_ = \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.u1.a  + \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.u1.b ;
assign { \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.u1.cout , \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.u1.s  } = _212_ + \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.u1.cin ;
assign _213_ = \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.u2.a  + \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.u2.b ;
assign { \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.u2.cout , \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.u2.s  } = _213_ + \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.u2.cin ;
assign ret_V_18_fu_450_p2 = { mul_ln731_reg_819[5], mul_ln731_reg_819[5], mul_ln731_reg_819, 2'h0 } | { op_0, 2'h0 };
always @(posedge ap_clk)
trunc_ln851_1_reg_851 <= 2'h0;
always @(posedge ap_clk)
shl_ln1299_reg_866 <= _036_;
always @(posedge ap_clk)
sext_ln850_reg_973 <= _035_;
always @(posedge ap_clk)
ret_V_9_reg_893 <= _032_;
always @(posedge ap_clk)
ret_V_25_reg_985 <= _027_;
always @(posedge ap_clk)
ret_V_24_reg_963 <= _026_;
always @(posedge ap_clk)
tmp_3_reg_968 <= _038_;
always @(posedge ap_clk)
ush_reg_741 <= _042_;
always @(posedge ap_clk)
ret_V_2_reg_746 <= _028_;
always @(posedge ap_clk)
ret_V_22_reg_751 <= _024_;
always @(posedge ap_clk)
ret_V_21_cast_reg_756 <= _022_;
always @(posedge ap_clk)
trunc_ln851_3_reg_763 <= _040_;
always @(posedge ap_clk)
ret_V_19_reg_903 <= _020_;
always @(posedge ap_clk)
ret_V_21_reg_908 <= _023_;
always @(posedge ap_clk)
_561_ <= _019_;
assign ret_V_18_reg_839[9:2] = _561_;
always @(posedge ap_clk)
ret_V_4_cast_reg_844 <= _029_;
always @(posedge ap_clk)
ret_V_20_reg_856 <= _021_;
always @(posedge ap_clk)
ret_V_8_reg_861 <= _031_;
always @(posedge ap_clk)
ret_V_12_reg_789 <= _017_;
always @(posedge ap_clk)
ret_V_5_reg_888 <= _030_;
always @(posedge ap_clk)
op_25_V_reg_898 <= _015_;
always @(posedge ap_clk)
op_23_V_reg_943 <= _014_;
always @(posedge ap_clk)
mul_ln728_reg_814 <= _012_;
always @(posedge ap_clk)
trunc_ln1118_reg_682 <= _039_;
always @(posedge ap_clk)
isNeg_reg_693 <= _011_;
always @(posedge ap_clk)
ret_V_reg_699 <= _033_;
always @(posedge ap_clk)
trunc_ln851_reg_706 <= _041_;
always @(posedge ap_clk)
sub_ln1367_reg_721 <= _037_;
always @(posedge ap_clk)
icmp_ln851_reg_726 <= _010_;
always @(posedge ap_clk)
r_reg_774 <= _016_;
always @(posedge ap_clk)
ret_V_17_reg_779 <= _018_;
always @(posedge ap_clk)
icmp_ln851_3_reg_784 <= _009_;
always @(posedge ap_clk)
mul_ln731_reg_819 <= _013_;
always @(posedge ap_clk)
icmp_ln851_2_reg_834 <= _008_;
always @(posedge ap_clk)
icmp_ln851_1_reg_876 <= _007_;
always @(posedge ap_clk)
sext_ln835_reg_881 <= _034_;
always @(posedge ap_clk)
ashr_ln1333_reg_871 <= _006_;
always @(posedge ap_clk)
ret_V_23_reg_804 <= _025_;
always @(posedge ap_clk)
add_ln69_4_reg_809 <= _003_;
always @(posedge ap_clk)
add_ln69_3_reg_995 <= _002_;
always @(posedge ap_clk)
add_ln69_reg_928 <= _004_;
always @(posedge ap_clk)
add_ln69_1_reg_933 <= _001_;
always @(posedge ap_clk)
add_ln691_reg_980 <= _000_;
always @(posedge ap_clk)
ap_CS_fsm <= _005_;
assign _043_ = _048_ ? 2'h2 : 2'h1;
assign _214_ = ap_CS_fsm == 1'h1;
function [24:0] _593_;
input [24:0] a;
input [624:0] b;
input [24:0] s;
case (s)
25'b0000000000000000000000001:
_593_ = b[24:0];
25'b0000000000000000000000010:
_593_ = b[49:25];
25'b0000000000000000000000100:
_593_ = b[74:50];
25'b0000000000000000000001000:
_593_ = b[99:75];
25'b0000000000000000000010000:
_593_ = b[124:100];
25'b0000000000000000000100000:
_593_ = b[149:125];
25'b0000000000000000001000000:
_593_ = b[174:150];
25'b0000000000000000010000000:
_593_ = b[199:175];
25'b0000000000000000100000000:
_593_ = b[224:200];
25'b0000000000000001000000000:
_593_ = b[249:225];
25'b0000000000000010000000000:
_593_ = b[274:250];
25'b0000000000000100000000000:
_593_ = b[299:275];
25'b0000000000001000000000000:
_593_ = b[324:300];
25'b0000000000010000000000000:
_593_ = b[349:325];
25'b0000000000100000000000000:
_593_ = b[374:350];
25'b0000000001000000000000000:
_593_ = b[399:375];
25'b0000000010000000000000000:
_593_ = b[424:400];
25'b0000000100000000000000000:
_593_ = b[449:425];
25'b0000001000000000000000000:
_593_ = b[474:450];
25'b0000010000000000000000000:
_593_ = b[499:475];
25'b0000100000000000000000000:
_593_ = b[524:500];
25'b0001000000000000000000000:
_593_ = b[549:525];
25'b0010000000000000000000000:
_593_ = b[574:550];
25'b0100000000000000000000000:
_593_ = b[599:575];
25'b1000000000000000000000000:
_593_ = b[624:600];
25'b0000000000000000000000000:
_593_ = a;
default:
_593_ = 25'bx;
endcase
endfunction
assign ap_NS_fsm = _593_(25'hxxxxxxx, { 23'h000000, _043_, 600'h000002000002000002000002000002000002000002000002000002000002000002000002000002000002000002000002000002000002000002000002000002000002000002000000000001 }, { _214_, _238_, _237_, _236_, _235_, _234_, _233_, _232_, _231_, _230_, _229_, _228_, _227_, _226_, _225_, _224_, _223_, _222_, _221_, _220_, _219_, _218_, _217_, _216_, _215_ });
assign _215_ = ap_CS_fsm == 25'h1000000;
assign _216_ = ap_CS_fsm == 24'h800000;
assign _217_ = ap_CS_fsm == 23'h400000;
assign _218_ = ap_CS_fsm == 22'h200000;
assign _219_ = ap_CS_fsm == 21'h100000;
assign _220_ = ap_CS_fsm == 20'h80000;
assign _221_ = ap_CS_fsm == 19'h40000;
assign _222_ = ap_CS_fsm == 18'h20000;
assign _223_ = ap_CS_fsm == 17'h10000;
assign _224_ = ap_CS_fsm == 16'h8000;
assign _225_ = ap_CS_fsm == 15'h4000;
assign _226_ = ap_CS_fsm == 14'h2000;
assign _227_ = ap_CS_fsm == 13'h1000;
assign _228_ = ap_CS_fsm == 12'h800;
assign _229_ = ap_CS_fsm == 11'h400;
assign _230_ = ap_CS_fsm == 10'h200;
assign _231_ = ap_CS_fsm == 9'h100;
assign _232_ = ap_CS_fsm == 8'h80;
assign _233_ = ap_CS_fsm == 7'h40;
assign _234_ = ap_CS_fsm == 6'h20;
assign _235_ = ap_CS_fsm == 5'h10;
assign _236_ = ap_CS_fsm == 4'h8;
assign _237_ = ap_CS_fsm == 3'h4;
assign _238_ = ap_CS_fsm == 2'h2;
assign op_28_ap_vld = ap_CS_fsm[24] ? 1'h1 : 1'h0;
assign ap_idle = _047_ ? 1'h1 : 1'h0;
assign _036_ = _046_ ? grp_fu_325_p2 : shl_ln1299_reg_866;
assign _035_ = ap_CS_fsm[18] ? { tmp_3_reg_968[18], tmp_3_reg_968 } : sext_ln850_reg_973;
assign _032_ = _045_ ? grp_fu_493_p2 : ret_V_9_reg_893;
assign _027_ = ap_CS_fsm[20] ? ret_V_25_fu_641_p3 : ret_V_25_reg_985;
assign _038_ = ap_CS_fsm[17] ? grp_fu_600_p2[19:1] : tmp_3_reg_968;
assign _026_ = ap_CS_fsm[17] ? grp_fu_600_p2 : ret_V_24_reg_963;
assign _040_ = ap_CS_fsm[2] ? grp_fu_297_p2[7:0] : trunc_ln851_3_reg_763;
assign _022_ = ap_CS_fsm[2] ? grp_fu_297_p2[9:8] : ret_V_21_cast_reg_756;
assign _024_ = ap_CS_fsm[2] ? grp_fu_297_p2 : ret_V_22_reg_751;
assign _028_ = ap_CS_fsm[2] ? grp_fu_276_p2 : ret_V_2_reg_746;
assign _042_ = ap_CS_fsm[2] ? ush_fu_303_p3 : ush_reg_741;
assign _023_ = ap_CS_fsm[11] ? ret_V_21_fu_549_p3 : ret_V_21_reg_908;
assign _020_ = ap_CS_fsm[11] ? ret_V_19_fu_530_p3 : ret_V_19_reg_903;
assign _031_ = ap_CS_fsm[8] ? grp_fu_415_p2[19:3] : ret_V_8_reg_861;
assign _021_ = ap_CS_fsm[8] ? grp_fu_415_p2 : ret_V_20_reg_856;
assign _029_ = ap_CS_fsm[8] ? ret_V_18_fu_450_p2[3:2] : ret_V_4_cast_reg_844;
assign _019_ = ap_CS_fsm[8] ? ret_V_18_fu_450_p2[9:2] : ret_V_18_reg_839[9:2];
assign _017_ = ap_CS_fsm[4] ? grp_fu_364_p2 : ret_V_12_reg_789;
assign _015_ = ap_CS_fsm[10] ? op_25_V_fu_512_p2 : op_25_V_reg_898;
assign _030_ = ap_CS_fsm[10] ? grp_fu_485_p2 : ret_V_5_reg_888;
assign _014_ = ap_CS_fsm[15] ? grp_fu_580_p2 : op_23_V_reg_943;
assign _012_ = ap_CS_fsm[6] ? grp_fu_201_p2 : mul_ln728_reg_814;
assign _041_ = ap_CS_fsm[0] ? 25'h0000000 : trunc_ln851_reg_706;
assign _033_ = ap_CS_fsm[0] ? { op_8[15:1], ret_V_16_fu_229_p2[25] } : ret_V_reg_699;
assign _011_ = ap_CS_fsm[0] ? op_9[3] : isNeg_reg_693;
assign _039_ = ap_CS_fsm[0] ? op_8[8:0] : trunc_ln1118_reg_682;
assign _010_ = ap_CS_fsm[1] ? icmp_ln851_fu_271_p2 : icmp_ln851_reg_726;
assign _037_ = ap_CS_fsm[1] ? grp_fu_215_p2 : sub_ln1367_reg_721;
assign _009_ = ap_CS_fsm[3] ? icmp_ln851_3_fu_359_p2 : icmp_ln851_3_reg_784;
assign _018_ = ap_CS_fsm[3] ? ret_V_17_fu_352_p3 : ret_V_17_reg_779;
assign _016_ = ap_CS_fsm[3] ? r_fu_335_p2 : r_reg_774;
assign _008_ = ap_CS_fsm[7] ? icmp_ln851_2_fu_425_p2 : icmp_ln851_2_reg_834;
assign _013_ = ap_CS_fsm[7] ? grp_fu_257_p2 : mul_ln731_reg_819;
assign _034_ = ap_CS_fsm[9] ? { ret_V_8_reg_861[16], ret_V_8_reg_861 } : sext_ln835_reg_881;
assign _007_ = ap_CS_fsm[9] ? icmp_ln851_1_fu_480_p2 : icmp_ln851_1_reg_876;
assign _006_ = _044_ ? grp_fu_330_p2 : ashr_ln1333_reg_871;
assign _003_ = ap_CS_fsm[5] ? grp_fu_375_p2 : add_ln69_4_reg_809;
assign _025_ = ap_CS_fsm[5] ? ret_V_23_fu_393_p3 : ret_V_23_reg_804;
assign _002_ = ap_CS_fsm[22] ? grp_fu_651_p2 : add_ln69_3_reg_995;
assign _001_ = ap_CS_fsm[13] ? grp_fu_571_p2 : add_ln69_1_reg_933;
assign _004_ = ap_CS_fsm[13] ? grp_fu_566_p2 : add_ln69_reg_928;
assign _000_ = ap_CS_fsm[19] ? grp_fu_619_p2 : add_ln691_reg_980;
assign _005_ = ap_rst ? 25'h0000001 : ap_NS_fsm;
assign icmp_ln851_1_fu_480_p2 = _052_ ? 1'h1 : 1'h0;
assign icmp_ln851_2_fu_425_p2 = _053_ ? 1'h1 : 1'h0;
assign icmp_ln851_3_fu_359_p2 = _054_ ? 1'h1 : 1'h0;
assign icmp_ln851_fu_271_p2 = _055_ ? 1'h1 : 1'h0;
assign op_16_V_fu_505_p3 = isNeg_reg_693 ? shl_ln1299_reg_866[0] : ashr_ln1333_reg_871[0];
assign ret_V_17_fu_352_p3 = op_8[15] ? select_ln850_fu_347_p3 : ret_V_reg_699;
assign ret_V_19_fu_530_p3 = ret_V_18_reg_839[9] ? select_ln850_1_fu_525_p3 : ret_V_4_cast_reg_844;
assign ret_V_21_fu_549_p3 = ret_V_20_reg_856[19] ? select_ln850_2_fu_544_p3 : sext_ln835_reg_881;
assign ret_V_23_fu_393_p3 = ret_V_22_reg_751[16] ? select_ln850_3_fu_388_p3 : ret_V_21_cast_reg_756;
assign ret_V_25_fu_641_p3 = ret_V_24_reg_963[19] ? select_ln850_4_fu_635_p3 : sext_ln850_reg_973;
assign select_ln850_1_fu_525_p3 = icmp_ln851_1_reg_876 ? ret_V_4_cast_reg_844 : ret_V_5_reg_888;
assign select_ln850_2_fu_544_p3 = icmp_ln851_2_reg_834 ? sext_ln835_reg_881 : ret_V_9_reg_893;
assign select_ln850_3_fu_388_p3 = icmp_ln851_3_reg_784 ? ret_V_21_cast_reg_756 : ret_V_12_reg_789;
assign select_ln850_4_fu_635_p3 = op_15[0] ? add_ln691_reg_980 : sext_ln850_reg_973;
assign select_ln850_fu_347_p3 = icmp_ln851_reg_726 ? ret_V_reg_699 : ret_V_2_reg_746;
assign ush_fu_303_p3 = isNeg_reg_693 ? sub_ln1367_reg_721 : op_9;
assign ap_CS_fsm_state1 = ap_CS_fsm[0];
assign ap_CS_fsm_state10 = ap_CS_fsm[9];
assign ap_CS_fsm_state11 = ap_CS_fsm[10];
assign ap_CS_fsm_state12 = ap_CS_fsm[11];
assign ap_CS_fsm_state13 = ap_CS_fsm[12];
assign ap_CS_fsm_state14 = ap_CS_fsm[13];
assign ap_CS_fsm_state15 = ap_CS_fsm[14];
assign ap_CS_fsm_state16 = ap_CS_fsm[15];
assign ap_CS_fsm_state17 = ap_CS_fsm[16];
assign ap_CS_fsm_state18 = ap_CS_fsm[17];
assign ap_CS_fsm_state19 = ap_CS_fsm[18];
assign ap_CS_fsm_state2 = ap_CS_fsm[1];
assign ap_CS_fsm_state20 = ap_CS_fsm[19];
assign ap_CS_fsm_state21 = ap_CS_fsm[20];
assign ap_CS_fsm_state22 = ap_CS_fsm[21];
assign ap_CS_fsm_state23 = ap_CS_fsm[22];
assign ap_CS_fsm_state24 = ap_CS_fsm[23];
assign ap_CS_fsm_state25 = ap_CS_fsm[24];
assign ap_CS_fsm_state3 = ap_CS_fsm[2];
assign ap_CS_fsm_state4 = ap_CS_fsm[3];
assign ap_CS_fsm_state5 = ap_CS_fsm[4];
assign ap_CS_fsm_state6 = ap_CS_fsm[5];
assign ap_CS_fsm_state7 = ap_CS_fsm[6];
assign ap_CS_fsm_state8 = ap_CS_fsm[7];
assign ap_CS_fsm_state9 = ap_CS_fsm[8];
assign ap_done = op_28_ap_vld;
assign ap_ready = op_28_ap_vld;
assign grp_fu_201_p1 = op_5;
assign grp_fu_201_p10 = { 12'h000, op_5 };
assign grp_fu_257_p0 = op_1[5:0];
assign grp_fu_257_p1 = op_2[5:0];
assign grp_fu_297_p0 = { 1'h0, op_2, 8'h00 };
assign grp_fu_297_p1 = { 7'h00, op_10, 8'h00 };
assign grp_fu_375_p0 = { ret_V_17_reg_779[15], ret_V_17_reg_779 };
assign grp_fu_375_p1 = { r_reg_774[3], r_reg_774[3], r_reg_774[3], r_reg_774[3], r_reg_774[3], r_reg_774[3], r_reg_774[3], r_reg_774[3], r_reg_774[3], r_reg_774[3], r_reg_774[3], r_reg_774[3], r_reg_774[3], r_reg_774 };
assign grp_fu_415_p0 = { 1'h0, mul_ln728_reg_814, 3'h0 };
assign grp_fu_415_p1 = { op_7[3], op_7[3], op_7[3], op_7[3], op_7[3], op_7[3], op_7[3], op_7[3], op_7[3], op_7[3], op_7[3], op_7[3], op_7[3], op_7[3], op_7[3], op_7[3], op_7 };
assign grp_fu_493_p0 = { ret_V_8_reg_861[16], ret_V_8_reg_861 };
assign grp_fu_566_p1 = { 16'h0000, ret_V_19_reg_903 };
assign grp_fu_571_p0 = { op_13[1], op_13[1], op_13 };
assign grp_fu_571_p1 = { 2'h0, ret_V_23_reg_804 };
assign grp_fu_580_p0 = { add_ln69_1_reg_933[3], add_ln69_1_reg_933[3], add_ln69_1_reg_933[3], add_ln69_1_reg_933[3], add_ln69_1_reg_933[3], add_ln69_1_reg_933[3], add_ln69_1_reg_933[3], add_ln69_1_reg_933[3], add_ln69_1_reg_933[3], add_ln69_1_reg_933[3], add_ln69_1_reg_933[3], add_ln69_1_reg_933[3], add_ln69_1_reg_933[3], add_ln69_1_reg_933[3], add_ln69_1_reg_933 };
assign grp_fu_600_p0 = { op_23_V_reg_943[17], op_23_V_reg_943, 1'h0 };
assign grp_fu_600_p1 = { op_15[1], op_15[1], op_15[1], op_15[1], op_15[1], op_15[1], op_15[1], op_15[1], op_15[1], op_15[1], op_15[1], op_15[1], op_15[1], op_15[1], op_15[1], op_15[1], op_15[1], op_15[1], op_15 };
assign grp_fu_619_p0 = { tmp_3_reg_968[18], tmp_3_reg_968 };
assign grp_fu_651_p0 = { 19'h00000, op_25_V_reg_898 };
assign grp_fu_659_p0 = { add_ln69_4_reg_809[16], add_ln69_4_reg_809[16], add_ln69_4_reg_809[16], add_ln69_4_reg_809 };
assign lhs_V_fu_438_p3 = { op_0, 2'h0 };
assign op_28 = { grp_fu_659_p2[19], grp_fu_659_p2[19], grp_fu_659_p2[19], grp_fu_659_p2[19], grp_fu_659_p2[19], grp_fu_659_p2[19], grp_fu_659_p2[19], grp_fu_659_p2[19], grp_fu_659_p2[19], grp_fu_659_p2[19], grp_fu_659_p2[19], grp_fu_659_p2[19], grp_fu_659_p2 };
assign op_4_V_fu_431_p3 = { mul_ln731_reg_819, 2'h0 };
assign op_6_V_fu_263_p3 = { op_2, 8'h00 };
assign p_Result_1_fu_518_p3 = ret_V_18_reg_839[9];
assign p_Result_2_fu_537_p3 = ret_V_20_reg_856[19];
assign p_Result_3_fu_381_p3 = ret_V_22_reg_751[16];
assign p_Result_4_fu_625_p3 = ret_V_24_reg_963[19];
assign p_Result_s_fu_340_p1 = op_8;
assign p_Result_s_fu_340_p3 = op_8[15];
assign ret_V_16_fu_229_p2[24:0] = 25'h0000000;
assign ret_V_16_fu_229_p2[40:26] = op_8[15:1];
assign rhs_2_fu_404_p3 = { mul_ln728_reg_814, 3'h0 };
assign rhs_3_fu_285_p3 = { op_10, 8'h00 };
assign rhs_fu_221_p1 = op_8;
assign rhs_fu_221_p3 = { op_8, 25'h0000000 };
assign sext_ln1192_1_fu_585_p0 = op_15;
assign sext_ln1192_fu_400_p0 = op_7;
assign sext_ln703_fu_446_p1 = { mul_ln731_reg_819[5], mul_ln731_reg_819[5], mul_ln731_reg_819, 2'h0 };
assign sext_ln835_fu_490_p1 = { ret_V_8_reg_861[16], ret_V_8_reg_861 };
assign sext_ln850_fu_616_p1 = { tmp_3_reg_968[18], tmp_3_reg_968 };
assign tmp_fu_589_p3 = { op_23_V_reg_943, 1'h0 };
assign trunc_ln1118_fu_193_p0 = op_8;
assign trunc_ln1118_fu_193_p1 = op_8[8:0];
assign trunc_ln1368_1_fu_502_p1 = ashr_ln1333_reg_871[0];
assign trunc_ln1368_fu_499_p1 = shl_ln1299_reg_866[0];
assign trunc_ln851_1_fu_466_p1 = ret_V_18_fu_450_p2[1:0];
assign trunc_ln851_2_fu_421_p0 = op_7;
assign trunc_ln851_2_fu_421_p1 = op_7[2:0];
assign trunc_ln851_3_fu_318_p1 = grp_fu_297_p2[7:0];
assign trunc_ln851_4_fu_632_p0 = op_15;
assign trunc_ln851_4_fu_632_p1 = op_15[0];
assign trunc_ln851_fu_245_p1 = 25'h0000000;
assign zext_ln1367_fu_322_p1 = { 5'h00, ush_reg_741 };
assign \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.ain_s0  = \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.a ;
assign \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.s  = { \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.fas_s2 , \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.sum_s1  };
assign \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.u2.a  = \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.ain_s1 ;
assign \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.u2.b  = \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.bin_s1 ;
assign \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.u2.cin  = \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.carry_s1 ;
assign \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.facout_s2  = \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.u2.cout ;
assign \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.fas_s2  = \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.u2.s ;
assign \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.u1.a  = \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.a [1:0];
assign \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.u1.b  = \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.bin_s0 [1:0];
assign \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.u1.cin  = 1'h1;
assign \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.facout_s1  = \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.u1.cout ;
assign \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.fas_s1  = \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.u1.s ;
assign \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.a  = \sub_4ns_4ns_4_2_1_U2.din0 ;
assign \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.b  = \sub_4ns_4ns_4_2_1_U2.din1 ;
assign \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.ce  = \sub_4ns_4ns_4_2_1_U2.ce ;
assign \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.clk  = \sub_4ns_4ns_4_2_1_U2.clk ;
assign \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.reset  = \sub_4ns_4ns_4_2_1_U2.reset ;
assign \sub_4ns_4ns_4_2_1_U2.dout  = \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.s ;
assign \sub_4ns_4ns_4_2_1_U2.ce  = 1'h1;
assign \sub_4ns_4ns_4_2_1_U2.clk  = ap_clk;
assign \sub_4ns_4ns_4_2_1_U2.din0  = 4'h0;
assign \sub_4ns_4ns_4_2_1_U2.din1  = op_9;
assign grp_fu_215_p2 = \sub_4ns_4ns_4_2_1_U2.dout ;
assign \sub_4ns_4ns_4_2_1_U2.reset  = ap_rst;
assign \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.ain_s0  = \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.a ;
assign \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.s  = { \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.fas_s2 , \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.sum_s1  };
assign \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.u2.a  = \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.ain_s1 ;
assign \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.u2.b  = \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.bin_s1 ;
assign \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.u2.cin  = \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.carry_s1 ;
assign \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.facout_s2  = \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.u2.cout ;
assign \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.fas_s2  = \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.u2.s ;
assign \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.u1.a  = \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.a [7:0];
assign \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.u1.b  = \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.bin_s0 [7:0];
assign \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.u1.cin  = 1'h1;
assign \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.facout_s1  = \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.u1.cout ;
assign \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.fas_s1  = \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.u1.s ;
assign \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.a  = \sub_17ns_17ns_17_2_1_U5.din0 ;
assign \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.b  = \sub_17ns_17ns_17_2_1_U5.din1 ;
assign \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.ce  = \sub_17ns_17ns_17_2_1_U5.ce ;
assign \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.clk  = \sub_17ns_17ns_17_2_1_U5.clk ;
assign \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.reset  = \sub_17ns_17ns_17_2_1_U5.reset ;
assign \sub_17ns_17ns_17_2_1_U5.dout  = \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.s ;
assign \sub_17ns_17ns_17_2_1_U5.ce  = 1'h1;
assign \sub_17ns_17ns_17_2_1_U5.clk  = ap_clk;
assign \sub_17ns_17ns_17_2_1_U5.din0  = { 1'h0, op_2, 8'h00 };
assign \sub_17ns_17ns_17_2_1_U5.din1  = { 7'h00, op_10, 8'h00 };
assign grp_fu_297_p2 = \sub_17ns_17ns_17_2_1_U5.dout ;
assign \sub_17ns_17ns_17_2_1_U5.reset  = ap_rst;
assign \shl_9ns_4ns_9_7_1_U6.din1_cast  = \shl_9ns_4ns_9_7_1_U6.din1 [3:0];
assign \shl_9ns_4ns_9_7_1_U6.din1_mask  = 4'h1;
assign \shl_9ns_4ns_9_7_1_U6.ce  = 1'h1;
assign \shl_9ns_4ns_9_7_1_U6.clk  = ap_clk;
assign \shl_9ns_4ns_9_7_1_U6.din0  = trunc_ln1118_reg_682;
assign \shl_9ns_4ns_9_7_1_U6.din1  = { 5'h00, ush_reg_741 };
assign grp_fu_325_p2 = \shl_9ns_4ns_9_7_1_U6.dout ;
assign \shl_9ns_4ns_9_7_1_U6.reset  = ap_rst;
assign \mul_6s_6s_6_7_1_U3.top_mul_6s_6s_6_7_1_Mul_DSP_1_U.p  = \mul_6s_6s_6_7_1_U3.top_mul_6s_6s_6_7_1_Mul_DSP_1_U.buff4 ;
assign \mul_6s_6s_6_7_1_U3.top_mul_6s_6s_6_7_1_Mul_DSP_1_U.a  = \mul_6s_6s_6_7_1_U3.din0 ;
assign \mul_6s_6s_6_7_1_U3.top_mul_6s_6s_6_7_1_Mul_DSP_1_U.b  = \mul_6s_6s_6_7_1_U3.din1 ;
assign \mul_6s_6s_6_7_1_U3.top_mul_6s_6s_6_7_1_Mul_DSP_1_U.ce  = \mul_6s_6s_6_7_1_U3.ce ;
assign \mul_6s_6s_6_7_1_U3.top_mul_6s_6s_6_7_1_Mul_DSP_1_U.clk  = \mul_6s_6s_6_7_1_U3.clk ;
assign \mul_6s_6s_6_7_1_U3.dout  = \mul_6s_6s_6_7_1_U3.top_mul_6s_6s_6_7_1_Mul_DSP_1_U.p ;
assign \mul_6s_6s_6_7_1_U3.ce  = 1'h1;
assign \mul_6s_6s_6_7_1_U3.clk  = ap_clk;
assign \mul_6s_6s_6_7_1_U3.din0  = op_1[5:0];
assign \mul_6s_6s_6_7_1_U3.din1  = op_2[5:0];
assign grp_fu_257_p2 = \mul_6s_6s_6_7_1_U3.dout ;
assign \mul_6s_6s_6_7_1_U3.reset  = ap_rst;
assign \mul_16s_4ns_16_7_1_U1.top_mul_16s_4ns_16_7_1_Mul_DSP_0_U.p  = \mul_16s_4ns_16_7_1_U1.top_mul_16s_4ns_16_7_1_Mul_DSP_0_U.buff4 ;
assign \mul_16s_4ns_16_7_1_U1.top_mul_16s_4ns_16_7_1_Mul_DSP_0_U.a  = \mul_16s_4ns_16_7_1_U1.din0 ;
assign \mul_16s_4ns_16_7_1_U1.top_mul_16s_4ns_16_7_1_Mul_DSP_0_U.b  = \mul_16s_4ns_16_7_1_U1.din1 ;
assign \mul_16s_4ns_16_7_1_U1.top_mul_16s_4ns_16_7_1_Mul_DSP_0_U.ce  = \mul_16s_4ns_16_7_1_U1.ce ;
assign \mul_16s_4ns_16_7_1_U1.top_mul_16s_4ns_16_7_1_Mul_DSP_0_U.clk  = \mul_16s_4ns_16_7_1_U1.clk ;
assign \mul_16s_4ns_16_7_1_U1.dout  = \mul_16s_4ns_16_7_1_U1.top_mul_16s_4ns_16_7_1_Mul_DSP_0_U.p ;
assign \mul_16s_4ns_16_7_1_U1.ce  = 1'h1;
assign \mul_16s_4ns_16_7_1_U1.clk  = ap_clk;
assign \mul_16s_4ns_16_7_1_U1.din0  = op_8;
assign \mul_16s_4ns_16_7_1_U1.din1  = op_5;
assign grp_fu_201_p2 = \mul_16s_4ns_16_7_1_U1.dout ;
assign \mul_16s_4ns_16_7_1_U1.reset  = ap_rst;
assign \ashr_9ns_4ns_9_7_1_U7.din1_cast  = \ashr_9ns_4ns_9_7_1_U7.din1 [3:0];
assign \ashr_9ns_4ns_9_7_1_U7.din1_mask  = 4'h1;
assign \ashr_9ns_4ns_9_7_1_U7.ce  = 1'h1;
assign \ashr_9ns_4ns_9_7_1_U7.clk  = ap_clk;
assign \ashr_9ns_4ns_9_7_1_U7.din0  = trunc_ln1118_reg_682;
assign \ashr_9ns_4ns_9_7_1_U7.din1  = { 5'h00, ush_reg_741 };
assign grp_fu_330_p2 = \ashr_9ns_4ns_9_7_1_U7.dout ;
assign \ashr_9ns_4ns_9_7_1_U7.reset  = ap_rst;
assign \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.ain_s0  = \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.a ;
assign \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.bin_s0  = \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.b ;
assign \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.s  = { \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.fas_s2 , \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.sum_s1  };
assign \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.u2.a  = \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.ain_s1 ;
assign \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.u2.b  = \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.bin_s1 ;
assign \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.u2.cin  = \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.carry_s1 ;
assign \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.facout_s2  = \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.u2.cout ;
assign \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.fas_s2  = \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.u2.s ;
assign \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.u1.a  = \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.a [1:0];
assign \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.u1.b  = \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.b [1:0];
assign \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.u1.cin  = 1'h0;
assign \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.facout_s1  = \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.u1.cout ;
assign \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.fas_s1  = \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.u1.s ;
assign \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.a  = \add_4s_4ns_4_2_1_U14.din0 ;
assign \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.b  = \add_4s_4ns_4_2_1_U14.din1 ;
assign \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.ce  = \add_4s_4ns_4_2_1_U14.ce ;
assign \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.clk  = \add_4s_4ns_4_2_1_U14.clk ;
assign \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.reset  = \add_4s_4ns_4_2_1_U14.reset ;
assign \add_4s_4ns_4_2_1_U14.dout  = \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.s ;
assign \add_4s_4ns_4_2_1_U14.ce  = 1'h1;
assign \add_4s_4ns_4_2_1_U14.clk  = ap_clk;
assign \add_4s_4ns_4_2_1_U14.din0  = { op_13[1], op_13[1], op_13 };
assign \add_4s_4ns_4_2_1_U14.din1  = { 2'h0, ret_V_23_reg_804 };
assign grp_fu_571_p2 = \add_4s_4ns_4_2_1_U14.dout ;
assign \add_4s_4ns_4_2_1_U14.reset  = ap_rst;
assign \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.ain_s0  = \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.a ;
assign \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.bin_s0  = \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.b ;
assign \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.s  = { \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.fas_s2 , \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.sum_s1  };
assign \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.u2.a  = \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.ain_s1 ;
assign \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.u2.b  = \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.bin_s1 ;
assign \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.u2.cin  = \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.carry_s1 ;
assign \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.facout_s2  = \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.u2.cout ;
assign \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.fas_s2  = \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.u2.s ;
assign \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.u1.a  = \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.a [0];
assign \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.u1.b  = \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.b [0];
assign \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.u1.cin  = 1'h0;
assign \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.facout_s1  = \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.u1.cout ;
assign \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.fas_s1  = \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.u1.s ;
assign \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.a  = \add_2ns_2ns_2_2_1_U8.din0 ;
assign \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.b  = \add_2ns_2ns_2_2_1_U8.din1 ;
assign \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.ce  = \add_2ns_2ns_2_2_1_U8.ce ;
assign \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.clk  = \add_2ns_2ns_2_2_1_U8.clk ;
assign \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.reset  = \add_2ns_2ns_2_2_1_U8.reset ;
assign \add_2ns_2ns_2_2_1_U8.dout  = \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.s ;
assign \add_2ns_2ns_2_2_1_U8.ce  = 1'h1;
assign \add_2ns_2ns_2_2_1_U8.clk  = ap_clk;
assign \add_2ns_2ns_2_2_1_U8.din0  = ret_V_21_cast_reg_756;
assign \add_2ns_2ns_2_2_1_U8.din1  = 2'h1;
assign grp_fu_364_p2 = \add_2ns_2ns_2_2_1_U8.dout ;
assign \add_2ns_2ns_2_2_1_U8.reset  = ap_rst;
assign \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.ain_s0  = \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.a ;
assign \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.bin_s0  = \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.b ;
assign \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.s  = { \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.fas_s2 , \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.sum_s1  };
assign \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.u2.a  = \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.ain_s1 ;
assign \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.u2.b  = \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.bin_s1 ;
assign \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.u2.cin  = \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.carry_s1 ;
assign \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.facout_s2  = \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.u2.cout ;
assign \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.fas_s2  = \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.u2.s ;
assign \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.u1.a  = \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.a [0];
assign \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.u1.b  = \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.b [0];
assign \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.u1.cin  = 1'h0;
assign \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.facout_s1  = \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.u1.cout ;
assign \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.fas_s1  = \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.u1.s ;
assign \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.a  = \add_2ns_2ns_2_2_1_U11.din0 ;
assign \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.b  = \add_2ns_2ns_2_2_1_U11.din1 ;
assign \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.ce  = \add_2ns_2ns_2_2_1_U11.ce ;
assign \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.clk  = \add_2ns_2ns_2_2_1_U11.clk ;
assign \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.reset  = \add_2ns_2ns_2_2_1_U11.reset ;
assign \add_2ns_2ns_2_2_1_U11.dout  = \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.s ;
assign \add_2ns_2ns_2_2_1_U11.ce  = 1'h1;
assign \add_2ns_2ns_2_2_1_U11.clk  = ap_clk;
assign \add_2ns_2ns_2_2_1_U11.din0  = ret_V_4_cast_reg_844;
assign \add_2ns_2ns_2_2_1_U11.din1  = 2'h1;
assign grp_fu_485_p2 = \add_2ns_2ns_2_2_1_U11.dout ;
assign \add_2ns_2ns_2_2_1_U11.reset  = ap_rst;
assign \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.ain_s0  = \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.a ;
assign \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.bin_s0  = \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.b ;
assign \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.s  = { \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.fas_s2 , \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.sum_s1  };
assign \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.u2.a  = \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.ain_s1 ;
assign \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.u2.b  = \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.bin_s1 ;
assign \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.u2.cin  = \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.carry_s1 ;
assign \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.facout_s2  = \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.u2.cout ;
assign \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.fas_s2  = \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.u2.s ;
assign \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.u1.a  = \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.a [9:0];
assign \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.u1.b  = \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.b [9:0];
assign \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.u1.cin  = 1'h0;
assign \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.facout_s1  = \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.u1.cout ;
assign \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.fas_s1  = \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.u1.s ;
assign \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.a  = \add_20s_20s_20_2_1_U16.din0 ;
assign \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.b  = \add_20s_20s_20_2_1_U16.din1 ;
assign \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.ce  = \add_20s_20s_20_2_1_U16.ce ;
assign \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.clk  = \add_20s_20s_20_2_1_U16.clk ;
assign \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.reset  = \add_20s_20s_20_2_1_U16.reset ;
assign \add_20s_20s_20_2_1_U16.dout  = \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.s ;
assign \add_20s_20s_20_2_1_U16.ce  = 1'h1;
assign \add_20s_20s_20_2_1_U16.clk  = ap_clk;
assign \add_20s_20s_20_2_1_U16.din0  = { op_23_V_reg_943[17], op_23_V_reg_943, 1'h0 };
assign \add_20s_20s_20_2_1_U16.din1  = { op_15[1], op_15[1], op_15[1], op_15[1], op_15[1], op_15[1], op_15[1], op_15[1], op_15[1], op_15[1], op_15[1], op_15[1], op_15[1], op_15[1], op_15[1], op_15[1], op_15[1], op_15[1], op_15 };
assign grp_fu_600_p2 = \add_20s_20s_20_2_1_U16.dout ;
assign \add_20s_20s_20_2_1_U16.reset  = ap_rst;
assign \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.ain_s0  = \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.a ;
assign \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.bin_s0  = \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.b ;
assign \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.s  = { \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.fas_s2 , \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.sum_s1  };
assign \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.u2.a  = \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.ain_s1 ;
assign \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.u2.b  = \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.bin_s1 ;
assign \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.u2.cin  = \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.carry_s1 ;
assign \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.facout_s2  = \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.u2.cout ;
assign \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.fas_s2  = \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.u2.s ;
assign \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.u1.a  = \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.a [9:0];
assign \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.u1.b  = \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.b [9:0];
assign \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.u1.cin  = 1'h0;
assign \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.facout_s1  = \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.u1.cout ;
assign \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.fas_s1  = \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.u1.s ;
assign \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.a  = \add_20s_20ns_20_2_1_U19.din0 ;
assign \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.b  = \add_20s_20ns_20_2_1_U19.din1 ;
assign \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.ce  = \add_20s_20ns_20_2_1_U19.ce ;
assign \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.clk  = \add_20s_20ns_20_2_1_U19.clk ;
assign \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.reset  = \add_20s_20ns_20_2_1_U19.reset ;
assign \add_20s_20ns_20_2_1_U19.dout  = \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.s ;
assign \add_20s_20ns_20_2_1_U19.ce  = 1'h1;
assign \add_20s_20ns_20_2_1_U19.clk  = ap_clk;
assign \add_20s_20ns_20_2_1_U19.din0  = { add_ln69_4_reg_809[16], add_ln69_4_reg_809[16], add_ln69_4_reg_809[16], add_ln69_4_reg_809 };
assign \add_20s_20ns_20_2_1_U19.din1  = add_ln69_3_reg_995;
assign grp_fu_659_p2 = \add_20s_20ns_20_2_1_U19.dout ;
assign \add_20s_20ns_20_2_1_U19.reset  = ap_rst;
assign \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.ain_s0  = \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.a ;
assign \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.bin_s0  = \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.b ;
assign \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.s  = { \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.fas_s2 , \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.sum_s1  };
assign \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.u2.a  = \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.ain_s1 ;
assign \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.u2.b  = \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.bin_s1 ;
assign \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.u2.cin  = \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.carry_s1 ;
assign \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.facout_s2  = \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.u2.cout ;
assign \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.fas_s2  = \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.u2.s ;
assign \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.u1.a  = \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.a [9:0];
assign \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.u1.b  = \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.b [9:0];
assign \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.u1.cin  = 1'h0;
assign \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.facout_s1  = \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.u1.cout ;
assign \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.fas_s1  = \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.u1.s ;
assign \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.a  = \add_20s_20ns_20_2_1_U17.din0 ;
assign \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.b  = \add_20s_20ns_20_2_1_U17.din1 ;
assign \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.ce  = \add_20s_20ns_20_2_1_U17.ce ;
assign \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.clk  = \add_20s_20ns_20_2_1_U17.clk ;
assign \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.reset  = \add_20s_20ns_20_2_1_U17.reset ;
assign \add_20s_20ns_20_2_1_U17.dout  = \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.s ;
assign \add_20s_20ns_20_2_1_U17.ce  = 1'h1;
assign \add_20s_20ns_20_2_1_U17.clk  = ap_clk;
assign \add_20s_20ns_20_2_1_U17.din0  = { tmp_3_reg_968[18], tmp_3_reg_968 };
assign \add_20s_20ns_20_2_1_U17.din1  = 20'h00001;
assign grp_fu_619_p2 = \add_20s_20ns_20_2_1_U17.dout ;
assign \add_20s_20ns_20_2_1_U17.reset  = ap_rst;
assign \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.ain_s0  = \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.a ;
assign \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.bin_s0  = \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.b ;
assign \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.s  = { \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.fas_s2 , \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.sum_s1  };
assign \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.u2.a  = \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.ain_s1 ;
assign \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.u2.b  = \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.bin_s1 ;
assign \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.u2.cin  = \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.carry_s1 ;
assign \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.facout_s2  = \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.u2.cout ;
assign \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.fas_s2  = \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.u2.s ;
assign \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.u1.a  = \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.a [9:0];
assign \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.u1.b  = \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.b [9:0];
assign \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.u1.cin  = 1'h0;
assign \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.facout_s1  = \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.u1.cout ;
assign \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.fas_s1  = \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.u1.s ;
assign \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.a  = \add_20ns_20s_20_2_1_U10.din0 ;
assign \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.b  = \add_20ns_20s_20_2_1_U10.din1 ;
assign \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.ce  = \add_20ns_20s_20_2_1_U10.ce ;
assign \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.clk  = \add_20ns_20s_20_2_1_U10.clk ;
assign \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.reset  = \add_20ns_20s_20_2_1_U10.reset ;
assign \add_20ns_20s_20_2_1_U10.dout  = \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.s ;
assign \add_20ns_20s_20_2_1_U10.ce  = 1'h1;
assign \add_20ns_20s_20_2_1_U10.clk  = ap_clk;
assign \add_20ns_20s_20_2_1_U10.din0  = { 1'h0, mul_ln728_reg_814, 3'h0 };
assign \add_20ns_20s_20_2_1_U10.din1  = { op_7[3], op_7[3], op_7[3], op_7[3], op_7[3], op_7[3], op_7[3], op_7[3], op_7[3], op_7[3], op_7[3], op_7[3], op_7[3], op_7[3], op_7[3], op_7[3], op_7 };
assign grp_fu_415_p2 = \add_20ns_20s_20_2_1_U10.dout ;
assign \add_20ns_20s_20_2_1_U10.reset  = ap_rst;
assign \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.ain_s0  = \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.a ;
assign \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.bin_s0  = \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.b ;
assign \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.s  = { \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.fas_s2 , \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.sum_s1  };
assign \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.u2.a  = \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.ain_s1 ;
assign \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.u2.b  = \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.bin_s1 ;
assign \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.u2.cin  = \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.carry_s1 ;
assign \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.facout_s2  = \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.u2.cout ;
assign \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.fas_s2  = \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.u2.s ;
assign \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.u1.a  = \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.a [9:0];
assign \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.u1.b  = \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.b [9:0];
assign \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.u1.cin  = 1'h0;
assign \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.facout_s1  = \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.u1.cout ;
assign \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.fas_s1  = \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.u1.s ;
assign \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.a  = \add_20ns_20ns_20_2_1_U18.din0 ;
assign \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.b  = \add_20ns_20ns_20_2_1_U18.din1 ;
assign \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.ce  = \add_20ns_20ns_20_2_1_U18.ce ;
assign \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.clk  = \add_20ns_20ns_20_2_1_U18.clk ;
assign \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.reset  = \add_20ns_20ns_20_2_1_U18.reset ;
assign \add_20ns_20ns_20_2_1_U18.dout  = \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.s ;
assign \add_20ns_20ns_20_2_1_U18.ce  = 1'h1;
assign \add_20ns_20ns_20_2_1_U18.clk  = ap_clk;
assign \add_20ns_20ns_20_2_1_U18.din0  = { 19'h00000, op_25_V_reg_898 };
assign \add_20ns_20ns_20_2_1_U18.din1  = ret_V_25_reg_985;
assign grp_fu_651_p2 = \add_20ns_20ns_20_2_1_U18.dout ;
assign \add_20ns_20ns_20_2_1_U18.reset  = ap_rst;
assign \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.ain_s0  = \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.a ;
assign \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.bin_s0  = \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.b ;
assign \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.s  = { \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.fas_s2 , \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.sum_s1  };
assign \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.u2.a  = \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.ain_s1 ;
assign \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.u2.b  = \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.bin_s1 ;
assign \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.u2.cin  = \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.carry_s1 ;
assign \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.facout_s2  = \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.u2.cout ;
assign \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.fas_s2  = \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.u2.s ;
assign \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.u1.a  = \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.a [8:0];
assign \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.u1.b  = \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.b [8:0];
assign \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.u1.cin  = 1'h0;
assign \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.facout_s1  = \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.u1.cout ;
assign \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.fas_s1  = \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.u1.s ;
assign \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.a  = \add_18s_18ns_18_2_1_U15.din0 ;
assign \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.b  = \add_18s_18ns_18_2_1_U15.din1 ;
assign \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.ce  = \add_18s_18ns_18_2_1_U15.ce ;
assign \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.clk  = \add_18s_18ns_18_2_1_U15.clk ;
assign \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.reset  = \add_18s_18ns_18_2_1_U15.reset ;
assign \add_18s_18ns_18_2_1_U15.dout  = \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.s ;
assign \add_18s_18ns_18_2_1_U15.ce  = 1'h1;
assign \add_18s_18ns_18_2_1_U15.clk  = ap_clk;
assign \add_18s_18ns_18_2_1_U15.din0  = { add_ln69_1_reg_933[3], add_ln69_1_reg_933[3], add_ln69_1_reg_933[3], add_ln69_1_reg_933[3], add_ln69_1_reg_933[3], add_ln69_1_reg_933[3], add_ln69_1_reg_933[3], add_ln69_1_reg_933[3], add_ln69_1_reg_933[3], add_ln69_1_reg_933[3], add_ln69_1_reg_933[3], add_ln69_1_reg_933[3], add_ln69_1_reg_933[3], add_ln69_1_reg_933[3], add_ln69_1_reg_933 };
assign \add_18s_18ns_18_2_1_U15.din1  = add_ln69_reg_928;
assign grp_fu_580_p2 = \add_18s_18ns_18_2_1_U15.dout ;
assign \add_18s_18ns_18_2_1_U15.reset  = ap_rst;
assign \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.ain_s0  = \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.a ;
assign \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.bin_s0  = \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.b ;
assign \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.s  = { \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.fas_s2 , \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.sum_s1  };
assign \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.u2.a  = \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.ain_s1 ;
assign \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.u2.b  = \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.bin_s1 ;
assign \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.u2.cin  = \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.carry_s1 ;
assign \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.facout_s2  = \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.u2.cout ;
assign \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.fas_s2  = \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.u2.s ;
assign \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.u1.a  = \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.a [8:0];
assign \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.u1.b  = \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.b [8:0];
assign \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.u1.cin  = 1'h0;
assign \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.facout_s1  = \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.u1.cout ;
assign \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.fas_s1  = \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.u1.s ;
assign \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.a  = \add_18s_18ns_18_2_1_U12.din0 ;
assign \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.b  = \add_18s_18ns_18_2_1_U12.din1 ;
assign \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.ce  = \add_18s_18ns_18_2_1_U12.ce ;
assign \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.clk  = \add_18s_18ns_18_2_1_U12.clk ;
assign \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.reset  = \add_18s_18ns_18_2_1_U12.reset ;
assign \add_18s_18ns_18_2_1_U12.dout  = \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.s ;
assign \add_18s_18ns_18_2_1_U12.ce  = 1'h1;
assign \add_18s_18ns_18_2_1_U12.clk  = ap_clk;
assign \add_18s_18ns_18_2_1_U12.din0  = { ret_V_8_reg_861[16], ret_V_8_reg_861 };
assign \add_18s_18ns_18_2_1_U12.din1  = 18'h00001;
assign grp_fu_493_p2 = \add_18s_18ns_18_2_1_U12.dout ;
assign \add_18s_18ns_18_2_1_U12.reset  = ap_rst;
assign \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.ain_s0  = \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.a ;
assign \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.bin_s0  = \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.b ;
assign \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.s  = { \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.fas_s2 , \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.sum_s1  };
assign \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.u2.a  = \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.ain_s1 ;
assign \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.u2.b  = \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.bin_s1 ;
assign \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.u2.cin  = \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.carry_s1 ;
assign \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.facout_s2  = \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.u2.cout ;
assign \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.fas_s2  = \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.u2.s ;
assign \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.u1.a  = \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.a [8:0];
assign \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.u1.b  = \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.b [8:0];
assign \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.u1.cin  = 1'h0;
assign \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.facout_s1  = \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.u1.cout ;
assign \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.fas_s1  = \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.u1.s ;
assign \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.a  = \add_18ns_18ns_18_2_1_U13.din0 ;
assign \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.b  = \add_18ns_18ns_18_2_1_U13.din1 ;
assign \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.ce  = \add_18ns_18ns_18_2_1_U13.ce ;
assign \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.clk  = \add_18ns_18ns_18_2_1_U13.clk ;
assign \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.reset  = \add_18ns_18ns_18_2_1_U13.reset ;
assign \add_18ns_18ns_18_2_1_U13.dout  = \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.s ;
assign \add_18ns_18ns_18_2_1_U13.ce  = 1'h1;
assign \add_18ns_18ns_18_2_1_U13.clk  = ap_clk;
assign \add_18ns_18ns_18_2_1_U13.din0  = ret_V_21_reg_908;
assign \add_18ns_18ns_18_2_1_U13.din1  = { 16'h0000, ret_V_19_reg_903 };
assign grp_fu_566_p2 = \add_18ns_18ns_18_2_1_U13.dout ;
assign \add_18ns_18ns_18_2_1_U13.reset  = ap_rst;
assign \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.ain_s0  = \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.a ;
assign \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.bin_s0  = \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.b ;
assign \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.s  = { \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.fas_s2 , \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.sum_s1  };
assign \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.u2.a  = \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.ain_s1 ;
assign \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.u2.b  = \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.bin_s1 ;
assign \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.u2.cin  = \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.carry_s1 ;
assign \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.facout_s2  = \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.u2.cout ;
assign \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.fas_s2  = \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.u2.s ;
assign \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.u1.a  = \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.a [7:0];
assign \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.u1.b  = \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.b [7:0];
assign \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.u1.cin  = 1'h0;
assign \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.facout_s1  = \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.u1.cout ;
assign \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.fas_s1  = \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.u1.s ;
assign \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.a  = \add_17s_17s_17_2_1_U9.din0 ;
assign \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.b  = \add_17s_17s_17_2_1_U9.din1 ;
assign \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.ce  = \add_17s_17s_17_2_1_U9.ce ;
assign \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.clk  = \add_17s_17s_17_2_1_U9.clk ;
assign \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.reset  = \add_17s_17s_17_2_1_U9.reset ;
assign \add_17s_17s_17_2_1_U9.dout  = \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.s ;
assign \add_17s_17s_17_2_1_U9.ce  = 1'h1;
assign \add_17s_17s_17_2_1_U9.clk  = ap_clk;
assign \add_17s_17s_17_2_1_U9.din0  = { ret_V_17_reg_779[15], ret_V_17_reg_779 };
assign \add_17s_17s_17_2_1_U9.din1  = { r_reg_774[3], r_reg_774[3], r_reg_774[3], r_reg_774[3], r_reg_774[3], r_reg_774[3], r_reg_774[3], r_reg_774[3], r_reg_774[3], r_reg_774[3], r_reg_774[3], r_reg_774[3], r_reg_774[3], r_reg_774 };
assign grp_fu_375_p2 = \add_17s_17s_17_2_1_U9.dout ;
assign \add_17s_17s_17_2_1_U9.reset  = ap_rst;
assign \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.ain_s0  = \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.a ;
assign \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.bin_s0  = \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.b ;
assign \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.s  = { \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.fas_s2 , \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.sum_s1  };
assign \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.u2.a  = \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.ain_s1 ;
assign \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.u2.b  = \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.bin_s1 ;
assign \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.u2.cin  = \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.carry_s1 ;
assign \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.facout_s2  = \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.u2.cout ;
assign \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.fas_s2  = \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.u2.s ;
assign \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.u1.a  = \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.a [7:0];
assign \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.u1.b  = \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.b [7:0];
assign \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.u1.cin  = 1'h0;
assign \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.facout_s1  = \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.u1.cout ;
assign \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.fas_s1  = \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.u1.s ;
assign \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.a  = \add_16ns_16ns_16_2_1_U4.din0 ;
assign \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.b  = \add_16ns_16ns_16_2_1_U4.din1 ;
assign \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.ce  = \add_16ns_16ns_16_2_1_U4.ce ;
assign \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.clk  = \add_16ns_16ns_16_2_1_U4.clk ;
assign \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.reset  = \add_16ns_16ns_16_2_1_U4.reset ;
assign \add_16ns_16ns_16_2_1_U4.dout  = \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.s ;
assign \add_16ns_16ns_16_2_1_U4.ce  = 1'h1;
assign \add_16ns_16ns_16_2_1_U4.clk  = ap_clk;
assign \add_16ns_16ns_16_2_1_U4.din0  = ret_V_reg_699;
assign \add_16ns_16ns_16_2_1_U4.din1  = 16'h0001;
assign grp_fu_276_p2 = \add_16ns_16ns_16_2_1_U4.dout ;
assign \add_16ns_16ns_16_2_1_U4.reset  = ap_rst;
endmodule


// Machine B:
// Processed by function `add_clk_enable_signal` in `verilog_tricks.py`.
// Processed by function `remove_reset_signal` in `verilog_tricks.py`.
module top_B (
  ap_clk,
  ap_start,
  ap_done,
  ap_idle,
  ap_ready,
  op_0,
  op_1,
  op_2,
  op_5,
  op_7,
  op_8,
  op_9,
  op_10,
  op_13,
  op_15,
  op_28,
  op_28_ap_vld,
clk_enable
);
input clk_enable;


input ap_clk;
wire ap_rst;
assign ap_rst = op_28_ap_vld;
input ap_start;
input [7:0] op_0;
input [15:0] op_1;
input [1:0] op_10;
input [1:0] op_13;
input [1:0] op_15;
input [7:0] op_2;
input [3:0] op_5;
input [3:0] op_7;
input [15:0] op_8;
input [3:0] op_9;
output ap_done;
output ap_idle;
output ap_ready;
output [31:0] op_28;
output op_28_ap_vld;


reg [7:0] \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.ain_s1 ;
reg [7:0] \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.bin_s1 ;
reg \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.carry_s1 ;
reg [7:0] \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.sum_s1 ;
reg [8:0] \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.ain_s1 ;
reg [8:0] \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.bin_s1 ;
reg \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.carry_s1 ;
reg [7:0] \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.sum_s1 ;
reg [8:0] \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.ain_s1 ;
reg [8:0] \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.bin_s1 ;
reg \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.carry_s1 ;
reg [8:0] \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.sum_s1 ;
reg [8:0] \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.ain_s1 ;
reg [8:0] \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.bin_s1 ;
reg \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.carry_s1 ;
reg [8:0] \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.sum_s1 ;
reg [8:0] \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.ain_s1 ;
reg [8:0] \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.bin_s1 ;
reg \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.carry_s1 ;
reg [8:0] \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.sum_s1 ;
reg [9:0] \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.ain_s1 ;
reg [9:0] \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.bin_s1 ;
reg \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.carry_s1 ;
reg [9:0] \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.sum_s1 ;
reg [9:0] \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.ain_s1 ;
reg [9:0] \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.bin_s1 ;
reg \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.carry_s1 ;
reg [9:0] \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.sum_s1 ;
reg [9:0] \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.ain_s1 ;
reg [9:0] \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.bin_s1 ;
reg \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.carry_s1 ;
reg [9:0] \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.sum_s1 ;
reg [9:0] \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.ain_s1 ;
reg [9:0] \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.bin_s1 ;
reg \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.carry_s1 ;
reg [9:0] \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.sum_s1 ;
reg [9:0] \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.ain_s1 ;
reg [9:0] \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.bin_s1 ;
reg \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.carry_s1 ;
reg [9:0] \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.sum_s1 ;
reg \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.ain_s1 ;
reg \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.bin_s1 ;
reg \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.carry_s1 ;
reg \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.sum_s1 ;
reg \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.ain_s1 ;
reg \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.bin_s1 ;
reg \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.carry_s1 ;
reg \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.sum_s1 ;
reg [1:0] \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.ain_s1 ;
reg [1:0] \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.bin_s1 ;
reg \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.carry_s1 ;
reg [1:0] \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.sum_s1 ;
reg [19:0] add_ln691_reg_980;
reg [3:0] add_ln69_1_reg_933;
reg [19:0] add_ln69_3_reg_995;
reg [16:0] add_ln69_4_reg_809;
reg [17:0] add_ln69_reg_928;
reg [24:0] ap_CS_fsm = 25'h0000001;
reg [3:0] \ashr_9ns_4ns_9_7_1_U7.din1_cast_array[0] ;
reg [3:0] \ashr_9ns_4ns_9_7_1_U7.din1_cast_array[1] ;
reg [3:0] \ashr_9ns_4ns_9_7_1_U7.din1_cast_array[2] ;
reg [3:0] \ashr_9ns_4ns_9_7_1_U7.din1_cast_array[3] ;
reg [3:0] \ashr_9ns_4ns_9_7_1_U7.din1_cast_array[4] ;
reg [3:0] \ashr_9ns_4ns_9_7_1_U7.din1_cast_array[5] ;
reg [8:0] \ashr_9ns_4ns_9_7_1_U7.dout_array[0] ;
reg [8:0] \ashr_9ns_4ns_9_7_1_U7.dout_array[1] ;
reg [8:0] \ashr_9ns_4ns_9_7_1_U7.dout_array[2] ;
reg [8:0] \ashr_9ns_4ns_9_7_1_U7.dout_array[3] ;
reg [8:0] \ashr_9ns_4ns_9_7_1_U7.dout_array[4] ;
reg [8:0] \ashr_9ns_4ns_9_7_1_U7.dout_array[5] ;
reg [8:0] ashr_ln1333_reg_871;
reg icmp_ln851_1_reg_876;
reg icmp_ln851_2_reg_834;
reg icmp_ln851_3_reg_784;
reg icmp_ln851_reg_726;
reg isNeg_reg_693;
reg [15:0] \mul_16s_4ns_16_7_1_U1.top_mul_16s_4ns_16_7_1_Mul_DSP_0_U.a_reg0 ;
reg [3:0] \mul_16s_4ns_16_7_1_U1.top_mul_16s_4ns_16_7_1_Mul_DSP_0_U.b_reg0 ;
reg [15:0] \mul_16s_4ns_16_7_1_U1.top_mul_16s_4ns_16_7_1_Mul_DSP_0_U.buff0 ;
reg [15:0] \mul_16s_4ns_16_7_1_U1.top_mul_16s_4ns_16_7_1_Mul_DSP_0_U.buff1 ;
reg [15:0] \mul_16s_4ns_16_7_1_U1.top_mul_16s_4ns_16_7_1_Mul_DSP_0_U.buff2 ;
reg [15:0] \mul_16s_4ns_16_7_1_U1.top_mul_16s_4ns_16_7_1_Mul_DSP_0_U.buff3 ;
reg [15:0] \mul_16s_4ns_16_7_1_U1.top_mul_16s_4ns_16_7_1_Mul_DSP_0_U.buff4 ;
reg [5:0] \mul_6s_6s_6_7_1_U3.top_mul_6s_6s_6_7_1_Mul_DSP_1_U.a_reg0 ;
reg [5:0] \mul_6s_6s_6_7_1_U3.top_mul_6s_6s_6_7_1_Mul_DSP_1_U.b_reg0 ;
reg [5:0] \mul_6s_6s_6_7_1_U3.top_mul_6s_6s_6_7_1_Mul_DSP_1_U.buff0 ;
reg [5:0] \mul_6s_6s_6_7_1_U3.top_mul_6s_6s_6_7_1_Mul_DSP_1_U.buff1 ;
reg [5:0] \mul_6s_6s_6_7_1_U3.top_mul_6s_6s_6_7_1_Mul_DSP_1_U.buff2 ;
reg [5:0] \mul_6s_6s_6_7_1_U3.top_mul_6s_6s_6_7_1_Mul_DSP_1_U.buff3 ;
reg [5:0] \mul_6s_6s_6_7_1_U3.top_mul_6s_6s_6_7_1_Mul_DSP_1_U.buff4 ;
reg [15:0] mul_ln728_reg_814;
reg [5:0] mul_ln731_reg_819;
reg [17:0] op_23_V_reg_943;
reg op_25_V_reg_898;
reg [3:0] r_reg_774;
reg [1:0] ret_V_12_reg_789;
reg [15:0] ret_V_17_reg_779;
reg [1:0] ret_V_19_reg_903;
reg [19:0] ret_V_20_reg_856;
reg [1:0] ret_V_21_cast_reg_756;
reg [17:0] ret_V_21_reg_908;
reg [16:0] ret_V_22_reg_751;
reg [1:0] ret_V_23_reg_804;
reg [19:0] ret_V_24_reg_963;
reg [19:0] ret_V_25_reg_985;
reg [15:0] ret_V_2_reg_746;
reg [1:0] ret_V_4_cast_reg_844;
reg [1:0] ret_V_5_reg_888;
reg [16:0] ret_V_8_reg_861;
reg [17:0] ret_V_9_reg_893;
reg [15:0] ret_V_reg_699;
reg [17:0] sext_ln835_reg_881;
reg [19:0] sext_ln850_reg_973;
reg [3:0] \shl_9ns_4ns_9_7_1_U6.din1_cast_array[0] ;
reg [3:0] \shl_9ns_4ns_9_7_1_U6.din1_cast_array[1] ;
reg [3:0] \shl_9ns_4ns_9_7_1_U6.din1_cast_array[2] ;
reg [3:0] \shl_9ns_4ns_9_7_1_U6.din1_cast_array[3] ;
reg [3:0] \shl_9ns_4ns_9_7_1_U6.din1_cast_array[4] ;
reg [3:0] \shl_9ns_4ns_9_7_1_U6.din1_cast_array[5] ;
reg [8:0] \shl_9ns_4ns_9_7_1_U6.dout_array[0] ;
reg [8:0] \shl_9ns_4ns_9_7_1_U6.dout_array[1] ;
reg [8:0] \shl_9ns_4ns_9_7_1_U6.dout_array[2] ;
reg [8:0] \shl_9ns_4ns_9_7_1_U6.dout_array[3] ;
reg [8:0] \shl_9ns_4ns_9_7_1_U6.dout_array[4] ;
reg [8:0] \shl_9ns_4ns_9_7_1_U6.dout_array[5] ;
reg [8:0] shl_ln1299_reg_866;
reg [8:0] \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.ain_s1 ;
reg [8:0] \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.bin_s1 ;
reg \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.carry_s1 ;
reg [7:0] \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.sum_s1 ;
reg [1:0] \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.ain_s1 ;
reg [1:0] \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.bin_s1 ;
reg \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.carry_s1 ;
reg [1:0] \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.sum_s1 ;
reg [3:0] sub_ln1367_reg_721;
reg [18:0] tmp_3_reg_968;
reg [8:0] trunc_ln1118_reg_682;
reg [1:0] trunc_ln851_1_reg_851;
reg [7:0] trunc_ln851_3_reg_763;
reg [24:0] trunc_ln851_reg_706;
reg [3:0] ush_reg_741;
reg [7:0] _561_;
wire [19:0] _000_;
wire [3:0] _001_;
wire [19:0] _002_;
wire [16:0] _003_;
wire [17:0] _004_;
wire [24:0] _005_;
wire [8:0] _006_;
wire _007_;
wire _008_;
wire _009_;
wire _010_;
wire _011_;
wire [15:0] _012_;
wire [5:0] _013_;
wire [17:0] _014_;
wire _015_;
wire [3:0] _016_;
wire [1:0] _017_;
wire [15:0] _018_;
wire [7:0] _019_;
wire [1:0] _020_;
wire [19:0] _021_;
wire [1:0] _022_;
wire [17:0] _023_;
wire [16:0] _024_;
wire [1:0] _025_;
wire [19:0] _026_;
wire [19:0] _027_;
wire [15:0] _028_;
wire [1:0] _029_;
wire [1:0] _030_;
wire [16:0] _031_;
wire [17:0] _032_;
wire [15:0] _033_;
wire [17:0] _034_;
wire [19:0] _035_;
wire [8:0] _036_;
wire [3:0] _037_;
wire [18:0] _038_;
wire [8:0] _039_;
wire [7:0] _040_;
wire [24:0] _041_;
wire [3:0] _042_;
wire [1:0] _043_;
wire _044_;
wire _045_;
wire _046_;
wire _047_;
wire _048_;
wire _049_;
wire _050_;
wire _051_;
wire _052_;
wire _053_;
wire _054_;
wire _055_;
wire [7:0] _056_;
wire [7:0] _057_;
wire _058_;
wire [7:0] _059_;
wire [8:0] _060_;
wire [8:0] _061_;
wire [8:0] _062_;
wire [8:0] _063_;
wire _064_;
wire [7:0] _065_;
wire [8:0] _066_;
wire [9:0] _067_;
wire [8:0] _068_;
wire [8:0] _069_;
wire _070_;
wire [8:0] _071_;
wire [9:0] _072_;
wire [9:0] _073_;
wire [8:0] _074_;
wire [8:0] _075_;
wire _076_;
wire [8:0] _077_;
wire [9:0] _078_;
wire [9:0] _079_;
wire [8:0] _080_;
wire [8:0] _081_;
wire _082_;
wire [8:0] _083_;
wire [9:0] _084_;
wire [9:0] _085_;
wire [9:0] _086_;
wire [9:0] _087_;
wire _088_;
wire [9:0] _089_;
wire [10:0] _090_;
wire [10:0] _091_;
wire [9:0] _092_;
wire [9:0] _093_;
wire _094_;
wire [9:0] _095_;
wire [10:0] _096_;
wire [10:0] _097_;
wire [9:0] _098_;
wire [9:0] _099_;
wire _100_;
wire [9:0] _101_;
wire [10:0] _102_;
wire [10:0] _103_;
wire [9:0] _104_;
wire [9:0] _105_;
wire _106_;
wire [9:0] _107_;
wire [10:0] _108_;
wire [10:0] _109_;
wire [9:0] _110_;
wire [9:0] _111_;
wire _112_;
wire [9:0] _113_;
wire [10:0] _114_;
wire [10:0] _115_;
wire _116_;
wire _117_;
wire _118_;
wire _119_;
wire [1:0] _120_;
wire [1:0] _121_;
wire _122_;
wire _123_;
wire _124_;
wire _125_;
wire [1:0] _126_;
wire [1:0] _127_;
wire [1:0] _128_;
wire [1:0] _129_;
wire _130_;
wire [1:0] _131_;
wire [2:0] _132_;
wire [2:0] _133_;
wire [3:0] _134_;
wire [3:0] _135_;
wire [3:0] _136_;
wire [3:0] _137_;
wire [3:0] _138_;
wire [3:0] _139_;
wire [8:0] _140_;
wire [8:0] _141_;
wire [8:0] _142_;
wire [8:0] _143_;
wire [8:0] _144_;
wire [8:0] _145_;
wire [3:0] _146_;
wire [8:0] _147_;
wire [3:0] _148_;
wire [8:0] _149_;
wire [3:0] _150_;
wire [8:0] _151_;
wire [3:0] _152_;
wire [8:0] _153_;
wire [3:0] _154_;
wire [8:0] _155_;
wire [3:0] _156_;
wire [8:0] _157_;
wire [8:0] _158_;
wire [8:0] _159_;
wire [8:0] _160_;
wire [15:0] _161_;
wire [3:0] _162_;
wire [15:0] _163_;
wire [15:0] _164_;
wire [15:0] _165_;
wire [15:0] _166_;
wire [15:0] _167_;
wire [5:0] _168_;
wire [5:0] _169_;
wire [5:0] _170_;
wire [5:0] _171_;
wire [5:0] _172_;
wire [5:0] _173_;
wire [5:0] _174_;
wire [3:0] _175_;
wire [3:0] _176_;
wire [3:0] _177_;
wire [3:0] _178_;
wire [3:0] _179_;
wire [3:0] _180_;
wire [8:0] _181_;
wire [8:0] _182_;
wire [8:0] _183_;
wire [8:0] _184_;
wire [8:0] _185_;
wire [8:0] _186_;
wire [3:0] _187_;
wire [8:0] _188_;
wire [3:0] _189_;
wire [8:0] _190_;
wire [3:0] _191_;
wire [8:0] _192_;
wire [3:0] _193_;
wire [8:0] _194_;
wire [3:0] _195_;
wire [8:0] _196_;
wire [3:0] _197_;
wire [8:0] _198_;
wire [8:0] _199_;
wire [8:0] _200_;
wire [8:0] _201_;
wire [8:0] _202_;
wire [8:0] _203_;
wire _204_;
wire [7:0] _205_;
wire [8:0] _206_;
wire [9:0] _207_;
wire [1:0] _208_;
wire [1:0] _209_;
wire _210_;
wire [1:0] _211_;
wire [2:0] _212_;
wire [2:0] _213_;
wire _214_;
wire _215_;
wire _216_;
wire _217_;
wire _218_;
wire _219_;
wire _220_;
wire _221_;
wire _222_;
wire _223_;
wire _224_;
wire _225_;
wire _226_;
wire _227_;
wire _228_;
wire _229_;
wire _230_;
wire _231_;
wire _232_;
wire _233_;
wire _234_;
wire _235_;
wire _236_;
wire _237_;
wire _238_;
wire \add_16ns_16ns_16_2_1_U4.ce ;
wire \add_16ns_16ns_16_2_1_U4.clk ;
wire [15:0] \add_16ns_16ns_16_2_1_U4.din0 ;
wire [15:0] \add_16ns_16ns_16_2_1_U4.din1 ;
wire [15:0] \add_16ns_16ns_16_2_1_U4.dout ;
wire \add_16ns_16ns_16_2_1_U4.reset ;
wire [15:0] \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.a ;
wire [15:0] \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.ain_s0 ;
wire [15:0] \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.b ;
wire [15:0] \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.bin_s0 ;
wire \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.ce ;
wire \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.clk ;
wire \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.facout_s1 ;
wire \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.facout_s2 ;
wire [7:0] \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.fas_s1 ;
wire [7:0] \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.fas_s2 ;
wire \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.reset ;
wire [15:0] \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.s ;
wire [7:0] \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.u1.a ;
wire [7:0] \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.u1.b ;
wire \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.u1.cin ;
wire \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.u1.cout ;
wire [7:0] \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.u1.s ;
wire [7:0] \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.u2.a ;
wire [7:0] \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.u2.b ;
wire \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.u2.cin ;
wire \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.u2.cout ;
wire [7:0] \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.u2.s ;
wire \add_17s_17s_17_2_1_U9.ce ;
wire \add_17s_17s_17_2_1_U9.clk ;
wire [16:0] \add_17s_17s_17_2_1_U9.din0 ;
wire [16:0] \add_17s_17s_17_2_1_U9.din1 ;
wire [16:0] \add_17s_17s_17_2_1_U9.dout ;
wire \add_17s_17s_17_2_1_U9.reset ;
wire [16:0] \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.a ;
wire [16:0] \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.ain_s0 ;
wire [16:0] \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.b ;
wire [16:0] \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.bin_s0 ;
wire \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.ce ;
wire \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.clk ;
wire \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.facout_s1 ;
wire \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.facout_s2 ;
wire [7:0] \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.fas_s1 ;
wire [8:0] \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.fas_s2 ;
wire \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.reset ;
wire [16:0] \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.s ;
wire [7:0] \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.u1.a ;
wire [7:0] \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.u1.b ;
wire \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.u1.cin ;
wire \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.u1.cout ;
wire [7:0] \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.u1.s ;
wire [8:0] \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.u2.a ;
wire [8:0] \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.u2.b ;
wire \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.u2.cin ;
wire \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.u2.cout ;
wire [8:0] \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.u2.s ;
wire \add_18ns_18ns_18_2_1_U13.ce ;
wire \add_18ns_18ns_18_2_1_U13.clk ;
wire [17:0] \add_18ns_18ns_18_2_1_U13.din0 ;
wire [17:0] \add_18ns_18ns_18_2_1_U13.din1 ;
wire [17:0] \add_18ns_18ns_18_2_1_U13.dout ;
wire \add_18ns_18ns_18_2_1_U13.reset ;
wire [17:0] \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.a ;
wire [17:0] \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.ain_s0 ;
wire [17:0] \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.b ;
wire [17:0] \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.bin_s0 ;
wire \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.ce ;
wire \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.clk ;
wire \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.facout_s1 ;
wire \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.facout_s2 ;
wire [8:0] \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.fas_s1 ;
wire [8:0] \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.fas_s2 ;
wire \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.reset ;
wire [17:0] \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.s ;
wire [8:0] \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.u1.a ;
wire [8:0] \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.u1.b ;
wire \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.u1.cin ;
wire \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.u1.cout ;
wire [8:0] \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.u1.s ;
wire [8:0] \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.u2.a ;
wire [8:0] \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.u2.b ;
wire \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.u2.cin ;
wire \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.u2.cout ;
wire [8:0] \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.u2.s ;
wire \add_18s_18ns_18_2_1_U12.ce ;
wire \add_18s_18ns_18_2_1_U12.clk ;
wire [17:0] \add_18s_18ns_18_2_1_U12.din0 ;
wire [17:0] \add_18s_18ns_18_2_1_U12.din1 ;
wire [17:0] \add_18s_18ns_18_2_1_U12.dout ;
wire \add_18s_18ns_18_2_1_U12.reset ;
wire [17:0] \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.a ;
wire [17:0] \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.ain_s0 ;
wire [17:0] \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.b ;
wire [17:0] \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.bin_s0 ;
wire \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.ce ;
wire \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.clk ;
wire \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.facout_s1 ;
wire \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.facout_s2 ;
wire [8:0] \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.fas_s1 ;
wire [8:0] \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.fas_s2 ;
wire \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.reset ;
wire [17:0] \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.s ;
wire [8:0] \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.u1.a ;
wire [8:0] \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.u1.b ;
wire \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.u1.cin ;
wire \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.u1.cout ;
wire [8:0] \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.u1.s ;
wire [8:0] \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.u2.a ;
wire [8:0] \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.u2.b ;
wire \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.u2.cin ;
wire \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.u2.cout ;
wire [8:0] \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.u2.s ;
wire \add_18s_18ns_18_2_1_U15.ce ;
wire \add_18s_18ns_18_2_1_U15.clk ;
wire [17:0] \add_18s_18ns_18_2_1_U15.din0 ;
wire [17:0] \add_18s_18ns_18_2_1_U15.din1 ;
wire [17:0] \add_18s_18ns_18_2_1_U15.dout ;
wire \add_18s_18ns_18_2_1_U15.reset ;
wire [17:0] \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.a ;
wire [17:0] \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.ain_s0 ;
wire [17:0] \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.b ;
wire [17:0] \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.bin_s0 ;
wire \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.ce ;
wire \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.clk ;
wire \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.facout_s1 ;
wire \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.facout_s2 ;
wire [8:0] \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.fas_s1 ;
wire [8:0] \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.fas_s2 ;
wire \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.reset ;
wire [17:0] \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.s ;
wire [8:0] \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.u1.a ;
wire [8:0] \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.u1.b ;
wire \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.u1.cin ;
wire \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.u1.cout ;
wire [8:0] \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.u1.s ;
wire [8:0] \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.u2.a ;
wire [8:0] \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.u2.b ;
wire \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.u2.cin ;
wire \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.u2.cout ;
wire [8:0] \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.u2.s ;
wire \add_20ns_20ns_20_2_1_U18.ce ;
wire \add_20ns_20ns_20_2_1_U18.clk ;
wire [19:0] \add_20ns_20ns_20_2_1_U18.din0 ;
wire [19:0] \add_20ns_20ns_20_2_1_U18.din1 ;
wire [19:0] \add_20ns_20ns_20_2_1_U18.dout ;
wire \add_20ns_20ns_20_2_1_U18.reset ;
wire [19:0] \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.a ;
wire [19:0] \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.ain_s0 ;
wire [19:0] \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.b ;
wire [19:0] \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.bin_s0 ;
wire \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.ce ;
wire \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.clk ;
wire \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.facout_s1 ;
wire \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.facout_s2 ;
wire [9:0] \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.fas_s1 ;
wire [9:0] \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.fas_s2 ;
wire \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.reset ;
wire [19:0] \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.s ;
wire [9:0] \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.u1.a ;
wire [9:0] \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.u1.b ;
wire \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.u1.cin ;
wire \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.u1.cout ;
wire [9:0] \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.u1.s ;
wire [9:0] \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.u2.a ;
wire [9:0] \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.u2.b ;
wire \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.u2.cin ;
wire \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.u2.cout ;
wire [9:0] \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.u2.s ;
wire \add_20ns_20s_20_2_1_U10.ce ;
wire \add_20ns_20s_20_2_1_U10.clk ;
wire [19:0] \add_20ns_20s_20_2_1_U10.din0 ;
wire [19:0] \add_20ns_20s_20_2_1_U10.din1 ;
wire [19:0] \add_20ns_20s_20_2_1_U10.dout ;
wire \add_20ns_20s_20_2_1_U10.reset ;
wire [19:0] \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.a ;
wire [19:0] \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.ain_s0 ;
wire [19:0] \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.b ;
wire [19:0] \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.bin_s0 ;
wire \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.ce ;
wire \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.clk ;
wire \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.facout_s1 ;
wire \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.facout_s2 ;
wire [9:0] \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.fas_s1 ;
wire [9:0] \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.fas_s2 ;
wire \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.reset ;
wire [19:0] \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.s ;
wire [9:0] \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.u1.a ;
wire [9:0] \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.u1.b ;
wire \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.u1.cin ;
wire \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.u1.cout ;
wire [9:0] \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.u1.s ;
wire [9:0] \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.u2.a ;
wire [9:0] \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.u2.b ;
wire \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.u2.cin ;
wire \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.u2.cout ;
wire [9:0] \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.u2.s ;
wire \add_20s_20ns_20_2_1_U17.ce ;
wire \add_20s_20ns_20_2_1_U17.clk ;
wire [19:0] \add_20s_20ns_20_2_1_U17.din0 ;
wire [19:0] \add_20s_20ns_20_2_1_U17.din1 ;
wire [19:0] \add_20s_20ns_20_2_1_U17.dout ;
wire \add_20s_20ns_20_2_1_U17.reset ;
wire [19:0] \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.a ;
wire [19:0] \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.ain_s0 ;
wire [19:0] \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.b ;
wire [19:0] \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.bin_s0 ;
wire \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.ce ;
wire \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.clk ;
wire \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.facout_s1 ;
wire \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.facout_s2 ;
wire [9:0] \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.fas_s1 ;
wire [9:0] \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.fas_s2 ;
wire \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.reset ;
wire [19:0] \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.s ;
wire [9:0] \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.u1.a ;
wire [9:0] \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.u1.b ;
wire \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.u1.cin ;
wire \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.u1.cout ;
wire [9:0] \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.u1.s ;
wire [9:0] \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.u2.a ;
wire [9:0] \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.u2.b ;
wire \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.u2.cin ;
wire \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.u2.cout ;
wire [9:0] \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.u2.s ;
wire \add_20s_20ns_20_2_1_U19.ce ;
wire \add_20s_20ns_20_2_1_U19.clk ;
wire [19:0] \add_20s_20ns_20_2_1_U19.din0 ;
wire [19:0] \add_20s_20ns_20_2_1_U19.din1 ;
wire [19:0] \add_20s_20ns_20_2_1_U19.dout ;
wire \add_20s_20ns_20_2_1_U19.reset ;
wire [19:0] \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.a ;
wire [19:0] \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.ain_s0 ;
wire [19:0] \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.b ;
wire [19:0] \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.bin_s0 ;
wire \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.ce ;
wire \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.clk ;
wire \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.facout_s1 ;
wire \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.facout_s2 ;
wire [9:0] \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.fas_s1 ;
wire [9:0] \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.fas_s2 ;
wire \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.reset ;
wire [19:0] \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.s ;
wire [9:0] \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.u1.a ;
wire [9:0] \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.u1.b ;
wire \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.u1.cin ;
wire \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.u1.cout ;
wire [9:0] \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.u1.s ;
wire [9:0] \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.u2.a ;
wire [9:0] \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.u2.b ;
wire \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.u2.cin ;
wire \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.u2.cout ;
wire [9:0] \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.u2.s ;
wire \add_20s_20s_20_2_1_U16.ce ;
wire \add_20s_20s_20_2_1_U16.clk ;
wire [19:0] \add_20s_20s_20_2_1_U16.din0 ;
wire [19:0] \add_20s_20s_20_2_1_U16.din1 ;
wire [19:0] \add_20s_20s_20_2_1_U16.dout ;
wire \add_20s_20s_20_2_1_U16.reset ;
wire [19:0] \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.a ;
wire [19:0] \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.ain_s0 ;
wire [19:0] \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.b ;
wire [19:0] \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.bin_s0 ;
wire \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.ce ;
wire \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.clk ;
wire \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.facout_s1 ;
wire \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.facout_s2 ;
wire [9:0] \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.fas_s1 ;
wire [9:0] \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.fas_s2 ;
wire \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.reset ;
wire [19:0] \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.s ;
wire [9:0] \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.u1.a ;
wire [9:0] \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.u1.b ;
wire \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.u1.cin ;
wire \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.u1.cout ;
wire [9:0] \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.u1.s ;
wire [9:0] \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.u2.a ;
wire [9:0] \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.u2.b ;
wire \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.u2.cin ;
wire \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.u2.cout ;
wire [9:0] \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.u2.s ;
wire \add_2ns_2ns_2_2_1_U11.ce ;
wire \add_2ns_2ns_2_2_1_U11.clk ;
wire [1:0] \add_2ns_2ns_2_2_1_U11.din0 ;
wire [1:0] \add_2ns_2ns_2_2_1_U11.din1 ;
wire [1:0] \add_2ns_2ns_2_2_1_U11.dout ;
wire \add_2ns_2ns_2_2_1_U11.reset ;
wire [1:0] \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.a ;
wire [1:0] \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.ain_s0 ;
wire [1:0] \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.b ;
wire [1:0] \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.bin_s0 ;
wire \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.ce ;
wire \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.clk ;
wire \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.facout_s1 ;
wire \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.facout_s2 ;
wire \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.fas_s1 ;
wire \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.fas_s2 ;
wire \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.reset ;
wire [1:0] \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.s ;
wire \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.u1.a ;
wire \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.u1.b ;
wire \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.u1.cin ;
wire \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.u1.cout ;
wire \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.u1.s ;
wire \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.u2.a ;
wire \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.u2.b ;
wire \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.u2.cin ;
wire \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.u2.cout ;
wire \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.u2.s ;
wire \add_2ns_2ns_2_2_1_U8.ce ;
wire \add_2ns_2ns_2_2_1_U8.clk ;
wire [1:0] \add_2ns_2ns_2_2_1_U8.din0 ;
wire [1:0] \add_2ns_2ns_2_2_1_U8.din1 ;
wire [1:0] \add_2ns_2ns_2_2_1_U8.dout ;
wire \add_2ns_2ns_2_2_1_U8.reset ;
wire [1:0] \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.a ;
wire [1:0] \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.ain_s0 ;
wire [1:0] \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.b ;
wire [1:0] \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.bin_s0 ;
wire \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.ce ;
wire \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.clk ;
wire \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.facout_s1 ;
wire \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.facout_s2 ;
wire \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.fas_s1 ;
wire \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.fas_s2 ;
wire \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.reset ;
wire [1:0] \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.s ;
wire \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.u1.a ;
wire \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.u1.b ;
wire \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.u1.cin ;
wire \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.u1.cout ;
wire \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.u1.s ;
wire \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.u2.a ;
wire \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.u2.b ;
wire \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.u2.cin ;
wire \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.u2.cout ;
wire \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.u2.s ;
wire \add_4s_4ns_4_2_1_U14.ce ;
wire \add_4s_4ns_4_2_1_U14.clk ;
wire [3:0] \add_4s_4ns_4_2_1_U14.din0 ;
wire [3:0] \add_4s_4ns_4_2_1_U14.din1 ;
wire [3:0] \add_4s_4ns_4_2_1_U14.dout ;
wire \add_4s_4ns_4_2_1_U14.reset ;
wire [3:0] \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.a ;
wire [3:0] \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.ain_s0 ;
wire [3:0] \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.b ;
wire [3:0] \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.bin_s0 ;
wire \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.ce ;
wire \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.clk ;
wire \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.facout_s1 ;
wire \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.facout_s2 ;
wire [1:0] \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.fas_s1 ;
wire [1:0] \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.fas_s2 ;
wire \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.reset ;
wire [3:0] \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.s ;
wire [1:0] \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.u1.a ;
wire [1:0] \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.u1.b ;
wire \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.u1.cin ;
wire \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.u1.cout ;
wire [1:0] \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.u1.s ;
wire [1:0] \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.u2.a ;
wire [1:0] \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.u2.b ;
wire \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.u2.cin ;
wire \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.u2.cout ;
wire [1:0] \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.u2.s ;
wire ap_CS_fsm_state1;
wire ap_CS_fsm_state10;
wire ap_CS_fsm_state11;
wire ap_CS_fsm_state12;
wire ap_CS_fsm_state13;
wire ap_CS_fsm_state14;
wire ap_CS_fsm_state15;
wire ap_CS_fsm_state16;
wire ap_CS_fsm_state17;
wire ap_CS_fsm_state18;
wire ap_CS_fsm_state19;
wire ap_CS_fsm_state2;
wire ap_CS_fsm_state20;
wire ap_CS_fsm_state21;
wire ap_CS_fsm_state22;
wire ap_CS_fsm_state23;
wire ap_CS_fsm_state24;
wire ap_CS_fsm_state25;
wire ap_CS_fsm_state3;
wire ap_CS_fsm_state4;
wire ap_CS_fsm_state5;
wire ap_CS_fsm_state6;
wire ap_CS_fsm_state7;
wire ap_CS_fsm_state8;
wire ap_CS_fsm_state9;
wire [24:0] ap_NS_fsm;
wire ap_clk;
wire ap_done;
wire ap_idle;
wire ap_ready;
wire ap_rst;
wire ap_start;
wire \ashr_9ns_4ns_9_7_1_U7.ce ;
wire \ashr_9ns_4ns_9_7_1_U7.clk ;
wire [8:0] \ashr_9ns_4ns_9_7_1_U7.din0 ;
wire [8:0] \ashr_9ns_4ns_9_7_1_U7.din1 ;
wire [3:0] \ashr_9ns_4ns_9_7_1_U7.din1_cast ;
wire [3:0] \ashr_9ns_4ns_9_7_1_U7.din1_mask ;
wire [8:0] \ashr_9ns_4ns_9_7_1_U7.dout ;
wire \ashr_9ns_4ns_9_7_1_U7.reset ;
wire [3:0] grp_fu_201_p1;
wire [15:0] grp_fu_201_p10;
wire [15:0] grp_fu_201_p2;
wire [3:0] grp_fu_215_p2;
wire [5:0] grp_fu_257_p0;
wire [5:0] grp_fu_257_p1;
wire [5:0] grp_fu_257_p2;
wire [15:0] grp_fu_276_p2;
wire [16:0] grp_fu_297_p0;
wire [16:0] grp_fu_297_p1;
wire [16:0] grp_fu_297_p2;
wire [8:0] grp_fu_325_p2;
wire [8:0] grp_fu_330_p2;
wire [1:0] grp_fu_364_p2;
wire [16:0] grp_fu_375_p0;
wire [16:0] grp_fu_375_p1;
wire [16:0] grp_fu_375_p2;
wire [19:0] grp_fu_415_p0;
wire [19:0] grp_fu_415_p1;
wire [19:0] grp_fu_415_p2;
wire [1:0] grp_fu_485_p2;
wire [17:0] grp_fu_493_p0;
wire [17:0] grp_fu_493_p2;
wire [17:0] grp_fu_566_p1;
wire [17:0] grp_fu_566_p2;
wire [3:0] grp_fu_571_p0;
wire [3:0] grp_fu_571_p1;
wire [3:0] grp_fu_571_p2;
wire [17:0] grp_fu_580_p0;
wire [17:0] grp_fu_580_p2;
wire [19:0] grp_fu_600_p0;
wire [19:0] grp_fu_600_p1;
wire [19:0] grp_fu_600_p2;
wire [19:0] grp_fu_619_p0;
wire [19:0] grp_fu_619_p2;
wire [19:0] grp_fu_651_p0;
wire [19:0] grp_fu_651_p2;
wire [19:0] grp_fu_659_p0;
wire [19:0] grp_fu_659_p2;
wire icmp_ln851_1_fu_480_p2;
wire icmp_ln851_2_fu_425_p2;
wire icmp_ln851_3_fu_359_p2;
wire icmp_ln851_fu_271_p2;
wire [9:0] lhs_V_fu_438_p3;
wire \mul_16s_4ns_16_7_1_U1.ce ;
wire \mul_16s_4ns_16_7_1_U1.clk ;
wire [15:0] \mul_16s_4ns_16_7_1_U1.din0 ;
wire [3:0] \mul_16s_4ns_16_7_1_U1.din1 ;
wire [15:0] \mul_16s_4ns_16_7_1_U1.dout ;
wire \mul_16s_4ns_16_7_1_U1.reset ;
wire [15:0] \mul_16s_4ns_16_7_1_U1.top_mul_16s_4ns_16_7_1_Mul_DSP_0_U.a ;
wire [3:0] \mul_16s_4ns_16_7_1_U1.top_mul_16s_4ns_16_7_1_Mul_DSP_0_U.b ;
wire \mul_16s_4ns_16_7_1_U1.top_mul_16s_4ns_16_7_1_Mul_DSP_0_U.ce ;
wire \mul_16s_4ns_16_7_1_U1.top_mul_16s_4ns_16_7_1_Mul_DSP_0_U.clk ;
wire [15:0] \mul_16s_4ns_16_7_1_U1.top_mul_16s_4ns_16_7_1_Mul_DSP_0_U.p ;
wire [15:0] \mul_16s_4ns_16_7_1_U1.top_mul_16s_4ns_16_7_1_Mul_DSP_0_U.tmp_product ;
wire \mul_6s_6s_6_7_1_U3.ce ;
wire \mul_6s_6s_6_7_1_U3.clk ;
wire [5:0] \mul_6s_6s_6_7_1_U3.din0 ;
wire [5:0] \mul_6s_6s_6_7_1_U3.din1 ;
wire [5:0] \mul_6s_6s_6_7_1_U3.dout ;
wire \mul_6s_6s_6_7_1_U3.reset ;
wire [5:0] \mul_6s_6s_6_7_1_U3.top_mul_6s_6s_6_7_1_Mul_DSP_1_U.a ;
wire [5:0] \mul_6s_6s_6_7_1_U3.top_mul_6s_6s_6_7_1_Mul_DSP_1_U.b ;
wire \mul_6s_6s_6_7_1_U3.top_mul_6s_6s_6_7_1_Mul_DSP_1_U.ce ;
wire \mul_6s_6s_6_7_1_U3.top_mul_6s_6s_6_7_1_Mul_DSP_1_U.clk ;
wire [5:0] \mul_6s_6s_6_7_1_U3.top_mul_6s_6s_6_7_1_Mul_DSP_1_U.p ;
wire [5:0] \mul_6s_6s_6_7_1_U3.top_mul_6s_6s_6_7_1_Mul_DSP_1_U.tmp_product ;
wire [7:0] op_0;
wire [15:0] op_1;
wire [1:0] op_10;
wire [1:0] op_13;
wire [1:0] op_15;
wire op_16_V_fu_505_p3;
wire [7:0] op_2;
wire op_25_V_fu_512_p2;
wire [31:0] op_28;
wire op_28_ap_vld;
wire [7:0] op_4_V_fu_431_p3;
wire [3:0] op_5;
wire [15:0] op_6_V_fu_263_p3;
wire [3:0] op_7;
wire [15:0] op_8;
wire [3:0] op_9;
wire p_Result_1_fu_518_p3;
wire p_Result_2_fu_537_p3;
wire p_Result_3_fu_381_p3;
wire p_Result_4_fu_625_p3;
wire [15:0] p_Result_s_fu_340_p1;
wire p_Result_s_fu_340_p3;
wire [3:0] r_fu_335_p2;
wire [40:0] ret_V_16_fu_229_p2;
wire [15:0] ret_V_17_fu_352_p3;
wire [9:0] ret_V_18_fu_450_p2;
wire [9:0] ret_V_18_reg_839;
wire [1:0] ret_V_19_fu_530_p3;
wire [17:0] ret_V_21_fu_549_p3;
wire [1:0] ret_V_23_fu_393_p3;
wire [19:0] ret_V_25_fu_641_p3;
wire [18:0] rhs_2_fu_404_p3;
wire [9:0] rhs_3_fu_285_p3;
wire [15:0] rhs_fu_221_p1;
wire [40:0] rhs_fu_221_p3;
wire [1:0] select_ln850_1_fu_525_p3;
wire [17:0] select_ln850_2_fu_544_p3;
wire [1:0] select_ln850_3_fu_388_p3;
wire [19:0] select_ln850_4_fu_635_p3;
wire [15:0] select_ln850_fu_347_p3;
wire [1:0] sext_ln1192_1_fu_585_p0;
wire [3:0] sext_ln1192_fu_400_p0;
wire [9:0] sext_ln703_fu_446_p1;
wire [17:0] sext_ln835_fu_490_p1;
wire [19:0] sext_ln850_fu_616_p1;
wire \shl_9ns_4ns_9_7_1_U6.ce ;
wire \shl_9ns_4ns_9_7_1_U6.clk ;
wire [8:0] \shl_9ns_4ns_9_7_1_U6.din0 ;
wire [8:0] \shl_9ns_4ns_9_7_1_U6.din1 ;
wire [3:0] \shl_9ns_4ns_9_7_1_U6.din1_cast ;
wire [3:0] \shl_9ns_4ns_9_7_1_U6.din1_mask ;
wire [8:0] \shl_9ns_4ns_9_7_1_U6.dout ;
wire \shl_9ns_4ns_9_7_1_U6.reset ;
wire \sub_17ns_17ns_17_2_1_U5.ce ;
wire \sub_17ns_17ns_17_2_1_U5.clk ;
wire [16:0] \sub_17ns_17ns_17_2_1_U5.din0 ;
wire [16:0] \sub_17ns_17ns_17_2_1_U5.din1 ;
wire [16:0] \sub_17ns_17ns_17_2_1_U5.dout ;
wire \sub_17ns_17ns_17_2_1_U5.reset ;
wire [16:0] \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.a ;
wire [16:0] \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.ain_s0 ;
wire [16:0] \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.b ;
wire [16:0] \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.bin_s0 ;
wire \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.ce ;
wire \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.clk ;
wire \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.facout_s1 ;
wire \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.facout_s2 ;
wire [7:0] \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.fas_s1 ;
wire [8:0] \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.fas_s2 ;
wire \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.reset ;
wire [16:0] \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.s ;
wire [7:0] \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.u1.a ;
wire [7:0] \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.u1.b ;
wire \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.u1.cin ;
wire \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.u1.cout ;
wire [7:0] \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.u1.s ;
wire [8:0] \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.u2.a ;
wire [8:0] \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.u2.b ;
wire \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.u2.cin ;
wire \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.u2.cout ;
wire [8:0] \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.u2.s ;
wire \sub_4ns_4ns_4_2_1_U2.ce ;
wire \sub_4ns_4ns_4_2_1_U2.clk ;
wire [3:0] \sub_4ns_4ns_4_2_1_U2.din0 ;
wire [3:0] \sub_4ns_4ns_4_2_1_U2.din1 ;
wire [3:0] \sub_4ns_4ns_4_2_1_U2.dout ;
wire \sub_4ns_4ns_4_2_1_U2.reset ;
wire [3:0] \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.a ;
wire [3:0] \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.ain_s0 ;
wire [3:0] \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.b ;
wire [3:0] \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.bin_s0 ;
wire \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.ce ;
wire \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.clk ;
wire \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.facout_s1 ;
wire \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.facout_s2 ;
wire [1:0] \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.fas_s1 ;
wire [1:0] \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.fas_s2 ;
wire \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.reset ;
wire [3:0] \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.s ;
wire [1:0] \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.u1.a ;
wire [1:0] \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.u1.b ;
wire \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.u1.cin ;
wire \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.u1.cout ;
wire [1:0] \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.u1.s ;
wire [1:0] \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.u2.a ;
wire [1:0] \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.u2.b ;
wire \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.u2.cin ;
wire \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.u2.cout ;
wire [1:0] \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.u2.s ;
wire [18:0] tmp_fu_589_p3;
wire [15:0] trunc_ln1118_fu_193_p0;
wire [8:0] trunc_ln1118_fu_193_p1;
wire trunc_ln1368_1_fu_502_p1;
wire trunc_ln1368_fu_499_p1;
wire [1:0] trunc_ln851_1_fu_466_p1;
wire [3:0] trunc_ln851_2_fu_421_p0;
wire [2:0] trunc_ln851_2_fu_421_p1;
wire [7:0] trunc_ln851_3_fu_318_p1;
wire [1:0] trunc_ln851_4_fu_632_p0;
wire trunc_ln851_4_fu_632_p1;
wire [24:0] trunc_ln851_fu_245_p1;
wire [3:0] ush_fu_303_p3;
wire [8:0] zext_ln1367_fu_322_p1;


assign _044_ = _049_ & ap_CS_fsm[9];
assign _045_ = ap_CS_fsm[10] & _050_;
assign _046_ = isNeg_reg_693 & ap_CS_fsm[9];
assign _047_ = _051_ & ap_CS_fsm[0];
assign _048_ = ap_start & ap_CS_fsm[0];
assign op_25_V_fu_512_p2 = ~ op_16_V_fu_505_p3;
assign r_fu_335_p2 = ~ op_9;
assign ret_V_16_fu_229_p2[25] = ~ op_8[0];
assign _049_ = ~ isNeg_reg_693;
assign _050_ = ~ icmp_ln851_2_reg_834;
assign _051_ = ~ ap_start;
assign _052_ = ! trunc_ln851_1_reg_851;
assign _053_ = ! op_7[2:0];
assign _054_ = ! trunc_ln851_3_reg_763;
assign _055_ = ! trunc_ln851_reg_706;
always @(posedge \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.clk )
\add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.bin_s1  <= _057_;
always @(posedge \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.clk )
\add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.ain_s1  <= _056_;
always @(posedge \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.clk )
\add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.sum_s1  <= _059_;
always @(posedge \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.clk )
\add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.carry_s1  <= _058_;
assign _057_ = \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.ce  ? \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.b [15:8] : \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.bin_s1 ;
assign _056_ = \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.ce  ? \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.a [15:8] : \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.ain_s1 ;
assign _058_ = \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.ce  ? \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.facout_s1  : \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.carry_s1 ;
assign _059_ = \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.ce  ? \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.fas_s1  : \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.sum_s1 ;
assign _060_ = \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.u1.a  + \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.u1.b ;
assign { \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.u1.cout , \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.u1.s  } = _060_ + \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.u1.cin ;
assign _061_ = \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.u2.a  + \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.u2.b ;
assign { \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.u2.cout , \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.u2.s  } = _061_ + \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.u2.cin ;
always @(posedge \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.clk )
\add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.bin_s1  <= _063_;
always @(posedge \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.clk )
\add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.ain_s1  <= _062_;
always @(posedge \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.clk )
\add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.sum_s1  <= _065_;
always @(posedge \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.clk )
\add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.carry_s1  <= _064_;
assign _063_ = \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.ce  ? \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.b [16:8] : \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.bin_s1 ;
assign _062_ = \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.ce  ? \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.a [16:8] : \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.ain_s1 ;
assign _064_ = \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.ce  ? \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.facout_s1  : \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.carry_s1 ;
assign _065_ = \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.ce  ? \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.fas_s1  : \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.sum_s1 ;
assign _066_ = \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.u1.a  + \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.u1.b ;
assign { \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.u1.cout , \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.u1.s  } = _066_ + \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.u1.cin ;
assign _067_ = \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.u2.a  + \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.u2.b ;
assign { \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.u2.cout , \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.u2.s  } = _067_ + \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.u2.cin ;
always @(posedge \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.clk )
\add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.bin_s1  <= _069_;
always @(posedge \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.clk )
\add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.ain_s1  <= _068_;
always @(posedge \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.clk )
\add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.sum_s1  <= _071_;
always @(posedge \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.clk )
\add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.carry_s1  <= _070_;
assign _069_ = \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.ce  ? \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.b [17:9] : \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.bin_s1 ;
assign _068_ = \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.ce  ? \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.a [17:9] : \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.ain_s1 ;
assign _070_ = \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.ce  ? \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.facout_s1  : \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.carry_s1 ;
assign _071_ = \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.ce  ? \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.fas_s1  : \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.sum_s1 ;
assign _072_ = \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.u1.a  + \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.u1.b ;
assign { \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.u1.cout , \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.u1.s  } = _072_ + \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.u1.cin ;
assign _073_ = \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.u2.a  + \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.u2.b ;
assign { \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.u2.cout , \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.u2.s  } = _073_ + \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.u2.cin ;
always @(posedge \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.clk )
\add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.bin_s1  <= _075_;
always @(posedge \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.clk )
\add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.ain_s1  <= _074_;
always @(posedge \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.clk )
\add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.sum_s1  <= _077_;
always @(posedge \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.clk )
\add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.carry_s1  <= _076_;
assign _075_ = \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.ce  ? \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.b [17:9] : \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.bin_s1 ;
assign _074_ = \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.ce  ? \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.a [17:9] : \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.ain_s1 ;
assign _076_ = \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.ce  ? \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.facout_s1  : \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.carry_s1 ;
assign _077_ = \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.ce  ? \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.fas_s1  : \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.sum_s1 ;
assign _078_ = \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.u1.a  + \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.u1.b ;
assign { \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.u1.cout , \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.u1.s  } = _078_ + \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.u1.cin ;
assign _079_ = \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.u2.a  + \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.u2.b ;
assign { \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.u2.cout , \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.u2.s  } = _079_ + \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.u2.cin ;
always @(posedge \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.clk )
\add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.bin_s1  <= _081_;
always @(posedge \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.clk )
\add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.ain_s1  <= _080_;
always @(posedge \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.clk )
\add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.sum_s1  <= _083_;
always @(posedge \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.clk )
\add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.carry_s1  <= _082_;
assign _081_ = \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.ce  ? \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.b [17:9] : \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.bin_s1 ;
assign _080_ = \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.ce  ? \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.a [17:9] : \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.ain_s1 ;
assign _082_ = \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.ce  ? \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.facout_s1  : \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.carry_s1 ;
assign _083_ = \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.ce  ? \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.fas_s1  : \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.sum_s1 ;
assign _084_ = \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.u1.a  + \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.u1.b ;
assign { \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.u1.cout , \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.u1.s  } = _084_ + \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.u1.cin ;
assign _085_ = \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.u2.a  + \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.u2.b ;
assign { \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.u2.cout , \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.u2.s  } = _085_ + \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.u2.cin ;
always @(posedge \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.clk )
\add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.bin_s1  <= _087_;
always @(posedge \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.clk )
\add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.ain_s1  <= _086_;
always @(posedge \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.clk )
\add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.sum_s1  <= _089_;
always @(posedge \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.clk )
\add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.carry_s1  <= _088_;
assign _087_ = \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.ce  ? \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.b [19:10] : \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.bin_s1 ;
assign _086_ = \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.ce  ? \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.a [19:10] : \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.ain_s1 ;
assign _088_ = \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.ce  ? \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.facout_s1  : \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.carry_s1 ;
assign _089_ = \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.ce  ? \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.fas_s1  : \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.sum_s1 ;
assign _090_ = \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.u1.a  + \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.u1.b ;
assign { \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.u1.cout , \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.u1.s  } = _090_ + \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.u1.cin ;
assign _091_ = \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.u2.a  + \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.u2.b ;
assign { \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.u2.cout , \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.u2.s  } = _091_ + \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.u2.cin ;
always @(posedge \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.clk )
\add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.bin_s1  <= _093_;
always @(posedge \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.clk )
\add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.ain_s1  <= _092_;
always @(posedge \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.clk )
\add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.sum_s1  <= _095_;
always @(posedge \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.clk )
\add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.carry_s1  <= _094_;
assign _093_ = \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.ce  ? \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.b [19:10] : \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.bin_s1 ;
assign _092_ = \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.ce  ? \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.a [19:10] : \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.ain_s1 ;
assign _094_ = \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.ce  ? \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.facout_s1  : \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.carry_s1 ;
assign _095_ = \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.ce  ? \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.fas_s1  : \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.sum_s1 ;
assign _096_ = \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.u1.a  + \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.u1.b ;
assign { \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.u1.cout , \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.u1.s  } = _096_ + \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.u1.cin ;
assign _097_ = \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.u2.a  + \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.u2.b ;
assign { \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.u2.cout , \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.u2.s  } = _097_ + \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.u2.cin ;
always @(posedge \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.clk )
\add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.bin_s1  <= _099_;
always @(posedge \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.clk )
\add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.ain_s1  <= _098_;
always @(posedge \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.clk )
\add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.sum_s1  <= _101_;
always @(posedge \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.clk )
\add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.carry_s1  <= _100_;
assign _099_ = \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.ce  ? \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.b [19:10] : \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.bin_s1 ;
assign _098_ = \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.ce  ? \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.a [19:10] : \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.ain_s1 ;
assign _100_ = \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.ce  ? \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.facout_s1  : \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.carry_s1 ;
assign _101_ = \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.ce  ? \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.fas_s1  : \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.sum_s1 ;
assign _102_ = \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.u1.a  + \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.u1.b ;
assign { \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.u1.cout , \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.u1.s  } = _102_ + \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.u1.cin ;
assign _103_ = \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.u2.a  + \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.u2.b ;
assign { \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.u2.cout , \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.u2.s  } = _103_ + \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.u2.cin ;
always @(posedge \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.clk )
\add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.bin_s1  <= _105_;
always @(posedge \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.clk )
\add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.ain_s1  <= _104_;
always @(posedge \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.clk )
\add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.sum_s1  <= _107_;
always @(posedge \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.clk )
\add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.carry_s1  <= _106_;
assign _105_ = \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.ce  ? \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.b [19:10] : \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.bin_s1 ;
assign _104_ = \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.ce  ? \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.a [19:10] : \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.ain_s1 ;
assign _106_ = \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.ce  ? \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.facout_s1  : \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.carry_s1 ;
assign _107_ = \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.ce  ? \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.fas_s1  : \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.sum_s1 ;
assign _108_ = \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.u1.a  + \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.u1.b ;
assign { \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.u1.cout , \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.u1.s  } = _108_ + \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.u1.cin ;
assign _109_ = \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.u2.a  + \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.u2.b ;
assign { \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.u2.cout , \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.u2.s  } = _109_ + \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.u2.cin ;
always @(posedge \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.clk )
\add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.bin_s1  <= _111_;
always @(posedge \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.clk )
\add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.ain_s1  <= _110_;
always @(posedge \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.clk )
\add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.sum_s1  <= _113_;
always @(posedge \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.clk )
\add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.carry_s1  <= _112_;
assign _111_ = \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.ce  ? \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.b [19:10] : \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.bin_s1 ;
assign _110_ = \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.ce  ? \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.a [19:10] : \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.ain_s1 ;
assign _112_ = \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.ce  ? \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.facout_s1  : \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.carry_s1 ;
assign _113_ = \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.ce  ? \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.fas_s1  : \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.sum_s1 ;
assign _114_ = \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.u1.a  + \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.u1.b ;
assign { \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.u1.cout , \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.u1.s  } = _114_ + \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.u1.cin ;
assign _115_ = \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.u2.a  + \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.u2.b ;
assign { \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.u2.cout , \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.u2.s  } = _115_ + \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.u2.cin ;
always @(posedge \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.clk )
\add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.bin_s1  <= _117_;
always @(posedge \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.clk )
\add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.ain_s1  <= _116_;
always @(posedge \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.clk )
\add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.sum_s1  <= _119_;
always @(posedge \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.clk )
\add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.carry_s1  <= _118_;
assign _117_ = \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.ce  ? \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.b [1] : \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.bin_s1 ;
assign _116_ = \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.ce  ? \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.a [1] : \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.ain_s1 ;
assign _118_ = \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.ce  ? \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.facout_s1  : \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.carry_s1 ;
assign _119_ = \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.ce  ? \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.fas_s1  : \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.sum_s1 ;
assign _120_ = \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.u1.a  + \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.u1.b ;
assign { \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.u1.cout , \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.u1.s  } = _120_ + \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.u1.cin ;
assign _121_ = \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.u2.a  + \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.u2.b ;
assign { \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.u2.cout , \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.u2.s  } = _121_ + \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.u2.cin ;
always @(posedge \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.clk )
\add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.bin_s1  <= _123_;
always @(posedge \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.clk )
\add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.ain_s1  <= _122_;
always @(posedge \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.clk )
\add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.sum_s1  <= _125_;
always @(posedge \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.clk )
\add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.carry_s1  <= _124_;
assign _123_ = \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.ce  ? \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.b [1] : \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.bin_s1 ;
assign _122_ = \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.ce  ? \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.a [1] : \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.ain_s1 ;
assign _124_ = \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.ce  ? \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.facout_s1  : \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.carry_s1 ;
assign _125_ = \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.ce  ? \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.fas_s1  : \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.sum_s1 ;
assign _126_ = \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.u1.a  + \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.u1.b ;
assign { \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.u1.cout , \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.u1.s  } = _126_ + \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.u1.cin ;
assign _127_ = \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.u2.a  + \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.u2.b ;
assign { \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.u2.cout , \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.u2.s  } = _127_ + \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.u2.cin ;
always @(posedge \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.clk )
\add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.bin_s1  <= _129_;
always @(posedge \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.clk )
\add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.ain_s1  <= _128_;
always @(posedge \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.clk )
\add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.sum_s1  <= _131_;
always @(posedge \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.clk )
\add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.carry_s1  <= _130_;
assign _129_ = \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.ce  ? \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.b [3:2] : \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.bin_s1 ;
assign _128_ = \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.ce  ? \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.a [3:2] : \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.ain_s1 ;
assign _130_ = \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.ce  ? \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.facout_s1  : \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.carry_s1 ;
assign _131_ = \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.ce  ? \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.fas_s1  : \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.sum_s1 ;
assign _132_ = \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.u1.a  + \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.u1.b ;
assign { \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.u1.cout , \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.u1.s  } = _132_ + \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.u1.cin ;
assign _133_ = \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.u2.a  + \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.u2.b ;
assign { \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.u2.cout , \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.u2.s  } = _133_ + \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.u2.cin ;
always @(posedge \ashr_9ns_4ns_9_7_1_U7.clk )
\ashr_9ns_4ns_9_7_1_U7.dout_array[5]  <= _145_;
always @(posedge \ashr_9ns_4ns_9_7_1_U7.clk )
\ashr_9ns_4ns_9_7_1_U7.din1_cast_array[5]  <= _139_;
always @(posedge \ashr_9ns_4ns_9_7_1_U7.clk )
\ashr_9ns_4ns_9_7_1_U7.dout_array[4]  <= _144_;
always @(posedge \ashr_9ns_4ns_9_7_1_U7.clk )
\ashr_9ns_4ns_9_7_1_U7.din1_cast_array[4]  <= _138_;
always @(posedge \ashr_9ns_4ns_9_7_1_U7.clk )
\ashr_9ns_4ns_9_7_1_U7.dout_array[3]  <= _143_;
always @(posedge \ashr_9ns_4ns_9_7_1_U7.clk )
\ashr_9ns_4ns_9_7_1_U7.din1_cast_array[3]  <= _137_;
always @(posedge \ashr_9ns_4ns_9_7_1_U7.clk )
\ashr_9ns_4ns_9_7_1_U7.dout_array[2]  <= _142_;
always @(posedge \ashr_9ns_4ns_9_7_1_U7.clk )
\ashr_9ns_4ns_9_7_1_U7.din1_cast_array[2]  <= _136_;
always @(posedge \ashr_9ns_4ns_9_7_1_U7.clk )
\ashr_9ns_4ns_9_7_1_U7.dout_array[1]  <= _141_;
always @(posedge \ashr_9ns_4ns_9_7_1_U7.clk )
\ashr_9ns_4ns_9_7_1_U7.din1_cast_array[1]  <= _135_;
always @(posedge \ashr_9ns_4ns_9_7_1_U7.clk )
\ashr_9ns_4ns_9_7_1_U7.dout_array[0]  <= _140_;
always @(posedge \ashr_9ns_4ns_9_7_1_U7.clk )
\ashr_9ns_4ns_9_7_1_U7.din1_cast_array[0]  <= _134_;
assign _146_ = \ashr_9ns_4ns_9_7_1_U7.ce  ? \ashr_9ns_4ns_9_7_1_U7.din1_cast_array[4]  : \ashr_9ns_4ns_9_7_1_U7.din1_cast_array[5] ;
assign _139_ = \ashr_9ns_4ns_9_7_1_U7.reset  ? 4'h0 : _146_;
assign _147_ = \ashr_9ns_4ns_9_7_1_U7.ce  ? _160_ : \ashr_9ns_4ns_9_7_1_U7.dout_array[5] ;
assign _145_ = \ashr_9ns_4ns_9_7_1_U7.reset  ? 9'h000 : _147_;
assign _148_ = \ashr_9ns_4ns_9_7_1_U7.ce  ? \ashr_9ns_4ns_9_7_1_U7.din1_cast_array[3]  : \ashr_9ns_4ns_9_7_1_U7.din1_cast_array[4] ;
assign _138_ = \ashr_9ns_4ns_9_7_1_U7.reset  ? 4'h0 : _148_;
assign _149_ = \ashr_9ns_4ns_9_7_1_U7.ce  ? _159_ : \ashr_9ns_4ns_9_7_1_U7.dout_array[4] ;
assign _144_ = \ashr_9ns_4ns_9_7_1_U7.reset  ? 9'h000 : _149_;
assign _150_ = \ashr_9ns_4ns_9_7_1_U7.ce  ? \ashr_9ns_4ns_9_7_1_U7.din1_cast_array[2]  : \ashr_9ns_4ns_9_7_1_U7.din1_cast_array[3] ;
assign _137_ = \ashr_9ns_4ns_9_7_1_U7.reset  ? 4'h0 : _150_;
assign _151_ = \ashr_9ns_4ns_9_7_1_U7.ce  ? _158_ : \ashr_9ns_4ns_9_7_1_U7.dout_array[3] ;
assign _143_ = \ashr_9ns_4ns_9_7_1_U7.reset  ? 9'h000 : _151_;
assign _152_ = \ashr_9ns_4ns_9_7_1_U7.ce  ? \ashr_9ns_4ns_9_7_1_U7.din1_cast_array[1]  : \ashr_9ns_4ns_9_7_1_U7.din1_cast_array[2] ;
assign _136_ = \ashr_9ns_4ns_9_7_1_U7.reset  ? 4'h0 : _152_;
assign _153_ = \ashr_9ns_4ns_9_7_1_U7.ce  ? \ashr_9ns_4ns_9_7_1_U7.dout_array[1]  : \ashr_9ns_4ns_9_7_1_U7.dout_array[2] ;
assign _142_ = \ashr_9ns_4ns_9_7_1_U7.reset  ? 9'h000 : _153_;
assign _154_ = \ashr_9ns_4ns_9_7_1_U7.ce  ? \ashr_9ns_4ns_9_7_1_U7.din1_cast_array[0]  : \ashr_9ns_4ns_9_7_1_U7.din1_cast_array[1] ;
assign _135_ = \ashr_9ns_4ns_9_7_1_U7.reset  ? 4'h0 : _154_;
assign _155_ = \ashr_9ns_4ns_9_7_1_U7.ce  ? \ashr_9ns_4ns_9_7_1_U7.dout_array[0]  : \ashr_9ns_4ns_9_7_1_U7.dout_array[1] ;
assign _141_ = \ashr_9ns_4ns_9_7_1_U7.reset  ? 9'h000 : _155_;
assign _156_ = \ashr_9ns_4ns_9_7_1_U7.ce  ? \ashr_9ns_4ns_9_7_1_U7.din1 [3:0] : \ashr_9ns_4ns_9_7_1_U7.din1_cast_array[0] ;
assign _134_ = \ashr_9ns_4ns_9_7_1_U7.reset  ? 4'h0 : _156_;
assign _157_ = \ashr_9ns_4ns_9_7_1_U7.ce  ? \ashr_9ns_4ns_9_7_1_U7.din0  : \ashr_9ns_4ns_9_7_1_U7.dout_array[0] ;
assign _140_ = \ashr_9ns_4ns_9_7_1_U7.reset  ? 9'h000 : _157_;
assign _158_ = $signed(\ashr_9ns_4ns_9_7_1_U7.dout_array[2] ) >>> { \ashr_9ns_4ns_9_7_1_U7.din1_cast_array[2] [3], 3'h0 };
assign _159_ = $signed(\ashr_9ns_4ns_9_7_1_U7.dout_array[3] ) >>> { \ashr_9ns_4ns_9_7_1_U7.din1_cast_array[3] [2], 2'h0 };
assign _160_ = $signed(\ashr_9ns_4ns_9_7_1_U7.dout_array[4] ) >>> { \ashr_9ns_4ns_9_7_1_U7.din1_cast_array[4] [1], 1'h0 };
assign \ashr_9ns_4ns_9_7_1_U7.dout  = $signed(\ashr_9ns_4ns_9_7_1_U7.dout_array[5] ) >>> \ashr_9ns_4ns_9_7_1_U7.din1_cast_array[5] [0];
assign \mul_16s_4ns_16_7_1_U1.top_mul_16s_4ns_16_7_1_Mul_DSP_0_U.tmp_product  = $signed(\mul_16s_4ns_16_7_1_U1.top_mul_16s_4ns_16_7_1_Mul_DSP_0_U.a_reg0 ) * $signed({ 1'h0, \mul_16s_4ns_16_7_1_U1.top_mul_16s_4ns_16_7_1_Mul_DSP_0_U.b_reg0  });
always @(posedge \mul_16s_4ns_16_7_1_U1.top_mul_16s_4ns_16_7_1_Mul_DSP_0_U.clk )
\mul_16s_4ns_16_7_1_U1.top_mul_16s_4ns_16_7_1_Mul_DSP_0_U.a_reg0  <= _161_;
always @(posedge \mul_16s_4ns_16_7_1_U1.top_mul_16s_4ns_16_7_1_Mul_DSP_0_U.clk )
\mul_16s_4ns_16_7_1_U1.top_mul_16s_4ns_16_7_1_Mul_DSP_0_U.b_reg0  <= _162_;
always @(posedge \mul_16s_4ns_16_7_1_U1.top_mul_16s_4ns_16_7_1_Mul_DSP_0_U.clk )
\mul_16s_4ns_16_7_1_U1.top_mul_16s_4ns_16_7_1_Mul_DSP_0_U.buff0  <= _163_;
always @(posedge \mul_16s_4ns_16_7_1_U1.top_mul_16s_4ns_16_7_1_Mul_DSP_0_U.clk )
\mul_16s_4ns_16_7_1_U1.top_mul_16s_4ns_16_7_1_Mul_DSP_0_U.buff1  <= _164_;
always @(posedge \mul_16s_4ns_16_7_1_U1.top_mul_16s_4ns_16_7_1_Mul_DSP_0_U.clk )
\mul_16s_4ns_16_7_1_U1.top_mul_16s_4ns_16_7_1_Mul_DSP_0_U.buff2  <= _165_;
always @(posedge \mul_16s_4ns_16_7_1_U1.top_mul_16s_4ns_16_7_1_Mul_DSP_0_U.clk )
\mul_16s_4ns_16_7_1_U1.top_mul_16s_4ns_16_7_1_Mul_DSP_0_U.buff3  <= _166_;
always @(posedge \mul_16s_4ns_16_7_1_U1.top_mul_16s_4ns_16_7_1_Mul_DSP_0_U.clk )
\mul_16s_4ns_16_7_1_U1.top_mul_16s_4ns_16_7_1_Mul_DSP_0_U.buff4  <= _167_;
assign _167_ = \mul_16s_4ns_16_7_1_U1.top_mul_16s_4ns_16_7_1_Mul_DSP_0_U.ce  ? \mul_16s_4ns_16_7_1_U1.top_mul_16s_4ns_16_7_1_Mul_DSP_0_U.buff3  : \mul_16s_4ns_16_7_1_U1.top_mul_16s_4ns_16_7_1_Mul_DSP_0_U.buff4 ;
assign _166_ = \mul_16s_4ns_16_7_1_U1.top_mul_16s_4ns_16_7_1_Mul_DSP_0_U.ce  ? \mul_16s_4ns_16_7_1_U1.top_mul_16s_4ns_16_7_1_Mul_DSP_0_U.buff2  : \mul_16s_4ns_16_7_1_U1.top_mul_16s_4ns_16_7_1_Mul_DSP_0_U.buff3 ;
assign _165_ = \mul_16s_4ns_16_7_1_U1.top_mul_16s_4ns_16_7_1_Mul_DSP_0_U.ce  ? \mul_16s_4ns_16_7_1_U1.top_mul_16s_4ns_16_7_1_Mul_DSP_0_U.buff1  : \mul_16s_4ns_16_7_1_U1.top_mul_16s_4ns_16_7_1_Mul_DSP_0_U.buff2 ;
assign _164_ = \mul_16s_4ns_16_7_1_U1.top_mul_16s_4ns_16_7_1_Mul_DSP_0_U.ce  ? \mul_16s_4ns_16_7_1_U1.top_mul_16s_4ns_16_7_1_Mul_DSP_0_U.buff0  : \mul_16s_4ns_16_7_1_U1.top_mul_16s_4ns_16_7_1_Mul_DSP_0_U.buff1 ;
assign _163_ = \mul_16s_4ns_16_7_1_U1.top_mul_16s_4ns_16_7_1_Mul_DSP_0_U.ce  ? \mul_16s_4ns_16_7_1_U1.top_mul_16s_4ns_16_7_1_Mul_DSP_0_U.tmp_product  : \mul_16s_4ns_16_7_1_U1.top_mul_16s_4ns_16_7_1_Mul_DSP_0_U.buff0 ;
assign _162_ = \mul_16s_4ns_16_7_1_U1.top_mul_16s_4ns_16_7_1_Mul_DSP_0_U.ce  ? \mul_16s_4ns_16_7_1_U1.top_mul_16s_4ns_16_7_1_Mul_DSP_0_U.b  : \mul_16s_4ns_16_7_1_U1.top_mul_16s_4ns_16_7_1_Mul_DSP_0_U.b_reg0 ;
assign _161_ = \mul_16s_4ns_16_7_1_U1.top_mul_16s_4ns_16_7_1_Mul_DSP_0_U.ce  ? \mul_16s_4ns_16_7_1_U1.top_mul_16s_4ns_16_7_1_Mul_DSP_0_U.a  : \mul_16s_4ns_16_7_1_U1.top_mul_16s_4ns_16_7_1_Mul_DSP_0_U.a_reg0 ;
assign \mul_6s_6s_6_7_1_U3.top_mul_6s_6s_6_7_1_Mul_DSP_1_U.tmp_product  = $signed(\mul_6s_6s_6_7_1_U3.top_mul_6s_6s_6_7_1_Mul_DSP_1_U.a_reg0 ) * $signed(\mul_6s_6s_6_7_1_U3.top_mul_6s_6s_6_7_1_Mul_DSP_1_U.b_reg0 );
always @(posedge \mul_6s_6s_6_7_1_U3.top_mul_6s_6s_6_7_1_Mul_DSP_1_U.clk )
\mul_6s_6s_6_7_1_U3.top_mul_6s_6s_6_7_1_Mul_DSP_1_U.a_reg0  <= _168_;
always @(posedge \mul_6s_6s_6_7_1_U3.top_mul_6s_6s_6_7_1_Mul_DSP_1_U.clk )
\mul_6s_6s_6_7_1_U3.top_mul_6s_6s_6_7_1_Mul_DSP_1_U.b_reg0  <= _169_;
always @(posedge \mul_6s_6s_6_7_1_U3.top_mul_6s_6s_6_7_1_Mul_DSP_1_U.clk )
\mul_6s_6s_6_7_1_U3.top_mul_6s_6s_6_7_1_Mul_DSP_1_U.buff0  <= _170_;
always @(posedge \mul_6s_6s_6_7_1_U3.top_mul_6s_6s_6_7_1_Mul_DSP_1_U.clk )
\mul_6s_6s_6_7_1_U3.top_mul_6s_6s_6_7_1_Mul_DSP_1_U.buff1  <= _171_;
always @(posedge \mul_6s_6s_6_7_1_U3.top_mul_6s_6s_6_7_1_Mul_DSP_1_U.clk )
\mul_6s_6s_6_7_1_U3.top_mul_6s_6s_6_7_1_Mul_DSP_1_U.buff2  <= _172_;
always @(posedge \mul_6s_6s_6_7_1_U3.top_mul_6s_6s_6_7_1_Mul_DSP_1_U.clk )
\mul_6s_6s_6_7_1_U3.top_mul_6s_6s_6_7_1_Mul_DSP_1_U.buff3  <= _173_;
always @(posedge \mul_6s_6s_6_7_1_U3.top_mul_6s_6s_6_7_1_Mul_DSP_1_U.clk )
\mul_6s_6s_6_7_1_U3.top_mul_6s_6s_6_7_1_Mul_DSP_1_U.buff4  <= _174_;
assign _174_ = \mul_6s_6s_6_7_1_U3.top_mul_6s_6s_6_7_1_Mul_DSP_1_U.ce  ? \mul_6s_6s_6_7_1_U3.top_mul_6s_6s_6_7_1_Mul_DSP_1_U.buff3  : \mul_6s_6s_6_7_1_U3.top_mul_6s_6s_6_7_1_Mul_DSP_1_U.buff4 ;
assign _173_ = \mul_6s_6s_6_7_1_U3.top_mul_6s_6s_6_7_1_Mul_DSP_1_U.ce  ? \mul_6s_6s_6_7_1_U3.top_mul_6s_6s_6_7_1_Mul_DSP_1_U.buff2  : \mul_6s_6s_6_7_1_U3.top_mul_6s_6s_6_7_1_Mul_DSP_1_U.buff3 ;
assign _172_ = \mul_6s_6s_6_7_1_U3.top_mul_6s_6s_6_7_1_Mul_DSP_1_U.ce  ? \mul_6s_6s_6_7_1_U3.top_mul_6s_6s_6_7_1_Mul_DSP_1_U.buff1  : \mul_6s_6s_6_7_1_U3.top_mul_6s_6s_6_7_1_Mul_DSP_1_U.buff2 ;
assign _171_ = \mul_6s_6s_6_7_1_U3.top_mul_6s_6s_6_7_1_Mul_DSP_1_U.ce  ? \mul_6s_6s_6_7_1_U3.top_mul_6s_6s_6_7_1_Mul_DSP_1_U.buff0  : \mul_6s_6s_6_7_1_U3.top_mul_6s_6s_6_7_1_Mul_DSP_1_U.buff1 ;
assign _170_ = \mul_6s_6s_6_7_1_U3.top_mul_6s_6s_6_7_1_Mul_DSP_1_U.ce  ? \mul_6s_6s_6_7_1_U3.top_mul_6s_6s_6_7_1_Mul_DSP_1_U.tmp_product  : \mul_6s_6s_6_7_1_U3.top_mul_6s_6s_6_7_1_Mul_DSP_1_U.buff0 ;
assign _169_ = \mul_6s_6s_6_7_1_U3.top_mul_6s_6s_6_7_1_Mul_DSP_1_U.ce  ? \mul_6s_6s_6_7_1_U3.top_mul_6s_6s_6_7_1_Mul_DSP_1_U.b  : \mul_6s_6s_6_7_1_U3.top_mul_6s_6s_6_7_1_Mul_DSP_1_U.b_reg0 ;
assign _168_ = \mul_6s_6s_6_7_1_U3.top_mul_6s_6s_6_7_1_Mul_DSP_1_U.ce  ? \mul_6s_6s_6_7_1_U3.top_mul_6s_6s_6_7_1_Mul_DSP_1_U.a  : \mul_6s_6s_6_7_1_U3.top_mul_6s_6s_6_7_1_Mul_DSP_1_U.a_reg0 ;
always @(posedge \shl_9ns_4ns_9_7_1_U6.clk )
\shl_9ns_4ns_9_7_1_U6.dout_array[5]  <= _186_;
always @(posedge \shl_9ns_4ns_9_7_1_U6.clk )
\shl_9ns_4ns_9_7_1_U6.din1_cast_array[5]  <= _180_;
always @(posedge \shl_9ns_4ns_9_7_1_U6.clk )
\shl_9ns_4ns_9_7_1_U6.dout_array[4]  <= _185_;
always @(posedge \shl_9ns_4ns_9_7_1_U6.clk )
\shl_9ns_4ns_9_7_1_U6.din1_cast_array[4]  <= _179_;
always @(posedge \shl_9ns_4ns_9_7_1_U6.clk )
\shl_9ns_4ns_9_7_1_U6.dout_array[3]  <= _184_;
always @(posedge \shl_9ns_4ns_9_7_1_U6.clk )
\shl_9ns_4ns_9_7_1_U6.din1_cast_array[3]  <= _178_;
always @(posedge \shl_9ns_4ns_9_7_1_U6.clk )
\shl_9ns_4ns_9_7_1_U6.dout_array[2]  <= _183_;
always @(posedge \shl_9ns_4ns_9_7_1_U6.clk )
\shl_9ns_4ns_9_7_1_U6.din1_cast_array[2]  <= _177_;
always @(posedge \shl_9ns_4ns_9_7_1_U6.clk )
\shl_9ns_4ns_9_7_1_U6.dout_array[1]  <= _182_;
always @(posedge \shl_9ns_4ns_9_7_1_U6.clk )
\shl_9ns_4ns_9_7_1_U6.din1_cast_array[1]  <= _176_;
always @(posedge \shl_9ns_4ns_9_7_1_U6.clk )
\shl_9ns_4ns_9_7_1_U6.dout_array[0]  <= _181_;
always @(posedge \shl_9ns_4ns_9_7_1_U6.clk )
\shl_9ns_4ns_9_7_1_U6.din1_cast_array[0]  <= _175_;
assign _187_ = \shl_9ns_4ns_9_7_1_U6.ce  ? \shl_9ns_4ns_9_7_1_U6.din1_cast_array[4]  : \shl_9ns_4ns_9_7_1_U6.din1_cast_array[5] ;
assign _180_ = \shl_9ns_4ns_9_7_1_U6.reset  ? 4'h0 : _187_;
assign _188_ = \shl_9ns_4ns_9_7_1_U6.ce  ? _201_ : \shl_9ns_4ns_9_7_1_U6.dout_array[5] ;
assign _186_ = \shl_9ns_4ns_9_7_1_U6.reset  ? 9'h000 : _188_;
assign _189_ = \shl_9ns_4ns_9_7_1_U6.ce  ? \shl_9ns_4ns_9_7_1_U6.din1_cast_array[3]  : \shl_9ns_4ns_9_7_1_U6.din1_cast_array[4] ;
assign _179_ = \shl_9ns_4ns_9_7_1_U6.reset  ? 4'h0 : _189_;
assign _190_ = \shl_9ns_4ns_9_7_1_U6.ce  ? _200_ : \shl_9ns_4ns_9_7_1_U6.dout_array[4] ;
assign _185_ = \shl_9ns_4ns_9_7_1_U6.reset  ? 9'h000 : _190_;
assign _191_ = \shl_9ns_4ns_9_7_1_U6.ce  ? \shl_9ns_4ns_9_7_1_U6.din1_cast_array[2]  : \shl_9ns_4ns_9_7_1_U6.din1_cast_array[3] ;
assign _178_ = \shl_9ns_4ns_9_7_1_U6.reset  ? 4'h0 : _191_;
assign _192_ = \shl_9ns_4ns_9_7_1_U6.ce  ? _199_ : \shl_9ns_4ns_9_7_1_U6.dout_array[3] ;
assign _184_ = \shl_9ns_4ns_9_7_1_U6.reset  ? 9'h000 : _192_;
assign _193_ = \shl_9ns_4ns_9_7_1_U6.ce  ? \shl_9ns_4ns_9_7_1_U6.din1_cast_array[1]  : \shl_9ns_4ns_9_7_1_U6.din1_cast_array[2] ;
assign _177_ = \shl_9ns_4ns_9_7_1_U6.reset  ? 4'h0 : _193_;
assign _194_ = \shl_9ns_4ns_9_7_1_U6.ce  ? \shl_9ns_4ns_9_7_1_U6.dout_array[1]  : \shl_9ns_4ns_9_7_1_U6.dout_array[2] ;
assign _183_ = \shl_9ns_4ns_9_7_1_U6.reset  ? 9'h000 : _194_;
assign _195_ = \shl_9ns_4ns_9_7_1_U6.ce  ? \shl_9ns_4ns_9_7_1_U6.din1_cast_array[0]  : \shl_9ns_4ns_9_7_1_U6.din1_cast_array[1] ;
assign _176_ = \shl_9ns_4ns_9_7_1_U6.reset  ? 4'h0 : _195_;
assign _196_ = \shl_9ns_4ns_9_7_1_U6.ce  ? \shl_9ns_4ns_9_7_1_U6.dout_array[0]  : \shl_9ns_4ns_9_7_1_U6.dout_array[1] ;
assign _182_ = \shl_9ns_4ns_9_7_1_U6.reset  ? 9'h000 : _196_;
assign _197_ = \shl_9ns_4ns_9_7_1_U6.ce  ? \shl_9ns_4ns_9_7_1_U6.din1 [3:0] : \shl_9ns_4ns_9_7_1_U6.din1_cast_array[0] ;
assign _175_ = \shl_9ns_4ns_9_7_1_U6.reset  ? 4'h0 : _197_;
assign _198_ = \shl_9ns_4ns_9_7_1_U6.ce  ? \shl_9ns_4ns_9_7_1_U6.din0  : \shl_9ns_4ns_9_7_1_U6.dout_array[0] ;
assign _181_ = \shl_9ns_4ns_9_7_1_U6.reset  ? 9'h000 : _198_;
assign _199_ = \shl_9ns_4ns_9_7_1_U6.dout_array[2]  << { \shl_9ns_4ns_9_7_1_U6.din1_cast_array[2] [3], 3'h0 };
assign _200_ = \shl_9ns_4ns_9_7_1_U6.dout_array[3]  << { \shl_9ns_4ns_9_7_1_U6.din1_cast_array[3] [2], 2'h0 };
assign _201_ = \shl_9ns_4ns_9_7_1_U6.dout_array[4]  << { \shl_9ns_4ns_9_7_1_U6.din1_cast_array[4] [1], 1'h0 };
assign \shl_9ns_4ns_9_7_1_U6.dout  = \shl_9ns_4ns_9_7_1_U6.dout_array[5]  << \shl_9ns_4ns_9_7_1_U6.din1_cast_array[5] [0];
assign \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.bin_s0  = ~ \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.b ;
always @(posedge \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.clk )
\sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.bin_s1  <= _203_;
always @(posedge \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.clk )
\sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.ain_s1  <= _202_;
always @(posedge \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.clk )
\sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.sum_s1  <= _205_;
always @(posedge \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.clk )
\sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.carry_s1  <= _204_;
assign _203_ = \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.ce  ? \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.bin_s0 [16:8] : \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.bin_s1 ;
assign _202_ = \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.ce  ? \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.a [16:8] : \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.ain_s1 ;
assign _204_ = \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.ce  ? \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.facout_s1  : \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.carry_s1 ;
assign _205_ = \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.ce  ? \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.fas_s1  : \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.sum_s1 ;
assign _206_ = \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.u1.a  + \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.u1.b ;
assign { \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.u1.cout , \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.u1.s  } = _206_ + \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.u1.cin ;
assign _207_ = \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.u2.a  + \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.u2.b ;
assign { \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.u2.cout , \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.u2.s  } = _207_ + \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.u2.cin ;
assign \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.bin_s0  = ~ \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.b ;
always @(posedge \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.clk )
\sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.bin_s1  <= _209_;
always @(posedge \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.clk )
\sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.ain_s1  <= _208_;
always @(posedge \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.clk )
\sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.sum_s1  <= _211_;
always @(posedge \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.clk )
\sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.carry_s1  <= _210_;
assign _209_ = \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.ce  ? \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.bin_s0 [3:2] : \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.bin_s1 ;
assign _208_ = \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.ce  ? \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.a [3:2] : \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.ain_s1 ;
assign _210_ = \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.ce  ? \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.facout_s1  : \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.carry_s1 ;
assign _211_ = \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.ce  ? \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.fas_s1  : \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.sum_s1 ;
assign _212_ = \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.u1.a  + \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.u1.b ;
assign { \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.u1.cout , \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.u1.s  } = _212_ + \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.u1.cin ;
assign _213_ = \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.u2.a  + \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.u2.b ;
assign { \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.u2.cout , \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.u2.s  } = _213_ + \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.u2.cin ;
assign ret_V_18_fu_450_p2 = { mul_ln731_reg_819[5], mul_ln731_reg_819[5], mul_ln731_reg_819, 2'h0 } | { op_0, 2'h0 };
always @(posedge ap_clk)
trunc_ln851_1_reg_851 <= 2'h0;
always @(posedge ap_clk)
shl_ln1299_reg_866 <= _036_;
always @(posedge ap_clk)
sext_ln850_reg_973 <= _035_;
always @(posedge ap_clk)
ret_V_9_reg_893 <= _032_;
always @(posedge ap_clk)
ret_V_25_reg_985 <= _027_;
always @(posedge ap_clk)
ret_V_24_reg_963 <= _026_;
always @(posedge ap_clk)
tmp_3_reg_968 <= _038_;
always @(posedge ap_clk)
ush_reg_741 <= _042_;
always @(posedge ap_clk)
ret_V_2_reg_746 <= _028_;
always @(posedge ap_clk)
ret_V_22_reg_751 <= _024_;
always @(posedge ap_clk)
ret_V_21_cast_reg_756 <= _022_;
always @(posedge ap_clk)
trunc_ln851_3_reg_763 <= _040_;
always @(posedge ap_clk)
ret_V_19_reg_903 <= _020_;
always @(posedge ap_clk)
ret_V_21_reg_908 <= _023_;
always @(posedge ap_clk)
_561_ <= _019_;
assign ret_V_18_reg_839[9:2] = _561_;
always @(posedge ap_clk)
ret_V_4_cast_reg_844 <= _029_;
always @(posedge ap_clk)
ret_V_20_reg_856 <= _021_;
always @(posedge ap_clk)
ret_V_8_reg_861 <= _031_;
always @(posedge ap_clk)
ret_V_12_reg_789 <= _017_;
always @(posedge ap_clk)
ret_V_5_reg_888 <= _030_;
always @(posedge ap_clk)
op_25_V_reg_898 <= _015_;
always @(posedge ap_clk)
op_23_V_reg_943 <= _014_;
always @(posedge ap_clk)
mul_ln728_reg_814 <= _012_;
always @(posedge ap_clk)
trunc_ln1118_reg_682 <= _039_;
always @(posedge ap_clk)
isNeg_reg_693 <= _011_;
always @(posedge ap_clk)
ret_V_reg_699 <= _033_;
always @(posedge ap_clk)
trunc_ln851_reg_706 <= _041_;
always @(posedge ap_clk)
sub_ln1367_reg_721 <= _037_;
always @(posedge ap_clk)
icmp_ln851_reg_726 <= _010_;
always @(posedge ap_clk)
r_reg_774 <= _016_;
always @(posedge ap_clk)
ret_V_17_reg_779 <= _018_;
always @(posedge ap_clk)
icmp_ln851_3_reg_784 <= _009_;
always @(posedge ap_clk)
mul_ln731_reg_819 <= _013_;
always @(posedge ap_clk)
icmp_ln851_2_reg_834 <= _008_;
always @(posedge ap_clk)
icmp_ln851_1_reg_876 <= _007_;
always @(posedge ap_clk)
sext_ln835_reg_881 <= _034_;
always @(posedge ap_clk)
ashr_ln1333_reg_871 <= _006_;
always @(posedge ap_clk)
ret_V_23_reg_804 <= _025_;
always @(posedge ap_clk)
add_ln69_4_reg_809 <= _003_;
always @(posedge ap_clk)
add_ln69_3_reg_995 <= _002_;
always @(posedge ap_clk)
add_ln69_reg_928 <= _004_;
always @(posedge ap_clk)
add_ln69_1_reg_933 <= _001_;
always @(posedge ap_clk)
add_ln691_reg_980 <= _000_;
always @(posedge ap_clk)
ap_CS_fsm <= _005_;
assign _043_ = _048_ ? 2'h2 : 2'h1;
assign _214_ = ap_CS_fsm == 1'h1;
function [24:0] _593_;
input [24:0] a;
input [624:0] b;
input [24:0] s;
case (s)
25'b0000000000000000000000001:
_593_ = b[24:0];
25'b0000000000000000000000010:
_593_ = b[49:25];
25'b0000000000000000000000100:
_593_ = b[74:50];
25'b0000000000000000000001000:
_593_ = b[99:75];
25'b0000000000000000000010000:
_593_ = b[124:100];
25'b0000000000000000000100000:
_593_ = b[149:125];
25'b0000000000000000001000000:
_593_ = b[174:150];
25'b0000000000000000010000000:
_593_ = b[199:175];
25'b0000000000000000100000000:
_593_ = b[224:200];
25'b0000000000000001000000000:
_593_ = b[249:225];
25'b0000000000000010000000000:
_593_ = b[274:250];
25'b0000000000000100000000000:
_593_ = b[299:275];
25'b0000000000001000000000000:
_593_ = b[324:300];
25'b0000000000010000000000000:
_593_ = b[349:325];
25'b0000000000100000000000000:
_593_ = b[374:350];
25'b0000000001000000000000000:
_593_ = b[399:375];
25'b0000000010000000000000000:
_593_ = b[424:400];
25'b0000000100000000000000000:
_593_ = b[449:425];
25'b0000001000000000000000000:
_593_ = b[474:450];
25'b0000010000000000000000000:
_593_ = b[499:475];
25'b0000100000000000000000000:
_593_ = b[524:500];
25'b0001000000000000000000000:
_593_ = b[549:525];
25'b0010000000000000000000000:
_593_ = b[574:550];
25'b0100000000000000000000000:
_593_ = b[599:575];
25'b1000000000000000000000000:
_593_ = b[624:600];
25'b0000000000000000000000000:
_593_ = a;
default:
_593_ = 25'bx;
endcase
endfunction
assign ap_NS_fsm = _593_(25'hxxxxxxx, { 23'h000000, _043_, 600'h000002000002000002000002000002000002000002000002000002000002000002000002000002000002000002000002000002000002000002000002000002000002000002000000000001 }, { _214_, _238_, _237_, _236_, _235_, _234_, _233_, _232_, _231_, _230_, _229_, _228_, _227_, _226_, _225_, _224_, _223_, _222_, _221_, _220_, _219_, _218_, _217_, _216_, _215_ });
assign _215_ = ap_CS_fsm == 25'h1000000;
assign _216_ = ap_CS_fsm == 24'h800000;
assign _217_ = ap_CS_fsm == 23'h400000;
assign _218_ = ap_CS_fsm == 22'h200000;
assign _219_ = ap_CS_fsm == 21'h100000;
assign _220_ = ap_CS_fsm == 20'h80000;
assign _221_ = ap_CS_fsm == 19'h40000;
assign _222_ = ap_CS_fsm == 18'h20000;
assign _223_ = ap_CS_fsm == 17'h10000;
assign _224_ = ap_CS_fsm == 16'h8000;
assign _225_ = ap_CS_fsm == 15'h4000;
assign _226_ = ap_CS_fsm == 14'h2000;
assign _227_ = ap_CS_fsm == 13'h1000;
assign _228_ = ap_CS_fsm == 12'h800;
assign _229_ = ap_CS_fsm == 11'h400;
assign _230_ = ap_CS_fsm == 10'h200;
assign _231_ = ap_CS_fsm == 9'h100;
assign _232_ = ap_CS_fsm == 8'h80;
assign _233_ = ap_CS_fsm == 7'h40;
assign _234_ = ap_CS_fsm == 6'h20;
assign _235_ = ap_CS_fsm == 5'h10;
assign _236_ = ap_CS_fsm == 4'h8;
assign _237_ = ap_CS_fsm == 3'h4;
assign _238_ = ap_CS_fsm == 2'h2;
assign op_28_ap_vld = ap_CS_fsm[24] ? 1'h1 : 1'h0;
assign ap_idle = _047_ ? 1'h1 : 1'h0;
assign _036_ = _046_ ? grp_fu_325_p2 : shl_ln1299_reg_866;
assign _035_ = ap_CS_fsm[18] ? { tmp_3_reg_968[18], tmp_3_reg_968 } : sext_ln850_reg_973;
assign _032_ = _045_ ? grp_fu_493_p2 : ret_V_9_reg_893;
assign _027_ = ap_CS_fsm[20] ? ret_V_25_fu_641_p3 : ret_V_25_reg_985;
assign _038_ = ap_CS_fsm[17] ? grp_fu_600_p2[19:1] : tmp_3_reg_968;
assign _026_ = ap_CS_fsm[17] ? grp_fu_600_p2 : ret_V_24_reg_963;
assign _040_ = ap_CS_fsm[2] ? grp_fu_297_p2[7:0] : trunc_ln851_3_reg_763;
assign _022_ = ap_CS_fsm[2] ? grp_fu_297_p2[9:8] : ret_V_21_cast_reg_756;
assign _024_ = ap_CS_fsm[2] ? grp_fu_297_p2 : ret_V_22_reg_751;
assign _028_ = ap_CS_fsm[2] ? grp_fu_276_p2 : ret_V_2_reg_746;
assign _042_ = ap_CS_fsm[2] ? ush_fu_303_p3 : ush_reg_741;
assign _023_ = ap_CS_fsm[11] ? ret_V_21_fu_549_p3 : ret_V_21_reg_908;
assign _020_ = ap_CS_fsm[11] ? ret_V_19_fu_530_p3 : ret_V_19_reg_903;
assign _031_ = ap_CS_fsm[8] ? grp_fu_415_p2[19:3] : ret_V_8_reg_861;
assign _021_ = ap_CS_fsm[8] ? grp_fu_415_p2 : ret_V_20_reg_856;
assign _029_ = ap_CS_fsm[8] ? ret_V_18_fu_450_p2[3:2] : ret_V_4_cast_reg_844;
assign _019_ = ap_CS_fsm[8] ? ret_V_18_fu_450_p2[9:2] : ret_V_18_reg_839[9:2];
assign _017_ = ap_CS_fsm[4] ? grp_fu_364_p2 : ret_V_12_reg_789;
assign _015_ = ap_CS_fsm[10] ? op_25_V_fu_512_p2 : op_25_V_reg_898;
assign _030_ = ap_CS_fsm[10] ? grp_fu_485_p2 : ret_V_5_reg_888;
assign _014_ = ap_CS_fsm[15] ? grp_fu_580_p2 : op_23_V_reg_943;
assign _012_ = ap_CS_fsm[6] ? grp_fu_201_p2 : mul_ln728_reg_814;
assign _041_ = ap_CS_fsm[0] ? 25'h0000000 : trunc_ln851_reg_706;
assign _033_ = ap_CS_fsm[0] ? { op_8[15:1], ret_V_16_fu_229_p2[25] } : ret_V_reg_699;
assign _011_ = ap_CS_fsm[0] ? op_9[3] : isNeg_reg_693;
assign _039_ = ap_CS_fsm[0] ? op_8[8:0] : trunc_ln1118_reg_682;
assign _010_ = ap_CS_fsm[1] ? icmp_ln851_fu_271_p2 : icmp_ln851_reg_726;
assign _037_ = ap_CS_fsm[1] ? grp_fu_215_p2 : sub_ln1367_reg_721;
assign _009_ = ap_CS_fsm[3] ? icmp_ln851_3_fu_359_p2 : icmp_ln851_3_reg_784;
assign _018_ = ap_CS_fsm[3] ? ret_V_17_fu_352_p3 : ret_V_17_reg_779;
assign _016_ = ap_CS_fsm[3] ? r_fu_335_p2 : r_reg_774;
assign _008_ = ap_CS_fsm[7] ? icmp_ln851_2_fu_425_p2 : icmp_ln851_2_reg_834;
assign _013_ = ap_CS_fsm[7] ? grp_fu_257_p2 : mul_ln731_reg_819;
assign _034_ = ap_CS_fsm[9] ? { ret_V_8_reg_861[16], ret_V_8_reg_861 } : sext_ln835_reg_881;
assign _007_ = ap_CS_fsm[9] ? icmp_ln851_1_fu_480_p2 : icmp_ln851_1_reg_876;
assign _006_ = _044_ ? grp_fu_330_p2 : ashr_ln1333_reg_871;
assign _003_ = ap_CS_fsm[5] ? grp_fu_375_p2 : add_ln69_4_reg_809;
assign _025_ = ap_CS_fsm[5] ? ret_V_23_fu_393_p3 : ret_V_23_reg_804;
assign _002_ = ap_CS_fsm[22] ? grp_fu_651_p2 : add_ln69_3_reg_995;
assign _001_ = ap_CS_fsm[13] ? grp_fu_571_p2 : add_ln69_1_reg_933;
assign _004_ = ap_CS_fsm[13] ? grp_fu_566_p2 : add_ln69_reg_928;
assign _000_ = ap_CS_fsm[19] ? grp_fu_619_p2 : add_ln691_reg_980;
assign _005_ = ap_rst ? 25'h0000001 : ap_NS_fsm;
assign icmp_ln851_1_fu_480_p2 = _052_ ? 1'h1 : 1'h0;
assign icmp_ln851_2_fu_425_p2 = _053_ ? 1'h1 : 1'h0;
assign icmp_ln851_3_fu_359_p2 = _054_ ? 1'h1 : 1'h0;
assign icmp_ln851_fu_271_p2 = _055_ ? 1'h1 : 1'h0;
assign op_16_V_fu_505_p3 = isNeg_reg_693 ? shl_ln1299_reg_866[0] : ashr_ln1333_reg_871[0];
assign ret_V_17_fu_352_p3 = op_8[15] ? select_ln850_fu_347_p3 : ret_V_reg_699;
assign ret_V_19_fu_530_p3 = ret_V_18_reg_839[9] ? select_ln850_1_fu_525_p3 : ret_V_4_cast_reg_844;
assign ret_V_21_fu_549_p3 = ret_V_20_reg_856[19] ? select_ln850_2_fu_544_p3 : sext_ln835_reg_881;
assign ret_V_23_fu_393_p3 = ret_V_22_reg_751[16] ? select_ln850_3_fu_388_p3 : ret_V_21_cast_reg_756;
assign ret_V_25_fu_641_p3 = ret_V_24_reg_963[19] ? select_ln850_4_fu_635_p3 : sext_ln850_reg_973;
assign select_ln850_1_fu_525_p3 = icmp_ln851_1_reg_876 ? ret_V_4_cast_reg_844 : ret_V_5_reg_888;
assign select_ln850_2_fu_544_p3 = icmp_ln851_2_reg_834 ? sext_ln835_reg_881 : ret_V_9_reg_893;
assign select_ln850_3_fu_388_p3 = icmp_ln851_3_reg_784 ? ret_V_21_cast_reg_756 : ret_V_12_reg_789;
assign select_ln850_4_fu_635_p3 = op_15[0] ? add_ln691_reg_980 : sext_ln850_reg_973;
assign select_ln850_fu_347_p3 = icmp_ln851_reg_726 ? ret_V_reg_699 : ret_V_2_reg_746;
assign ush_fu_303_p3 = isNeg_reg_693 ? sub_ln1367_reg_721 : op_9;
assign ap_CS_fsm_state1 = ap_CS_fsm[0];
assign ap_CS_fsm_state10 = ap_CS_fsm[9];
assign ap_CS_fsm_state11 = ap_CS_fsm[10];
assign ap_CS_fsm_state12 = ap_CS_fsm[11];
assign ap_CS_fsm_state13 = ap_CS_fsm[12];
assign ap_CS_fsm_state14 = ap_CS_fsm[13];
assign ap_CS_fsm_state15 = ap_CS_fsm[14];
assign ap_CS_fsm_state16 = ap_CS_fsm[15];
assign ap_CS_fsm_state17 = ap_CS_fsm[16];
assign ap_CS_fsm_state18 = ap_CS_fsm[17];
assign ap_CS_fsm_state19 = ap_CS_fsm[18];
assign ap_CS_fsm_state2 = ap_CS_fsm[1];
assign ap_CS_fsm_state20 = ap_CS_fsm[19];
assign ap_CS_fsm_state21 = ap_CS_fsm[20];
assign ap_CS_fsm_state22 = ap_CS_fsm[21];
assign ap_CS_fsm_state23 = ap_CS_fsm[22];
assign ap_CS_fsm_state24 = ap_CS_fsm[23];
assign ap_CS_fsm_state25 = ap_CS_fsm[24];
assign ap_CS_fsm_state3 = ap_CS_fsm[2];
assign ap_CS_fsm_state4 = ap_CS_fsm[3];
assign ap_CS_fsm_state5 = ap_CS_fsm[4];
assign ap_CS_fsm_state6 = ap_CS_fsm[5];
assign ap_CS_fsm_state7 = ap_CS_fsm[6];
assign ap_CS_fsm_state8 = ap_CS_fsm[7];
assign ap_CS_fsm_state9 = ap_CS_fsm[8];
assign ap_done = op_28_ap_vld;
assign ap_ready = op_28_ap_vld;
assign grp_fu_201_p1 = op_5;
assign grp_fu_201_p10 = { 12'h000, op_5 };
assign grp_fu_257_p0 = op_1[5:0];
assign grp_fu_257_p1 = op_2[5:0];
assign grp_fu_297_p0 = { 1'h0, op_2, 8'h00 };
assign grp_fu_297_p1 = { 7'h00, op_10, 8'h00 };
assign grp_fu_375_p0 = { ret_V_17_reg_779[15], ret_V_17_reg_779 };
assign grp_fu_375_p1 = { r_reg_774[3], r_reg_774[3], r_reg_774[3], r_reg_774[3], r_reg_774[3], r_reg_774[3], r_reg_774[3], r_reg_774[3], r_reg_774[3], r_reg_774[3], r_reg_774[3], r_reg_774[3], r_reg_774[3], r_reg_774 };
assign grp_fu_415_p0 = { 1'h0, mul_ln728_reg_814, 3'h0 };
assign grp_fu_415_p1 = { op_7[3], op_7[3], op_7[3], op_7[3], op_7[3], op_7[3], op_7[3], op_7[3], op_7[3], op_7[3], op_7[3], op_7[3], op_7[3], op_7[3], op_7[3], op_7[3], op_7 };
assign grp_fu_493_p0 = { ret_V_8_reg_861[16], ret_V_8_reg_861 };
assign grp_fu_566_p1 = { 16'h0000, ret_V_19_reg_903 };
assign grp_fu_571_p0 = { op_13[1], op_13[1], op_13 };
assign grp_fu_571_p1 = { 2'h0, ret_V_23_reg_804 };
assign grp_fu_580_p0 = { add_ln69_1_reg_933[3], add_ln69_1_reg_933[3], add_ln69_1_reg_933[3], add_ln69_1_reg_933[3], add_ln69_1_reg_933[3], add_ln69_1_reg_933[3], add_ln69_1_reg_933[3], add_ln69_1_reg_933[3], add_ln69_1_reg_933[3], add_ln69_1_reg_933[3], add_ln69_1_reg_933[3], add_ln69_1_reg_933[3], add_ln69_1_reg_933[3], add_ln69_1_reg_933[3], add_ln69_1_reg_933 };
assign grp_fu_600_p0 = { op_23_V_reg_943[17], op_23_V_reg_943, 1'h0 };
assign grp_fu_600_p1 = { op_15[1], op_15[1], op_15[1], op_15[1], op_15[1], op_15[1], op_15[1], op_15[1], op_15[1], op_15[1], op_15[1], op_15[1], op_15[1], op_15[1], op_15[1], op_15[1], op_15[1], op_15[1], op_15 };
assign grp_fu_619_p0 = { tmp_3_reg_968[18], tmp_3_reg_968 };
assign grp_fu_651_p0 = { 19'h00000, op_25_V_reg_898 };
assign grp_fu_659_p0 = { add_ln69_4_reg_809[16], add_ln69_4_reg_809[16], add_ln69_4_reg_809[16], add_ln69_4_reg_809 };
assign lhs_V_fu_438_p3 = { op_0, 2'h0 };
assign op_28 = { grp_fu_659_p2[19], grp_fu_659_p2[19], grp_fu_659_p2[19], grp_fu_659_p2[19], grp_fu_659_p2[19], grp_fu_659_p2[19], grp_fu_659_p2[19], grp_fu_659_p2[19], grp_fu_659_p2[19], grp_fu_659_p2[19], grp_fu_659_p2[19], grp_fu_659_p2[19], grp_fu_659_p2 };
assign op_4_V_fu_431_p3 = { mul_ln731_reg_819, 2'h0 };
assign op_6_V_fu_263_p3 = { op_2, 8'h00 };
assign p_Result_1_fu_518_p3 = ret_V_18_reg_839[9];
assign p_Result_2_fu_537_p3 = ret_V_20_reg_856[19];
assign p_Result_3_fu_381_p3 = ret_V_22_reg_751[16];
assign p_Result_4_fu_625_p3 = ret_V_24_reg_963[19];
assign p_Result_s_fu_340_p1 = op_8;
assign p_Result_s_fu_340_p3 = op_8[15];
assign ret_V_16_fu_229_p2[24:0] = 25'h0000000;
assign ret_V_16_fu_229_p2[40:26] = op_8[15:1];
assign rhs_2_fu_404_p3 = { mul_ln728_reg_814, 3'h0 };
assign rhs_3_fu_285_p3 = { op_10, 8'h00 };
assign rhs_fu_221_p1 = op_8;
assign rhs_fu_221_p3 = { op_8, 25'h0000000 };
assign sext_ln1192_1_fu_585_p0 = op_15;
assign sext_ln1192_fu_400_p0 = op_7;
assign sext_ln703_fu_446_p1 = { mul_ln731_reg_819[5], mul_ln731_reg_819[5], mul_ln731_reg_819, 2'h0 };
assign sext_ln835_fu_490_p1 = { ret_V_8_reg_861[16], ret_V_8_reg_861 };
assign sext_ln850_fu_616_p1 = { tmp_3_reg_968[18], tmp_3_reg_968 };
assign tmp_fu_589_p3 = { op_23_V_reg_943, 1'h0 };
assign trunc_ln1118_fu_193_p0 = op_8;
assign trunc_ln1118_fu_193_p1 = op_8[8:0];
assign trunc_ln1368_1_fu_502_p1 = ashr_ln1333_reg_871[0];
assign trunc_ln1368_fu_499_p1 = shl_ln1299_reg_866[0];
assign trunc_ln851_1_fu_466_p1 = ret_V_18_fu_450_p2[1:0];
assign trunc_ln851_2_fu_421_p0 = op_7;
assign trunc_ln851_2_fu_421_p1 = op_7[2:0];
assign trunc_ln851_3_fu_318_p1 = grp_fu_297_p2[7:0];
assign trunc_ln851_4_fu_632_p0 = op_15;
assign trunc_ln851_4_fu_632_p1 = op_15[0];
assign trunc_ln851_fu_245_p1 = 25'h0000000;
assign zext_ln1367_fu_322_p1 = { 5'h00, ush_reg_741 };
assign \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.ain_s0  = \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.a ;
assign \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.s  = { \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.fas_s2 , \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.sum_s1  };
assign \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.u2.a  = \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.ain_s1 ;
assign \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.u2.b  = \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.bin_s1 ;
assign \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.u2.cin  = \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.carry_s1 ;
assign \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.facout_s2  = \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.u2.cout ;
assign \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.fas_s2  = \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.u2.s ;
assign \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.u1.a  = \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.a [1:0];
assign \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.u1.b  = \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.bin_s0 [1:0];
assign \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.u1.cin  = 1'h1;
assign \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.facout_s1  = \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.u1.cout ;
assign \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.fas_s1  = \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.u1.s ;
assign \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.a  = \sub_4ns_4ns_4_2_1_U2.din0 ;
assign \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.b  = \sub_4ns_4ns_4_2_1_U2.din1 ;
assign \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.ce  = \sub_4ns_4ns_4_2_1_U2.ce ;
assign \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.clk  = \sub_4ns_4ns_4_2_1_U2.clk ;
assign \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.reset  = \sub_4ns_4ns_4_2_1_U2.reset ;
assign \sub_4ns_4ns_4_2_1_U2.dout  = \sub_4ns_4ns_4_2_1_U2.top_sub_4ns_4ns_4_2_1_Adder_0_U.s ;
assign \sub_4ns_4ns_4_2_1_U2.ce  = 1'h1;
assign \sub_4ns_4ns_4_2_1_U2.clk  = ap_clk;
assign \sub_4ns_4ns_4_2_1_U2.din0  = 4'h0;
assign \sub_4ns_4ns_4_2_1_U2.din1  = op_9;
assign grp_fu_215_p2 = \sub_4ns_4ns_4_2_1_U2.dout ;
assign \sub_4ns_4ns_4_2_1_U2.reset  = ap_rst;
assign \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.ain_s0  = \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.a ;
assign \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.s  = { \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.fas_s2 , \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.sum_s1  };
assign \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.u2.a  = \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.ain_s1 ;
assign \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.u2.b  = \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.bin_s1 ;
assign \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.u2.cin  = \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.carry_s1 ;
assign \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.facout_s2  = \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.u2.cout ;
assign \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.fas_s2  = \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.u2.s ;
assign \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.u1.a  = \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.a [7:0];
assign \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.u1.b  = \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.bin_s0 [7:0];
assign \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.u1.cin  = 1'h1;
assign \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.facout_s1  = \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.u1.cout ;
assign \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.fas_s1  = \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.u1.s ;
assign \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.a  = \sub_17ns_17ns_17_2_1_U5.din0 ;
assign \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.b  = \sub_17ns_17ns_17_2_1_U5.din1 ;
assign \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.ce  = \sub_17ns_17ns_17_2_1_U5.ce ;
assign \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.clk  = \sub_17ns_17ns_17_2_1_U5.clk ;
assign \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.reset  = \sub_17ns_17ns_17_2_1_U5.reset ;
assign \sub_17ns_17ns_17_2_1_U5.dout  = \sub_17ns_17ns_17_2_1_U5.top_sub_17ns_17ns_17_2_1_Adder_2_U.s ;
assign \sub_17ns_17ns_17_2_1_U5.ce  = 1'h1;
assign \sub_17ns_17ns_17_2_1_U5.clk  = ap_clk;
assign \sub_17ns_17ns_17_2_1_U5.din0  = { 1'h0, op_2, 8'h00 };
assign \sub_17ns_17ns_17_2_1_U5.din1  = { 7'h00, op_10, 8'h00 };
assign grp_fu_297_p2 = \sub_17ns_17ns_17_2_1_U5.dout ;
assign \sub_17ns_17ns_17_2_1_U5.reset  = ap_rst;
assign \shl_9ns_4ns_9_7_1_U6.din1_cast  = \shl_9ns_4ns_9_7_1_U6.din1 [3:0];
assign \shl_9ns_4ns_9_7_1_U6.din1_mask  = 4'h1;
assign \shl_9ns_4ns_9_7_1_U6.ce  = 1'h1;
assign \shl_9ns_4ns_9_7_1_U6.clk  = ap_clk;
assign \shl_9ns_4ns_9_7_1_U6.din0  = trunc_ln1118_reg_682;
assign \shl_9ns_4ns_9_7_1_U6.din1  = { 5'h00, ush_reg_741 };
assign grp_fu_325_p2 = \shl_9ns_4ns_9_7_1_U6.dout ;
assign \shl_9ns_4ns_9_7_1_U6.reset  = ap_rst;
assign \mul_6s_6s_6_7_1_U3.top_mul_6s_6s_6_7_1_Mul_DSP_1_U.p  = \mul_6s_6s_6_7_1_U3.top_mul_6s_6s_6_7_1_Mul_DSP_1_U.buff4 ;
assign \mul_6s_6s_6_7_1_U3.top_mul_6s_6s_6_7_1_Mul_DSP_1_U.a  = \mul_6s_6s_6_7_1_U3.din0 ;
assign \mul_6s_6s_6_7_1_U3.top_mul_6s_6s_6_7_1_Mul_DSP_1_U.b  = \mul_6s_6s_6_7_1_U3.din1 ;
assign \mul_6s_6s_6_7_1_U3.top_mul_6s_6s_6_7_1_Mul_DSP_1_U.ce  = \mul_6s_6s_6_7_1_U3.ce ;
assign \mul_6s_6s_6_7_1_U3.top_mul_6s_6s_6_7_1_Mul_DSP_1_U.clk  = \mul_6s_6s_6_7_1_U3.clk ;
assign \mul_6s_6s_6_7_1_U3.dout  = \mul_6s_6s_6_7_1_U3.top_mul_6s_6s_6_7_1_Mul_DSP_1_U.p ;
assign \mul_6s_6s_6_7_1_U3.ce  = 1'h1;
assign \mul_6s_6s_6_7_1_U3.clk  = ap_clk;
assign \mul_6s_6s_6_7_1_U3.din0  = op_1[5:0];
assign \mul_6s_6s_6_7_1_U3.din1  = op_2[5:0];
assign grp_fu_257_p2 = \mul_6s_6s_6_7_1_U3.dout ;
assign \mul_6s_6s_6_7_1_U3.reset  = ap_rst;
assign \mul_16s_4ns_16_7_1_U1.top_mul_16s_4ns_16_7_1_Mul_DSP_0_U.p  = \mul_16s_4ns_16_7_1_U1.top_mul_16s_4ns_16_7_1_Mul_DSP_0_U.buff4 ;
assign \mul_16s_4ns_16_7_1_U1.top_mul_16s_4ns_16_7_1_Mul_DSP_0_U.a  = \mul_16s_4ns_16_7_1_U1.din0 ;
assign \mul_16s_4ns_16_7_1_U1.top_mul_16s_4ns_16_7_1_Mul_DSP_0_U.b  = \mul_16s_4ns_16_7_1_U1.din1 ;
assign \mul_16s_4ns_16_7_1_U1.top_mul_16s_4ns_16_7_1_Mul_DSP_0_U.ce  = \mul_16s_4ns_16_7_1_U1.ce ;
assign \mul_16s_4ns_16_7_1_U1.top_mul_16s_4ns_16_7_1_Mul_DSP_0_U.clk  = \mul_16s_4ns_16_7_1_U1.clk ;
assign \mul_16s_4ns_16_7_1_U1.dout  = \mul_16s_4ns_16_7_1_U1.top_mul_16s_4ns_16_7_1_Mul_DSP_0_U.p ;
assign \mul_16s_4ns_16_7_1_U1.ce  = 1'h1;
assign \mul_16s_4ns_16_7_1_U1.clk  = ap_clk;
assign \mul_16s_4ns_16_7_1_U1.din0  = op_8;
assign \mul_16s_4ns_16_7_1_U1.din1  = op_5;
assign grp_fu_201_p2 = \mul_16s_4ns_16_7_1_U1.dout ;
assign \mul_16s_4ns_16_7_1_U1.reset  = ap_rst;
assign \ashr_9ns_4ns_9_7_1_U7.din1_cast  = \ashr_9ns_4ns_9_7_1_U7.din1 [3:0];
assign \ashr_9ns_4ns_9_7_1_U7.din1_mask  = 4'h1;
assign \ashr_9ns_4ns_9_7_1_U7.ce  = 1'h1;
assign \ashr_9ns_4ns_9_7_1_U7.clk  = ap_clk;
assign \ashr_9ns_4ns_9_7_1_U7.din0  = trunc_ln1118_reg_682;
assign \ashr_9ns_4ns_9_7_1_U7.din1  = { 5'h00, ush_reg_741 };
assign grp_fu_330_p2 = \ashr_9ns_4ns_9_7_1_U7.dout ;
assign \ashr_9ns_4ns_9_7_1_U7.reset  = ap_rst;
assign \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.ain_s0  = \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.a ;
assign \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.bin_s0  = \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.b ;
assign \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.s  = { \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.fas_s2 , \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.sum_s1  };
assign \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.u2.a  = \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.ain_s1 ;
assign \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.u2.b  = \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.bin_s1 ;
assign \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.u2.cin  = \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.carry_s1 ;
assign \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.facout_s2  = \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.u2.cout ;
assign \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.fas_s2  = \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.u2.s ;
assign \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.u1.a  = \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.a [1:0];
assign \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.u1.b  = \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.b [1:0];
assign \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.u1.cin  = 1'h0;
assign \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.facout_s1  = \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.u1.cout ;
assign \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.fas_s1  = \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.u1.s ;
assign \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.a  = \add_4s_4ns_4_2_1_U14.din0 ;
assign \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.b  = \add_4s_4ns_4_2_1_U14.din1 ;
assign \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.ce  = \add_4s_4ns_4_2_1_U14.ce ;
assign \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.clk  = \add_4s_4ns_4_2_1_U14.clk ;
assign \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.reset  = \add_4s_4ns_4_2_1_U14.reset ;
assign \add_4s_4ns_4_2_1_U14.dout  = \add_4s_4ns_4_2_1_U14.top_add_4s_4ns_4_2_1_Adder_8_U.s ;
assign \add_4s_4ns_4_2_1_U14.ce  = 1'h1;
assign \add_4s_4ns_4_2_1_U14.clk  = ap_clk;
assign \add_4s_4ns_4_2_1_U14.din0  = { op_13[1], op_13[1], op_13 };
assign \add_4s_4ns_4_2_1_U14.din1  = { 2'h0, ret_V_23_reg_804 };
assign grp_fu_571_p2 = \add_4s_4ns_4_2_1_U14.dout ;
assign \add_4s_4ns_4_2_1_U14.reset  = ap_rst;
assign \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.ain_s0  = \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.a ;
assign \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.bin_s0  = \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.b ;
assign \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.s  = { \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.fas_s2 , \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.sum_s1  };
assign \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.u2.a  = \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.ain_s1 ;
assign \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.u2.b  = \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.bin_s1 ;
assign \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.u2.cin  = \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.carry_s1 ;
assign \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.facout_s2  = \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.u2.cout ;
assign \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.fas_s2  = \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.u2.s ;
assign \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.u1.a  = \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.a [0];
assign \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.u1.b  = \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.b [0];
assign \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.u1.cin  = 1'h0;
assign \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.facout_s1  = \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.u1.cout ;
assign \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.fas_s1  = \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.u1.s ;
assign \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.a  = \add_2ns_2ns_2_2_1_U8.din0 ;
assign \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.b  = \add_2ns_2ns_2_2_1_U8.din1 ;
assign \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.ce  = \add_2ns_2ns_2_2_1_U8.ce ;
assign \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.clk  = \add_2ns_2ns_2_2_1_U8.clk ;
assign \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.reset  = \add_2ns_2ns_2_2_1_U8.reset ;
assign \add_2ns_2ns_2_2_1_U8.dout  = \add_2ns_2ns_2_2_1_U8.top_add_2ns_2ns_2_2_1_Adder_3_U.s ;
assign \add_2ns_2ns_2_2_1_U8.ce  = 1'h1;
assign \add_2ns_2ns_2_2_1_U8.clk  = ap_clk;
assign \add_2ns_2ns_2_2_1_U8.din0  = ret_V_21_cast_reg_756;
assign \add_2ns_2ns_2_2_1_U8.din1  = 2'h1;
assign grp_fu_364_p2 = \add_2ns_2ns_2_2_1_U8.dout ;
assign \add_2ns_2ns_2_2_1_U8.reset  = ap_rst;
assign \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.ain_s0  = \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.a ;
assign \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.bin_s0  = \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.b ;
assign \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.s  = { \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.fas_s2 , \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.sum_s1  };
assign \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.u2.a  = \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.ain_s1 ;
assign \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.u2.b  = \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.bin_s1 ;
assign \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.u2.cin  = \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.carry_s1 ;
assign \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.facout_s2  = \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.u2.cout ;
assign \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.fas_s2  = \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.u2.s ;
assign \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.u1.a  = \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.a [0];
assign \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.u1.b  = \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.b [0];
assign \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.u1.cin  = 1'h0;
assign \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.facout_s1  = \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.u1.cout ;
assign \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.fas_s1  = \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.u1.s ;
assign \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.a  = \add_2ns_2ns_2_2_1_U11.din0 ;
assign \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.b  = \add_2ns_2ns_2_2_1_U11.din1 ;
assign \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.ce  = \add_2ns_2ns_2_2_1_U11.ce ;
assign \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.clk  = \add_2ns_2ns_2_2_1_U11.clk ;
assign \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.reset  = \add_2ns_2ns_2_2_1_U11.reset ;
assign \add_2ns_2ns_2_2_1_U11.dout  = \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_3_U.s ;
assign \add_2ns_2ns_2_2_1_U11.ce  = 1'h1;
assign \add_2ns_2ns_2_2_1_U11.clk  = ap_clk;
assign \add_2ns_2ns_2_2_1_U11.din0  = ret_V_4_cast_reg_844;
assign \add_2ns_2ns_2_2_1_U11.din1  = 2'h1;
assign grp_fu_485_p2 = \add_2ns_2ns_2_2_1_U11.dout ;
assign \add_2ns_2ns_2_2_1_U11.reset  = ap_rst;
assign \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.ain_s0  = \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.a ;
assign \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.bin_s0  = \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.b ;
assign \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.s  = { \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.fas_s2 , \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.sum_s1  };
assign \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.u2.a  = \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.ain_s1 ;
assign \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.u2.b  = \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.bin_s1 ;
assign \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.u2.cin  = \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.carry_s1 ;
assign \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.facout_s2  = \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.u2.cout ;
assign \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.fas_s2  = \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.u2.s ;
assign \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.u1.a  = \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.a [9:0];
assign \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.u1.b  = \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.b [9:0];
assign \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.u1.cin  = 1'h0;
assign \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.facout_s1  = \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.u1.cout ;
assign \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.fas_s1  = \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.u1.s ;
assign \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.a  = \add_20s_20s_20_2_1_U16.din0 ;
assign \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.b  = \add_20s_20s_20_2_1_U16.din1 ;
assign \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.ce  = \add_20s_20s_20_2_1_U16.ce ;
assign \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.clk  = \add_20s_20s_20_2_1_U16.clk ;
assign \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.reset  = \add_20s_20s_20_2_1_U16.reset ;
assign \add_20s_20s_20_2_1_U16.dout  = \add_20s_20s_20_2_1_U16.top_add_20s_20s_20_2_1_Adder_9_U.s ;
assign \add_20s_20s_20_2_1_U16.ce  = 1'h1;
assign \add_20s_20s_20_2_1_U16.clk  = ap_clk;
assign \add_20s_20s_20_2_1_U16.din0  = { op_23_V_reg_943[17], op_23_V_reg_943, 1'h0 };
assign \add_20s_20s_20_2_1_U16.din1  = { op_15[1], op_15[1], op_15[1], op_15[1], op_15[1], op_15[1], op_15[1], op_15[1], op_15[1], op_15[1], op_15[1], op_15[1], op_15[1], op_15[1], op_15[1], op_15[1], op_15[1], op_15[1], op_15 };
assign grp_fu_600_p2 = \add_20s_20s_20_2_1_U16.dout ;
assign \add_20s_20s_20_2_1_U16.reset  = ap_rst;
assign \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.ain_s0  = \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.a ;
assign \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.bin_s0  = \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.b ;
assign \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.s  = { \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.fas_s2 , \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.sum_s1  };
assign \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.u2.a  = \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.ain_s1 ;
assign \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.u2.b  = \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.bin_s1 ;
assign \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.u2.cin  = \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.carry_s1 ;
assign \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.facout_s2  = \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.u2.cout ;
assign \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.fas_s2  = \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.u2.s ;
assign \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.u1.a  = \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.a [9:0];
assign \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.u1.b  = \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.b [9:0];
assign \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.u1.cin  = 1'h0;
assign \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.facout_s1  = \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.u1.cout ;
assign \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.fas_s1  = \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.u1.s ;
assign \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.a  = \add_20s_20ns_20_2_1_U19.din0 ;
assign \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.b  = \add_20s_20ns_20_2_1_U19.din1 ;
assign \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.ce  = \add_20s_20ns_20_2_1_U19.ce ;
assign \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.clk  = \add_20s_20ns_20_2_1_U19.clk ;
assign \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.reset  = \add_20s_20ns_20_2_1_U19.reset ;
assign \add_20s_20ns_20_2_1_U19.dout  = \add_20s_20ns_20_2_1_U19.top_add_20s_20ns_20_2_1_Adder_10_U.s ;
assign \add_20s_20ns_20_2_1_U19.ce  = 1'h1;
assign \add_20s_20ns_20_2_1_U19.clk  = ap_clk;
assign \add_20s_20ns_20_2_1_U19.din0  = { add_ln69_4_reg_809[16], add_ln69_4_reg_809[16], add_ln69_4_reg_809[16], add_ln69_4_reg_809 };
assign \add_20s_20ns_20_2_1_U19.din1  = add_ln69_3_reg_995;
assign grp_fu_659_p2 = \add_20s_20ns_20_2_1_U19.dout ;
assign \add_20s_20ns_20_2_1_U19.reset  = ap_rst;
assign \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.ain_s0  = \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.a ;
assign \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.bin_s0  = \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.b ;
assign \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.s  = { \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.fas_s2 , \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.sum_s1  };
assign \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.u2.a  = \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.ain_s1 ;
assign \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.u2.b  = \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.bin_s1 ;
assign \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.u2.cin  = \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.carry_s1 ;
assign \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.facout_s2  = \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.u2.cout ;
assign \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.fas_s2  = \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.u2.s ;
assign \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.u1.a  = \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.a [9:0];
assign \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.u1.b  = \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.b [9:0];
assign \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.u1.cin  = 1'h0;
assign \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.facout_s1  = \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.u1.cout ;
assign \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.fas_s1  = \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.u1.s ;
assign \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.a  = \add_20s_20ns_20_2_1_U17.din0 ;
assign \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.b  = \add_20s_20ns_20_2_1_U17.din1 ;
assign \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.ce  = \add_20s_20ns_20_2_1_U17.ce ;
assign \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.clk  = \add_20s_20ns_20_2_1_U17.clk ;
assign \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.reset  = \add_20s_20ns_20_2_1_U17.reset ;
assign \add_20s_20ns_20_2_1_U17.dout  = \add_20s_20ns_20_2_1_U17.top_add_20s_20ns_20_2_1_Adder_10_U.s ;
assign \add_20s_20ns_20_2_1_U17.ce  = 1'h1;
assign \add_20s_20ns_20_2_1_U17.clk  = ap_clk;
assign \add_20s_20ns_20_2_1_U17.din0  = { tmp_3_reg_968[18], tmp_3_reg_968 };
assign \add_20s_20ns_20_2_1_U17.din1  = 20'h00001;
assign grp_fu_619_p2 = \add_20s_20ns_20_2_1_U17.dout ;
assign \add_20s_20ns_20_2_1_U17.reset  = ap_rst;
assign \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.ain_s0  = \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.a ;
assign \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.bin_s0  = \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.b ;
assign \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.s  = { \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.fas_s2 , \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.sum_s1  };
assign \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.u2.a  = \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.ain_s1 ;
assign \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.u2.b  = \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.bin_s1 ;
assign \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.u2.cin  = \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.carry_s1 ;
assign \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.facout_s2  = \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.u2.cout ;
assign \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.fas_s2  = \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.u2.s ;
assign \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.u1.a  = \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.a [9:0];
assign \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.u1.b  = \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.b [9:0];
assign \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.u1.cin  = 1'h0;
assign \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.facout_s1  = \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.u1.cout ;
assign \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.fas_s1  = \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.u1.s ;
assign \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.a  = \add_20ns_20s_20_2_1_U10.din0 ;
assign \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.b  = \add_20ns_20s_20_2_1_U10.din1 ;
assign \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.ce  = \add_20ns_20s_20_2_1_U10.ce ;
assign \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.clk  = \add_20ns_20s_20_2_1_U10.clk ;
assign \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.reset  = \add_20ns_20s_20_2_1_U10.reset ;
assign \add_20ns_20s_20_2_1_U10.dout  = \add_20ns_20s_20_2_1_U10.top_add_20ns_20s_20_2_1_Adder_5_U.s ;
assign \add_20ns_20s_20_2_1_U10.ce  = 1'h1;
assign \add_20ns_20s_20_2_1_U10.clk  = ap_clk;
assign \add_20ns_20s_20_2_1_U10.din0  = { 1'h0, mul_ln728_reg_814, 3'h0 };
assign \add_20ns_20s_20_2_1_U10.din1  = { op_7[3], op_7[3], op_7[3], op_7[3], op_7[3], op_7[3], op_7[3], op_7[3], op_7[3], op_7[3], op_7[3], op_7[3], op_7[3], op_7[3], op_7[3], op_7[3], op_7 };
assign grp_fu_415_p2 = \add_20ns_20s_20_2_1_U10.dout ;
assign \add_20ns_20s_20_2_1_U10.reset  = ap_rst;
assign \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.ain_s0  = \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.a ;
assign \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.bin_s0  = \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.b ;
assign \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.s  = { \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.fas_s2 , \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.sum_s1  };
assign \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.u2.a  = \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.ain_s1 ;
assign \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.u2.b  = \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.bin_s1 ;
assign \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.u2.cin  = \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.carry_s1 ;
assign \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.facout_s2  = \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.u2.cout ;
assign \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.fas_s2  = \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.u2.s ;
assign \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.u1.a  = \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.a [9:0];
assign \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.u1.b  = \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.b [9:0];
assign \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.u1.cin  = 1'h0;
assign \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.facout_s1  = \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.u1.cout ;
assign \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.fas_s1  = \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.u1.s ;
assign \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.a  = \add_20ns_20ns_20_2_1_U18.din0 ;
assign \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.b  = \add_20ns_20ns_20_2_1_U18.din1 ;
assign \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.ce  = \add_20ns_20ns_20_2_1_U18.ce ;
assign \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.clk  = \add_20ns_20ns_20_2_1_U18.clk ;
assign \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.reset  = \add_20ns_20ns_20_2_1_U18.reset ;
assign \add_20ns_20ns_20_2_1_U18.dout  = \add_20ns_20ns_20_2_1_U18.top_add_20ns_20ns_20_2_1_Adder_11_U.s ;
assign \add_20ns_20ns_20_2_1_U18.ce  = 1'h1;
assign \add_20ns_20ns_20_2_1_U18.clk  = ap_clk;
assign \add_20ns_20ns_20_2_1_U18.din0  = { 19'h00000, op_25_V_reg_898 };
assign \add_20ns_20ns_20_2_1_U18.din1  = ret_V_25_reg_985;
assign grp_fu_651_p2 = \add_20ns_20ns_20_2_1_U18.dout ;
assign \add_20ns_20ns_20_2_1_U18.reset  = ap_rst;
assign \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.ain_s0  = \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.a ;
assign \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.bin_s0  = \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.b ;
assign \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.s  = { \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.fas_s2 , \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.sum_s1  };
assign \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.u2.a  = \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.ain_s1 ;
assign \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.u2.b  = \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.bin_s1 ;
assign \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.u2.cin  = \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.carry_s1 ;
assign \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.facout_s2  = \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.u2.cout ;
assign \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.fas_s2  = \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.u2.s ;
assign \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.u1.a  = \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.a [8:0];
assign \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.u1.b  = \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.b [8:0];
assign \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.u1.cin  = 1'h0;
assign \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.facout_s1  = \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.u1.cout ;
assign \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.fas_s1  = \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.u1.s ;
assign \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.a  = \add_18s_18ns_18_2_1_U15.din0 ;
assign \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.b  = \add_18s_18ns_18_2_1_U15.din1 ;
assign \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.ce  = \add_18s_18ns_18_2_1_U15.ce ;
assign \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.clk  = \add_18s_18ns_18_2_1_U15.clk ;
assign \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.reset  = \add_18s_18ns_18_2_1_U15.reset ;
assign \add_18s_18ns_18_2_1_U15.dout  = \add_18s_18ns_18_2_1_U15.top_add_18s_18ns_18_2_1_Adder_6_U.s ;
assign \add_18s_18ns_18_2_1_U15.ce  = 1'h1;
assign \add_18s_18ns_18_2_1_U15.clk  = ap_clk;
assign \add_18s_18ns_18_2_1_U15.din0  = { add_ln69_1_reg_933[3], add_ln69_1_reg_933[3], add_ln69_1_reg_933[3], add_ln69_1_reg_933[3], add_ln69_1_reg_933[3], add_ln69_1_reg_933[3], add_ln69_1_reg_933[3], add_ln69_1_reg_933[3], add_ln69_1_reg_933[3], add_ln69_1_reg_933[3], add_ln69_1_reg_933[3], add_ln69_1_reg_933[3], add_ln69_1_reg_933[3], add_ln69_1_reg_933[3], add_ln69_1_reg_933 };
assign \add_18s_18ns_18_2_1_U15.din1  = add_ln69_reg_928;
assign grp_fu_580_p2 = \add_18s_18ns_18_2_1_U15.dout ;
assign \add_18s_18ns_18_2_1_U15.reset  = ap_rst;
assign \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.ain_s0  = \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.a ;
assign \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.bin_s0  = \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.b ;
assign \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.s  = { \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.fas_s2 , \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.sum_s1  };
assign \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.u2.a  = \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.ain_s1 ;
assign \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.u2.b  = \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.bin_s1 ;
assign \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.u2.cin  = \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.carry_s1 ;
assign \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.facout_s2  = \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.u2.cout ;
assign \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.fas_s2  = \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.u2.s ;
assign \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.u1.a  = \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.a [8:0];
assign \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.u1.b  = \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.b [8:0];
assign \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.u1.cin  = 1'h0;
assign \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.facout_s1  = \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.u1.cout ;
assign \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.fas_s1  = \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.u1.s ;
assign \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.a  = \add_18s_18ns_18_2_1_U12.din0 ;
assign \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.b  = \add_18s_18ns_18_2_1_U12.din1 ;
assign \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.ce  = \add_18s_18ns_18_2_1_U12.ce ;
assign \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.clk  = \add_18s_18ns_18_2_1_U12.clk ;
assign \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.reset  = \add_18s_18ns_18_2_1_U12.reset ;
assign \add_18s_18ns_18_2_1_U12.dout  = \add_18s_18ns_18_2_1_U12.top_add_18s_18ns_18_2_1_Adder_6_U.s ;
assign \add_18s_18ns_18_2_1_U12.ce  = 1'h1;
assign \add_18s_18ns_18_2_1_U12.clk  = ap_clk;
assign \add_18s_18ns_18_2_1_U12.din0  = { ret_V_8_reg_861[16], ret_V_8_reg_861 };
assign \add_18s_18ns_18_2_1_U12.din1  = 18'h00001;
assign grp_fu_493_p2 = \add_18s_18ns_18_2_1_U12.dout ;
assign \add_18s_18ns_18_2_1_U12.reset  = ap_rst;
assign \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.ain_s0  = \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.a ;
assign \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.bin_s0  = \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.b ;
assign \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.s  = { \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.fas_s2 , \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.sum_s1  };
assign \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.u2.a  = \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.ain_s1 ;
assign \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.u2.b  = \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.bin_s1 ;
assign \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.u2.cin  = \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.carry_s1 ;
assign \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.facout_s2  = \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.u2.cout ;
assign \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.fas_s2  = \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.u2.s ;
assign \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.u1.a  = \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.a [8:0];
assign \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.u1.b  = \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.b [8:0];
assign \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.u1.cin  = 1'h0;
assign \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.facout_s1  = \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.u1.cout ;
assign \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.fas_s1  = \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.u1.s ;
assign \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.a  = \add_18ns_18ns_18_2_1_U13.din0 ;
assign \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.b  = \add_18ns_18ns_18_2_1_U13.din1 ;
assign \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.ce  = \add_18ns_18ns_18_2_1_U13.ce ;
assign \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.clk  = \add_18ns_18ns_18_2_1_U13.clk ;
assign \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.reset  = \add_18ns_18ns_18_2_1_U13.reset ;
assign \add_18ns_18ns_18_2_1_U13.dout  = \add_18ns_18ns_18_2_1_U13.top_add_18ns_18ns_18_2_1_Adder_7_U.s ;
assign \add_18ns_18ns_18_2_1_U13.ce  = 1'h1;
assign \add_18ns_18ns_18_2_1_U13.clk  = ap_clk;
assign \add_18ns_18ns_18_2_1_U13.din0  = ret_V_21_reg_908;
assign \add_18ns_18ns_18_2_1_U13.din1  = { 16'h0000, ret_V_19_reg_903 };
assign grp_fu_566_p2 = \add_18ns_18ns_18_2_1_U13.dout ;
assign \add_18ns_18ns_18_2_1_U13.reset  = ap_rst;
assign \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.ain_s0  = \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.a ;
assign \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.bin_s0  = \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.b ;
assign \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.s  = { \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.fas_s2 , \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.sum_s1  };
assign \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.u2.a  = \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.ain_s1 ;
assign \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.u2.b  = \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.bin_s1 ;
assign \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.u2.cin  = \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.carry_s1 ;
assign \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.facout_s2  = \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.u2.cout ;
assign \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.fas_s2  = \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.u2.s ;
assign \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.u1.a  = \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.a [7:0];
assign \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.u1.b  = \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.b [7:0];
assign \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.u1.cin  = 1'h0;
assign \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.facout_s1  = \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.u1.cout ;
assign \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.fas_s1  = \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.u1.s ;
assign \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.a  = \add_17s_17s_17_2_1_U9.din0 ;
assign \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.b  = \add_17s_17s_17_2_1_U9.din1 ;
assign \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.ce  = \add_17s_17s_17_2_1_U9.ce ;
assign \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.clk  = \add_17s_17s_17_2_1_U9.clk ;
assign \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.reset  = \add_17s_17s_17_2_1_U9.reset ;
assign \add_17s_17s_17_2_1_U9.dout  = \add_17s_17s_17_2_1_U9.top_add_17s_17s_17_2_1_Adder_4_U.s ;
assign \add_17s_17s_17_2_1_U9.ce  = 1'h1;
assign \add_17s_17s_17_2_1_U9.clk  = ap_clk;
assign \add_17s_17s_17_2_1_U9.din0  = { ret_V_17_reg_779[15], ret_V_17_reg_779 };
assign \add_17s_17s_17_2_1_U9.din1  = { r_reg_774[3], r_reg_774[3], r_reg_774[3], r_reg_774[3], r_reg_774[3], r_reg_774[3], r_reg_774[3], r_reg_774[3], r_reg_774[3], r_reg_774[3], r_reg_774[3], r_reg_774[3], r_reg_774[3], r_reg_774 };
assign grp_fu_375_p2 = \add_17s_17s_17_2_1_U9.dout ;
assign \add_17s_17s_17_2_1_U9.reset  = ap_rst;
assign \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.ain_s0  = \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.a ;
assign \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.bin_s0  = \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.b ;
assign \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.s  = { \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.fas_s2 , \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.sum_s1  };
assign \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.u2.a  = \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.ain_s1 ;
assign \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.u2.b  = \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.bin_s1 ;
assign \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.u2.cin  = \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.carry_s1 ;
assign \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.facout_s2  = \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.u2.cout ;
assign \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.fas_s2  = \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.u2.s ;
assign \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.u1.a  = \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.a [7:0];
assign \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.u1.b  = \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.b [7:0];
assign \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.u1.cin  = 1'h0;
assign \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.facout_s1  = \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.u1.cout ;
assign \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.fas_s1  = \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.u1.s ;
assign \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.a  = \add_16ns_16ns_16_2_1_U4.din0 ;
assign \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.b  = \add_16ns_16ns_16_2_1_U4.din1 ;
assign \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.ce  = \add_16ns_16ns_16_2_1_U4.ce ;
assign \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.clk  = \add_16ns_16ns_16_2_1_U4.clk ;
assign \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.reset  = \add_16ns_16ns_16_2_1_U4.reset ;
assign \add_16ns_16ns_16_2_1_U4.dout  = \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_1_U.s ;
assign \add_16ns_16ns_16_2_1_U4.ce  = 1'h1;
assign \add_16ns_16ns_16_2_1_U4.clk  = ap_clk;
assign \add_16ns_16ns_16_2_1_U4.din0  = ret_V_reg_699;
assign \add_16ns_16ns_16_2_1_U4.din1  = 16'h0001;
assign grp_fu_276_p2 = \add_16ns_16ns_16_2_1_U4.dout ;
assign \add_16ns_16ns_16_2_1_U4.reset  = ap_rst;
endmodule


// Product machine:
module top_A_times_top_B (ap_start, op_0, op_1, op_10, op_13, op_15, op_2, op_5, op_7, op_8, op_9, ap_clk, unsafe_signal);
input ap_start;
input [7:0] op_0;
input [15:0] op_1;
input [1:0] op_10;
input [1:0] op_13;
input [1:0] op_15;
input [7:0] op_2;
input [3:0] op_5;
input [3:0] op_7;
input [15:0] op_8;
input [3:0] op_9;
input ap_clk;
output unsafe_signal;
reg _setup;
initial _setup = 1'b0;
always @ (posedge ap_clk) _setup <= 1'b1;
reg ap_start_internal;
always @ (posedge ap_clk) if (!_setup) ap_start_internal <= ap_start;
reg [7:0] op_0_internal;
always @ (posedge ap_clk) if (!_setup) op_0_internal <= op_0;
reg [15:0] op_1_internal;
always @ (posedge ap_clk) if (!_setup) op_1_internal <= op_1;
reg [1:0] op_10_internal;
always @ (posedge ap_clk) if (!_setup) op_10_internal <= op_10;
reg [1:0] op_13_internal;
always @ (posedge ap_clk) if (!_setup) op_13_internal <= op_13;
reg [1:0] op_15_internal;
always @ (posedge ap_clk) if (!_setup) op_15_internal <= op_15;
reg [7:0] op_2_internal;
always @ (posedge ap_clk) if (!_setup) op_2_internal <= op_2;
reg [3:0] op_5_internal;
always @ (posedge ap_clk) if (!_setup) op_5_internal <= op_5;
reg [3:0] op_7_internal;
always @ (posedge ap_clk) if (!_setup) op_7_internal <= op_7;
reg [15:0] op_8_internal;
always @ (posedge ap_clk) if (!_setup) op_8_internal <= op_8;
reg [3:0] op_9_internal;
always @ (posedge ap_clk) if (!_setup) op_9_internal <= op_9;
wire ap_done_A;
wire ap_done_B;
wire ap_done_eq;
assign ap_done_eq = ap_done_A == ap_done_B;
wire ap_idle_A;
wire ap_idle_B;
wire ap_idle_eq;
assign ap_idle_eq = ap_idle_A == ap_idle_B;
wire ap_ready_A;
wire ap_ready_B;
wire ap_ready_eq;
assign ap_ready_eq = ap_ready_A == ap_ready_B;
wire [31:0] op_28_A;
wire [31:0] op_28_B;
wire op_28_eq;
assign op_28_eq = op_28_A == op_28_B;
wire op_28_ap_vld_A;
wire op_28_ap_vld_B;
wire clk_enable_A;
wire clk_enable_B;
assign clk_enable_A = _setup & (~op_28_ap_vld_A | op_28_ap_vld_B);
assign clk_enable_B = _setup;
wire divergent;
assign divergent = ~(ap_done_eq & ap_idle_eq & ap_ready_eq & op_28_eq);
assign unsafe_signal = op_28_ap_vld_A & op_28_ap_vld_B & divergent;
top_A instance_A (
    .ap_clk(ap_clk),
    .clk_enable(clk_enable_A),
    .ap_start(ap_start_internal),
    .op_0(op_0_internal),
    .op_1(op_1_internal),
    .op_10(op_10_internal),
    .op_13(op_13_internal),
    .op_15(op_15_internal),
    .op_2(op_2_internal),
    .op_5(op_5_internal),
    .op_7(op_7_internal),
    .op_8(op_8_internal),
    .op_9(op_9_internal),
    .ap_done(ap_done_A),
    .ap_idle(ap_idle_A),
    .ap_ready(ap_ready_A),
    .op_28(op_28_A),
    .op_28_ap_vld(op_28_ap_vld_A)
);
top_B instance_B (
    .ap_clk(ap_clk),
    .clk_enable(clk_enable_B),
    .ap_start(ap_start_internal),
    .op_0(op_0_internal),
    .op_1(op_1_internal),
    .op_10(op_10_internal),
    .op_13(op_13_internal),
    .op_15(op_15_internal),
    .op_2(op_2_internal),
    .op_5(op_5_internal),
    .op_7(op_7_internal),
    .op_8(op_8_internal),
    .op_9(op_9_internal),
    .ap_done(ap_done_B),
    .ap_idle(ap_idle_B),
    .ap_ready(ap_ready_B),
    .op_28(op_28_B),
    .op_28_ap_vld(op_28_ap_vld_B)
);
endmodule
