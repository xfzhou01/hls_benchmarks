// Processed by function `construct_kairos` in `verilog_tricks.py`.
// Machine A:
// Processed by function `add_clk_enable_signal` in `verilog_tricks.py`.
// Processed by function `remove_reset_signal` in `verilog_tricks.py`.
module top_A (
  ap_clk,
  ap_start,
  ap_done,
  ap_idle,
  ap_ready,
  op_0,
  op_2,
  op_3,
  op_5,
  op_10,
  op_11,
  op_12,
  op_13,
  op_14,
  op_15,
  op_17,
  op_18,
  op_19,
  op_31,
  op_31_ap_vld,
clk_enable
);
input clk_enable;


input ap_clk;
wire ap_rst;
assign ap_rst = op_31_ap_vld;
input ap_start;
input [3:0] op_0;
input [1:0] op_10;
input op_11;
input [31:0] op_12;
input [31:0] op_13;
input [7:0] op_14;
input [3:0] op_15;
input [31:0] op_17;
input op_18;
input op_19;
input [1:0] op_2;
input [3:0] op_3;
input [3:0] op_5;
output ap_done;
output ap_idle;
output ap_ready;
output [31:0] op_31;
output op_31_ap_vld;


reg [11:0] \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.ain_s1 ;
reg [11:0] \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.bin_s1 ;
reg \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.carry_s1 ;
reg [11:0] \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.sum_s1 ;
reg \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.ain_s1 ;
reg \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.bin_s1 ;
reg \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.carry_s1 ;
reg \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.sum_s1 ;
reg \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_0_U.ain_s1 ;
reg \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_0_U.bin_s1 ;
reg \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_0_U.carry_s1 ;
reg \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_0_U.sum_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s1 ;
reg \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.carry_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.sum_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s1 ;
reg \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.carry_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.sum_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s1 ;
reg \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.carry_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.sum_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s1 ;
reg \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.carry_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.sum_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s1 ;
reg \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.carry_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.sum_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s1 ;
reg \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.carry_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.sum_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s1 ;
reg \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.carry_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.sum_s1 ;
reg [16:0] \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.ain_s1 ;
reg [16:0] \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.bin_s1 ;
reg \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.carry_s1 ;
reg [15:0] \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.sum_s1 ;
reg [16:0] \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.ain_s1 ;
reg [16:0] \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.bin_s1 ;
reg \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.carry_s1 ;
reg [16:0] \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.sum_s1 ;
reg [17:0] \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.ain_s1 ;
reg [17:0] \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.bin_s1 ;
reg \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.carry_s1 ;
reg [16:0] \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.sum_s1 ;
reg [19:0] \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.ain_s1 ;
reg [19:0] \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.bin_s1 ;
reg \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.carry_s1 ;
reg [19:0] \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.sum_s1 ;
reg [26:0] \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.ain_s1 ;
reg [26:0] \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.bin_s1 ;
reg \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.carry_s1 ;
reg [26:0] \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.sum_s1 ;
reg [2:0] \add_6s_6ns_6_2_1_U4.top_add_6s_6ns_6_2_1_Adder_2_U.ain_s1 ;
reg [2:0] \add_6s_6ns_6_2_1_U4.top_add_6s_6ns_6_2_1_Adder_2_U.bin_s1 ;
reg \add_6s_6ns_6_2_1_U4.top_add_6s_6ns_6_2_1_Adder_2_U.carry_s1 ;
reg [2:0] \add_6s_6ns_6_2_1_U4.top_add_6s_6ns_6_2_1_Adder_2_U.sum_s1 ;
reg [2:0] \add_6s_6s_6_2_1_U2.top_add_6s_6s_6_2_1_Adder_1_U.ain_s1 ;
reg [2:0] \add_6s_6s_6_2_1_U2.top_add_6s_6s_6_2_1_Adder_1_U.bin_s1 ;
reg \add_6s_6s_6_2_1_U2.top_add_6s_6s_6_2_1_Adder_1_U.carry_s1 ;
reg [2:0] \add_6s_6s_6_2_1_U2.top_add_6s_6s_6_2_1_Adder_1_U.sum_s1 ;
reg [31:0] add_ln691_1_reg_913;
reg [31:0] add_ln691_2_reg_950;
reg [31:0] add_ln691_3_reg_987;
reg [31:0] add_ln691_4_reg_1034;
reg [23:0] add_ln691_reg_876;
reg [1:0] add_ln69_1_reg_829;
reg [5:0] add_ln69_reg_824;
reg [38:0] ap_CS_fsm = 39'h0000000001;
reg icmp_ln1494_reg_779;
reg icmp_ln1499_reg_757;
reg icmp_ln851_1_reg_854;
reg icmp_ln851_2_reg_896;
reg icmp_ln851_3_reg_933;
reg icmp_ln851_4_reg_1017;
reg icmp_ln851_reg_789;
reg [5:0] op_23_V_reg_839;
reg [31:0] op_28_V_reg_1002;
reg [1:0] ret_V_13_reg_799;
reg [32:0] ret_V_14_reg_859;
reg [34:0] ret_V_15_reg_901;
reg [39:0] ret_V_16_reg_938;
reg [33:0] ret_V_17_reg_975;
reg [31:0] ret_V_18_cast_reg_943;
reg [31:0] ret_V_18_reg_992;
reg [53:0] ret_V_19_reg_1022;
reg [31:0] ret_V_20_cast_reg_980;
reg [31:0] ret_V_20_reg_1039;
reg [31:0] ret_V_21_reg_1049;
reg [31:0] ret_V_22_cast_reg_1027;
reg [31:0] ret_V_7_cast_reg_906;
reg [1:0] ret_V_cast_reg_767;
reg [1:0] ret_V_reg_794;
reg [31:0] select_ln1192_1_reg_1054;
reg [31:0] select_ln1192_reg_1044;
reg [31:0] select_ln353_1_reg_918;
reg [31:0] select_ln353_2_reg_955;
reg [23:0] select_ln353_reg_881;
reg [31:0] select_ln69_1_reg_997;
reg [1:0] select_ln69_reg_804;
reg [23:0] sext_ln850_reg_869;
reg signbit_reg_784;
reg [22:0] tmp_reg_864;
reg [2:0] trunc_ln851_reg_774;
reg [3:0] _453_;
wire [31:0] _000_;
wire [31:0] _001_;
wire [31:0] _002_;
wire [31:0] _003_;
wire [23:0] _004_;
wire [1:0] _005_;
wire [5:0] _006_;
wire [38:0] _007_;
wire _008_;
wire _009_;
wire _010_;
wire _011_;
wire _012_;
wire _013_;
wire _014_;
wire [5:0] _015_;
wire [31:0] _016_;
wire [3:0] _017_;
wire [1:0] _018_;
wire [32:0] _019_;
wire [34:0] _020_;
wire [39:0] _021_;
wire [33:0] _022_;
wire [31:0] _023_;
wire [31:0] _024_;
wire [53:0] _025_;
wire [31:0] _026_;
wire [31:0] _027_;
wire [31:0] _028_;
wire [31:0] _029_;
wire [31:0] _030_;
wire [1:0] _031_;
wire [1:0] _032_;
wire [31:0] _033_;
wire [31:0] _034_;
wire [31:0] _035_;
wire [31:0] _036_;
wire [23:0] _037_;
wire [31:0] _038_;
wire [1:0] _039_;
wire [23:0] _040_;
wire _041_;
wire [22:0] _042_;
wire [1:0] _043_;
wire _044_;
wire _045_;
wire _046_;
wire _047_;
wire _048_;
wire _049_;
wire _050_;
wire _051_;
wire _052_;
wire [11:0] _053_;
wire [11:0] _054_;
wire _055_;
wire [11:0] _056_;
wire [12:0] _057_;
wire [12:0] _058_;
wire _059_;
wire _060_;
wire _061_;
wire _062_;
wire [1:0] _063_;
wire [1:0] _064_;
wire _065_;
wire _066_;
wire _067_;
wire _068_;
wire [1:0] _069_;
wire [1:0] _070_;
wire [15:0] _071_;
wire [15:0] _072_;
wire _073_;
wire [15:0] _074_;
wire [16:0] _075_;
wire [16:0] _076_;
wire [15:0] _077_;
wire [15:0] _078_;
wire _079_;
wire [15:0] _080_;
wire [16:0] _081_;
wire [16:0] _082_;
wire [15:0] _083_;
wire [15:0] _084_;
wire _085_;
wire [15:0] _086_;
wire [16:0] _087_;
wire [16:0] _088_;
wire [15:0] _089_;
wire [15:0] _090_;
wire _091_;
wire [15:0] _092_;
wire [16:0] _093_;
wire [16:0] _094_;
wire [15:0] _095_;
wire [15:0] _096_;
wire _097_;
wire [15:0] _098_;
wire [16:0] _099_;
wire [16:0] _100_;
wire [15:0] _101_;
wire [15:0] _102_;
wire _103_;
wire [15:0] _104_;
wire [16:0] _105_;
wire [16:0] _106_;
wire [15:0] _107_;
wire [15:0] _108_;
wire _109_;
wire [15:0] _110_;
wire [16:0] _111_;
wire [16:0] _112_;
wire [16:0] _113_;
wire [16:0] _114_;
wire _115_;
wire [15:0] _116_;
wire [16:0] _117_;
wire [17:0] _118_;
wire [16:0] _119_;
wire [16:0] _120_;
wire _121_;
wire [16:0] _122_;
wire [17:0] _123_;
wire [17:0] _124_;
wire [17:0] _125_;
wire [17:0] _126_;
wire _127_;
wire [16:0] _128_;
wire [17:0] _129_;
wire [18:0] _130_;
wire [19:0] _131_;
wire [19:0] _132_;
wire _133_;
wire [19:0] _134_;
wire [20:0] _135_;
wire [20:0] _136_;
wire [26:0] _137_;
wire [26:0] _138_;
wire _139_;
wire [26:0] _140_;
wire [27:0] _141_;
wire [27:0] _142_;
wire [2:0] _143_;
wire [2:0] _144_;
wire _145_;
wire [2:0] _146_;
wire [3:0] _147_;
wire [3:0] _148_;
wire [2:0] _149_;
wire [2:0] _150_;
wire _151_;
wire [2:0] _152_;
wire [3:0] _153_;
wire [3:0] _154_;
wire _155_;
wire _156_;
wire _157_;
wire _158_;
wire _159_;
wire _160_;
wire _161_;
wire _162_;
wire _163_;
wire _164_;
wire _165_;
wire _166_;
wire _167_;
wire _168_;
wire _169_;
wire _170_;
wire _171_;
wire _172_;
wire _173_;
wire _174_;
wire _175_;
wire _176_;
wire _177_;
wire _178_;
wire _179_;
wire _180_;
wire _181_;
wire _182_;
wire _183_;
wire _184_;
wire _185_;
wire _186_;
wire _187_;
wire _188_;
wire _189_;
wire _190_;
wire _191_;
wire _192_;
wire _193_;
wire _194_;
wire _195_;
wire _196_;
wire _197_;
wire _198_;
wire _199_;
wire \add_24s_24ns_24_2_1_U6.ce ;
wire \add_24s_24ns_24_2_1_U6.clk ;
wire [23:0] \add_24s_24ns_24_2_1_U6.din0 ;
wire [23:0] \add_24s_24ns_24_2_1_U6.din1 ;
wire [23:0] \add_24s_24ns_24_2_1_U6.dout ;
wire \add_24s_24ns_24_2_1_U6.reset ;
wire [23:0] \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.a ;
wire [23:0] \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.ain_s0 ;
wire [23:0] \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.b ;
wire [23:0] \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.bin_s0 ;
wire \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.ce ;
wire \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.clk ;
wire \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.facout_s1 ;
wire \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.facout_s2 ;
wire [11:0] \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.fas_s1 ;
wire [11:0] \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.fas_s2 ;
wire \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.reset ;
wire [23:0] \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.s ;
wire [11:0] \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.u1.a ;
wire [11:0] \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.u1.b ;
wire \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.u1.cin ;
wire \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.u1.cout ;
wire [11:0] \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.u1.s ;
wire [11:0] \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.u2.a ;
wire [11:0] \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.u2.b ;
wire \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.u2.cin ;
wire \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.u2.cout ;
wire [11:0] \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.u2.s ;
wire \add_2ns_2ns_2_2_1_U1.ce ;
wire \add_2ns_2ns_2_2_1_U1.clk ;
wire [1:0] \add_2ns_2ns_2_2_1_U1.din0 ;
wire [1:0] \add_2ns_2ns_2_2_1_U1.din1 ;
wire [1:0] \add_2ns_2ns_2_2_1_U1.dout ;
wire \add_2ns_2ns_2_2_1_U1.reset ;
wire [1:0] \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.a ;
wire [1:0] \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.ain_s0 ;
wire [1:0] \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.b ;
wire [1:0] \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.bin_s0 ;
wire \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.ce ;
wire \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.clk ;
wire \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.facout_s1 ;
wire \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.facout_s2 ;
wire \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.fas_s1 ;
wire \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.fas_s2 ;
wire \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.reset ;
wire [1:0] \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.s ;
wire \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.u1.a ;
wire \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.u1.b ;
wire \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.u1.cin ;
wire \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.u1.cout ;
wire \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.u1.s ;
wire \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.u2.a ;
wire \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.u2.b ;
wire \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.u2.cin ;
wire \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.u2.cout ;
wire \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.u2.s ;
wire \add_2ns_2ns_2_2_1_U3.ce ;
wire \add_2ns_2ns_2_2_1_U3.clk ;
wire [1:0] \add_2ns_2ns_2_2_1_U3.din0 ;
wire [1:0] \add_2ns_2ns_2_2_1_U3.din1 ;
wire [1:0] \add_2ns_2ns_2_2_1_U3.dout ;
wire \add_2ns_2ns_2_2_1_U3.reset ;
wire [1:0] \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_0_U.a ;
wire [1:0] \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_0_U.ain_s0 ;
wire [1:0] \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_0_U.b ;
wire [1:0] \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_0_U.bin_s0 ;
wire \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_0_U.ce ;
wire \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_0_U.clk ;
wire \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_0_U.facout_s1 ;
wire \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_0_U.facout_s2 ;
wire \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_0_U.fas_s1 ;
wire \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_0_U.fas_s2 ;
wire \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_0_U.reset ;
wire [1:0] \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_0_U.s ;
wire \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_0_U.u1.a ;
wire \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_0_U.u1.b ;
wire \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_0_U.u1.cin ;
wire \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_0_U.u1.cout ;
wire \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_0_U.u1.s ;
wire \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_0_U.u2.a ;
wire \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_0_U.u2.b ;
wire \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_0_U.u2.cin ;
wire \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_0_U.u2.cout ;
wire \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_0_U.u2.s ;
wire \add_32ns_32ns_32_2_1_U10.ce ;
wire \add_32ns_32ns_32_2_1_U10.clk ;
wire [31:0] \add_32ns_32ns_32_2_1_U10.din0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U10.din1 ;
wire [31:0] \add_32ns_32ns_32_2_1_U10.dout ;
wire \add_32ns_32ns_32_2_1_U10.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.a ;
wire [31:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.b ;
wire [31:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s0 ;
wire \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.ce ;
wire \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.clk ;
wire \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s1 ;
wire \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s2 ;
wire [15:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s1 ;
wire [15:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s2 ;
wire \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.b ;
wire \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cin ;
wire \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.b ;
wire \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cin ;
wire \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.s ;
wire \add_32ns_32ns_32_2_1_U12.ce ;
wire \add_32ns_32ns_32_2_1_U12.clk ;
wire [31:0] \add_32ns_32ns_32_2_1_U12.din0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U12.din1 ;
wire [31:0] \add_32ns_32ns_32_2_1_U12.dout ;
wire \add_32ns_32ns_32_2_1_U12.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.a ;
wire [31:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.b ;
wire [31:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s0 ;
wire \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.ce ;
wire \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.clk ;
wire \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s1 ;
wire \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s2 ;
wire [15:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s1 ;
wire [15:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s2 ;
wire \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.b ;
wire \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cin ;
wire \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.b ;
wire \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cin ;
wire \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.s ;
wire \add_32ns_32ns_32_2_1_U13.ce ;
wire \add_32ns_32ns_32_2_1_U13.clk ;
wire [31:0] \add_32ns_32ns_32_2_1_U13.din0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U13.din1 ;
wire [31:0] \add_32ns_32ns_32_2_1_U13.dout ;
wire \add_32ns_32ns_32_2_1_U13.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.a ;
wire [31:0] \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.b ;
wire [31:0] \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s0 ;
wire \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.ce ;
wire \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.clk ;
wire \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s1 ;
wire \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s2 ;
wire [15:0] \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s1 ;
wire [15:0] \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s2 ;
wire \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.b ;
wire \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cin ;
wire \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.b ;
wire \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cin ;
wire \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.s ;
wire \add_32ns_32ns_32_2_1_U15.ce ;
wire \add_32ns_32ns_32_2_1_U15.clk ;
wire [31:0] \add_32ns_32ns_32_2_1_U15.din0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U15.din1 ;
wire [31:0] \add_32ns_32ns_32_2_1_U15.dout ;
wire \add_32ns_32ns_32_2_1_U15.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.a ;
wire [31:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.b ;
wire [31:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s0 ;
wire \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.ce ;
wire \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.clk ;
wire \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s1 ;
wire \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s2 ;
wire [15:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s1 ;
wire [15:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s2 ;
wire \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.b ;
wire \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cin ;
wire \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.b ;
wire \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cin ;
wire \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.s ;
wire \add_32ns_32ns_32_2_1_U16.ce ;
wire \add_32ns_32ns_32_2_1_U16.clk ;
wire [31:0] \add_32ns_32ns_32_2_1_U16.din0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U16.din1 ;
wire [31:0] \add_32ns_32ns_32_2_1_U16.dout ;
wire \add_32ns_32ns_32_2_1_U16.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.a ;
wire [31:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.b ;
wire [31:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s0 ;
wire \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.ce ;
wire \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.clk ;
wire \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s1 ;
wire \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s2 ;
wire [15:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s1 ;
wire [15:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s2 ;
wire \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.b ;
wire \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cin ;
wire \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.b ;
wire \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cin ;
wire \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.s ;
wire \add_32ns_32ns_32_2_1_U17.ce ;
wire \add_32ns_32ns_32_2_1_U17.clk ;
wire [31:0] \add_32ns_32ns_32_2_1_U17.din0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U17.din1 ;
wire [31:0] \add_32ns_32ns_32_2_1_U17.dout ;
wire \add_32ns_32ns_32_2_1_U17.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.a ;
wire [31:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.b ;
wire [31:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s0 ;
wire \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.ce ;
wire \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.clk ;
wire \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s1 ;
wire \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s2 ;
wire [15:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s1 ;
wire [15:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s2 ;
wire \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.b ;
wire \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cin ;
wire \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.b ;
wire \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cin ;
wire \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.s ;
wire \add_32ns_32ns_32_2_1_U8.ce ;
wire \add_32ns_32ns_32_2_1_U8.clk ;
wire [31:0] \add_32ns_32ns_32_2_1_U8.din0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U8.din1 ;
wire [31:0] \add_32ns_32ns_32_2_1_U8.dout ;
wire \add_32ns_32ns_32_2_1_U8.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.a ;
wire [31:0] \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.b ;
wire [31:0] \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s0 ;
wire \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.ce ;
wire \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.clk ;
wire \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s1 ;
wire \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s2 ;
wire [15:0] \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s1 ;
wire [15:0] \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s2 ;
wire \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.b ;
wire \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cin ;
wire \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.b ;
wire \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cin ;
wire \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.s ;
wire \add_33s_33s_33_2_1_U5.ce ;
wire \add_33s_33s_33_2_1_U5.clk ;
wire [32:0] \add_33s_33s_33_2_1_U5.din0 ;
wire [32:0] \add_33s_33s_33_2_1_U5.din1 ;
wire [32:0] \add_33s_33s_33_2_1_U5.dout ;
wire \add_33s_33s_33_2_1_U5.reset ;
wire [32:0] \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.a ;
wire [32:0] \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.ain_s0 ;
wire [32:0] \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.b ;
wire [32:0] \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.bin_s0 ;
wire \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.ce ;
wire \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.clk ;
wire \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.facout_s1 ;
wire \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.facout_s2 ;
wire [15:0] \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.fas_s1 ;
wire [16:0] \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.fas_s2 ;
wire \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.reset ;
wire [32:0] \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.s ;
wire [15:0] \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.u1.a ;
wire [15:0] \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.u1.b ;
wire \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.u1.cin ;
wire \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.u1.cout ;
wire [15:0] \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.u1.s ;
wire [16:0] \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.u2.a ;
wire [16:0] \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.u2.b ;
wire \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.u2.cin ;
wire \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.u2.cout ;
wire [16:0] \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.u2.s ;
wire \add_34s_34s_34_2_1_U11.ce ;
wire \add_34s_34s_34_2_1_U11.clk ;
wire [33:0] \add_34s_34s_34_2_1_U11.din0 ;
wire [33:0] \add_34s_34s_34_2_1_U11.din1 ;
wire [33:0] \add_34s_34s_34_2_1_U11.dout ;
wire \add_34s_34s_34_2_1_U11.reset ;
wire [33:0] \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.a ;
wire [33:0] \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.ain_s0 ;
wire [33:0] \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.b ;
wire [33:0] \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.bin_s0 ;
wire \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.ce ;
wire \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.clk ;
wire \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.facout_s1 ;
wire \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.facout_s2 ;
wire [16:0] \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.fas_s1 ;
wire [16:0] \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.fas_s2 ;
wire \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.reset ;
wire [33:0] \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.s ;
wire [16:0] \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.u1.a ;
wire [16:0] \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.u1.b ;
wire \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.u1.cin ;
wire \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.u1.cout ;
wire [16:0] \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.u1.s ;
wire [16:0] \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.u2.a ;
wire [16:0] \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.u2.b ;
wire \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.u2.cin ;
wire \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.u2.cout ;
wire [16:0] \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.u2.s ;
wire \add_35s_35s_35_2_1_U7.ce ;
wire \add_35s_35s_35_2_1_U7.clk ;
wire [34:0] \add_35s_35s_35_2_1_U7.din0 ;
wire [34:0] \add_35s_35s_35_2_1_U7.din1 ;
wire [34:0] \add_35s_35s_35_2_1_U7.dout ;
wire \add_35s_35s_35_2_1_U7.reset ;
wire [34:0] \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.a ;
wire [34:0] \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.ain_s0 ;
wire [34:0] \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.b ;
wire [34:0] \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.bin_s0 ;
wire \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.ce ;
wire \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.clk ;
wire \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.facout_s1 ;
wire \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.facout_s2 ;
wire [16:0] \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.fas_s1 ;
wire [17:0] \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.fas_s2 ;
wire \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.reset ;
wire [34:0] \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.s ;
wire [16:0] \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.u1.a ;
wire [16:0] \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.u1.b ;
wire \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.u1.cin ;
wire \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.u1.cout ;
wire [16:0] \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.u1.s ;
wire [17:0] \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.u2.a ;
wire [17:0] \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.u2.b ;
wire \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.u2.cin ;
wire \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.u2.cout ;
wire [17:0] \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.u2.s ;
wire \add_40s_40s_40_2_1_U9.ce ;
wire \add_40s_40s_40_2_1_U9.clk ;
wire [39:0] \add_40s_40s_40_2_1_U9.din0 ;
wire [39:0] \add_40s_40s_40_2_1_U9.din1 ;
wire [39:0] \add_40s_40s_40_2_1_U9.dout ;
wire \add_40s_40s_40_2_1_U9.reset ;
wire [39:0] \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.a ;
wire [39:0] \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.ain_s0 ;
wire [39:0] \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.b ;
wire [39:0] \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.bin_s0 ;
wire \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.ce ;
wire \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.clk ;
wire \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.facout_s1 ;
wire \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.facout_s2 ;
wire [19:0] \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.fas_s1 ;
wire [19:0] \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.fas_s2 ;
wire \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.reset ;
wire [39:0] \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.s ;
wire [19:0] \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.u1.a ;
wire [19:0] \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.u1.b ;
wire \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.u1.cin ;
wire \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.u1.cout ;
wire [19:0] \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.u1.s ;
wire [19:0] \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.u2.a ;
wire [19:0] \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.u2.b ;
wire \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.u2.cin ;
wire \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.u2.cout ;
wire [19:0] \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.u2.s ;
wire \add_54s_54s_54_2_1_U14.ce ;
wire \add_54s_54s_54_2_1_U14.clk ;
wire [53:0] \add_54s_54s_54_2_1_U14.din0 ;
wire [53:0] \add_54s_54s_54_2_1_U14.din1 ;
wire [53:0] \add_54s_54s_54_2_1_U14.dout ;
wire \add_54s_54s_54_2_1_U14.reset ;
wire [53:0] \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.a ;
wire [53:0] \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.ain_s0 ;
wire [53:0] \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.b ;
wire [53:0] \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.bin_s0 ;
wire \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.ce ;
wire \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.clk ;
wire \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.facout_s1 ;
wire \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.facout_s2 ;
wire [26:0] \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.fas_s1 ;
wire [26:0] \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.fas_s2 ;
wire \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.reset ;
wire [53:0] \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.s ;
wire [26:0] \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.u1.a ;
wire [26:0] \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.u1.b ;
wire \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.u1.cin ;
wire \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.u1.cout ;
wire [26:0] \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.u1.s ;
wire [26:0] \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.u2.a ;
wire [26:0] \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.u2.b ;
wire \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.u2.cin ;
wire \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.u2.cout ;
wire [26:0] \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.u2.s ;
wire \add_6s_6ns_6_2_1_U4.ce ;
wire \add_6s_6ns_6_2_1_U4.clk ;
wire [5:0] \add_6s_6ns_6_2_1_U4.din0 ;
wire [5:0] \add_6s_6ns_6_2_1_U4.din1 ;
wire [5:0] \add_6s_6ns_6_2_1_U4.dout ;
wire \add_6s_6ns_6_2_1_U4.reset ;
wire [5:0] \add_6s_6ns_6_2_1_U4.top_add_6s_6ns_6_2_1_Adder_2_U.a ;
wire [5:0] \add_6s_6ns_6_2_1_U4.top_add_6s_6ns_6_2_1_Adder_2_U.ain_s0 ;
wire [5:0] \add_6s_6ns_6_2_1_U4.top_add_6s_6ns_6_2_1_Adder_2_U.b ;
wire [5:0] \add_6s_6ns_6_2_1_U4.top_add_6s_6ns_6_2_1_Adder_2_U.bin_s0 ;
wire \add_6s_6ns_6_2_1_U4.top_add_6s_6ns_6_2_1_Adder_2_U.ce ;
wire \add_6s_6ns_6_2_1_U4.top_add_6s_6ns_6_2_1_Adder_2_U.clk ;
wire \add_6s_6ns_6_2_1_U4.top_add_6s_6ns_6_2_1_Adder_2_U.facout_s1 ;
wire \add_6s_6ns_6_2_1_U4.top_add_6s_6ns_6_2_1_Adder_2_U.facout_s2 ;
wire [2:0] \add_6s_6ns_6_2_1_U4.top_add_6s_6ns_6_2_1_Adder_2_U.fas_s1 ;
wire [2:0] \add_6s_6ns_6_2_1_U4.top_add_6s_6ns_6_2_1_Adder_2_U.fas_s2 ;
wire \add_6s_6ns_6_2_1_U4.top_add_6s_6ns_6_2_1_Adder_2_U.reset ;
wire [5:0] \add_6s_6ns_6_2_1_U4.top_add_6s_6ns_6_2_1_Adder_2_U.s ;
wire [2:0] \add_6s_6ns_6_2_1_U4.top_add_6s_6ns_6_2_1_Adder_2_U.u1.a ;
wire [2:0] \add_6s_6ns_6_2_1_U4.top_add_6s_6ns_6_2_1_Adder_2_U.u1.b ;
wire \add_6s_6ns_6_2_1_U4.top_add_6s_6ns_6_2_1_Adder_2_U.u1.cin ;
wire \add_6s_6ns_6_2_1_U4.top_add_6s_6ns_6_2_1_Adder_2_U.u1.cout ;
wire [2:0] \add_6s_6ns_6_2_1_U4.top_add_6s_6ns_6_2_1_Adder_2_U.u1.s ;
wire [2:0] \add_6s_6ns_6_2_1_U4.top_add_6s_6ns_6_2_1_Adder_2_U.u2.a ;
wire [2:0] \add_6s_6ns_6_2_1_U4.top_add_6s_6ns_6_2_1_Adder_2_U.u2.b ;
wire \add_6s_6ns_6_2_1_U4.top_add_6s_6ns_6_2_1_Adder_2_U.u2.cin ;
wire \add_6s_6ns_6_2_1_U4.top_add_6s_6ns_6_2_1_Adder_2_U.u2.cout ;
wire [2:0] \add_6s_6ns_6_2_1_U4.top_add_6s_6ns_6_2_1_Adder_2_U.u2.s ;
wire \add_6s_6s_6_2_1_U2.ce ;
wire \add_6s_6s_6_2_1_U2.clk ;
wire [5:0] \add_6s_6s_6_2_1_U2.din0 ;
wire [5:0] \add_6s_6s_6_2_1_U2.din1 ;
wire [5:0] \add_6s_6s_6_2_1_U2.dout ;
wire \add_6s_6s_6_2_1_U2.reset ;
wire [5:0] \add_6s_6s_6_2_1_U2.top_add_6s_6s_6_2_1_Adder_1_U.a ;
wire [5:0] \add_6s_6s_6_2_1_U2.top_add_6s_6s_6_2_1_Adder_1_U.ain_s0 ;
wire [5:0] \add_6s_6s_6_2_1_U2.top_add_6s_6s_6_2_1_Adder_1_U.b ;
wire [5:0] \add_6s_6s_6_2_1_U2.top_add_6s_6s_6_2_1_Adder_1_U.bin_s0 ;
wire \add_6s_6s_6_2_1_U2.top_add_6s_6s_6_2_1_Adder_1_U.ce ;
wire \add_6s_6s_6_2_1_U2.top_add_6s_6s_6_2_1_Adder_1_U.clk ;
wire \add_6s_6s_6_2_1_U2.top_add_6s_6s_6_2_1_Adder_1_U.facout_s1 ;
wire \add_6s_6s_6_2_1_U2.top_add_6s_6s_6_2_1_Adder_1_U.facout_s2 ;
wire [2:0] \add_6s_6s_6_2_1_U2.top_add_6s_6s_6_2_1_Adder_1_U.fas_s1 ;
wire [2:0] \add_6s_6s_6_2_1_U2.top_add_6s_6s_6_2_1_Adder_1_U.fas_s2 ;
wire \add_6s_6s_6_2_1_U2.top_add_6s_6s_6_2_1_Adder_1_U.reset ;
wire [5:0] \add_6s_6s_6_2_1_U2.top_add_6s_6s_6_2_1_Adder_1_U.s ;
wire [2:0] \add_6s_6s_6_2_1_U2.top_add_6s_6s_6_2_1_Adder_1_U.u1.a ;
wire [2:0] \add_6s_6s_6_2_1_U2.top_add_6s_6s_6_2_1_Adder_1_U.u1.b ;
wire \add_6s_6s_6_2_1_U2.top_add_6s_6s_6_2_1_Adder_1_U.u1.cin ;
wire \add_6s_6s_6_2_1_U2.top_add_6s_6s_6_2_1_Adder_1_U.u1.cout ;
wire [2:0] \add_6s_6s_6_2_1_U2.top_add_6s_6s_6_2_1_Adder_1_U.u1.s ;
wire [2:0] \add_6s_6s_6_2_1_U2.top_add_6s_6s_6_2_1_Adder_1_U.u2.a ;
wire [2:0] \add_6s_6s_6_2_1_U2.top_add_6s_6s_6_2_1_Adder_1_U.u2.b ;
wire \add_6s_6s_6_2_1_U2.top_add_6s_6s_6_2_1_Adder_1_U.u2.cin ;
wire \add_6s_6s_6_2_1_U2.top_add_6s_6s_6_2_1_Adder_1_U.u2.cout ;
wire [2:0] \add_6s_6s_6_2_1_U2.top_add_6s_6s_6_2_1_Adder_1_U.u2.s ;
wire ap_CS_fsm_state1;
wire ap_CS_fsm_state10;
wire ap_CS_fsm_state11;
wire ap_CS_fsm_state12;
wire ap_CS_fsm_state13;
wire ap_CS_fsm_state14;
wire ap_CS_fsm_state15;
wire ap_CS_fsm_state16;
wire ap_CS_fsm_state17;
wire ap_CS_fsm_state18;
wire ap_CS_fsm_state19;
wire ap_CS_fsm_state2;
wire ap_CS_fsm_state20;
wire ap_CS_fsm_state21;
wire ap_CS_fsm_state22;
wire ap_CS_fsm_state23;
wire ap_CS_fsm_state24;
wire ap_CS_fsm_state25;
wire ap_CS_fsm_state26;
wire ap_CS_fsm_state27;
wire ap_CS_fsm_state28;
wire ap_CS_fsm_state29;
wire ap_CS_fsm_state3;
wire ap_CS_fsm_state30;
wire ap_CS_fsm_state31;
wire ap_CS_fsm_state32;
wire ap_CS_fsm_state33;
wire ap_CS_fsm_state34;
wire ap_CS_fsm_state35;
wire ap_CS_fsm_state36;
wire ap_CS_fsm_state37;
wire ap_CS_fsm_state38;
wire ap_CS_fsm_state39;
wire ap_CS_fsm_state4;
wire ap_CS_fsm_state5;
wire ap_CS_fsm_state6;
wire ap_CS_fsm_state7;
wire ap_CS_fsm_state8;
wire ap_CS_fsm_state9;
wire [38:0] ap_NS_fsm;
wire ap_clk;
wire ap_done;
wire ap_idle;
wire ap_ready;
wire ap_rst;
wire ap_start;
wire [1:0] grp_fu_320_p2;
wire [5:0] grp_fu_369_p0;
wire [5:0] grp_fu_369_p1;
wire [5:0] grp_fu_369_p2;
wire [1:0] grp_fu_375_p0;
wire [1:0] grp_fu_375_p2;
wire [5:0] grp_fu_383_p0;
wire [5:0] grp_fu_383_p2;
wire [32:0] grp_fu_403_p0;
wire [32:0] grp_fu_403_p1;
wire [32:0] grp_fu_403_p2;
wire [23:0] grp_fu_432_p0;
wire [23:0] grp_fu_432_p2;
wire [34:0] grp_fu_472_p0;
wire [34:0] grp_fu_472_p1;
wire [34:0] grp_fu_472_p2;
wire [31:0] grp_fu_498_p2;
wire [39:0] grp_fu_537_p0;
wire [39:0] grp_fu_537_p1;
wire [39:0] grp_fu_537_p2;
wire [31:0] grp_fu_563_p2;
wire [33:0] grp_fu_602_p0;
wire [33:0] grp_fu_602_p1;
wire [33:0] grp_fu_602_p2;
wire [31:0] grp_fu_618_p2;
wire [31:0] grp_fu_663_p2;
wire [53:0] grp_fu_682_p0;
wire [53:0] grp_fu_682_p1;
wire [53:0] grp_fu_682_p2;
wire [31:0] grp_fu_708_p2;
wire [31:0] grp_fu_740_p2;
wire [31:0] grp_fu_752_p2;
wire icmp_ln1494_fu_303_p2;
wire icmp_ln1499_fu_253_p2;
wire icmp_ln851_1_fu_413_p2;
wire icmp_ln851_2_fu_482_p2;
wire icmp_ln851_3_fu_547_p2;
wire icmp_ln851_4_fu_692_p2;
wire icmp_ln851_fu_315_p2;
wire [3:0] op_0;
wire [1:0] op_10;
wire op_11;
wire [31:0] op_12;
wire [31:0] op_13;
wire [7:0] op_14;
wire [3:0] op_15;
wire op_16_V_fu_627_p2;
wire [31:0] op_17;
wire op_18;
wire op_19;
wire [1:0] op_2;
wire [4:0] op_20_V_fu_352_p3;
wire [3:0] op_3;
wire [31:0] op_31;
wire op_31_ap_vld;
wire [7:0] op_4_V_fu_233_p3;
wire [3:0] op_5;
wire p_Result_1_fu_438_p3;
wire p_Result_2_fu_503_p3;
wire p_Result_3_fu_568_p3;
wire p_Result_4_fu_632_p3;
wire p_Result_5_fu_713_p3;
wire p_Result_s_fu_325_p3;
wire [6:0] ret_V_12_fu_271_p2;
wire [6:0] ret_V_12_reg_762;
wire [1:0] ret_V_13_fu_337_p3;
wire [31:0] ret_V_18_fu_648_p3;
wire [31:0] ret_V_20_fu_725_p3;
wire [15:0] rhs_2_fu_392_p3;
wire [38:0] rhs_3_fu_526_p3;
wire [32:0] rhs_4_fu_591_p3;
wire [52:0] rhs_6_fu_671_p3;
wire [6:0] rhs_fu_263_p3;
wire [31:0] select_ln1192_1_fu_744_p3;
wire [31:0] select_ln1192_fu_732_p3;
wire [31:0] select_ln353_1_fu_515_p3;
wire [31:0] select_ln353_2_fu_580_p3;
wire [23:0] select_ln353_fu_450_p3;
wire [31:0] select_ln69_1_fu_655_p3;
wire [1:0] select_ln69_fu_344_p3;
wire [23:0] select_ln850_1_fu_445_p3;
wire [31:0] select_ln850_2_fu_510_p3;
wire [31:0] select_ln850_3_fu_575_p3;
wire [31:0] select_ln850_4_fu_642_p3;
wire [31:0] select_ln850_5_fu_720_p3;
wire [1:0] select_ln850_fu_332_p3;
wire [31:0] sext_ln1192_fu_388_p0;
wire [7:0] sext_ln1494_fu_299_p1;
wire [3:0] sext_ln1499_fu_249_p0;
wire [4:0] sext_ln1499_fu_249_p1;
wire [31:0] sext_ln703_1_fu_457_p0;
wire [7:0] sext_ln703_2_fu_522_p0;
wire [3:0] sext_ln703_3_fu_587_p0;
wire [31:0] sext_ln703_4_fu_667_p0;
wire [3:0] sext_ln703_fu_259_p0;
wire [6:0] sext_ln703_fu_259_p1;
wire [23:0] sext_ln850_fu_429_p1;
wire [3:0] shl_ln728_2_fu_291_p1;
wire [6:0] shl_ln728_2_fu_291_p3;
wire [4:0] shl_ln_fu_241_p3;
wire signbit_fu_309_p2;
wire [25:0] tmp_3_fu_461_p3;
wire trunc_ln1195_fu_623_p1;
wire [31:0] trunc_ln851_1_fu_409_p0;
wire [9:0] trunc_ln851_1_fu_409_p1;
wire [31:0] trunc_ln851_2_fu_478_p0;
wire [1:0] trunc_ln851_2_fu_478_p1;
wire [7:0] trunc_ln851_3_fu_543_p0;
wire [6:0] trunc_ln851_3_fu_543_p1;
wire [3:0] trunc_ln851_4_fu_639_p0;
wire trunc_ln851_4_fu_639_p1;
wire [31:0] trunc_ln851_5_fu_688_p0;
wire [20:0] trunc_ln851_5_fu_688_p1;
wire [2:0] trunc_ln851_fu_287_p1;


assign _044_ = ap_CS_fsm[16] & icmp_ln851_2_reg_896;
assign _045_ = icmp_ln851_3_reg_933 & ap_CS_fsm[21];
assign _046_ = icmp_ln851_4_reg_1017 & ap_CS_fsm[33];
assign _047_ = ap_CS_fsm[11] & icmp_ln851_1_reg_854;
assign _048_ = _050_ & ap_CS_fsm[0];
assign _049_ = ap_start & ap_CS_fsm[0];
assign ret_V_12_fu_271_p2 = { op_3[3], op_3[3], op_3[3], op_3 } & { op_5, 3'h0 };
assign _050_ = ~ ap_start;
assign _051_ = ! trunc_ln851_reg_774;
assign _052_ = { op_3[3], op_3 } == { op_2, 3'h0 };
always @(posedge \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.clk )
\add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.bin_s1  <= _054_;
always @(posedge \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.clk )
\add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.ain_s1  <= _053_;
always @(posedge \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.clk )
\add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.sum_s1  <= _056_;
always @(posedge \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.clk )
\add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.carry_s1  <= _055_;
assign _054_ = \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.ce  ? \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.b [23:12] : \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.bin_s1 ;
assign _053_ = \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.ce  ? \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.a [23:12] : \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.ain_s1 ;
assign _055_ = \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.ce  ? \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.facout_s1  : \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.carry_s1 ;
assign _056_ = \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.ce  ? \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.fas_s1  : \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.sum_s1 ;
assign _057_ = \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.u1.a  + \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.u1.b ;
assign { \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.u1.cout , \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.u1.s  } = _057_ + \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.u1.cin ;
assign _058_ = \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.u2.a  + \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.u2.b ;
assign { \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.u2.cout , \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.u2.s  } = _058_ + \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.u2.cin ;
always @(posedge \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.clk )
\add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.bin_s1  <= _060_;
always @(posedge \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.clk )
\add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.ain_s1  <= _059_;
always @(posedge \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.clk )
\add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.sum_s1  <= _062_;
always @(posedge \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.clk )
\add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.carry_s1  <= _061_;
assign _060_ = \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.ce  ? \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.b [1] : \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.bin_s1 ;
assign _059_ = \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.ce  ? \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.a [1] : \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.ain_s1 ;
assign _061_ = \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.ce  ? \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.facout_s1  : \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.carry_s1 ;
assign _062_ = \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.ce  ? \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.fas_s1  : \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.sum_s1 ;
assign _063_ = \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.u1.a  + \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.u1.b ;
assign { \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.u1.cout , \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.u1.s  } = _063_ + \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.u1.cin ;
assign _064_ = \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.u2.a  + \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.u2.b ;
assign { \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.u2.cout , \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.u2.s  } = _064_ + \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.u2.cin ;
always @(posedge \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_0_U.clk )
\add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_0_U.bin_s1  <= _066_;
always @(posedge \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_0_U.clk )
\add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_0_U.ain_s1  <= _065_;
always @(posedge \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_0_U.clk )
\add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_0_U.sum_s1  <= _068_;
always @(posedge \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_0_U.clk )
\add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_0_U.carry_s1  <= _067_;
assign _066_ = \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_0_U.ce  ? \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_0_U.b [1] : \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_0_U.bin_s1 ;
assign _065_ = \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_0_U.ce  ? \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_0_U.a [1] : \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_0_U.ain_s1 ;
assign _067_ = \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_0_U.ce  ? \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_0_U.facout_s1  : \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_0_U.carry_s1 ;
assign _068_ = \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_0_U.ce  ? \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_0_U.fas_s1  : \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_0_U.sum_s1 ;
assign _069_ = \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_0_U.u1.a  + \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_0_U.u1.b ;
assign { \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_0_U.u1.cout , \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_0_U.u1.s  } = _069_ + \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_0_U.u1.cin ;
assign _070_ = \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_0_U.u2.a  + \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_0_U.u2.b ;
assign { \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_0_U.u2.cout , \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_0_U.u2.s  } = _070_ + \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_0_U.u2.cin ;
always @(posedge \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.clk )
\add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s1  <= _072_;
always @(posedge \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.clk )
\add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s1  <= _071_;
always @(posedge \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.clk )
\add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.sum_s1  <= _074_;
always @(posedge \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.clk )
\add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.carry_s1  <= _073_;
assign _072_ = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  ? \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.b [31:16] : \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s1 ;
assign _071_ = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  ? \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.a [31:16] : \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s1 ;
assign _073_ = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  ? \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s1  : \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.carry_s1 ;
assign _074_ = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  ? \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s1  : \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.sum_s1 ;
assign _075_ = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.a  + \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.b ;
assign { \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cout , \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.s  } = _075_ + \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cin ;
assign _076_ = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.a  + \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.b ;
assign { \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cout , \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.s  } = _076_ + \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cin ;
always @(posedge \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.clk )
\add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s1  <= _078_;
always @(posedge \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.clk )
\add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s1  <= _077_;
always @(posedge \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.clk )
\add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.sum_s1  <= _080_;
always @(posedge \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.clk )
\add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.carry_s1  <= _079_;
assign _078_ = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  ? \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.b [31:16] : \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s1 ;
assign _077_ = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  ? \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.a [31:16] : \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s1 ;
assign _079_ = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  ? \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s1  : \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.carry_s1 ;
assign _080_ = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  ? \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s1  : \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.sum_s1 ;
assign _081_ = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.a  + \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.b ;
assign { \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cout , \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.s  } = _081_ + \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cin ;
assign _082_ = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.a  + \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.b ;
assign { \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cout , \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.s  } = _082_ + \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cin ;
always @(posedge \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.clk )
\add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s1  <= _084_;
always @(posedge \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.clk )
\add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s1  <= _083_;
always @(posedge \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.clk )
\add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.sum_s1  <= _086_;
always @(posedge \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.clk )
\add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.carry_s1  <= _085_;
assign _084_ = \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  ? \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.b [31:16] : \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s1 ;
assign _083_ = \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  ? \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.a [31:16] : \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s1 ;
assign _085_ = \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  ? \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s1  : \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.carry_s1 ;
assign _086_ = \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  ? \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s1  : \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.sum_s1 ;
assign _087_ = \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.a  + \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.b ;
assign { \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cout , \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.s  } = _087_ + \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cin ;
assign _088_ = \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.a  + \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.b ;
assign { \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cout , \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.s  } = _088_ + \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cin ;
always @(posedge \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.clk )
\add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s1  <= _090_;
always @(posedge \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.clk )
\add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s1  <= _089_;
always @(posedge \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.clk )
\add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.sum_s1  <= _092_;
always @(posedge \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.clk )
\add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.carry_s1  <= _091_;
assign _090_ = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  ? \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.b [31:16] : \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s1 ;
assign _089_ = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  ? \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.a [31:16] : \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s1 ;
assign _091_ = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  ? \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s1  : \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.carry_s1 ;
assign _092_ = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  ? \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s1  : \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.sum_s1 ;
assign _093_ = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.a  + \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.b ;
assign { \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cout , \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.s  } = _093_ + \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cin ;
assign _094_ = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.a  + \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.b ;
assign { \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cout , \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.s  } = _094_ + \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cin ;
always @(posedge \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.clk )
\add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s1  <= _096_;
always @(posedge \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.clk )
\add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s1  <= _095_;
always @(posedge \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.clk )
\add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.sum_s1  <= _098_;
always @(posedge \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.clk )
\add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.carry_s1  <= _097_;
assign _096_ = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  ? \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.b [31:16] : \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s1 ;
assign _095_ = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  ? \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.a [31:16] : \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s1 ;
assign _097_ = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  ? \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s1  : \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.carry_s1 ;
assign _098_ = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  ? \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s1  : \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.sum_s1 ;
assign _099_ = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.a  + \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.b ;
assign { \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cout , \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.s  } = _099_ + \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cin ;
assign _100_ = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.a  + \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.b ;
assign { \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cout , \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.s  } = _100_ + \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cin ;
always @(posedge \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.clk )
\add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s1  <= _102_;
always @(posedge \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.clk )
\add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s1  <= _101_;
always @(posedge \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.clk )
\add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.sum_s1  <= _104_;
always @(posedge \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.clk )
\add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.carry_s1  <= _103_;
assign _102_ = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  ? \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.b [31:16] : \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s1 ;
assign _101_ = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  ? \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.a [31:16] : \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s1 ;
assign _103_ = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  ? \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s1  : \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.carry_s1 ;
assign _104_ = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  ? \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s1  : \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.sum_s1 ;
assign _105_ = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.a  + \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.b ;
assign { \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cout , \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.s  } = _105_ + \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cin ;
assign _106_ = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.a  + \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.b ;
assign { \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cout , \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.s  } = _106_ + \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cin ;
always @(posedge \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.clk )
\add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s1  <= _108_;
always @(posedge \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.clk )
\add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s1  <= _107_;
always @(posedge \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.clk )
\add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.sum_s1  <= _110_;
always @(posedge \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.clk )
\add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.carry_s1  <= _109_;
assign _108_ = \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  ? \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.b [31:16] : \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s1 ;
assign _107_ = \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  ? \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.a [31:16] : \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s1 ;
assign _109_ = \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  ? \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s1  : \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.carry_s1 ;
assign _110_ = \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  ? \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s1  : \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.sum_s1 ;
assign _111_ = \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.a  + \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.b ;
assign { \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cout , \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.s  } = _111_ + \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cin ;
assign _112_ = \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.a  + \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.b ;
assign { \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cout , \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.s  } = _112_ + \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cin ;
always @(posedge \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.clk )
\add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.bin_s1  <= _114_;
always @(posedge \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.clk )
\add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.ain_s1  <= _113_;
always @(posedge \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.clk )
\add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.sum_s1  <= _116_;
always @(posedge \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.clk )
\add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.carry_s1  <= _115_;
assign _114_ = \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.ce  ? \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.b [32:16] : \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.bin_s1 ;
assign _113_ = \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.ce  ? \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.a [32:16] : \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.ain_s1 ;
assign _115_ = \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.ce  ? \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.facout_s1  : \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.carry_s1 ;
assign _116_ = \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.ce  ? \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.fas_s1  : \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.sum_s1 ;
assign _117_ = \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.u1.a  + \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.u1.b ;
assign { \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.u1.cout , \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.u1.s  } = _117_ + \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.u1.cin ;
assign _118_ = \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.u2.a  + \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.u2.b ;
assign { \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.u2.cout , \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.u2.s  } = _118_ + \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.u2.cin ;
always @(posedge \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.clk )
\add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.bin_s1  <= _120_;
always @(posedge \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.clk )
\add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.ain_s1  <= _119_;
always @(posedge \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.clk )
\add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.sum_s1  <= _122_;
always @(posedge \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.clk )
\add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.carry_s1  <= _121_;
assign _120_ = \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.ce  ? \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.b [33:17] : \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.bin_s1 ;
assign _119_ = \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.ce  ? \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.a [33:17] : \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.ain_s1 ;
assign _121_ = \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.ce  ? \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.facout_s1  : \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.carry_s1 ;
assign _122_ = \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.ce  ? \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.fas_s1  : \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.sum_s1 ;
assign _123_ = \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.u1.a  + \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.u1.b ;
assign { \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.u1.cout , \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.u1.s  } = _123_ + \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.u1.cin ;
assign _124_ = \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.u2.a  + \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.u2.b ;
assign { \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.u2.cout , \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.u2.s  } = _124_ + \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.u2.cin ;
always @(posedge \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.clk )
\add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.bin_s1  <= _126_;
always @(posedge \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.clk )
\add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.ain_s1  <= _125_;
always @(posedge \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.clk )
\add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.sum_s1  <= _128_;
always @(posedge \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.clk )
\add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.carry_s1  <= _127_;
assign _126_ = \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.ce  ? \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.b [34:17] : \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.bin_s1 ;
assign _125_ = \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.ce  ? \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.a [34:17] : \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.ain_s1 ;
assign _127_ = \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.ce  ? \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.facout_s1  : \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.carry_s1 ;
assign _128_ = \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.ce  ? \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.fas_s1  : \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.sum_s1 ;
assign _129_ = \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.u1.a  + \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.u1.b ;
assign { \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.u1.cout , \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.u1.s  } = _129_ + \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.u1.cin ;
assign _130_ = \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.u2.a  + \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.u2.b ;
assign { \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.u2.cout , \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.u2.s  } = _130_ + \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.u2.cin ;
always @(posedge \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.clk )
\add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.bin_s1  <= _132_;
always @(posedge \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.clk )
\add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.ain_s1  <= _131_;
always @(posedge \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.clk )
\add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.sum_s1  <= _134_;
always @(posedge \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.clk )
\add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.carry_s1  <= _133_;
assign _132_ = \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.ce  ? \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.b [39:20] : \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.bin_s1 ;
assign _131_ = \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.ce  ? \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.a [39:20] : \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.ain_s1 ;
assign _133_ = \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.ce  ? \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.facout_s1  : \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.carry_s1 ;
assign _134_ = \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.ce  ? \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.fas_s1  : \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.sum_s1 ;
assign _135_ = \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.u1.a  + \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.u1.b ;
assign { \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.u1.cout , \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.u1.s  } = _135_ + \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.u1.cin ;
assign _136_ = \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.u2.a  + \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.u2.b ;
assign { \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.u2.cout , \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.u2.s  } = _136_ + \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.u2.cin ;
always @(posedge \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.clk )
\add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.bin_s1  <= _138_;
always @(posedge \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.clk )
\add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.ain_s1  <= _137_;
always @(posedge \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.clk )
\add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.sum_s1  <= _140_;
always @(posedge \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.clk )
\add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.carry_s1  <= _139_;
assign _138_ = \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.ce  ? \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.b [53:27] : \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.bin_s1 ;
assign _137_ = \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.ce  ? \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.a [53:27] : \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.ain_s1 ;
assign _139_ = \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.ce  ? \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.facout_s1  : \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.carry_s1 ;
assign _140_ = \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.ce  ? \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.fas_s1  : \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.sum_s1 ;
assign _141_ = \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.u1.a  + \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.u1.b ;
assign { \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.u1.cout , \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.u1.s  } = _141_ + \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.u1.cin ;
assign _142_ = \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.u2.a  + \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.u2.b ;
assign { \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.u2.cout , \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.u2.s  } = _142_ + \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.u2.cin ;
always @(posedge \add_6s_6ns_6_2_1_U4.top_add_6s_6ns_6_2_1_Adder_2_U.clk )
\add_6s_6ns_6_2_1_U4.top_add_6s_6ns_6_2_1_Adder_2_U.bin_s1  <= _144_;
always @(posedge \add_6s_6ns_6_2_1_U4.top_add_6s_6ns_6_2_1_Adder_2_U.clk )
\add_6s_6ns_6_2_1_U4.top_add_6s_6ns_6_2_1_Adder_2_U.ain_s1  <= _143_;
always @(posedge \add_6s_6ns_6_2_1_U4.top_add_6s_6ns_6_2_1_Adder_2_U.clk )
\add_6s_6ns_6_2_1_U4.top_add_6s_6ns_6_2_1_Adder_2_U.sum_s1  <= _146_;
always @(posedge \add_6s_6ns_6_2_1_U4.top_add_6s_6ns_6_2_1_Adder_2_U.clk )
\add_6s_6ns_6_2_1_U4.top_add_6s_6ns_6_2_1_Adder_2_U.carry_s1  <= _145_;
assign _144_ = \add_6s_6ns_6_2_1_U4.top_add_6s_6ns_6_2_1_Adder_2_U.ce  ? \add_6s_6ns_6_2_1_U4.top_add_6s_6ns_6_2_1_Adder_2_U.b [5:3] : \add_6s_6ns_6_2_1_U4.top_add_6s_6ns_6_2_1_Adder_2_U.bin_s1 ;
assign _143_ = \add_6s_6ns_6_2_1_U4.top_add_6s_6ns_6_2_1_Adder_2_U.ce  ? \add_6s_6ns_6_2_1_U4.top_add_6s_6ns_6_2_1_Adder_2_U.a [5:3] : \add_6s_6ns_6_2_1_U4.top_add_6s_6ns_6_2_1_Adder_2_U.ain_s1 ;
assign _145_ = \add_6s_6ns_6_2_1_U4.top_add_6s_6ns_6_2_1_Adder_2_U.ce  ? \add_6s_6ns_6_2_1_U4.top_add_6s_6ns_6_2_1_Adder_2_U.facout_s1  : \add_6s_6ns_6_2_1_U4.top_add_6s_6ns_6_2_1_Adder_2_U.carry_s1 ;
assign _146_ = \add_6s_6ns_6_2_1_U4.top_add_6s_6ns_6_2_1_Adder_2_U.ce  ? \add_6s_6ns_6_2_1_U4.top_add_6s_6ns_6_2_1_Adder_2_U.fas_s1  : \add_6s_6ns_6_2_1_U4.top_add_6s_6ns_6_2_1_Adder_2_U.sum_s1 ;
assign _147_ = \add_6s_6ns_6_2_1_U4.top_add_6s_6ns_6_2_1_Adder_2_U.u1.a  + \add_6s_6ns_6_2_1_U4.top_add_6s_6ns_6_2_1_Adder_2_U.u1.b ;
assign { \add_6s_6ns_6_2_1_U4.top_add_6s_6ns_6_2_1_Adder_2_U.u1.cout , \add_6s_6ns_6_2_1_U4.top_add_6s_6ns_6_2_1_Adder_2_U.u1.s  } = _147_ + \add_6s_6ns_6_2_1_U4.top_add_6s_6ns_6_2_1_Adder_2_U.u1.cin ;
assign _148_ = \add_6s_6ns_6_2_1_U4.top_add_6s_6ns_6_2_1_Adder_2_U.u2.a  + \add_6s_6ns_6_2_1_U4.top_add_6s_6ns_6_2_1_Adder_2_U.u2.b ;
assign { \add_6s_6ns_6_2_1_U4.top_add_6s_6ns_6_2_1_Adder_2_U.u2.cout , \add_6s_6ns_6_2_1_U4.top_add_6s_6ns_6_2_1_Adder_2_U.u2.s  } = _148_ + \add_6s_6ns_6_2_1_U4.top_add_6s_6ns_6_2_1_Adder_2_U.u2.cin ;
always @(posedge \add_6s_6s_6_2_1_U2.top_add_6s_6s_6_2_1_Adder_1_U.clk )
\add_6s_6s_6_2_1_U2.top_add_6s_6s_6_2_1_Adder_1_U.bin_s1  <= _150_;
always @(posedge \add_6s_6s_6_2_1_U2.top_add_6s_6s_6_2_1_Adder_1_U.clk )
\add_6s_6s_6_2_1_U2.top_add_6s_6s_6_2_1_Adder_1_U.ain_s1  <= _149_;
always @(posedge \add_6s_6s_6_2_1_U2.top_add_6s_6s_6_2_1_Adder_1_U.clk )
\add_6s_6s_6_2_1_U2.top_add_6s_6s_6_2_1_Adder_1_U.sum_s1  <= _152_;
always @(posedge \add_6s_6s_6_2_1_U2.top_add_6s_6s_6_2_1_Adder_1_U.clk )
\add_6s_6s_6_2_1_U2.top_add_6s_6s_6_2_1_Adder_1_U.carry_s1  <= _151_;
assign _150_ = \add_6s_6s_6_2_1_U2.top_add_6s_6s_6_2_1_Adder_1_U.ce  ? \add_6s_6s_6_2_1_U2.top_add_6s_6s_6_2_1_Adder_1_U.b [5:3] : \add_6s_6s_6_2_1_U2.top_add_6s_6s_6_2_1_Adder_1_U.bin_s1 ;
assign _149_ = \add_6s_6s_6_2_1_U2.top_add_6s_6s_6_2_1_Adder_1_U.ce  ? \add_6s_6s_6_2_1_U2.top_add_6s_6s_6_2_1_Adder_1_U.a [5:3] : \add_6s_6s_6_2_1_U2.top_add_6s_6s_6_2_1_Adder_1_U.ain_s1 ;
assign _151_ = \add_6s_6s_6_2_1_U2.top_add_6s_6s_6_2_1_Adder_1_U.ce  ? \add_6s_6s_6_2_1_U2.top_add_6s_6s_6_2_1_Adder_1_U.facout_s1  : \add_6s_6s_6_2_1_U2.top_add_6s_6s_6_2_1_Adder_1_U.carry_s1 ;
assign _152_ = \add_6s_6s_6_2_1_U2.top_add_6s_6s_6_2_1_Adder_1_U.ce  ? \add_6s_6s_6_2_1_U2.top_add_6s_6s_6_2_1_Adder_1_U.fas_s1  : \add_6s_6s_6_2_1_U2.top_add_6s_6s_6_2_1_Adder_1_U.sum_s1 ;
assign _153_ = \add_6s_6s_6_2_1_U2.top_add_6s_6s_6_2_1_Adder_1_U.u1.a  + \add_6s_6s_6_2_1_U2.top_add_6s_6s_6_2_1_Adder_1_U.u1.b ;
assign { \add_6s_6s_6_2_1_U2.top_add_6s_6s_6_2_1_Adder_1_U.u1.cout , \add_6s_6s_6_2_1_U2.top_add_6s_6s_6_2_1_Adder_1_U.u1.s  } = _153_ + \add_6s_6s_6_2_1_U2.top_add_6s_6s_6_2_1_Adder_1_U.u1.cin ;
assign _154_ = \add_6s_6s_6_2_1_U2.top_add_6s_6s_6_2_1_Adder_1_U.u2.a  + \add_6s_6s_6_2_1_U2.top_add_6s_6s_6_2_1_Adder_1_U.u2.b ;
assign { \add_6s_6s_6_2_1_U2.top_add_6s_6s_6_2_1_Adder_1_U.u2.cout , \add_6s_6s_6_2_1_U2.top_add_6s_6s_6_2_1_Adder_1_U.u2.s  } = _154_ + \add_6s_6s_6_2_1_U2.top_add_6s_6s_6_2_1_Adder_1_U.u2.cin ;
assign _155_ = $signed({ op_3, 3'h0 }) > $signed({ op_2, 6'h00 });
assign _156_ = { op_2, 3'h0 } != { op_3[3], op_3 };
assign _157_ = | op_12[9:0];
assign _158_ = | op_13[1:0];
assign _159_ = | op_14[6:0];
assign _160_ = | op_17[20:0];
assign op_16_V_fu_627_p2 = op_10[0] | signbit_reg_784;
always @(posedge ap_clk)
trunc_ln851_reg_774 <= 3'h0;
always @(posedge ap_clk)
sext_ln850_reg_869 <= _040_;
always @(posedge ap_clk)
select_ln353_reg_881 <= _037_;
always @(posedge ap_clk)
select_ln353_2_reg_955 <= _036_;
always @(posedge ap_clk)
select_ln353_1_reg_918 <= _035_;
always @(posedge ap_clk)
ret_V_reg_794 <= _032_;
always @(posedge ap_clk)
ret_V_21_reg_1049 <= _028_;
always @(posedge ap_clk)
select_ln1192_1_reg_1054 <= _033_;
always @(posedge ap_clk)
ret_V_20_reg_1039 <= _027_;
always @(posedge ap_clk)
select_ln1192_reg_1044 <= _034_;
always @(posedge ap_clk)
ret_V_19_reg_1022 <= _025_;
always @(posedge ap_clk)
ret_V_22_cast_reg_1027 <= _029_;
always @(posedge ap_clk)
ret_V_18_reg_992 <= _024_;
always @(posedge ap_clk)
select_ln69_1_reg_997 <= _038_;
always @(posedge ap_clk)
ret_V_17_reg_975 <= _022_;
always @(posedge ap_clk)
ret_V_20_cast_reg_980 <= _026_;
always @(posedge ap_clk)
ret_V_16_reg_938 <= _021_;
always @(posedge ap_clk)
ret_V_18_cast_reg_943 <= _023_;
always @(posedge ap_clk)
ret_V_15_reg_901 <= _020_;
always @(posedge ap_clk)
ret_V_7_cast_reg_906 <= _030_;
always @(posedge ap_clk)
ret_V_14_reg_859 <= _019_;
always @(posedge ap_clk)
tmp_reg_864 <= _042_;
always @(posedge ap_clk)
ret_V_13_reg_799 <= _018_;
always @(posedge ap_clk)
select_ln69_reg_804 <= _039_;
always @(posedge ap_clk)
op_28_V_reg_1002 <= _016_;
always @(posedge ap_clk)
op_23_V_reg_839 <= _015_;
always @(posedge ap_clk)
icmp_ln851_reg_789 <= _014_;
always @(posedge ap_clk)
icmp_ln851_4_reg_1017 <= _013_;
always @(posedge ap_clk)
icmp_ln851_3_reg_933 <= _012_;
always @(posedge ap_clk)
icmp_ln851_2_reg_896 <= _011_;
always @(posedge ap_clk)
icmp_ln851_1_reg_854 <= _010_;
always @(posedge ap_clk)
icmp_ln1499_reg_757 <= _009_;
always @(posedge ap_clk)
_453_ <= _017_;
assign ret_V_12_reg_762[6:3] = _453_;
always @(posedge ap_clk)
ret_V_cast_reg_767 <= _031_;
always @(posedge ap_clk)
icmp_ln1494_reg_779 <= _008_;
always @(posedge ap_clk)
signbit_reg_784 <= _041_;
always @(posedge ap_clk)
add_ln69_reg_824 <= _006_;
always @(posedge ap_clk)
add_ln69_1_reg_829 <= _005_;
always @(posedge ap_clk)
add_ln691_reg_876 <= _004_;
always @(posedge ap_clk)
add_ln691_4_reg_1034 <= _003_;
always @(posedge ap_clk)
add_ln691_3_reg_987 <= _002_;
always @(posedge ap_clk)
add_ln691_2_reg_950 <= _001_;
always @(posedge ap_clk)
add_ln691_1_reg_913 <= _000_;
always @(posedge ap_clk)
ap_CS_fsm <= _007_;
assign _043_ = _049_ ? 2'h2 : 2'h1;
assign _161_ = ap_CS_fsm == 1'h1;
function [38:0] _467_;
input [38:0] a;
input [1520:0] b;
input [38:0] s;
case (s)
39'b000000000000000000000000000000000000001:
_467_ = b[38:0];
39'b000000000000000000000000000000000000010:
_467_ = b[77:39];
39'b000000000000000000000000000000000000100:
_467_ = b[116:78];
39'b000000000000000000000000000000000001000:
_467_ = b[155:117];
39'b000000000000000000000000000000000010000:
_467_ = b[194:156];
39'b000000000000000000000000000000000100000:
_467_ = b[233:195];
39'b000000000000000000000000000000001000000:
_467_ = b[272:234];
39'b000000000000000000000000000000010000000:
_467_ = b[311:273];
39'b000000000000000000000000000000100000000:
_467_ = b[350:312];
39'b000000000000000000000000000001000000000:
_467_ = b[389:351];
39'b000000000000000000000000000010000000000:
_467_ = b[428:390];
39'b000000000000000000000000000100000000000:
_467_ = b[467:429];
39'b000000000000000000000000001000000000000:
_467_ = b[506:468];
39'b000000000000000000000000010000000000000:
_467_ = b[545:507];
39'b000000000000000000000000100000000000000:
_467_ = b[584:546];
39'b000000000000000000000001000000000000000:
_467_ = b[623:585];
39'b000000000000000000000010000000000000000:
_467_ = b[662:624];
39'b000000000000000000000100000000000000000:
_467_ = b[701:663];
39'b000000000000000000001000000000000000000:
_467_ = b[740:702];
39'b000000000000000000010000000000000000000:
_467_ = b[779:741];
39'b000000000000000000100000000000000000000:
_467_ = b[818:780];
39'b000000000000000001000000000000000000000:
_467_ = b[857:819];
39'b000000000000000010000000000000000000000:
_467_ = b[896:858];
39'b000000000000000100000000000000000000000:
_467_ = b[935:897];
39'b000000000000001000000000000000000000000:
_467_ = b[974:936];
39'b000000000000010000000000000000000000000:
_467_ = b[1013:975];
39'b000000000000100000000000000000000000000:
_467_ = b[1052:1014];
39'b000000000001000000000000000000000000000:
_467_ = b[1091:1053];
39'b000000000010000000000000000000000000000:
_467_ = b[1130:1092];
39'b000000000100000000000000000000000000000:
_467_ = b[1169:1131];
39'b000000001000000000000000000000000000000:
_467_ = b[1208:1170];
39'b000000010000000000000000000000000000000:
_467_ = b[1247:1209];
39'b000000100000000000000000000000000000000:
_467_ = b[1286:1248];
39'b000001000000000000000000000000000000000:
_467_ = b[1325:1287];
39'b000010000000000000000000000000000000000:
_467_ = b[1364:1326];
39'b000100000000000000000000000000000000000:
_467_ = b[1403:1365];
39'b001000000000000000000000000000000000000:
_467_ = b[1442:1404];
39'b010000000000000000000000000000000000000:
_467_ = b[1481:1443];
39'b100000000000000000000000000000000000000:
_467_ = b[1520:1482];
39'b000000000000000000000000000000000000000:
_467_ = a;
default:
_467_ = 39'bx;
endcase
endfunction
assign ap_NS_fsm = _467_(39'hxxxxxxxxxx, { 37'h0000000000, _043_, 1482'h00000000020000000008000000002000000000800000000200000000080000000020000000008000000002000000000800000000200000000080000000020000000008000000002000000000800000000200000000080000000020000000008000000002000000000800000000200000000080000000020000000008000000002000000000800000000200000000080000000020000000008000000002000000000800000000200000000080000000020000000000000000001 }, { _161_, _199_, _198_, _197_, _196_, _195_, _194_, _193_, _192_, _191_, _190_, _189_, _188_, _187_, _186_, _185_, _184_, _183_, _182_, _181_, _180_, _179_, _178_, _177_, _176_, _175_, _174_, _173_, _172_, _171_, _170_, _169_, _168_, _167_, _166_, _165_, _164_, _163_, _162_ });
assign _162_ = ap_CS_fsm == 39'h4000000000;
assign _163_ = ap_CS_fsm == 38'h2000000000;
assign _164_ = ap_CS_fsm == 37'h1000000000;
assign _165_ = ap_CS_fsm == 36'h800000000;
assign _166_ = ap_CS_fsm == 35'h400000000;
assign _167_ = ap_CS_fsm == 34'h200000000;
assign _168_ = ap_CS_fsm == 33'h100000000;
assign _169_ = ap_CS_fsm == 32'd2147483648;
assign _170_ = ap_CS_fsm == 31'h40000000;
assign _171_ = ap_CS_fsm == 30'h20000000;
assign _172_ = ap_CS_fsm == 29'h10000000;
assign _173_ = ap_CS_fsm == 28'h8000000;
assign _174_ = ap_CS_fsm == 27'h4000000;
assign _175_ = ap_CS_fsm == 26'h2000000;
assign _176_ = ap_CS_fsm == 25'h1000000;
assign _177_ = ap_CS_fsm == 24'h800000;
assign _178_ = ap_CS_fsm == 23'h400000;
assign _179_ = ap_CS_fsm == 22'h200000;
assign _180_ = ap_CS_fsm == 21'h100000;
assign _181_ = ap_CS_fsm == 20'h80000;
assign _182_ = ap_CS_fsm == 19'h40000;
assign _183_ = ap_CS_fsm == 18'h20000;
assign _184_ = ap_CS_fsm == 17'h10000;
assign _185_ = ap_CS_fsm == 16'h8000;
assign _186_ = ap_CS_fsm == 15'h4000;
assign _187_ = ap_CS_fsm == 14'h2000;
assign _188_ = ap_CS_fsm == 13'h1000;
assign _189_ = ap_CS_fsm == 12'h800;
assign _190_ = ap_CS_fsm == 11'h400;
assign _191_ = ap_CS_fsm == 10'h200;
assign _192_ = ap_CS_fsm == 9'h100;
assign _193_ = ap_CS_fsm == 8'h80;
assign _194_ = ap_CS_fsm == 7'h40;
assign _195_ = ap_CS_fsm == 6'h20;
assign _196_ = ap_CS_fsm == 5'h10;
assign _197_ = ap_CS_fsm == 4'h8;
assign _198_ = ap_CS_fsm == 3'h4;
assign _199_ = ap_CS_fsm == 2'h2;
assign op_31_ap_vld = ap_CS_fsm[38] ? 1'h1 : 1'h0;
assign ap_idle = _048_ ? 1'h1 : 1'h0;
assign _040_ = ap_CS_fsm[10] ? { tmp_reg_864[22], tmp_reg_864 } : sext_ln850_reg_869;
assign _037_ = ap_CS_fsm[12] ? select_ln353_fu_450_p3 : select_ln353_reg_881;
assign _036_ = ap_CS_fsm[22] ? select_ln353_2_fu_580_p3 : select_ln353_2_reg_955;
assign _035_ = ap_CS_fsm[17] ? select_ln353_1_fu_515_p3 : select_ln353_1_reg_918;
assign _032_ = ap_CS_fsm[2] ? grp_fu_320_p2 : ret_V_reg_794;
assign _033_ = ap_CS_fsm[36] ? select_ln1192_1_fu_744_p3 : select_ln1192_1_reg_1054;
assign _028_ = ap_CS_fsm[36] ? grp_fu_740_p2 : ret_V_21_reg_1049;
assign _034_ = ap_CS_fsm[34] ? select_ln1192_fu_732_p3 : select_ln1192_reg_1044;
assign _027_ = ap_CS_fsm[34] ? ret_V_20_fu_725_p3 : ret_V_20_reg_1039;
assign _029_ = ap_CS_fsm[31] ? grp_fu_682_p2[52:21] : ret_V_22_cast_reg_1027;
assign _025_ = ap_CS_fsm[31] ? grp_fu_682_p2 : ret_V_19_reg_1022;
assign _038_ = ap_CS_fsm[27] ? select_ln69_1_fu_655_p3 : select_ln69_1_reg_997;
assign _024_ = ap_CS_fsm[27] ? ret_V_18_fu_648_p3 : ret_V_18_reg_992;
assign _026_ = ap_CS_fsm[24] ? grp_fu_602_p2[32:1] : ret_V_20_cast_reg_980;
assign _022_ = ap_CS_fsm[24] ? grp_fu_602_p2 : ret_V_17_reg_975;
assign _023_ = ap_CS_fsm[19] ? grp_fu_537_p2[38:7] : ret_V_18_cast_reg_943;
assign _021_ = ap_CS_fsm[19] ? grp_fu_537_p2 : ret_V_16_reg_938;
assign _030_ = ap_CS_fsm[14] ? grp_fu_472_p2[33:2] : ret_V_7_cast_reg_906;
assign _020_ = ap_CS_fsm[14] ? grp_fu_472_p2 : ret_V_15_reg_901;
assign _042_ = ap_CS_fsm[9] ? grp_fu_403_p2[32:10] : tmp_reg_864;
assign _019_ = ap_CS_fsm[9] ? grp_fu_403_p2 : ret_V_14_reg_859;
assign _039_ = ap_CS_fsm[3] ? select_ln69_fu_344_p3 : select_ln69_reg_804;
assign _018_ = ap_CS_fsm[3] ? ret_V_13_fu_337_p3 : ret_V_13_reg_799;
assign _016_ = ap_CS_fsm[29] ? grp_fu_663_p2 : op_28_V_reg_1002;
assign _015_ = ap_CS_fsm[7] ? grp_fu_383_p2 : op_23_V_reg_839;
assign _014_ = ap_CS_fsm[1] ? icmp_ln851_fu_315_p2 : icmp_ln851_reg_789;
assign _013_ = ap_CS_fsm[30] ? icmp_ln851_4_fu_692_p2 : icmp_ln851_4_reg_1017;
assign _012_ = ap_CS_fsm[18] ? icmp_ln851_3_fu_547_p2 : icmp_ln851_3_reg_933;
assign _011_ = ap_CS_fsm[13] ? icmp_ln851_2_fu_482_p2 : icmp_ln851_2_reg_896;
assign _010_ = ap_CS_fsm[8] ? icmp_ln851_1_fu_413_p2 : icmp_ln851_1_reg_854;
assign _041_ = ap_CS_fsm[0] ? signbit_fu_309_p2 : signbit_reg_784;
assign _008_ = ap_CS_fsm[0] ? icmp_ln1494_fu_303_p2 : icmp_ln1494_reg_779;
assign _031_ = ap_CS_fsm[0] ? ret_V_12_fu_271_p2[4:3] : ret_V_cast_reg_767;
assign _017_ = ap_CS_fsm[0] ? ret_V_12_fu_271_p2[6:3] : ret_V_12_reg_762[6:3];
assign _009_ = ap_CS_fsm[0] ? icmp_ln1499_fu_253_p2 : icmp_ln1499_reg_757;
assign _005_ = ap_CS_fsm[5] ? grp_fu_375_p2 : add_ln69_1_reg_829;
assign _006_ = ap_CS_fsm[5] ? grp_fu_369_p2 : add_ln69_reg_824;
assign _004_ = _047_ ? grp_fu_432_p2 : add_ln691_reg_876;
assign _003_ = _046_ ? grp_fu_708_p2 : add_ln691_4_reg_1034;
assign _002_ = ap_CS_fsm[26] ? grp_fu_618_p2 : add_ln691_3_reg_987;
assign _001_ = _045_ ? grp_fu_563_p2 : add_ln691_2_reg_950;
assign _000_ = _044_ ? grp_fu_498_p2 : add_ln691_1_reg_913;
assign _007_ = ap_rst ? 39'h0000000001 : ap_NS_fsm;
assign icmp_ln1494_fu_303_p2 = _155_ ? 1'h1 : 1'h0;
assign icmp_ln1499_fu_253_p2 = _156_ ? 1'h1 : 1'h0;
assign icmp_ln851_1_fu_413_p2 = _157_ ? 1'h1 : 1'h0;
assign icmp_ln851_2_fu_482_p2 = _158_ ? 1'h1 : 1'h0;
assign icmp_ln851_3_fu_547_p2 = _159_ ? 1'h1 : 1'h0;
assign icmp_ln851_4_fu_692_p2 = _160_ ? 1'h1 : 1'h0;
assign icmp_ln851_fu_315_p2 = _051_ ? 1'h1 : 1'h0;
assign ret_V_13_fu_337_p3 = ret_V_12_reg_762[6] ? select_ln850_fu_332_p3 : ret_V_cast_reg_767;
assign ret_V_18_fu_648_p3 = ret_V_17_reg_975[33] ? select_ln850_4_fu_642_p3 : ret_V_20_cast_reg_980;
assign ret_V_20_fu_725_p3 = ret_V_19_reg_1022[53] ? select_ln850_5_fu_720_p3 : ret_V_22_cast_reg_1027;
assign select_ln1192_1_fu_744_p3 = op_19 ? 32'd4294967295 : 32'd0;
assign select_ln1192_fu_732_p3 = op_18 ? 32'd4294967295 : 32'd0;
assign select_ln353_1_fu_515_p3 = ret_V_15_reg_901[34] ? select_ln850_2_fu_510_p3 : ret_V_7_cast_reg_906;
assign select_ln353_2_fu_580_p3 = ret_V_16_reg_938[39] ? select_ln850_3_fu_575_p3 : ret_V_18_cast_reg_943;
assign select_ln353_fu_450_p3 = ret_V_14_reg_859[32] ? select_ln850_1_fu_445_p3 : sext_ln850_reg_869;
assign select_ln69_1_fu_655_p3 = op_16_V_fu_627_p2 ? 32'd4294967295 : 32'd0;
assign select_ln69_fu_344_p3 = op_11 ? 2'h3 : 2'h0;
assign select_ln850_1_fu_445_p3 = icmp_ln851_1_reg_854 ? add_ln691_reg_876 : sext_ln850_reg_869;
assign select_ln850_2_fu_510_p3 = icmp_ln851_2_reg_896 ? add_ln691_1_reg_913 : ret_V_7_cast_reg_906;
assign select_ln850_3_fu_575_p3 = icmp_ln851_3_reg_933 ? add_ln691_2_reg_950 : ret_V_18_cast_reg_943;
assign select_ln850_4_fu_642_p3 = op_15[0] ? add_ln691_3_reg_987 : ret_V_20_cast_reg_980;
assign select_ln850_5_fu_720_p3 = icmp_ln851_4_reg_1017 ? add_ln691_4_reg_1034 : ret_V_22_cast_reg_1027;
assign select_ln850_fu_332_p3 = icmp_ln851_reg_789 ? ret_V_cast_reg_767 : ret_V_reg_794;
assign signbit_fu_309_p2 = _052_ ? 1'h1 : 1'h0;
assign ap_CS_fsm_state1 = ap_CS_fsm[0];
assign ap_CS_fsm_state10 = ap_CS_fsm[9];
assign ap_CS_fsm_state11 = ap_CS_fsm[10];
assign ap_CS_fsm_state12 = ap_CS_fsm[11];
assign ap_CS_fsm_state13 = ap_CS_fsm[12];
assign ap_CS_fsm_state14 = ap_CS_fsm[13];
assign ap_CS_fsm_state15 = ap_CS_fsm[14];
assign ap_CS_fsm_state16 = ap_CS_fsm[15];
assign ap_CS_fsm_state17 = ap_CS_fsm[16];
assign ap_CS_fsm_state18 = ap_CS_fsm[17];
assign ap_CS_fsm_state19 = ap_CS_fsm[18];
assign ap_CS_fsm_state2 = ap_CS_fsm[1];
assign ap_CS_fsm_state20 = ap_CS_fsm[19];
assign ap_CS_fsm_state21 = ap_CS_fsm[20];
assign ap_CS_fsm_state22 = ap_CS_fsm[21];
assign ap_CS_fsm_state23 = ap_CS_fsm[22];
assign ap_CS_fsm_state24 = ap_CS_fsm[23];
assign ap_CS_fsm_state25 = ap_CS_fsm[24];
assign ap_CS_fsm_state26 = ap_CS_fsm[25];
assign ap_CS_fsm_state27 = ap_CS_fsm[26];
assign ap_CS_fsm_state28 = ap_CS_fsm[27];
assign ap_CS_fsm_state29 = ap_CS_fsm[28];
assign ap_CS_fsm_state3 = ap_CS_fsm[2];
assign ap_CS_fsm_state30 = ap_CS_fsm[29];
assign ap_CS_fsm_state31 = ap_CS_fsm[30];
assign ap_CS_fsm_state32 = ap_CS_fsm[31];
assign ap_CS_fsm_state33 = ap_CS_fsm[32];
assign ap_CS_fsm_state34 = ap_CS_fsm[33];
assign ap_CS_fsm_state35 = ap_CS_fsm[34];
assign ap_CS_fsm_state36 = ap_CS_fsm[35];
assign ap_CS_fsm_state37 = ap_CS_fsm[36];
assign ap_CS_fsm_state38 = ap_CS_fsm[37];
assign ap_CS_fsm_state39 = ap_CS_fsm[38];
assign ap_CS_fsm_state4 = ap_CS_fsm[3];
assign ap_CS_fsm_state5 = ap_CS_fsm[4];
assign ap_CS_fsm_state6 = ap_CS_fsm[5];
assign ap_CS_fsm_state7 = ap_CS_fsm[6];
assign ap_CS_fsm_state8 = ap_CS_fsm[7];
assign ap_CS_fsm_state9 = ap_CS_fsm[8];
assign ap_done = op_31_ap_vld;
assign ap_ready = op_31_ap_vld;
assign grp_fu_369_p0 = { op_0[3], op_0, icmp_ln1499_reg_757 };
assign grp_fu_369_p1 = { ret_V_13_reg_799[1], ret_V_13_reg_799[1], ret_V_13_reg_799[1], ret_V_13_reg_799[1], ret_V_13_reg_799 };
assign grp_fu_375_p0 = { 1'h0, icmp_ln1494_reg_779 };
assign grp_fu_383_p0 = { add_ln69_1_reg_829[1], add_ln69_1_reg_829[1], add_ln69_1_reg_829[1], add_ln69_1_reg_829[1], add_ln69_1_reg_829 };
assign grp_fu_403_p0 = { op_23_V_reg_839[5], op_23_V_reg_839[5], op_23_V_reg_839[5], op_23_V_reg_839[5], op_23_V_reg_839[5], op_23_V_reg_839[5], op_23_V_reg_839[5], op_23_V_reg_839[5], op_23_V_reg_839[5], op_23_V_reg_839[5], op_23_V_reg_839[5], op_23_V_reg_839[5], op_23_V_reg_839[5], op_23_V_reg_839[5], op_23_V_reg_839[5], op_23_V_reg_839[5], op_23_V_reg_839[5], op_23_V_reg_839, 10'h000 };
assign grp_fu_403_p1 = { op_12[31], op_12 };
assign grp_fu_432_p0 = { tmp_reg_864[22], tmp_reg_864 };
assign grp_fu_472_p0 = { select_ln353_reg_881[23], select_ln353_reg_881[23], select_ln353_reg_881[23], select_ln353_reg_881[23], select_ln353_reg_881[23], select_ln353_reg_881[23], select_ln353_reg_881[23], select_ln353_reg_881[23], select_ln353_reg_881[23], select_ln353_reg_881, 2'h0 };
assign grp_fu_472_p1 = { op_13[31], op_13[31], op_13[31], op_13 };
assign grp_fu_537_p0 = { select_ln353_1_reg_918[31], select_ln353_1_reg_918, 7'h00 };
assign grp_fu_537_p1 = { op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14 };
assign grp_fu_602_p0 = { select_ln353_2_reg_955[31], select_ln353_2_reg_955, 1'h0 };
assign grp_fu_602_p1 = { op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15 };
assign grp_fu_682_p0 = { op_28_V_reg_1002[31], op_28_V_reg_1002, 21'h000000 };
assign grp_fu_682_p1 = { op_17[31], op_17[31], op_17[31], op_17[31], op_17[31], op_17[31], op_17[31], op_17[31], op_17[31], op_17[31], op_17[31], op_17[31], op_17[31], op_17[31], op_17[31], op_17[31], op_17[31], op_17[31], op_17[31], op_17[31], op_17[31], op_17[31], op_17 };
assign op_20_V_fu_352_p3 = { op_0, icmp_ln1499_reg_757 };
assign op_31 = grp_fu_752_p2;
assign op_4_V_fu_233_p3 = { op_2, 6'h00 };
assign p_Result_1_fu_438_p3 = ret_V_14_reg_859[32];
assign p_Result_2_fu_503_p3 = ret_V_15_reg_901[34];
assign p_Result_3_fu_568_p3 = ret_V_16_reg_938[39];
assign p_Result_4_fu_632_p3 = ret_V_17_reg_975[33];
assign p_Result_5_fu_713_p3 = ret_V_19_reg_1022[53];
assign p_Result_s_fu_325_p3 = ret_V_12_reg_762[6];
assign rhs_2_fu_392_p3 = { op_23_V_reg_839, 10'h000 };
assign rhs_3_fu_526_p3 = { select_ln353_1_reg_918, 7'h00 };
assign rhs_4_fu_591_p3 = { select_ln353_2_reg_955, 1'h0 };
assign rhs_6_fu_671_p3 = { op_28_V_reg_1002, 21'h000000 };
assign rhs_fu_263_p3 = { op_5, 3'h0 };
assign sext_ln1192_fu_388_p0 = op_12;
assign sext_ln1494_fu_299_p1 = { op_3[3], op_3, 3'h0 };
assign sext_ln1499_fu_249_p0 = op_3;
assign sext_ln1499_fu_249_p1 = { op_3[3], op_3 };
assign sext_ln703_1_fu_457_p0 = op_13;
assign sext_ln703_2_fu_522_p0 = op_14;
assign sext_ln703_3_fu_587_p0 = op_15;
assign sext_ln703_4_fu_667_p0 = op_17;
assign sext_ln703_fu_259_p0 = op_3;
assign sext_ln703_fu_259_p1 = { op_3[3], op_3[3], op_3[3], op_3 };
assign sext_ln850_fu_429_p1 = { tmp_reg_864[22], tmp_reg_864 };
assign shl_ln728_2_fu_291_p1 = op_3;
assign shl_ln728_2_fu_291_p3 = { op_3, 3'h0 };
assign shl_ln_fu_241_p3 = { op_2, 3'h0 };
assign tmp_3_fu_461_p3 = { select_ln353_reg_881, 2'h0 };
assign trunc_ln1195_fu_623_p1 = op_10[0];
assign trunc_ln851_1_fu_409_p0 = op_12;
assign trunc_ln851_1_fu_409_p1 = op_12[9:0];
assign trunc_ln851_2_fu_478_p0 = op_13;
assign trunc_ln851_2_fu_478_p1 = op_13[1:0];
assign trunc_ln851_3_fu_543_p0 = op_14;
assign trunc_ln851_3_fu_543_p1 = op_14[6:0];
assign trunc_ln851_4_fu_639_p0 = op_15;
assign trunc_ln851_4_fu_639_p1 = op_15[0];
assign trunc_ln851_5_fu_688_p0 = op_17;
assign trunc_ln851_5_fu_688_p1 = op_17[20:0];
assign trunc_ln851_fu_287_p1 = ret_V_12_fu_271_p2[2:0];
assign \add_6s_6s_6_2_1_U2.top_add_6s_6s_6_2_1_Adder_1_U.ain_s0  = \add_6s_6s_6_2_1_U2.top_add_6s_6s_6_2_1_Adder_1_U.a ;
assign \add_6s_6s_6_2_1_U2.top_add_6s_6s_6_2_1_Adder_1_U.bin_s0  = \add_6s_6s_6_2_1_U2.top_add_6s_6s_6_2_1_Adder_1_U.b ;
assign \add_6s_6s_6_2_1_U2.top_add_6s_6s_6_2_1_Adder_1_U.s  = { \add_6s_6s_6_2_1_U2.top_add_6s_6s_6_2_1_Adder_1_U.fas_s2 , \add_6s_6s_6_2_1_U2.top_add_6s_6s_6_2_1_Adder_1_U.sum_s1  };
assign \add_6s_6s_6_2_1_U2.top_add_6s_6s_6_2_1_Adder_1_U.u2.a  = \add_6s_6s_6_2_1_U2.top_add_6s_6s_6_2_1_Adder_1_U.ain_s1 ;
assign \add_6s_6s_6_2_1_U2.top_add_6s_6s_6_2_1_Adder_1_U.u2.b  = \add_6s_6s_6_2_1_U2.top_add_6s_6s_6_2_1_Adder_1_U.bin_s1 ;
assign \add_6s_6s_6_2_1_U2.top_add_6s_6s_6_2_1_Adder_1_U.u2.cin  = \add_6s_6s_6_2_1_U2.top_add_6s_6s_6_2_1_Adder_1_U.carry_s1 ;
assign \add_6s_6s_6_2_1_U2.top_add_6s_6s_6_2_1_Adder_1_U.facout_s2  = \add_6s_6s_6_2_1_U2.top_add_6s_6s_6_2_1_Adder_1_U.u2.cout ;
assign \add_6s_6s_6_2_1_U2.top_add_6s_6s_6_2_1_Adder_1_U.fas_s2  = \add_6s_6s_6_2_1_U2.top_add_6s_6s_6_2_1_Adder_1_U.u2.s ;
assign \add_6s_6s_6_2_1_U2.top_add_6s_6s_6_2_1_Adder_1_U.u1.a  = \add_6s_6s_6_2_1_U2.top_add_6s_6s_6_2_1_Adder_1_U.a [2:0];
assign \add_6s_6s_6_2_1_U2.top_add_6s_6s_6_2_1_Adder_1_U.u1.b  = \add_6s_6s_6_2_1_U2.top_add_6s_6s_6_2_1_Adder_1_U.b [2:0];
assign \add_6s_6s_6_2_1_U2.top_add_6s_6s_6_2_1_Adder_1_U.u1.cin  = 1'h0;
assign \add_6s_6s_6_2_1_U2.top_add_6s_6s_6_2_1_Adder_1_U.facout_s1  = \add_6s_6s_6_2_1_U2.top_add_6s_6s_6_2_1_Adder_1_U.u1.cout ;
assign \add_6s_6s_6_2_1_U2.top_add_6s_6s_6_2_1_Adder_1_U.fas_s1  = \add_6s_6s_6_2_1_U2.top_add_6s_6s_6_2_1_Adder_1_U.u1.s ;
assign \add_6s_6s_6_2_1_U2.top_add_6s_6s_6_2_1_Adder_1_U.a  = \add_6s_6s_6_2_1_U2.din0 ;
assign \add_6s_6s_6_2_1_U2.top_add_6s_6s_6_2_1_Adder_1_U.b  = \add_6s_6s_6_2_1_U2.din1 ;
assign \add_6s_6s_6_2_1_U2.top_add_6s_6s_6_2_1_Adder_1_U.ce  = \add_6s_6s_6_2_1_U2.ce ;
assign \add_6s_6s_6_2_1_U2.top_add_6s_6s_6_2_1_Adder_1_U.clk  = \add_6s_6s_6_2_1_U2.clk ;
assign \add_6s_6s_6_2_1_U2.top_add_6s_6s_6_2_1_Adder_1_U.reset  = \add_6s_6s_6_2_1_U2.reset ;
assign \add_6s_6s_6_2_1_U2.dout  = \add_6s_6s_6_2_1_U2.top_add_6s_6s_6_2_1_Adder_1_U.s ;
assign \add_6s_6s_6_2_1_U2.ce  = 1'h1;
assign \add_6s_6s_6_2_1_U2.clk  = ap_clk;
assign \add_6s_6s_6_2_1_U2.din0  = { op_0[3], op_0, icmp_ln1499_reg_757 };
assign \add_6s_6s_6_2_1_U2.din1  = { ret_V_13_reg_799[1], ret_V_13_reg_799[1], ret_V_13_reg_799[1], ret_V_13_reg_799[1], ret_V_13_reg_799 };
assign grp_fu_369_p2 = \add_6s_6s_6_2_1_U2.dout ;
assign \add_6s_6s_6_2_1_U2.reset  = ap_rst;
assign \add_6s_6ns_6_2_1_U4.top_add_6s_6ns_6_2_1_Adder_2_U.ain_s0  = \add_6s_6ns_6_2_1_U4.top_add_6s_6ns_6_2_1_Adder_2_U.a ;
assign \add_6s_6ns_6_2_1_U4.top_add_6s_6ns_6_2_1_Adder_2_U.bin_s0  = \add_6s_6ns_6_2_1_U4.top_add_6s_6ns_6_2_1_Adder_2_U.b ;
assign \add_6s_6ns_6_2_1_U4.top_add_6s_6ns_6_2_1_Adder_2_U.s  = { \add_6s_6ns_6_2_1_U4.top_add_6s_6ns_6_2_1_Adder_2_U.fas_s2 , \add_6s_6ns_6_2_1_U4.top_add_6s_6ns_6_2_1_Adder_2_U.sum_s1  };
assign \add_6s_6ns_6_2_1_U4.top_add_6s_6ns_6_2_1_Adder_2_U.u2.a  = \add_6s_6ns_6_2_1_U4.top_add_6s_6ns_6_2_1_Adder_2_U.ain_s1 ;
assign \add_6s_6ns_6_2_1_U4.top_add_6s_6ns_6_2_1_Adder_2_U.u2.b  = \add_6s_6ns_6_2_1_U4.top_add_6s_6ns_6_2_1_Adder_2_U.bin_s1 ;
assign \add_6s_6ns_6_2_1_U4.top_add_6s_6ns_6_2_1_Adder_2_U.u2.cin  = \add_6s_6ns_6_2_1_U4.top_add_6s_6ns_6_2_1_Adder_2_U.carry_s1 ;
assign \add_6s_6ns_6_2_1_U4.top_add_6s_6ns_6_2_1_Adder_2_U.facout_s2  = \add_6s_6ns_6_2_1_U4.top_add_6s_6ns_6_2_1_Adder_2_U.u2.cout ;
assign \add_6s_6ns_6_2_1_U4.top_add_6s_6ns_6_2_1_Adder_2_U.fas_s2  = \add_6s_6ns_6_2_1_U4.top_add_6s_6ns_6_2_1_Adder_2_U.u2.s ;
assign \add_6s_6ns_6_2_1_U4.top_add_6s_6ns_6_2_1_Adder_2_U.u1.a  = \add_6s_6ns_6_2_1_U4.top_add_6s_6ns_6_2_1_Adder_2_U.a [2:0];
assign \add_6s_6ns_6_2_1_U4.top_add_6s_6ns_6_2_1_Adder_2_U.u1.b  = \add_6s_6ns_6_2_1_U4.top_add_6s_6ns_6_2_1_Adder_2_U.b [2:0];
assign \add_6s_6ns_6_2_1_U4.top_add_6s_6ns_6_2_1_Adder_2_U.u1.cin  = 1'h0;
assign \add_6s_6ns_6_2_1_U4.top_add_6s_6ns_6_2_1_Adder_2_U.facout_s1  = \add_6s_6ns_6_2_1_U4.top_add_6s_6ns_6_2_1_Adder_2_U.u1.cout ;
assign \add_6s_6ns_6_2_1_U4.top_add_6s_6ns_6_2_1_Adder_2_U.fas_s1  = \add_6s_6ns_6_2_1_U4.top_add_6s_6ns_6_2_1_Adder_2_U.u1.s ;
assign \add_6s_6ns_6_2_1_U4.top_add_6s_6ns_6_2_1_Adder_2_U.a  = \add_6s_6ns_6_2_1_U4.din0 ;
assign \add_6s_6ns_6_2_1_U4.top_add_6s_6ns_6_2_1_Adder_2_U.b  = \add_6s_6ns_6_2_1_U4.din1 ;
assign \add_6s_6ns_6_2_1_U4.top_add_6s_6ns_6_2_1_Adder_2_U.ce  = \add_6s_6ns_6_2_1_U4.ce ;
assign \add_6s_6ns_6_2_1_U4.top_add_6s_6ns_6_2_1_Adder_2_U.clk  = \add_6s_6ns_6_2_1_U4.clk ;
assign \add_6s_6ns_6_2_1_U4.top_add_6s_6ns_6_2_1_Adder_2_U.reset  = \add_6s_6ns_6_2_1_U4.reset ;
assign \add_6s_6ns_6_2_1_U4.dout  = \add_6s_6ns_6_2_1_U4.top_add_6s_6ns_6_2_1_Adder_2_U.s ;
assign \add_6s_6ns_6_2_1_U4.ce  = 1'h1;
assign \add_6s_6ns_6_2_1_U4.clk  = ap_clk;
assign \add_6s_6ns_6_2_1_U4.din0  = { add_ln69_1_reg_829[1], add_ln69_1_reg_829[1], add_ln69_1_reg_829[1], add_ln69_1_reg_829[1], add_ln69_1_reg_829 };
assign \add_6s_6ns_6_2_1_U4.din1  = add_ln69_reg_824;
assign grp_fu_383_p2 = \add_6s_6ns_6_2_1_U4.dout ;
assign \add_6s_6ns_6_2_1_U4.reset  = ap_rst;
assign \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.ain_s0  = \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.a ;
assign \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.bin_s0  = \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.b ;
assign \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.s  = { \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.fas_s2 , \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.sum_s1  };
assign \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.u2.a  = \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.ain_s1 ;
assign \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.u2.b  = \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.bin_s1 ;
assign \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.u2.cin  = \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.carry_s1 ;
assign \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.facout_s2  = \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.u2.cout ;
assign \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.fas_s2  = \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.u2.s ;
assign \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.u1.a  = \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.a [26:0];
assign \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.u1.b  = \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.b [26:0];
assign \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.u1.cin  = 1'h0;
assign \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.facout_s1  = \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.u1.cout ;
assign \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.fas_s1  = \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.u1.s ;
assign \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.a  = \add_54s_54s_54_2_1_U14.din0 ;
assign \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.b  = \add_54s_54s_54_2_1_U14.din1 ;
assign \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.ce  = \add_54s_54s_54_2_1_U14.ce ;
assign \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.clk  = \add_54s_54s_54_2_1_U14.clk ;
assign \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.reset  = \add_54s_54s_54_2_1_U14.reset ;
assign \add_54s_54s_54_2_1_U14.dout  = \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.s ;
assign \add_54s_54s_54_2_1_U14.ce  = 1'h1;
assign \add_54s_54s_54_2_1_U14.clk  = ap_clk;
assign \add_54s_54s_54_2_1_U14.din0  = { op_28_V_reg_1002[31], op_28_V_reg_1002, 21'h000000 };
assign \add_54s_54s_54_2_1_U14.din1  = { op_17[31], op_17[31], op_17[31], op_17[31], op_17[31], op_17[31], op_17[31], op_17[31], op_17[31], op_17[31], op_17[31], op_17[31], op_17[31], op_17[31], op_17[31], op_17[31], op_17[31], op_17[31], op_17[31], op_17[31], op_17[31], op_17[31], op_17 };
assign grp_fu_682_p2 = \add_54s_54s_54_2_1_U14.dout ;
assign \add_54s_54s_54_2_1_U14.reset  = ap_rst;
assign \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.ain_s0  = \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.a ;
assign \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.bin_s0  = \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.b ;
assign \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.s  = { \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.fas_s2 , \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.sum_s1  };
assign \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.u2.a  = \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.ain_s1 ;
assign \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.u2.b  = \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.bin_s1 ;
assign \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.u2.cin  = \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.carry_s1 ;
assign \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.facout_s2  = \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.u2.cout ;
assign \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.fas_s2  = \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.u2.s ;
assign \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.u1.a  = \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.a [19:0];
assign \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.u1.b  = \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.b [19:0];
assign \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.u1.cin  = 1'h0;
assign \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.facout_s1  = \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.u1.cout ;
assign \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.fas_s1  = \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.u1.s ;
assign \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.a  = \add_40s_40s_40_2_1_U9.din0 ;
assign \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.b  = \add_40s_40s_40_2_1_U9.din1 ;
assign \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.ce  = \add_40s_40s_40_2_1_U9.ce ;
assign \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.clk  = \add_40s_40s_40_2_1_U9.clk ;
assign \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.reset  = \add_40s_40s_40_2_1_U9.reset ;
assign \add_40s_40s_40_2_1_U9.dout  = \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.s ;
assign \add_40s_40s_40_2_1_U9.ce  = 1'h1;
assign \add_40s_40s_40_2_1_U9.clk  = ap_clk;
assign \add_40s_40s_40_2_1_U9.din0  = { select_ln353_1_reg_918[31], select_ln353_1_reg_918, 7'h00 };
assign \add_40s_40s_40_2_1_U9.din1  = { op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14 };
assign grp_fu_537_p2 = \add_40s_40s_40_2_1_U9.dout ;
assign \add_40s_40s_40_2_1_U9.reset  = ap_rst;
assign \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.ain_s0  = \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.a ;
assign \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.bin_s0  = \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.b ;
assign \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.s  = { \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.fas_s2 , \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.sum_s1  };
assign \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.u2.a  = \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.ain_s1 ;
assign \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.u2.b  = \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.bin_s1 ;
assign \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.u2.cin  = \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.carry_s1 ;
assign \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.facout_s2  = \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.u2.cout ;
assign \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.fas_s2  = \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.u2.s ;
assign \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.u1.a  = \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.a [16:0];
assign \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.u1.b  = \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.b [16:0];
assign \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.u1.cin  = 1'h0;
assign \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.facout_s1  = \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.u1.cout ;
assign \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.fas_s1  = \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.u1.s ;
assign \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.a  = \add_35s_35s_35_2_1_U7.din0 ;
assign \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.b  = \add_35s_35s_35_2_1_U7.din1 ;
assign \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.ce  = \add_35s_35s_35_2_1_U7.ce ;
assign \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.clk  = \add_35s_35s_35_2_1_U7.clk ;
assign \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.reset  = \add_35s_35s_35_2_1_U7.reset ;
assign \add_35s_35s_35_2_1_U7.dout  = \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.s ;
assign \add_35s_35s_35_2_1_U7.ce  = 1'h1;
assign \add_35s_35s_35_2_1_U7.clk  = ap_clk;
assign \add_35s_35s_35_2_1_U7.din0  = { select_ln353_reg_881[23], select_ln353_reg_881[23], select_ln353_reg_881[23], select_ln353_reg_881[23], select_ln353_reg_881[23], select_ln353_reg_881[23], select_ln353_reg_881[23], select_ln353_reg_881[23], select_ln353_reg_881[23], select_ln353_reg_881, 2'h0 };
assign \add_35s_35s_35_2_1_U7.din1  = { op_13[31], op_13[31], op_13[31], op_13 };
assign grp_fu_472_p2 = \add_35s_35s_35_2_1_U7.dout ;
assign \add_35s_35s_35_2_1_U7.reset  = ap_rst;
assign \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.ain_s0  = \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.a ;
assign \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.bin_s0  = \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.b ;
assign \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.s  = { \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.fas_s2 , \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.sum_s1  };
assign \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.u2.a  = \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.ain_s1 ;
assign \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.u2.b  = \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.bin_s1 ;
assign \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.u2.cin  = \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.carry_s1 ;
assign \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.facout_s2  = \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.u2.cout ;
assign \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.fas_s2  = \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.u2.s ;
assign \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.u1.a  = \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.a [16:0];
assign \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.u1.b  = \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.b [16:0];
assign \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.u1.cin  = 1'h0;
assign \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.facout_s1  = \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.u1.cout ;
assign \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.fas_s1  = \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.u1.s ;
assign \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.a  = \add_34s_34s_34_2_1_U11.din0 ;
assign \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.b  = \add_34s_34s_34_2_1_U11.din1 ;
assign \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.ce  = \add_34s_34s_34_2_1_U11.ce ;
assign \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.clk  = \add_34s_34s_34_2_1_U11.clk ;
assign \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.reset  = \add_34s_34s_34_2_1_U11.reset ;
assign \add_34s_34s_34_2_1_U11.dout  = \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.s ;
assign \add_34s_34s_34_2_1_U11.ce  = 1'h1;
assign \add_34s_34s_34_2_1_U11.clk  = ap_clk;
assign \add_34s_34s_34_2_1_U11.din0  = { select_ln353_2_reg_955[31], select_ln353_2_reg_955, 1'h0 };
assign \add_34s_34s_34_2_1_U11.din1  = { op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15 };
assign grp_fu_602_p2 = \add_34s_34s_34_2_1_U11.dout ;
assign \add_34s_34s_34_2_1_U11.reset  = ap_rst;
assign \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.ain_s0  = \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.a ;
assign \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.bin_s0  = \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.b ;
assign \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.s  = { \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.fas_s2 , \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.sum_s1  };
assign \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.u2.a  = \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.ain_s1 ;
assign \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.u2.b  = \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.bin_s1 ;
assign \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.u2.cin  = \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.carry_s1 ;
assign \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.facout_s2  = \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.u2.cout ;
assign \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.fas_s2  = \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.u2.s ;
assign \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.u1.a  = \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.a [15:0];
assign \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.u1.b  = \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.b [15:0];
assign \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.u1.cin  = 1'h0;
assign \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.facout_s1  = \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.u1.cout ;
assign \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.fas_s1  = \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.u1.s ;
assign \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.a  = \add_33s_33s_33_2_1_U5.din0 ;
assign \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.b  = \add_33s_33s_33_2_1_U5.din1 ;
assign \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.ce  = \add_33s_33s_33_2_1_U5.ce ;
assign \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.clk  = \add_33s_33s_33_2_1_U5.clk ;
assign \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.reset  = \add_33s_33s_33_2_1_U5.reset ;
assign \add_33s_33s_33_2_1_U5.dout  = \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.s ;
assign \add_33s_33s_33_2_1_U5.ce  = 1'h1;
assign \add_33s_33s_33_2_1_U5.clk  = ap_clk;
assign \add_33s_33s_33_2_1_U5.din0  = { op_23_V_reg_839[5], op_23_V_reg_839[5], op_23_V_reg_839[5], op_23_V_reg_839[5], op_23_V_reg_839[5], op_23_V_reg_839[5], op_23_V_reg_839[5], op_23_V_reg_839[5], op_23_V_reg_839[5], op_23_V_reg_839[5], op_23_V_reg_839[5], op_23_V_reg_839[5], op_23_V_reg_839[5], op_23_V_reg_839[5], op_23_V_reg_839[5], op_23_V_reg_839[5], op_23_V_reg_839[5], op_23_V_reg_839, 10'h000 };
assign \add_33s_33s_33_2_1_U5.din1  = { op_12[31], op_12 };
assign grp_fu_403_p2 = \add_33s_33s_33_2_1_U5.dout ;
assign \add_33s_33s_33_2_1_U5.reset  = ap_rst;
assign \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s0  = \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.a ;
assign \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s0  = \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.b ;
assign \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.s  = { \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s2 , \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.sum_s1  };
assign \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.a  = \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s1 ;
assign \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.b  = \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s1 ;
assign \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cin  = \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.carry_s1 ;
assign \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s2  = \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cout ;
assign \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s2  = \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.s ;
assign \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.a  = \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.a [15:0];
assign \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.b  = \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.b [15:0];
assign \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cin  = 1'h0;
assign \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s1  = \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cout ;
assign \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s1  = \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.s ;
assign \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.a  = \add_32ns_32ns_32_2_1_U8.din0 ;
assign \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.b  = \add_32ns_32ns_32_2_1_U8.din1 ;
assign \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  = \add_32ns_32ns_32_2_1_U8.ce ;
assign \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.clk  = \add_32ns_32ns_32_2_1_U8.clk ;
assign \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.reset  = \add_32ns_32ns_32_2_1_U8.reset ;
assign \add_32ns_32ns_32_2_1_U8.dout  = \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.s ;
assign \add_32ns_32ns_32_2_1_U8.ce  = 1'h1;
assign \add_32ns_32ns_32_2_1_U8.clk  = ap_clk;
assign \add_32ns_32ns_32_2_1_U8.din0  = ret_V_7_cast_reg_906;
assign \add_32ns_32ns_32_2_1_U8.din1  = 32'd1;
assign grp_fu_498_p2 = \add_32ns_32ns_32_2_1_U8.dout ;
assign \add_32ns_32ns_32_2_1_U8.reset  = ap_rst;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s0  = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.a ;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s0  = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.b ;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.s  = { \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s2 , \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.sum_s1  };
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.a  = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s1 ;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.b  = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s1 ;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cin  = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.carry_s1 ;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s2  = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cout ;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s2  = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.s ;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.a  = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.a [15:0];
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.b  = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.b [15:0];
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cin  = 1'h0;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s1  = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cout ;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s1  = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.s ;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.a  = \add_32ns_32ns_32_2_1_U17.din0 ;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.b  = \add_32ns_32ns_32_2_1_U17.din1 ;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  = \add_32ns_32ns_32_2_1_U17.ce ;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.clk  = \add_32ns_32ns_32_2_1_U17.clk ;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.reset  = \add_32ns_32ns_32_2_1_U17.reset ;
assign \add_32ns_32ns_32_2_1_U17.dout  = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.s ;
assign \add_32ns_32ns_32_2_1_U17.ce  = 1'h1;
assign \add_32ns_32ns_32_2_1_U17.clk  = ap_clk;
assign \add_32ns_32ns_32_2_1_U17.din0  = ret_V_21_reg_1049;
assign \add_32ns_32ns_32_2_1_U17.din1  = select_ln1192_1_reg_1054;
assign grp_fu_752_p2 = \add_32ns_32ns_32_2_1_U17.dout ;
assign \add_32ns_32ns_32_2_1_U17.reset  = ap_rst;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s0  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.a ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s0  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.b ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.s  = { \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s2 , \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.sum_s1  };
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.a  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s1 ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.b  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s1 ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cin  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.carry_s1 ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s2  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cout ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s2  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.s ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.a  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.a [15:0];
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.b  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.b [15:0];
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cin  = 1'h0;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s1  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cout ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s1  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.s ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.a  = \add_32ns_32ns_32_2_1_U16.din0 ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.b  = \add_32ns_32ns_32_2_1_U16.din1 ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  = \add_32ns_32ns_32_2_1_U16.ce ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.clk  = \add_32ns_32ns_32_2_1_U16.clk ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.reset  = \add_32ns_32ns_32_2_1_U16.reset ;
assign \add_32ns_32ns_32_2_1_U16.dout  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.s ;
assign \add_32ns_32ns_32_2_1_U16.ce  = 1'h1;
assign \add_32ns_32ns_32_2_1_U16.clk  = ap_clk;
assign \add_32ns_32ns_32_2_1_U16.din0  = ret_V_20_reg_1039;
assign \add_32ns_32ns_32_2_1_U16.din1  = select_ln1192_reg_1044;
assign grp_fu_740_p2 = \add_32ns_32ns_32_2_1_U16.dout ;
assign \add_32ns_32ns_32_2_1_U16.reset  = ap_rst;
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s0  = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.a ;
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s0  = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.b ;
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.s  = { \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s2 , \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.sum_s1  };
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.a  = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s1 ;
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.b  = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s1 ;
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cin  = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.carry_s1 ;
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s2  = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cout ;
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s2  = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.s ;
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.a  = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.a [15:0];
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.b  = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.b [15:0];
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cin  = 1'h0;
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s1  = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cout ;
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s1  = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.s ;
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.a  = \add_32ns_32ns_32_2_1_U15.din0 ;
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.b  = \add_32ns_32ns_32_2_1_U15.din1 ;
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  = \add_32ns_32ns_32_2_1_U15.ce ;
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.clk  = \add_32ns_32ns_32_2_1_U15.clk ;
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.reset  = \add_32ns_32ns_32_2_1_U15.reset ;
assign \add_32ns_32ns_32_2_1_U15.dout  = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.s ;
assign \add_32ns_32ns_32_2_1_U15.ce  = 1'h1;
assign \add_32ns_32ns_32_2_1_U15.clk  = ap_clk;
assign \add_32ns_32ns_32_2_1_U15.din0  = ret_V_22_cast_reg_1027;
assign \add_32ns_32ns_32_2_1_U15.din1  = 32'd1;
assign grp_fu_708_p2 = \add_32ns_32ns_32_2_1_U15.dout ;
assign \add_32ns_32ns_32_2_1_U15.reset  = ap_rst;
assign \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s0  = \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.a ;
assign \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s0  = \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.b ;
assign \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.s  = { \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s2 , \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.sum_s1  };
assign \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.a  = \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s1 ;
assign \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.b  = \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s1 ;
assign \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cin  = \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.carry_s1 ;
assign \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s2  = \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cout ;
assign \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s2  = \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.s ;
assign \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.a  = \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.a [15:0];
assign \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.b  = \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.b [15:0];
assign \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cin  = 1'h0;
assign \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s1  = \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cout ;
assign \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s1  = \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.s ;
assign \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.a  = \add_32ns_32ns_32_2_1_U13.din0 ;
assign \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.b  = \add_32ns_32ns_32_2_1_U13.din1 ;
assign \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  = \add_32ns_32ns_32_2_1_U13.ce ;
assign \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.clk  = \add_32ns_32ns_32_2_1_U13.clk ;
assign \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.reset  = \add_32ns_32ns_32_2_1_U13.reset ;
assign \add_32ns_32ns_32_2_1_U13.dout  = \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.s ;
assign \add_32ns_32ns_32_2_1_U13.ce  = 1'h1;
assign \add_32ns_32ns_32_2_1_U13.clk  = ap_clk;
assign \add_32ns_32ns_32_2_1_U13.din0  = ret_V_18_reg_992;
assign \add_32ns_32ns_32_2_1_U13.din1  = select_ln69_1_reg_997;
assign grp_fu_663_p2 = \add_32ns_32ns_32_2_1_U13.dout ;
assign \add_32ns_32ns_32_2_1_U13.reset  = ap_rst;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s0  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.a ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s0  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.b ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.s  = { \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s2 , \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.sum_s1  };
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.a  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s1 ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.b  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s1 ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cin  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.carry_s1 ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s2  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cout ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s2  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.s ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.a  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.a [15:0];
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.b  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.b [15:0];
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cin  = 1'h0;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s1  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cout ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s1  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.s ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.a  = \add_32ns_32ns_32_2_1_U12.din0 ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.b  = \add_32ns_32ns_32_2_1_U12.din1 ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  = \add_32ns_32ns_32_2_1_U12.ce ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.clk  = \add_32ns_32ns_32_2_1_U12.clk ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.reset  = \add_32ns_32ns_32_2_1_U12.reset ;
assign \add_32ns_32ns_32_2_1_U12.dout  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.s ;
assign \add_32ns_32ns_32_2_1_U12.ce  = 1'h1;
assign \add_32ns_32ns_32_2_1_U12.clk  = ap_clk;
assign \add_32ns_32ns_32_2_1_U12.din0  = ret_V_20_cast_reg_980;
assign \add_32ns_32ns_32_2_1_U12.din1  = 32'd1;
assign grp_fu_618_p2 = \add_32ns_32ns_32_2_1_U12.dout ;
assign \add_32ns_32ns_32_2_1_U12.reset  = ap_rst;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s0  = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.a ;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s0  = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.b ;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.s  = { \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s2 , \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.sum_s1  };
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.a  = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s1 ;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.b  = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s1 ;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cin  = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.carry_s1 ;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s2  = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cout ;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s2  = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.s ;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.a  = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.a [15:0];
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.b  = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.b [15:0];
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cin  = 1'h0;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s1  = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cout ;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s1  = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.s ;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.a  = \add_32ns_32ns_32_2_1_U10.din0 ;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.b  = \add_32ns_32ns_32_2_1_U10.din1 ;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  = \add_32ns_32ns_32_2_1_U10.ce ;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.clk  = \add_32ns_32ns_32_2_1_U10.clk ;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.reset  = \add_32ns_32ns_32_2_1_U10.reset ;
assign \add_32ns_32ns_32_2_1_U10.dout  = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.s ;
assign \add_32ns_32ns_32_2_1_U10.ce  = 1'h1;
assign \add_32ns_32ns_32_2_1_U10.clk  = ap_clk;
assign \add_32ns_32ns_32_2_1_U10.din0  = ret_V_18_cast_reg_943;
assign \add_32ns_32ns_32_2_1_U10.din1  = 32'd1;
assign grp_fu_563_p2 = \add_32ns_32ns_32_2_1_U10.dout ;
assign \add_32ns_32ns_32_2_1_U10.reset  = ap_rst;
assign \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_0_U.ain_s0  = \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_0_U.a ;
assign \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_0_U.bin_s0  = \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_0_U.b ;
assign \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_0_U.s  = { \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_0_U.fas_s2 , \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_0_U.sum_s1  };
assign \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_0_U.u2.a  = \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_0_U.ain_s1 ;
assign \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_0_U.u2.b  = \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_0_U.bin_s1 ;
assign \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_0_U.u2.cin  = \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_0_U.carry_s1 ;
assign \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_0_U.facout_s2  = \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_0_U.u2.cout ;
assign \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_0_U.fas_s2  = \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_0_U.u2.s ;
assign \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_0_U.u1.a  = \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_0_U.a [0];
assign \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_0_U.u1.b  = \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_0_U.b [0];
assign \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_0_U.u1.cin  = 1'h0;
assign \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_0_U.facout_s1  = \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_0_U.u1.cout ;
assign \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_0_U.fas_s1  = \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_0_U.u1.s ;
assign \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_0_U.a  = \add_2ns_2ns_2_2_1_U3.din0 ;
assign \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_0_U.b  = \add_2ns_2ns_2_2_1_U3.din1 ;
assign \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_0_U.ce  = \add_2ns_2ns_2_2_1_U3.ce ;
assign \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_0_U.clk  = \add_2ns_2ns_2_2_1_U3.clk ;
assign \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_0_U.reset  = \add_2ns_2ns_2_2_1_U3.reset ;
assign \add_2ns_2ns_2_2_1_U3.dout  = \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_0_U.s ;
assign \add_2ns_2ns_2_2_1_U3.ce  = 1'h1;
assign \add_2ns_2ns_2_2_1_U3.clk  = ap_clk;
assign \add_2ns_2ns_2_2_1_U3.din0  = { 1'h0, icmp_ln1494_reg_779 };
assign \add_2ns_2ns_2_2_1_U3.din1  = select_ln69_reg_804;
assign grp_fu_375_p2 = \add_2ns_2ns_2_2_1_U3.dout ;
assign \add_2ns_2ns_2_2_1_U3.reset  = ap_rst;
assign \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.ain_s0  = \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.a ;
assign \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.bin_s0  = \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.b ;
assign \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.s  = { \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.fas_s2 , \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.sum_s1  };
assign \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.u2.a  = \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.ain_s1 ;
assign \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.u2.b  = \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.bin_s1 ;
assign \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.u2.cin  = \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.carry_s1 ;
assign \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.facout_s2  = \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.u2.cout ;
assign \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.fas_s2  = \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.u2.s ;
assign \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.u1.a  = \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.a [0];
assign \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.u1.b  = \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.b [0];
assign \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.u1.cin  = 1'h0;
assign \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.facout_s1  = \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.u1.cout ;
assign \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.fas_s1  = \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.u1.s ;
assign \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.a  = \add_2ns_2ns_2_2_1_U1.din0 ;
assign \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.b  = \add_2ns_2ns_2_2_1_U1.din1 ;
assign \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.ce  = \add_2ns_2ns_2_2_1_U1.ce ;
assign \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.clk  = \add_2ns_2ns_2_2_1_U1.clk ;
assign \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.reset  = \add_2ns_2ns_2_2_1_U1.reset ;
assign \add_2ns_2ns_2_2_1_U1.dout  = \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.s ;
assign \add_2ns_2ns_2_2_1_U1.ce  = 1'h1;
assign \add_2ns_2ns_2_2_1_U1.clk  = ap_clk;
assign \add_2ns_2ns_2_2_1_U1.din0  = ret_V_cast_reg_767;
assign \add_2ns_2ns_2_2_1_U1.din1  = 2'h1;
assign grp_fu_320_p2 = \add_2ns_2ns_2_2_1_U1.dout ;
assign \add_2ns_2ns_2_2_1_U1.reset  = ap_rst;
assign \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.ain_s0  = \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.a ;
assign \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.bin_s0  = \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.b ;
assign \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.s  = { \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.fas_s2 , \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.sum_s1  };
assign \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.u2.a  = \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.ain_s1 ;
assign \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.u2.b  = \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.bin_s1 ;
assign \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.u2.cin  = \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.carry_s1 ;
assign \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.facout_s2  = \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.u2.cout ;
assign \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.fas_s2  = \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.u2.s ;
assign \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.u1.a  = \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.a [11:0];
assign \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.u1.b  = \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.b [11:0];
assign \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.u1.cin  = 1'h0;
assign \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.facout_s1  = \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.u1.cout ;
assign \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.fas_s1  = \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.u1.s ;
assign \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.a  = \add_24s_24ns_24_2_1_U6.din0 ;
assign \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.b  = \add_24s_24ns_24_2_1_U6.din1 ;
assign \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.ce  = \add_24s_24ns_24_2_1_U6.ce ;
assign \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.clk  = \add_24s_24ns_24_2_1_U6.clk ;
assign \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.reset  = \add_24s_24ns_24_2_1_U6.reset ;
assign \add_24s_24ns_24_2_1_U6.dout  = \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.s ;
assign \add_24s_24ns_24_2_1_U6.ce  = 1'h1;
assign \add_24s_24ns_24_2_1_U6.clk  = ap_clk;
assign \add_24s_24ns_24_2_1_U6.din0  = { tmp_reg_864[22], tmp_reg_864 };
assign \add_24s_24ns_24_2_1_U6.din1  = 24'h000001;
assign grp_fu_432_p2 = \add_24s_24ns_24_2_1_U6.dout ;
assign \add_24s_24ns_24_2_1_U6.reset  = ap_rst;
endmodule


// Machine B:
// Processed by function `add_clk_enable_signal` in `verilog_tricks.py`.
// Processed by function `remove_reset_signal` in `verilog_tricks.py`.
module top_B (
  ap_clk,
  ap_start,
  ap_done,
  ap_idle,
  ap_ready,
  op_0,
  op_2,
  op_3,
  op_5,
  op_10,
  op_11,
  op_12,
  op_13,
  op_14,
  op_15,
  op_17,
  op_18,
  op_19,
  op_31,
  op_31_ap_vld,
clk_enable
);
input clk_enable;


input ap_clk;
wire ap_rst;
assign ap_rst = op_31_ap_vld;
input ap_start;
input [3:0] op_0;
input [1:0] op_10;
input op_11;
input [31:0] op_12;
input [31:0] op_13;
input [7:0] op_14;
input [3:0] op_15;
input [31:0] op_17;
input op_18;
input op_19;
input [1:0] op_2;
input [3:0] op_3;
input [3:0] op_5;
output ap_done;
output ap_idle;
output ap_ready;
output [31:0] op_31;
output op_31_ap_vld;


reg [11:0] \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.ain_s1 ;
reg [11:0] \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.bin_s1 ;
reg \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.carry_s1 ;
reg [11:0] \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.sum_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s1 ;
reg \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.carry_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.sum_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s1 ;
reg \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.carry_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.sum_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s1 ;
reg \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.carry_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.sum_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s1 ;
reg \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.carry_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.sum_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s1 ;
reg \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.carry_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.sum_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s1 ;
reg \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.carry_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.sum_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s1 ;
reg \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.carry_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.sum_s1 ;
reg [16:0] \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.ain_s1 ;
reg [16:0] \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.bin_s1 ;
reg \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.carry_s1 ;
reg [15:0] \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.sum_s1 ;
reg [16:0] \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.ain_s1 ;
reg [16:0] \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.bin_s1 ;
reg \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.carry_s1 ;
reg [16:0] \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.sum_s1 ;
reg [17:0] \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.ain_s1 ;
reg [17:0] \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.bin_s1 ;
reg \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.carry_s1 ;
reg [16:0] \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.sum_s1 ;
reg [19:0] \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.ain_s1 ;
reg [19:0] \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.bin_s1 ;
reg \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.carry_s1 ;
reg [19:0] \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.sum_s1 ;
reg [26:0] \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.ain_s1 ;
reg [26:0] \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.bin_s1 ;
reg \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.carry_s1 ;
reg [26:0] \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.sum_s1 ;
reg [31:0] add_ln691_1_reg_881;
reg [31:0] add_ln691_2_reg_918;
reg [31:0] add_ln691_3_reg_955;
reg [31:0] add_ln691_4_reg_1002;
reg [23:0] add_ln691_reg_844;
reg [1:0] add_ln69_1_reg_802;
reg [5:0] add_ln69_reg_797;
reg [34:0] ap_CS_fsm = 35'h000000001;
reg icmp_ln1494_reg_782;
reg icmp_ln1499_reg_760;
reg icmp_ln851_1_reg_822;
reg icmp_ln851_2_reg_864;
reg icmp_ln851_3_reg_901;
reg icmp_ln851_4_reg_985;
reg icmp_ln851_reg_777;
reg [5:0] op_23_V_reg_807;
reg [31:0] op_28_V_reg_970;
reg [32:0] ret_V_14_reg_827;
reg [34:0] ret_V_15_reg_869;
reg [39:0] ret_V_16_reg_906;
reg [33:0] ret_V_17_reg_943;
reg [31:0] ret_V_18_cast_reg_911;
reg [31:0] ret_V_18_reg_960;
reg [53:0] ret_V_19_reg_990;
reg [31:0] ret_V_20_cast_reg_948;
reg [31:0] ret_V_20_reg_1007;
reg [31:0] ret_V_21_reg_1017;
reg [31:0] ret_V_22_cast_reg_995;
reg [31:0] ret_V_7_cast_reg_874;
reg [1:0] ret_V_cast_reg_770;
reg [1:0] ret_V_reg_792;
reg [31:0] select_ln1192_1_reg_1022;
reg [31:0] select_ln1192_reg_1012;
reg [31:0] select_ln353_1_reg_886;
reg [31:0] select_ln353_2_reg_923;
reg [23:0] select_ln353_reg_849;
reg [31:0] select_ln69_1_reg_965;
reg [23:0] sext_ln850_reg_837;
reg signbit_reg_787;
reg [22:0] tmp_reg_832;
reg [3:0] _379_;
wire [31:0] _000_;
wire [31:0] _001_;
wire [31:0] _002_;
wire [31:0] _003_;
wire [23:0] _004_;
wire [1:0] _005_;
wire [5:0] _006_;
wire [34:0] _007_;
wire _008_;
wire _009_;
wire _010_;
wire _011_;
wire _012_;
wire _013_;
wire _014_;
wire [5:0] _015_;
wire [31:0] _016_;
wire [3:0] _017_;
wire [32:0] _018_;
wire [34:0] _019_;
wire [39:0] _020_;
wire [33:0] _021_;
wire [31:0] _022_;
wire [31:0] _023_;
wire [53:0] _024_;
wire [31:0] _025_;
wire [31:0] _026_;
wire [31:0] _027_;
wire [31:0] _028_;
wire [31:0] _029_;
wire [1:0] _030_;
wire [1:0] _031_;
wire [31:0] _032_;
wire [31:0] _033_;
wire [31:0] _034_;
wire [31:0] _035_;
wire [23:0] _036_;
wire [31:0] _037_;
wire [23:0] _038_;
wire _039_;
wire [22:0] _040_;
wire [1:0] _041_;
wire _042_;
wire _043_;
wire _044_;
wire _045_;
wire _046_;
wire _047_;
wire _048_;
wire _049_;
wire _050_;
wire _051_;
wire _052_;
wire [11:0] _053_;
wire [11:0] _054_;
wire _055_;
wire [11:0] _056_;
wire [12:0] _057_;
wire [12:0] _058_;
wire [15:0] _059_;
wire [15:0] _060_;
wire _061_;
wire [15:0] _062_;
wire [16:0] _063_;
wire [16:0] _064_;
wire [15:0] _065_;
wire [15:0] _066_;
wire _067_;
wire [15:0] _068_;
wire [16:0] _069_;
wire [16:0] _070_;
wire [15:0] _071_;
wire [15:0] _072_;
wire _073_;
wire [15:0] _074_;
wire [16:0] _075_;
wire [16:0] _076_;
wire [15:0] _077_;
wire [15:0] _078_;
wire _079_;
wire [15:0] _080_;
wire [16:0] _081_;
wire [16:0] _082_;
wire [15:0] _083_;
wire [15:0] _084_;
wire _085_;
wire [15:0] _086_;
wire [16:0] _087_;
wire [16:0] _088_;
wire [15:0] _089_;
wire [15:0] _090_;
wire _091_;
wire [15:0] _092_;
wire [16:0] _093_;
wire [16:0] _094_;
wire [15:0] _095_;
wire [15:0] _096_;
wire _097_;
wire [15:0] _098_;
wire [16:0] _099_;
wire [16:0] _100_;
wire [16:0] _101_;
wire [16:0] _102_;
wire _103_;
wire [15:0] _104_;
wire [16:0] _105_;
wire [17:0] _106_;
wire [16:0] _107_;
wire [16:0] _108_;
wire _109_;
wire [16:0] _110_;
wire [17:0] _111_;
wire [17:0] _112_;
wire [17:0] _113_;
wire [17:0] _114_;
wire _115_;
wire [16:0] _116_;
wire [17:0] _117_;
wire [18:0] _118_;
wire [19:0] _119_;
wire [19:0] _120_;
wire _121_;
wire [19:0] _122_;
wire [20:0] _123_;
wire [20:0] _124_;
wire [26:0] _125_;
wire [26:0] _126_;
wire _127_;
wire [26:0] _128_;
wire [27:0] _129_;
wire [27:0] _130_;
wire _131_;
wire _132_;
wire _133_;
wire _134_;
wire _135_;
wire _136_;
wire _137_;
wire _138_;
wire _139_;
wire _140_;
wire _141_;
wire _142_;
wire _143_;
wire _144_;
wire _145_;
wire _146_;
wire _147_;
wire _148_;
wire _149_;
wire _150_;
wire _151_;
wire _152_;
wire _153_;
wire _154_;
wire _155_;
wire _156_;
wire _157_;
wire _158_;
wire _159_;
wire _160_;
wire _161_;
wire _162_;
wire _163_;
wire _164_;
wire _165_;
wire _166_;
wire _167_;
wire _168_;
wire _169_;
wire _170_;
wire _171_;
wire \add_24s_24ns_24_2_1_U6.ce ;
wire \add_24s_24ns_24_2_1_U6.clk ;
wire [23:0] \add_24s_24ns_24_2_1_U6.din0 ;
wire [23:0] \add_24s_24ns_24_2_1_U6.din1 ;
wire [23:0] \add_24s_24ns_24_2_1_U6.dout ;
wire \add_24s_24ns_24_2_1_U6.reset ;
wire [23:0] \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.a ;
wire [23:0] \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.ain_s0 ;
wire [23:0] \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.b ;
wire [23:0] \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.bin_s0 ;
wire \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.ce ;
wire \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.clk ;
wire \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.facout_s1 ;
wire \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.facout_s2 ;
wire [11:0] \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.fas_s1 ;
wire [11:0] \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.fas_s2 ;
wire \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.reset ;
wire [23:0] \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.s ;
wire [11:0] \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.u1.a ;
wire [11:0] \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.u1.b ;
wire \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.u1.cin ;
wire \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.u1.cout ;
wire [11:0] \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.u1.s ;
wire [11:0] \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.u2.a ;
wire [11:0] \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.u2.b ;
wire \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.u2.cin ;
wire \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.u2.cout ;
wire [11:0] \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.u2.s ;
wire [1:0] \add_2ns_2ns_2_1_1_U1.din0 ;
wire [1:0] \add_2ns_2ns_2_1_1_U1.din1 ;
wire [1:0] \add_2ns_2ns_2_1_1_U1.dout ;
wire [1:0] \add_2ns_2ns_2_1_1_U1.top_add_2ns_2ns_2_1_1_Adder_0_U.a ;
wire [1:0] \add_2ns_2ns_2_1_1_U1.top_add_2ns_2ns_2_1_1_Adder_0_U.b ;
wire [1:0] \add_2ns_2ns_2_1_1_U1.top_add_2ns_2ns_2_1_1_Adder_0_U.s ;
wire [1:0] \add_2ns_2ns_2_1_1_U3.din0 ;
wire [1:0] \add_2ns_2ns_2_1_1_U3.din1 ;
wire [1:0] \add_2ns_2ns_2_1_1_U3.dout ;
wire [1:0] \add_2ns_2ns_2_1_1_U3.top_add_2ns_2ns_2_1_1_Adder_0_U.a ;
wire [1:0] \add_2ns_2ns_2_1_1_U3.top_add_2ns_2ns_2_1_1_Adder_0_U.b ;
wire [1:0] \add_2ns_2ns_2_1_1_U3.top_add_2ns_2ns_2_1_1_Adder_0_U.s ;
wire \add_32ns_32ns_32_2_1_U10.ce ;
wire \add_32ns_32ns_32_2_1_U10.clk ;
wire [31:0] \add_32ns_32ns_32_2_1_U10.din0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U10.din1 ;
wire [31:0] \add_32ns_32ns_32_2_1_U10.dout ;
wire \add_32ns_32ns_32_2_1_U10.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.a ;
wire [31:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.b ;
wire [31:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s0 ;
wire \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.ce ;
wire \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.clk ;
wire \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s1 ;
wire \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s2 ;
wire [15:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s1 ;
wire [15:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s2 ;
wire \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.b ;
wire \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cin ;
wire \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.b ;
wire \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cin ;
wire \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.s ;
wire \add_32ns_32ns_32_2_1_U12.ce ;
wire \add_32ns_32ns_32_2_1_U12.clk ;
wire [31:0] \add_32ns_32ns_32_2_1_U12.din0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U12.din1 ;
wire [31:0] \add_32ns_32ns_32_2_1_U12.dout ;
wire \add_32ns_32ns_32_2_1_U12.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.a ;
wire [31:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.b ;
wire [31:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s0 ;
wire \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.ce ;
wire \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.clk ;
wire \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s1 ;
wire \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s2 ;
wire [15:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s1 ;
wire [15:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s2 ;
wire \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.b ;
wire \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cin ;
wire \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.b ;
wire \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cin ;
wire \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.s ;
wire \add_32ns_32ns_32_2_1_U13.ce ;
wire \add_32ns_32ns_32_2_1_U13.clk ;
wire [31:0] \add_32ns_32ns_32_2_1_U13.din0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U13.din1 ;
wire [31:0] \add_32ns_32ns_32_2_1_U13.dout ;
wire \add_32ns_32ns_32_2_1_U13.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.a ;
wire [31:0] \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.b ;
wire [31:0] \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s0 ;
wire \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.ce ;
wire \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.clk ;
wire \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s1 ;
wire \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s2 ;
wire [15:0] \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s1 ;
wire [15:0] \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s2 ;
wire \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.b ;
wire \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cin ;
wire \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.b ;
wire \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cin ;
wire \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.s ;
wire \add_32ns_32ns_32_2_1_U15.ce ;
wire \add_32ns_32ns_32_2_1_U15.clk ;
wire [31:0] \add_32ns_32ns_32_2_1_U15.din0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U15.din1 ;
wire [31:0] \add_32ns_32ns_32_2_1_U15.dout ;
wire \add_32ns_32ns_32_2_1_U15.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.a ;
wire [31:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.b ;
wire [31:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s0 ;
wire \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.ce ;
wire \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.clk ;
wire \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s1 ;
wire \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s2 ;
wire [15:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s1 ;
wire [15:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s2 ;
wire \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.b ;
wire \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cin ;
wire \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.b ;
wire \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cin ;
wire \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.s ;
wire \add_32ns_32ns_32_2_1_U16.ce ;
wire \add_32ns_32ns_32_2_1_U16.clk ;
wire [31:0] \add_32ns_32ns_32_2_1_U16.din0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U16.din1 ;
wire [31:0] \add_32ns_32ns_32_2_1_U16.dout ;
wire \add_32ns_32ns_32_2_1_U16.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.a ;
wire [31:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.b ;
wire [31:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s0 ;
wire \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.ce ;
wire \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.clk ;
wire \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s1 ;
wire \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s2 ;
wire [15:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s1 ;
wire [15:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s2 ;
wire \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.b ;
wire \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cin ;
wire \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.b ;
wire \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cin ;
wire \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.s ;
wire \add_32ns_32ns_32_2_1_U17.ce ;
wire \add_32ns_32ns_32_2_1_U17.clk ;
wire [31:0] \add_32ns_32ns_32_2_1_U17.din0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U17.din1 ;
wire [31:0] \add_32ns_32ns_32_2_1_U17.dout ;
wire \add_32ns_32ns_32_2_1_U17.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.a ;
wire [31:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.b ;
wire [31:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s0 ;
wire \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.ce ;
wire \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.clk ;
wire \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s1 ;
wire \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s2 ;
wire [15:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s1 ;
wire [15:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s2 ;
wire \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.b ;
wire \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cin ;
wire \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.b ;
wire \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cin ;
wire \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.s ;
wire \add_32ns_32ns_32_2_1_U8.ce ;
wire \add_32ns_32ns_32_2_1_U8.clk ;
wire [31:0] \add_32ns_32ns_32_2_1_U8.din0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U8.din1 ;
wire [31:0] \add_32ns_32ns_32_2_1_U8.dout ;
wire \add_32ns_32ns_32_2_1_U8.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.a ;
wire [31:0] \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.b ;
wire [31:0] \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s0 ;
wire \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.ce ;
wire \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.clk ;
wire \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s1 ;
wire \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s2 ;
wire [15:0] \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s1 ;
wire [15:0] \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s2 ;
wire \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.b ;
wire \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cin ;
wire \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.b ;
wire \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cin ;
wire \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.s ;
wire \add_33s_33s_33_2_1_U5.ce ;
wire \add_33s_33s_33_2_1_U5.clk ;
wire [32:0] \add_33s_33s_33_2_1_U5.din0 ;
wire [32:0] \add_33s_33s_33_2_1_U5.din1 ;
wire [32:0] \add_33s_33s_33_2_1_U5.dout ;
wire \add_33s_33s_33_2_1_U5.reset ;
wire [32:0] \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.a ;
wire [32:0] \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.ain_s0 ;
wire [32:0] \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.b ;
wire [32:0] \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.bin_s0 ;
wire \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.ce ;
wire \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.clk ;
wire \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.facout_s1 ;
wire \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.facout_s2 ;
wire [15:0] \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.fas_s1 ;
wire [16:0] \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.fas_s2 ;
wire \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.reset ;
wire [32:0] \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.s ;
wire [15:0] \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.u1.a ;
wire [15:0] \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.u1.b ;
wire \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.u1.cin ;
wire \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.u1.cout ;
wire [15:0] \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.u1.s ;
wire [16:0] \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.u2.a ;
wire [16:0] \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.u2.b ;
wire \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.u2.cin ;
wire \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.u2.cout ;
wire [16:0] \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.u2.s ;
wire \add_34s_34s_34_2_1_U11.ce ;
wire \add_34s_34s_34_2_1_U11.clk ;
wire [33:0] \add_34s_34s_34_2_1_U11.din0 ;
wire [33:0] \add_34s_34s_34_2_1_U11.din1 ;
wire [33:0] \add_34s_34s_34_2_1_U11.dout ;
wire \add_34s_34s_34_2_1_U11.reset ;
wire [33:0] \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.a ;
wire [33:0] \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.ain_s0 ;
wire [33:0] \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.b ;
wire [33:0] \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.bin_s0 ;
wire \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.ce ;
wire \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.clk ;
wire \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.facout_s1 ;
wire \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.facout_s2 ;
wire [16:0] \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.fas_s1 ;
wire [16:0] \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.fas_s2 ;
wire \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.reset ;
wire [33:0] \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.s ;
wire [16:0] \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.u1.a ;
wire [16:0] \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.u1.b ;
wire \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.u1.cin ;
wire \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.u1.cout ;
wire [16:0] \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.u1.s ;
wire [16:0] \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.u2.a ;
wire [16:0] \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.u2.b ;
wire \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.u2.cin ;
wire \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.u2.cout ;
wire [16:0] \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.u2.s ;
wire \add_35s_35s_35_2_1_U7.ce ;
wire \add_35s_35s_35_2_1_U7.clk ;
wire [34:0] \add_35s_35s_35_2_1_U7.din0 ;
wire [34:0] \add_35s_35s_35_2_1_U7.din1 ;
wire [34:0] \add_35s_35s_35_2_1_U7.dout ;
wire \add_35s_35s_35_2_1_U7.reset ;
wire [34:0] \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.a ;
wire [34:0] \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.ain_s0 ;
wire [34:0] \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.b ;
wire [34:0] \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.bin_s0 ;
wire \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.ce ;
wire \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.clk ;
wire \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.facout_s1 ;
wire \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.facout_s2 ;
wire [16:0] \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.fas_s1 ;
wire [17:0] \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.fas_s2 ;
wire \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.reset ;
wire [34:0] \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.s ;
wire [16:0] \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.u1.a ;
wire [16:0] \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.u1.b ;
wire \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.u1.cin ;
wire \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.u1.cout ;
wire [16:0] \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.u1.s ;
wire [17:0] \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.u2.a ;
wire [17:0] \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.u2.b ;
wire \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.u2.cin ;
wire \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.u2.cout ;
wire [17:0] \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.u2.s ;
wire \add_40s_40s_40_2_1_U9.ce ;
wire \add_40s_40s_40_2_1_U9.clk ;
wire [39:0] \add_40s_40s_40_2_1_U9.din0 ;
wire [39:0] \add_40s_40s_40_2_1_U9.din1 ;
wire [39:0] \add_40s_40s_40_2_1_U9.dout ;
wire \add_40s_40s_40_2_1_U9.reset ;
wire [39:0] \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.a ;
wire [39:0] \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.ain_s0 ;
wire [39:0] \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.b ;
wire [39:0] \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.bin_s0 ;
wire \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.ce ;
wire \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.clk ;
wire \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.facout_s1 ;
wire \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.facout_s2 ;
wire [19:0] \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.fas_s1 ;
wire [19:0] \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.fas_s2 ;
wire \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.reset ;
wire [39:0] \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.s ;
wire [19:0] \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.u1.a ;
wire [19:0] \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.u1.b ;
wire \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.u1.cin ;
wire \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.u1.cout ;
wire [19:0] \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.u1.s ;
wire [19:0] \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.u2.a ;
wire [19:0] \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.u2.b ;
wire \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.u2.cin ;
wire \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.u2.cout ;
wire [19:0] \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.u2.s ;
wire \add_54s_54s_54_2_1_U14.ce ;
wire \add_54s_54s_54_2_1_U14.clk ;
wire [53:0] \add_54s_54s_54_2_1_U14.din0 ;
wire [53:0] \add_54s_54s_54_2_1_U14.din1 ;
wire [53:0] \add_54s_54s_54_2_1_U14.dout ;
wire \add_54s_54s_54_2_1_U14.reset ;
wire [53:0] \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.a ;
wire [53:0] \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.ain_s0 ;
wire [53:0] \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.b ;
wire [53:0] \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.bin_s0 ;
wire \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.ce ;
wire \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.clk ;
wire \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.facout_s1 ;
wire \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.facout_s2 ;
wire [26:0] \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.fas_s1 ;
wire [26:0] \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.fas_s2 ;
wire \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.reset ;
wire [53:0] \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.s ;
wire [26:0] \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.u1.a ;
wire [26:0] \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.u1.b ;
wire \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.u1.cin ;
wire \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.u1.cout ;
wire [26:0] \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.u1.s ;
wire [26:0] \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.u2.a ;
wire [26:0] \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.u2.b ;
wire \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.u2.cin ;
wire \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.u2.cout ;
wire [26:0] \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.u2.s ;
wire [5:0] \add_6s_6ns_6_1_1_U4.din0 ;
wire [5:0] \add_6s_6ns_6_1_1_U4.din1 ;
wire [5:0] \add_6s_6ns_6_1_1_U4.dout ;
wire [5:0] \add_6s_6ns_6_1_1_U4.top_add_6s_6ns_6_1_1_Adder_2_U.a ;
wire [5:0] \add_6s_6ns_6_1_1_U4.top_add_6s_6ns_6_1_1_Adder_2_U.b ;
wire [5:0] \add_6s_6ns_6_1_1_U4.top_add_6s_6ns_6_1_1_Adder_2_U.s ;
wire [5:0] \add_6s_6s_6_1_1_U2.din0 ;
wire [5:0] \add_6s_6s_6_1_1_U2.din1 ;
wire [5:0] \add_6s_6s_6_1_1_U2.dout ;
wire [5:0] \add_6s_6s_6_1_1_U2.top_add_6s_6s_6_1_1_Adder_1_U.a ;
wire [5:0] \add_6s_6s_6_1_1_U2.top_add_6s_6s_6_1_1_Adder_1_U.b ;
wire [5:0] \add_6s_6s_6_1_1_U2.top_add_6s_6s_6_1_1_Adder_1_U.s ;
wire [1:0] add_ln69_1_fu_377_p0;
wire [1:0] add_ln69_1_fu_377_p1;
wire [1:0] add_ln69_1_fu_377_p2;
wire [5:0] add_ln69_fu_371_p0;
wire [5:0] add_ln69_fu_371_p1;
wire [5:0] add_ln69_fu_371_p2;
wire ap_CS_fsm_state1;
wire ap_CS_fsm_state10;
wire ap_CS_fsm_state11;
wire ap_CS_fsm_state12;
wire ap_CS_fsm_state13;
wire ap_CS_fsm_state14;
wire ap_CS_fsm_state15;
wire ap_CS_fsm_state16;
wire ap_CS_fsm_state17;
wire ap_CS_fsm_state18;
wire ap_CS_fsm_state19;
wire ap_CS_fsm_state2;
wire ap_CS_fsm_state20;
wire ap_CS_fsm_state21;
wire ap_CS_fsm_state22;
wire ap_CS_fsm_state23;
wire ap_CS_fsm_state24;
wire ap_CS_fsm_state25;
wire ap_CS_fsm_state26;
wire ap_CS_fsm_state27;
wire ap_CS_fsm_state28;
wire ap_CS_fsm_state29;
wire ap_CS_fsm_state3;
wire ap_CS_fsm_state30;
wire ap_CS_fsm_state31;
wire ap_CS_fsm_state32;
wire ap_CS_fsm_state33;
wire ap_CS_fsm_state34;
wire ap_CS_fsm_state35;
wire ap_CS_fsm_state4;
wire ap_CS_fsm_state5;
wire ap_CS_fsm_state6;
wire ap_CS_fsm_state7;
wire ap_CS_fsm_state8;
wire ap_CS_fsm_state9;
wire [34:0] ap_NS_fsm;
wire ap_clk;
wire ap_done;
wire ap_idle;
wire ap_ready;
wire ap_rst;
wire ap_start;
wire [32:0] grp_fu_406_p0;
wire [32:0] grp_fu_406_p1;
wire [32:0] grp_fu_406_p2;
wire [23:0] grp_fu_435_p0;
wire [23:0] grp_fu_435_p2;
wire [34:0] grp_fu_475_p0;
wire [34:0] grp_fu_475_p1;
wire [34:0] grp_fu_475_p2;
wire [31:0] grp_fu_501_p2;
wire [39:0] grp_fu_540_p0;
wire [39:0] grp_fu_540_p1;
wire [39:0] grp_fu_540_p2;
wire [31:0] grp_fu_566_p2;
wire [33:0] grp_fu_605_p0;
wire [33:0] grp_fu_605_p1;
wire [33:0] grp_fu_605_p2;
wire [31:0] grp_fu_621_p2;
wire [31:0] grp_fu_666_p2;
wire [53:0] grp_fu_685_p0;
wire [53:0] grp_fu_685_p1;
wire [53:0] grp_fu_685_p2;
wire [31:0] grp_fu_711_p2;
wire [31:0] grp_fu_743_p2;
wire [31:0] grp_fu_755_p2;
wire icmp_ln1494_fu_309_p2;
wire icmp_ln1499_fu_253_p2;
wire icmp_ln851_1_fu_416_p2;
wire icmp_ln851_2_fu_485_p2;
wire icmp_ln851_3_fu_550_p2;
wire icmp_ln851_4_fu_695_p2;
wire icmp_ln851_fu_291_p2;
wire [3:0] op_0;
wire [1:0] op_10;
wire op_11;
wire [31:0] op_12;
wire [31:0] op_13;
wire [7:0] op_14;
wire [3:0] op_15;
wire op_16_V_fu_630_p2;
wire [31:0] op_17;
wire op_18;
wire op_19;
wire [1:0] op_2;
wire [4:0] op_20_V_fu_345_p3;
wire [5:0] op_23_V_fu_386_p0;
wire [5:0] op_23_V_fu_386_p2;
wire [3:0] op_3;
wire [31:0] op_31;
wire op_31_ap_vld;
wire [7:0] op_4_V_fu_233_p3;
wire [3:0] op_5;
wire p_Result_1_fu_441_p3;
wire p_Result_2_fu_506_p3;
wire p_Result_3_fu_571_p3;
wire p_Result_4_fu_635_p3;
wire p_Result_5_fu_716_p3;
wire p_Result_s_fu_326_p3;
wire [6:0] ret_V_12_fu_271_p2;
wire [6:0] ret_V_12_reg_765;
wire [1:0] ret_V_13_fu_338_p3;
wire [31:0] ret_V_18_fu_651_p3;
wire [31:0] ret_V_20_fu_728_p3;
wire [1:0] ret_V_fu_321_p2;
wire [15:0] rhs_2_fu_395_p3;
wire [38:0] rhs_3_fu_529_p3;
wire [32:0] rhs_4_fu_594_p3;
wire [52:0] rhs_6_fu_674_p3;
wire [6:0] rhs_fu_263_p3;
wire [31:0] select_ln1192_1_fu_747_p3;
wire [31:0] select_ln1192_fu_735_p3;
wire [31:0] select_ln353_1_fu_518_p3;
wire [31:0] select_ln353_2_fu_583_p3;
wire [23:0] select_ln353_fu_453_p3;
wire [31:0] select_ln69_1_fu_658_p3;
wire [23:0] select_ln850_1_fu_448_p3;
wire [31:0] select_ln850_2_fu_513_p3;
wire [31:0] select_ln850_3_fu_578_p3;
wire [31:0] select_ln850_4_fu_645_p3;
wire [31:0] select_ln850_5_fu_723_p3;
wire [1:0] select_ln850_fu_333_p3;
wire [31:0] sext_ln1192_fu_391_p0;
wire [7:0] sext_ln1494_fu_305_p1;
wire [3:0] sext_ln1499_fu_249_p0;
wire [4:0] sext_ln1499_fu_249_p1;
wire [31:0] sext_ln703_1_fu_460_p0;
wire [7:0] sext_ln703_2_fu_525_p0;
wire [3:0] sext_ln703_3_fu_590_p0;
wire [31:0] sext_ln703_4_fu_670_p0;
wire [3:0] sext_ln703_fu_259_p0;
wire [6:0] sext_ln703_fu_259_p1;
wire [23:0] sext_ln850_fu_432_p1;
wire [3:0] shl_ln728_2_fu_297_p1;
wire [6:0] shl_ln728_2_fu_297_p3;
wire [4:0] shl_ln_fu_241_p3;
wire signbit_fu_315_p2;
wire [25:0] tmp_3_fu_464_p3;
wire trunc_ln1195_fu_626_p1;
wire [31:0] trunc_ln851_1_fu_412_p0;
wire [9:0] trunc_ln851_1_fu_412_p1;
wire [31:0] trunc_ln851_2_fu_481_p0;
wire [1:0] trunc_ln851_2_fu_481_p1;
wire [7:0] trunc_ln851_3_fu_546_p0;
wire [6:0] trunc_ln851_3_fu_546_p1;
wire [3:0] trunc_ln851_4_fu_642_p0;
wire trunc_ln851_4_fu_642_p1;
wire [31:0] trunc_ln851_5_fu_691_p0;
wire [20:0] trunc_ln851_5_fu_691_p1;
wire [2:0] trunc_ln851_fu_287_p1;


assign _042_ = ap_CS_fsm[12] & icmp_ln851_2_reg_864;
assign _043_ = ap_CS_fsm[17] & icmp_ln851_3_reg_901;
assign _044_ = icmp_ln851_4_reg_985 & ap_CS_fsm[29];
assign _045_ = ap_CS_fsm[7] & icmp_ln851_1_reg_822;
assign _046_ = _049_ & ap_CS_fsm[1];
assign _047_ = _050_ & ap_CS_fsm[0];
assign _048_ = ap_start & ap_CS_fsm[0];
assign ret_V_12_fu_271_p2 = { op_3[3], op_3[3], op_3[3], op_3 } & { op_5, 3'h0 };
assign _049_ = ~ icmp_ln851_reg_777;
assign _050_ = ~ ap_start;
assign _051_ = ! ret_V_12_fu_271_p2[2:0];
assign _052_ = { op_3[3], op_3 } == { op_2, 3'h0 };
always @(posedge \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.clk )
\add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.bin_s1  <= _054_;
always @(posedge \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.clk )
\add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.ain_s1  <= _053_;
always @(posedge \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.clk )
\add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.sum_s1  <= _056_;
always @(posedge \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.clk )
\add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.carry_s1  <= _055_;
assign _054_ = \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.ce  ? \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.b [23:12] : \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.bin_s1 ;
assign _053_ = \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.ce  ? \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.a [23:12] : \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.ain_s1 ;
assign _055_ = \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.ce  ? \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.facout_s1  : \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.carry_s1 ;
assign _056_ = \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.ce  ? \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.fas_s1  : \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.sum_s1 ;
assign _057_ = \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.u1.a  + \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.u1.b ;
assign { \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.u1.cout , \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.u1.s  } = _057_ + \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.u1.cin ;
assign _058_ = \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.u2.a  + \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.u2.b ;
assign { \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.u2.cout , \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.u2.s  } = _058_ + \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.u2.cin ;
assign \add_2ns_2ns_2_1_1_U1.top_add_2ns_2ns_2_1_1_Adder_0_U.s  = \add_2ns_2ns_2_1_1_U1.top_add_2ns_2ns_2_1_1_Adder_0_U.a  + \add_2ns_2ns_2_1_1_U1.top_add_2ns_2ns_2_1_1_Adder_0_U.b ;
assign \add_2ns_2ns_2_1_1_U3.top_add_2ns_2ns_2_1_1_Adder_0_U.s  = \add_2ns_2ns_2_1_1_U3.top_add_2ns_2ns_2_1_1_Adder_0_U.a  + \add_2ns_2ns_2_1_1_U3.top_add_2ns_2ns_2_1_1_Adder_0_U.b ;
always @(posedge \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.clk )
\add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s1  <= _060_;
always @(posedge \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.clk )
\add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s1  <= _059_;
always @(posedge \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.clk )
\add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.sum_s1  <= _062_;
always @(posedge \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.clk )
\add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.carry_s1  <= _061_;
assign _060_ = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  ? \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.b [31:16] : \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s1 ;
assign _059_ = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  ? \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.a [31:16] : \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s1 ;
assign _061_ = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  ? \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s1  : \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.carry_s1 ;
assign _062_ = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  ? \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s1  : \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.sum_s1 ;
assign _063_ = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.a  + \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.b ;
assign { \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cout , \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.s  } = _063_ + \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cin ;
assign _064_ = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.a  + \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.b ;
assign { \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cout , \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.s  } = _064_ + \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cin ;
always @(posedge \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.clk )
\add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s1  <= _066_;
always @(posedge \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.clk )
\add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s1  <= _065_;
always @(posedge \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.clk )
\add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.sum_s1  <= _068_;
always @(posedge \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.clk )
\add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.carry_s1  <= _067_;
assign _066_ = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  ? \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.b [31:16] : \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s1 ;
assign _065_ = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  ? \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.a [31:16] : \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s1 ;
assign _067_ = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  ? \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s1  : \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.carry_s1 ;
assign _068_ = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  ? \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s1  : \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.sum_s1 ;
assign _069_ = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.a  + \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.b ;
assign { \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cout , \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.s  } = _069_ + \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cin ;
assign _070_ = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.a  + \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.b ;
assign { \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cout , \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.s  } = _070_ + \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cin ;
always @(posedge \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.clk )
\add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s1  <= _072_;
always @(posedge \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.clk )
\add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s1  <= _071_;
always @(posedge \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.clk )
\add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.sum_s1  <= _074_;
always @(posedge \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.clk )
\add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.carry_s1  <= _073_;
assign _072_ = \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  ? \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.b [31:16] : \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s1 ;
assign _071_ = \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  ? \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.a [31:16] : \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s1 ;
assign _073_ = \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  ? \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s1  : \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.carry_s1 ;
assign _074_ = \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  ? \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s1  : \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.sum_s1 ;
assign _075_ = \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.a  + \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.b ;
assign { \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cout , \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.s  } = _075_ + \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cin ;
assign _076_ = \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.a  + \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.b ;
assign { \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cout , \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.s  } = _076_ + \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cin ;
always @(posedge \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.clk )
\add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s1  <= _078_;
always @(posedge \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.clk )
\add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s1  <= _077_;
always @(posedge \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.clk )
\add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.sum_s1  <= _080_;
always @(posedge \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.clk )
\add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.carry_s1  <= _079_;
assign _078_ = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  ? \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.b [31:16] : \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s1 ;
assign _077_ = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  ? \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.a [31:16] : \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s1 ;
assign _079_ = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  ? \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s1  : \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.carry_s1 ;
assign _080_ = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  ? \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s1  : \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.sum_s1 ;
assign _081_ = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.a  + \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.b ;
assign { \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cout , \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.s  } = _081_ + \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cin ;
assign _082_ = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.a  + \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.b ;
assign { \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cout , \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.s  } = _082_ + \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cin ;
always @(posedge \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.clk )
\add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s1  <= _084_;
always @(posedge \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.clk )
\add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s1  <= _083_;
always @(posedge \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.clk )
\add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.sum_s1  <= _086_;
always @(posedge \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.clk )
\add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.carry_s1  <= _085_;
assign _084_ = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  ? \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.b [31:16] : \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s1 ;
assign _083_ = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  ? \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.a [31:16] : \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s1 ;
assign _085_ = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  ? \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s1  : \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.carry_s1 ;
assign _086_ = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  ? \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s1  : \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.sum_s1 ;
assign _087_ = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.a  + \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.b ;
assign { \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cout , \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.s  } = _087_ + \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cin ;
assign _088_ = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.a  + \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.b ;
assign { \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cout , \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.s  } = _088_ + \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cin ;
always @(posedge \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.clk )
\add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s1  <= _090_;
always @(posedge \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.clk )
\add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s1  <= _089_;
always @(posedge \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.clk )
\add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.sum_s1  <= _092_;
always @(posedge \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.clk )
\add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.carry_s1  <= _091_;
assign _090_ = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  ? \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.b [31:16] : \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s1 ;
assign _089_ = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  ? \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.a [31:16] : \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s1 ;
assign _091_ = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  ? \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s1  : \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.carry_s1 ;
assign _092_ = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  ? \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s1  : \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.sum_s1 ;
assign _093_ = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.a  + \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.b ;
assign { \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cout , \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.s  } = _093_ + \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cin ;
assign _094_ = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.a  + \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.b ;
assign { \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cout , \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.s  } = _094_ + \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cin ;
always @(posedge \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.clk )
\add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s1  <= _096_;
always @(posedge \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.clk )
\add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s1  <= _095_;
always @(posedge \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.clk )
\add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.sum_s1  <= _098_;
always @(posedge \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.clk )
\add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.carry_s1  <= _097_;
assign _096_ = \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  ? \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.b [31:16] : \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s1 ;
assign _095_ = \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  ? \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.a [31:16] : \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s1 ;
assign _097_ = \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  ? \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s1  : \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.carry_s1 ;
assign _098_ = \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  ? \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s1  : \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.sum_s1 ;
assign _099_ = \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.a  + \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.b ;
assign { \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cout , \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.s  } = _099_ + \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cin ;
assign _100_ = \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.a  + \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.b ;
assign { \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cout , \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.s  } = _100_ + \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cin ;
always @(posedge \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.clk )
\add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.bin_s1  <= _102_;
always @(posedge \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.clk )
\add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.ain_s1  <= _101_;
always @(posedge \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.clk )
\add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.sum_s1  <= _104_;
always @(posedge \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.clk )
\add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.carry_s1  <= _103_;
assign _102_ = \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.ce  ? \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.b [32:16] : \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.bin_s1 ;
assign _101_ = \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.ce  ? \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.a [32:16] : \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.ain_s1 ;
assign _103_ = \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.ce  ? \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.facout_s1  : \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.carry_s1 ;
assign _104_ = \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.ce  ? \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.fas_s1  : \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.sum_s1 ;
assign _105_ = \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.u1.a  + \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.u1.b ;
assign { \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.u1.cout , \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.u1.s  } = _105_ + \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.u1.cin ;
assign _106_ = \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.u2.a  + \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.u2.b ;
assign { \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.u2.cout , \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.u2.s  } = _106_ + \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.u2.cin ;
always @(posedge \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.clk )
\add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.bin_s1  <= _108_;
always @(posedge \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.clk )
\add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.ain_s1  <= _107_;
always @(posedge \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.clk )
\add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.sum_s1  <= _110_;
always @(posedge \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.clk )
\add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.carry_s1  <= _109_;
assign _108_ = \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.ce  ? \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.b [33:17] : \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.bin_s1 ;
assign _107_ = \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.ce  ? \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.a [33:17] : \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.ain_s1 ;
assign _109_ = \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.ce  ? \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.facout_s1  : \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.carry_s1 ;
assign _110_ = \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.ce  ? \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.fas_s1  : \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.sum_s1 ;
assign _111_ = \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.u1.a  + \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.u1.b ;
assign { \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.u1.cout , \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.u1.s  } = _111_ + \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.u1.cin ;
assign _112_ = \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.u2.a  + \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.u2.b ;
assign { \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.u2.cout , \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.u2.s  } = _112_ + \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.u2.cin ;
always @(posedge \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.clk )
\add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.bin_s1  <= _114_;
always @(posedge \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.clk )
\add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.ain_s1  <= _113_;
always @(posedge \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.clk )
\add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.sum_s1  <= _116_;
always @(posedge \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.clk )
\add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.carry_s1  <= _115_;
assign _114_ = \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.ce  ? \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.b [34:17] : \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.bin_s1 ;
assign _113_ = \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.ce  ? \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.a [34:17] : \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.ain_s1 ;
assign _115_ = \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.ce  ? \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.facout_s1  : \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.carry_s1 ;
assign _116_ = \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.ce  ? \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.fas_s1  : \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.sum_s1 ;
assign _117_ = \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.u1.a  + \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.u1.b ;
assign { \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.u1.cout , \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.u1.s  } = _117_ + \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.u1.cin ;
assign _118_ = \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.u2.a  + \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.u2.b ;
assign { \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.u2.cout , \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.u2.s  } = _118_ + \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.u2.cin ;
always @(posedge \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.clk )
\add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.bin_s1  <= _120_;
always @(posedge \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.clk )
\add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.ain_s1  <= _119_;
always @(posedge \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.clk )
\add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.sum_s1  <= _122_;
always @(posedge \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.clk )
\add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.carry_s1  <= _121_;
assign _120_ = \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.ce  ? \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.b [39:20] : \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.bin_s1 ;
assign _119_ = \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.ce  ? \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.a [39:20] : \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.ain_s1 ;
assign _121_ = \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.ce  ? \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.facout_s1  : \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.carry_s1 ;
assign _122_ = \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.ce  ? \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.fas_s1  : \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.sum_s1 ;
assign _123_ = \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.u1.a  + \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.u1.b ;
assign { \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.u1.cout , \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.u1.s  } = _123_ + \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.u1.cin ;
assign _124_ = \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.u2.a  + \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.u2.b ;
assign { \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.u2.cout , \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.u2.s  } = _124_ + \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.u2.cin ;
always @(posedge \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.clk )
\add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.bin_s1  <= _126_;
always @(posedge \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.clk )
\add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.ain_s1  <= _125_;
always @(posedge \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.clk )
\add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.sum_s1  <= _128_;
always @(posedge \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.clk )
\add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.carry_s1  <= _127_;
assign _126_ = \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.ce  ? \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.b [53:27] : \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.bin_s1 ;
assign _125_ = \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.ce  ? \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.a [53:27] : \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.ain_s1 ;
assign _127_ = \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.ce  ? \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.facout_s1  : \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.carry_s1 ;
assign _128_ = \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.ce  ? \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.fas_s1  : \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.sum_s1 ;
assign _129_ = \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.u1.a  + \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.u1.b ;
assign { \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.u1.cout , \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.u1.s  } = _129_ + \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.u1.cin ;
assign _130_ = \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.u2.a  + \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.u2.b ;
assign { \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.u2.cout , \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.u2.s  } = _130_ + \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.u2.cin ;
assign \add_6s_6ns_6_1_1_U4.top_add_6s_6ns_6_1_1_Adder_2_U.s  = \add_6s_6ns_6_1_1_U4.top_add_6s_6ns_6_1_1_Adder_2_U.a  + \add_6s_6ns_6_1_1_U4.top_add_6s_6ns_6_1_1_Adder_2_U.b ;
assign \add_6s_6s_6_1_1_U2.top_add_6s_6s_6_1_1_Adder_1_U.s  = \add_6s_6s_6_1_1_U2.top_add_6s_6s_6_1_1_Adder_1_U.a  + \add_6s_6s_6_1_1_U2.top_add_6s_6s_6_1_1_Adder_1_U.b ;
assign _131_ = $signed({ op_3, 3'h0 }) > $signed({ op_2, 6'h00 });
assign _132_ = { op_2, 3'h0 } != { op_3[3], op_3 };
assign _133_ = | op_12[9:0];
assign _134_ = | op_13[1:0];
assign _135_ = | op_14[6:0];
assign _136_ = | op_17[20:0];
assign op_16_V_fu_630_p2 = op_10[0] | signbit_reg_787;
always @(posedge ap_clk)
sext_ln850_reg_837 <= _038_;
always @(posedge ap_clk)
select_ln353_reg_849 <= _036_;
always @(posedge ap_clk)
select_ln353_2_reg_923 <= _035_;
always @(posedge ap_clk)
select_ln353_1_reg_886 <= _034_;
always @(posedge ap_clk)
ret_V_reg_792 <= _031_;
always @(posedge ap_clk)
ret_V_21_reg_1017 <= _027_;
always @(posedge ap_clk)
select_ln1192_1_reg_1022 <= _032_;
always @(posedge ap_clk)
ret_V_20_reg_1007 <= _026_;
always @(posedge ap_clk)
select_ln1192_reg_1012 <= _033_;
always @(posedge ap_clk)
ret_V_19_reg_990 <= _024_;
always @(posedge ap_clk)
ret_V_22_cast_reg_995 <= _028_;
always @(posedge ap_clk)
ret_V_18_reg_960 <= _023_;
always @(posedge ap_clk)
select_ln69_1_reg_965 <= _037_;
always @(posedge ap_clk)
ret_V_17_reg_943 <= _021_;
always @(posedge ap_clk)
ret_V_20_cast_reg_948 <= _025_;
always @(posedge ap_clk)
ret_V_16_reg_906 <= _020_;
always @(posedge ap_clk)
ret_V_18_cast_reg_911 <= _022_;
always @(posedge ap_clk)
ret_V_15_reg_869 <= _019_;
always @(posedge ap_clk)
ret_V_7_cast_reg_874 <= _029_;
always @(posedge ap_clk)
ret_V_14_reg_827 <= _018_;
always @(posedge ap_clk)
tmp_reg_832 <= _040_;
always @(posedge ap_clk)
op_28_V_reg_970 <= _016_;
always @(posedge ap_clk)
op_23_V_reg_807 <= _015_;
always @(posedge ap_clk)
icmp_ln851_4_reg_985 <= _013_;
always @(posedge ap_clk)
icmp_ln851_3_reg_901 <= _012_;
always @(posedge ap_clk)
icmp_ln851_2_reg_864 <= _011_;
always @(posedge ap_clk)
icmp_ln851_1_reg_822 <= _010_;
always @(posedge ap_clk)
icmp_ln1499_reg_760 <= _009_;
always @(posedge ap_clk)
_379_ <= _017_;
assign ret_V_12_reg_765[6:3] = _379_;
always @(posedge ap_clk)
ret_V_cast_reg_770 <= _030_;
always @(posedge ap_clk)
icmp_ln851_reg_777 <= _014_;
always @(posedge ap_clk)
icmp_ln1494_reg_782 <= _008_;
always @(posedge ap_clk)
signbit_reg_787 <= _039_;
always @(posedge ap_clk)
add_ln69_reg_797 <= _006_;
always @(posedge ap_clk)
add_ln69_1_reg_802 <= _005_;
always @(posedge ap_clk)
add_ln691_reg_844 <= _004_;
always @(posedge ap_clk)
add_ln691_4_reg_1002 <= _003_;
always @(posedge ap_clk)
add_ln691_3_reg_955 <= _002_;
always @(posedge ap_clk)
add_ln691_2_reg_918 <= _001_;
always @(posedge ap_clk)
add_ln691_1_reg_881 <= _000_;
always @(posedge ap_clk)
ap_CS_fsm <= _007_;
assign _041_ = _048_ ? 2'h2 : 2'h1;
assign _137_ = ap_CS_fsm == 1'h1;
function [34:0] _394_;
input [34:0] a;
input [1224:0] b;
input [34:0] s;
case (s)
35'b00000000000000000000000000000000001:
_394_ = b[34:0];
35'b00000000000000000000000000000000010:
_394_ = b[69:35];
35'b00000000000000000000000000000000100:
_394_ = b[104:70];
35'b00000000000000000000000000000001000:
_394_ = b[139:105];
35'b00000000000000000000000000000010000:
_394_ = b[174:140];
35'b00000000000000000000000000000100000:
_394_ = b[209:175];
35'b00000000000000000000000000001000000:
_394_ = b[244:210];
35'b00000000000000000000000000010000000:
_394_ = b[279:245];
35'b00000000000000000000000000100000000:
_394_ = b[314:280];
35'b00000000000000000000000001000000000:
_394_ = b[349:315];
35'b00000000000000000000000010000000000:
_394_ = b[384:350];
35'b00000000000000000000000100000000000:
_394_ = b[419:385];
35'b00000000000000000000001000000000000:
_394_ = b[454:420];
35'b00000000000000000000010000000000000:
_394_ = b[489:455];
35'b00000000000000000000100000000000000:
_394_ = b[524:490];
35'b00000000000000000001000000000000000:
_394_ = b[559:525];
35'b00000000000000000010000000000000000:
_394_ = b[594:560];
35'b00000000000000000100000000000000000:
_394_ = b[629:595];
35'b00000000000000001000000000000000000:
_394_ = b[664:630];
35'b00000000000000010000000000000000000:
_394_ = b[699:665];
35'b00000000000000100000000000000000000:
_394_ = b[734:700];
35'b00000000000001000000000000000000000:
_394_ = b[769:735];
35'b00000000000010000000000000000000000:
_394_ = b[804:770];
35'b00000000000100000000000000000000000:
_394_ = b[839:805];
35'b00000000001000000000000000000000000:
_394_ = b[874:840];
35'b00000000010000000000000000000000000:
_394_ = b[909:875];
35'b00000000100000000000000000000000000:
_394_ = b[944:910];
35'b00000001000000000000000000000000000:
_394_ = b[979:945];
35'b00000010000000000000000000000000000:
_394_ = b[1014:980];
35'b00000100000000000000000000000000000:
_394_ = b[1049:1015];
35'b00001000000000000000000000000000000:
_394_ = b[1084:1050];
35'b00010000000000000000000000000000000:
_394_ = b[1119:1085];
35'b00100000000000000000000000000000000:
_394_ = b[1154:1120];
35'b01000000000000000000000000000000000:
_394_ = b[1189:1155];
35'b10000000000000000000000000000000000:
_394_ = b[1224:1190];
35'b00000000000000000000000000000000000:
_394_ = a;
default:
_394_ = 35'bx;
endcase
endfunction
assign ap_NS_fsm = _394_(35'hxxxxxxxxx, { 33'h000000000, _041_, 1190'h0000000020000000080000000200000000800000002000000008000000020000000080000000200000000800000002000000008000000020000000080000000200000000800000002000000008000000020000000080000000200000000800000002000000008000000020000000080000000200000000800000002000000008000000020000000080000000200000000000000001 }, { _137_, _171_, _170_, _169_, _168_, _167_, _166_, _165_, _164_, _163_, _162_, _161_, _160_, _159_, _158_, _157_, _156_, _155_, _154_, _153_, _152_, _151_, _150_, _149_, _148_, _147_, _146_, _145_, _144_, _143_, _142_, _141_, _140_, _139_, _138_ });
assign _138_ = ap_CS_fsm == 35'h400000000;
assign _139_ = ap_CS_fsm == 34'h200000000;
assign _140_ = ap_CS_fsm == 33'h100000000;
assign _141_ = ap_CS_fsm == 32'd2147483648;
assign _142_ = ap_CS_fsm == 31'h40000000;
assign _143_ = ap_CS_fsm == 30'h20000000;
assign _144_ = ap_CS_fsm == 29'h10000000;
assign _145_ = ap_CS_fsm == 28'h8000000;
assign _146_ = ap_CS_fsm == 27'h4000000;
assign _147_ = ap_CS_fsm == 26'h2000000;
assign _148_ = ap_CS_fsm == 25'h1000000;
assign _149_ = ap_CS_fsm == 24'h800000;
assign _150_ = ap_CS_fsm == 23'h400000;
assign _151_ = ap_CS_fsm == 22'h200000;
assign _152_ = ap_CS_fsm == 21'h100000;
assign _153_ = ap_CS_fsm == 20'h80000;
assign _154_ = ap_CS_fsm == 19'h40000;
assign _155_ = ap_CS_fsm == 18'h20000;
assign _156_ = ap_CS_fsm == 17'h10000;
assign _157_ = ap_CS_fsm == 16'h8000;
assign _158_ = ap_CS_fsm == 15'h4000;
assign _159_ = ap_CS_fsm == 14'h2000;
assign _160_ = ap_CS_fsm == 13'h1000;
assign _161_ = ap_CS_fsm == 12'h800;
assign _162_ = ap_CS_fsm == 11'h400;
assign _163_ = ap_CS_fsm == 10'h200;
assign _164_ = ap_CS_fsm == 9'h100;
assign _165_ = ap_CS_fsm == 8'h80;
assign _166_ = ap_CS_fsm == 7'h40;
assign _167_ = ap_CS_fsm == 6'h20;
assign _168_ = ap_CS_fsm == 5'h10;
assign _169_ = ap_CS_fsm == 4'h8;
assign _170_ = ap_CS_fsm == 3'h4;
assign _171_ = ap_CS_fsm == 2'h2;
assign op_31_ap_vld = ap_CS_fsm[34] ? 1'h1 : 1'h0;
assign ap_idle = _047_ ? 1'h1 : 1'h0;
assign _038_ = ap_CS_fsm[6] ? { tmp_reg_832[22], tmp_reg_832 } : sext_ln850_reg_837;
assign _036_ = ap_CS_fsm[8] ? select_ln353_fu_453_p3 : select_ln353_reg_849;
assign _035_ = ap_CS_fsm[18] ? select_ln353_2_fu_583_p3 : select_ln353_2_reg_923;
assign _034_ = ap_CS_fsm[13] ? select_ln353_1_fu_518_p3 : select_ln353_1_reg_886;
assign _031_ = _046_ ? ret_V_fu_321_p2 : ret_V_reg_792;
assign _032_ = ap_CS_fsm[32] ? select_ln1192_1_fu_747_p3 : select_ln1192_1_reg_1022;
assign _027_ = ap_CS_fsm[32] ? grp_fu_743_p2 : ret_V_21_reg_1017;
assign _033_ = ap_CS_fsm[30] ? select_ln1192_fu_735_p3 : select_ln1192_reg_1012;
assign _026_ = ap_CS_fsm[30] ? ret_V_20_fu_728_p3 : ret_V_20_reg_1007;
assign _028_ = ap_CS_fsm[27] ? grp_fu_685_p2[52:21] : ret_V_22_cast_reg_995;
assign _024_ = ap_CS_fsm[27] ? grp_fu_685_p2 : ret_V_19_reg_990;
assign _037_ = ap_CS_fsm[23] ? select_ln69_1_fu_658_p3 : select_ln69_1_reg_965;
assign _023_ = ap_CS_fsm[23] ? ret_V_18_fu_651_p3 : ret_V_18_reg_960;
assign _025_ = ap_CS_fsm[20] ? grp_fu_605_p2[32:1] : ret_V_20_cast_reg_948;
assign _021_ = ap_CS_fsm[20] ? grp_fu_605_p2 : ret_V_17_reg_943;
assign _022_ = ap_CS_fsm[15] ? grp_fu_540_p2[38:7] : ret_V_18_cast_reg_911;
assign _020_ = ap_CS_fsm[15] ? grp_fu_540_p2 : ret_V_16_reg_906;
assign _029_ = ap_CS_fsm[10] ? grp_fu_475_p2[33:2] : ret_V_7_cast_reg_874;
assign _019_ = ap_CS_fsm[10] ? grp_fu_475_p2 : ret_V_15_reg_869;
assign _040_ = ap_CS_fsm[5] ? grp_fu_406_p2[32:10] : tmp_reg_832;
assign _018_ = ap_CS_fsm[5] ? grp_fu_406_p2 : ret_V_14_reg_827;
assign _016_ = ap_CS_fsm[25] ? grp_fu_666_p2 : op_28_V_reg_970;
assign _015_ = ap_CS_fsm[3] ? op_23_V_fu_386_p2 : op_23_V_reg_807;
assign _013_ = ap_CS_fsm[26] ? icmp_ln851_4_fu_695_p2 : icmp_ln851_4_reg_985;
assign _012_ = ap_CS_fsm[14] ? icmp_ln851_3_fu_550_p2 : icmp_ln851_3_reg_901;
assign _011_ = ap_CS_fsm[9] ? icmp_ln851_2_fu_485_p2 : icmp_ln851_2_reg_864;
assign _010_ = ap_CS_fsm[4] ? icmp_ln851_1_fu_416_p2 : icmp_ln851_1_reg_822;
assign _039_ = ap_CS_fsm[0] ? signbit_fu_315_p2 : signbit_reg_787;
assign _008_ = ap_CS_fsm[0] ? icmp_ln1494_fu_309_p2 : icmp_ln1494_reg_782;
assign _014_ = ap_CS_fsm[0] ? icmp_ln851_fu_291_p2 : icmp_ln851_reg_777;
assign _030_ = ap_CS_fsm[0] ? ret_V_12_fu_271_p2[4:3] : ret_V_cast_reg_770;
assign _017_ = ap_CS_fsm[0] ? ret_V_12_fu_271_p2[6:3] : ret_V_12_reg_765[6:3];
assign _009_ = ap_CS_fsm[0] ? icmp_ln1499_fu_253_p2 : icmp_ln1499_reg_760;
assign _005_ = ap_CS_fsm[2] ? add_ln69_1_fu_377_p2 : add_ln69_1_reg_802;
assign _006_ = ap_CS_fsm[2] ? add_ln69_fu_371_p2 : add_ln69_reg_797;
assign _004_ = _045_ ? grp_fu_435_p2 : add_ln691_reg_844;
assign _003_ = _044_ ? grp_fu_711_p2 : add_ln691_4_reg_1002;
assign _002_ = ap_CS_fsm[22] ? grp_fu_621_p2 : add_ln691_3_reg_955;
assign _001_ = _043_ ? grp_fu_566_p2 : add_ln691_2_reg_918;
assign _000_ = _042_ ? grp_fu_501_p2 : add_ln691_1_reg_881;
assign _007_ = ap_rst ? 35'h000000001 : ap_NS_fsm;
assign add_ln69_1_fu_377_p1 = op_11 ? 2'h3 : 2'h0;
assign icmp_ln1494_fu_309_p2 = _131_ ? 1'h1 : 1'h0;
assign icmp_ln1499_fu_253_p2 = _132_ ? 1'h1 : 1'h0;
assign icmp_ln851_1_fu_416_p2 = _133_ ? 1'h1 : 1'h0;
assign icmp_ln851_2_fu_485_p2 = _134_ ? 1'h1 : 1'h0;
assign icmp_ln851_3_fu_550_p2 = _135_ ? 1'h1 : 1'h0;
assign icmp_ln851_4_fu_695_p2 = _136_ ? 1'h1 : 1'h0;
assign icmp_ln851_fu_291_p2 = _051_ ? 1'h1 : 1'h0;
assign ret_V_13_fu_338_p3 = ret_V_12_reg_765[6] ? select_ln850_fu_333_p3 : ret_V_cast_reg_770;
assign ret_V_18_fu_651_p3 = ret_V_17_reg_943[33] ? select_ln850_4_fu_645_p3 : ret_V_20_cast_reg_948;
assign ret_V_20_fu_728_p3 = ret_V_19_reg_990[53] ? select_ln850_5_fu_723_p3 : ret_V_22_cast_reg_995;
assign select_ln1192_1_fu_747_p3 = op_19 ? 32'd4294967295 : 32'd0;
assign select_ln1192_fu_735_p3 = op_18 ? 32'd4294967295 : 32'd0;
assign select_ln353_1_fu_518_p3 = ret_V_15_reg_869[34] ? select_ln850_2_fu_513_p3 : ret_V_7_cast_reg_874;
assign select_ln353_2_fu_583_p3 = ret_V_16_reg_906[39] ? select_ln850_3_fu_578_p3 : ret_V_18_cast_reg_911;
assign select_ln353_fu_453_p3 = ret_V_14_reg_827[32] ? select_ln850_1_fu_448_p3 : sext_ln850_reg_837;
assign select_ln69_1_fu_658_p3 = op_16_V_fu_630_p2 ? 32'd4294967295 : 32'd0;
assign select_ln850_1_fu_448_p3 = icmp_ln851_1_reg_822 ? add_ln691_reg_844 : sext_ln850_reg_837;
assign select_ln850_2_fu_513_p3 = icmp_ln851_2_reg_864 ? add_ln691_1_reg_881 : ret_V_7_cast_reg_874;
assign select_ln850_3_fu_578_p3 = icmp_ln851_3_reg_901 ? add_ln691_2_reg_918 : ret_V_18_cast_reg_911;
assign select_ln850_4_fu_645_p3 = op_15[0] ? add_ln691_3_reg_955 : ret_V_20_cast_reg_948;
assign select_ln850_5_fu_723_p3 = icmp_ln851_4_reg_985 ? add_ln691_4_reg_1002 : ret_V_22_cast_reg_995;
assign select_ln850_fu_333_p3 = icmp_ln851_reg_777 ? ret_V_cast_reg_770 : ret_V_reg_792;
assign signbit_fu_315_p2 = _052_ ? 1'h1 : 1'h0;
assign add_ln69_1_fu_377_p0 = { 1'h0, icmp_ln1494_reg_782 };
assign add_ln69_fu_371_p0 = { op_0[3], op_0, icmp_ln1499_reg_760 };
assign add_ln69_fu_371_p1 = { ret_V_13_fu_338_p3[1], ret_V_13_fu_338_p3[1], ret_V_13_fu_338_p3[1], ret_V_13_fu_338_p3[1], ret_V_13_fu_338_p3 };
assign ap_CS_fsm_state1 = ap_CS_fsm[0];
assign ap_CS_fsm_state10 = ap_CS_fsm[9];
assign ap_CS_fsm_state11 = ap_CS_fsm[10];
assign ap_CS_fsm_state12 = ap_CS_fsm[11];
assign ap_CS_fsm_state13 = ap_CS_fsm[12];
assign ap_CS_fsm_state14 = ap_CS_fsm[13];
assign ap_CS_fsm_state15 = ap_CS_fsm[14];
assign ap_CS_fsm_state16 = ap_CS_fsm[15];
assign ap_CS_fsm_state17 = ap_CS_fsm[16];
assign ap_CS_fsm_state18 = ap_CS_fsm[17];
assign ap_CS_fsm_state19 = ap_CS_fsm[18];
assign ap_CS_fsm_state2 = ap_CS_fsm[1];
assign ap_CS_fsm_state20 = ap_CS_fsm[19];
assign ap_CS_fsm_state21 = ap_CS_fsm[20];
assign ap_CS_fsm_state22 = ap_CS_fsm[21];
assign ap_CS_fsm_state23 = ap_CS_fsm[22];
assign ap_CS_fsm_state24 = ap_CS_fsm[23];
assign ap_CS_fsm_state25 = ap_CS_fsm[24];
assign ap_CS_fsm_state26 = ap_CS_fsm[25];
assign ap_CS_fsm_state27 = ap_CS_fsm[26];
assign ap_CS_fsm_state28 = ap_CS_fsm[27];
assign ap_CS_fsm_state29 = ap_CS_fsm[28];
assign ap_CS_fsm_state3 = ap_CS_fsm[2];
assign ap_CS_fsm_state30 = ap_CS_fsm[29];
assign ap_CS_fsm_state31 = ap_CS_fsm[30];
assign ap_CS_fsm_state32 = ap_CS_fsm[31];
assign ap_CS_fsm_state33 = ap_CS_fsm[32];
assign ap_CS_fsm_state34 = ap_CS_fsm[33];
assign ap_CS_fsm_state35 = ap_CS_fsm[34];
assign ap_CS_fsm_state4 = ap_CS_fsm[3];
assign ap_CS_fsm_state5 = ap_CS_fsm[4];
assign ap_CS_fsm_state6 = ap_CS_fsm[5];
assign ap_CS_fsm_state7 = ap_CS_fsm[6];
assign ap_CS_fsm_state8 = ap_CS_fsm[7];
assign ap_CS_fsm_state9 = ap_CS_fsm[8];
assign ap_done = op_31_ap_vld;
assign ap_ready = op_31_ap_vld;
assign grp_fu_406_p0 = { op_23_V_reg_807[5], op_23_V_reg_807[5], op_23_V_reg_807[5], op_23_V_reg_807[5], op_23_V_reg_807[5], op_23_V_reg_807[5], op_23_V_reg_807[5], op_23_V_reg_807[5], op_23_V_reg_807[5], op_23_V_reg_807[5], op_23_V_reg_807[5], op_23_V_reg_807[5], op_23_V_reg_807[5], op_23_V_reg_807[5], op_23_V_reg_807[5], op_23_V_reg_807[5], op_23_V_reg_807[5], op_23_V_reg_807, 10'h000 };
assign grp_fu_406_p1 = { op_12[31], op_12 };
assign grp_fu_435_p0 = { tmp_reg_832[22], tmp_reg_832 };
assign grp_fu_475_p0 = { select_ln353_reg_849[23], select_ln353_reg_849[23], select_ln353_reg_849[23], select_ln353_reg_849[23], select_ln353_reg_849[23], select_ln353_reg_849[23], select_ln353_reg_849[23], select_ln353_reg_849[23], select_ln353_reg_849[23], select_ln353_reg_849, 2'h0 };
assign grp_fu_475_p1 = { op_13[31], op_13[31], op_13[31], op_13 };
assign grp_fu_540_p0 = { select_ln353_1_reg_886[31], select_ln353_1_reg_886, 7'h00 };
assign grp_fu_540_p1 = { op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14 };
assign grp_fu_605_p0 = { select_ln353_2_reg_923[31], select_ln353_2_reg_923, 1'h0 };
assign grp_fu_605_p1 = { op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15 };
assign grp_fu_685_p0 = { op_28_V_reg_970[31], op_28_V_reg_970, 21'h000000 };
assign grp_fu_685_p1 = { op_17[31], op_17[31], op_17[31], op_17[31], op_17[31], op_17[31], op_17[31], op_17[31], op_17[31], op_17[31], op_17[31], op_17[31], op_17[31], op_17[31], op_17[31], op_17[31], op_17[31], op_17[31], op_17[31], op_17[31], op_17[31], op_17[31], op_17 };
assign op_20_V_fu_345_p3 = { op_0, icmp_ln1499_reg_760 };
assign op_23_V_fu_386_p0 = { add_ln69_1_reg_802[1], add_ln69_1_reg_802[1], add_ln69_1_reg_802[1], add_ln69_1_reg_802[1], add_ln69_1_reg_802 };
assign op_31 = grp_fu_755_p2;
assign op_4_V_fu_233_p3 = { op_2, 6'h00 };
assign p_Result_1_fu_441_p3 = ret_V_14_reg_827[32];
assign p_Result_2_fu_506_p3 = ret_V_15_reg_869[34];
assign p_Result_3_fu_571_p3 = ret_V_16_reg_906[39];
assign p_Result_4_fu_635_p3 = ret_V_17_reg_943[33];
assign p_Result_5_fu_716_p3 = ret_V_19_reg_990[53];
assign p_Result_s_fu_326_p3 = ret_V_12_reg_765[6];
assign rhs_2_fu_395_p3 = { op_23_V_reg_807, 10'h000 };
assign rhs_3_fu_529_p3 = { select_ln353_1_reg_886, 7'h00 };
assign rhs_4_fu_594_p3 = { select_ln353_2_reg_923, 1'h0 };
assign rhs_6_fu_674_p3 = { op_28_V_reg_970, 21'h000000 };
assign rhs_fu_263_p3 = { op_5, 3'h0 };
assign sext_ln1192_fu_391_p0 = op_12;
assign sext_ln1494_fu_305_p1 = { op_3[3], op_3, 3'h0 };
assign sext_ln1499_fu_249_p0 = op_3;
assign sext_ln1499_fu_249_p1 = { op_3[3], op_3 };
assign sext_ln703_1_fu_460_p0 = op_13;
assign sext_ln703_2_fu_525_p0 = op_14;
assign sext_ln703_3_fu_590_p0 = op_15;
assign sext_ln703_4_fu_670_p0 = op_17;
assign sext_ln703_fu_259_p0 = op_3;
assign sext_ln703_fu_259_p1 = { op_3[3], op_3[3], op_3[3], op_3 };
assign sext_ln850_fu_432_p1 = { tmp_reg_832[22], tmp_reg_832 };
assign shl_ln728_2_fu_297_p1 = op_3;
assign shl_ln728_2_fu_297_p3 = { op_3, 3'h0 };
assign shl_ln_fu_241_p3 = { op_2, 3'h0 };
assign tmp_3_fu_464_p3 = { select_ln353_reg_849, 2'h0 };
assign trunc_ln1195_fu_626_p1 = op_10[0];
assign trunc_ln851_1_fu_412_p0 = op_12;
assign trunc_ln851_1_fu_412_p1 = op_12[9:0];
assign trunc_ln851_2_fu_481_p0 = op_13;
assign trunc_ln851_2_fu_481_p1 = op_13[1:0];
assign trunc_ln851_3_fu_546_p0 = op_14;
assign trunc_ln851_3_fu_546_p1 = op_14[6:0];
assign trunc_ln851_4_fu_642_p0 = op_15;
assign trunc_ln851_4_fu_642_p1 = op_15[0];
assign trunc_ln851_5_fu_691_p0 = op_17;
assign trunc_ln851_5_fu_691_p1 = op_17[20:0];
assign trunc_ln851_fu_287_p1 = ret_V_12_fu_271_p2[2:0];
assign \add_6s_6s_6_1_1_U2.top_add_6s_6s_6_1_1_Adder_1_U.a  = \add_6s_6s_6_1_1_U2.din0 ;
assign \add_6s_6s_6_1_1_U2.top_add_6s_6s_6_1_1_Adder_1_U.b  = \add_6s_6s_6_1_1_U2.din1 ;
assign \add_6s_6s_6_1_1_U2.dout  = \add_6s_6s_6_1_1_U2.top_add_6s_6s_6_1_1_Adder_1_U.s ;
assign \add_6s_6s_6_1_1_U2.din0  = { op_0[3], op_0, icmp_ln1499_reg_760 };
assign \add_6s_6s_6_1_1_U2.din1  = { ret_V_13_fu_338_p3[1], ret_V_13_fu_338_p3[1], ret_V_13_fu_338_p3[1], ret_V_13_fu_338_p3[1], ret_V_13_fu_338_p3 };
assign add_ln69_fu_371_p2 = \add_6s_6s_6_1_1_U2.dout ;
assign \add_6s_6ns_6_1_1_U4.top_add_6s_6ns_6_1_1_Adder_2_U.a  = \add_6s_6ns_6_1_1_U4.din0 ;
assign \add_6s_6ns_6_1_1_U4.top_add_6s_6ns_6_1_1_Adder_2_U.b  = \add_6s_6ns_6_1_1_U4.din1 ;
assign \add_6s_6ns_6_1_1_U4.dout  = \add_6s_6ns_6_1_1_U4.top_add_6s_6ns_6_1_1_Adder_2_U.s ;
assign \add_6s_6ns_6_1_1_U4.din0  = { add_ln69_1_reg_802[1], add_ln69_1_reg_802[1], add_ln69_1_reg_802[1], add_ln69_1_reg_802[1], add_ln69_1_reg_802 };
assign \add_6s_6ns_6_1_1_U4.din1  = add_ln69_reg_797;
assign op_23_V_fu_386_p2 = \add_6s_6ns_6_1_1_U4.dout ;
assign \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.ain_s0  = \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.a ;
assign \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.bin_s0  = \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.b ;
assign \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.s  = { \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.fas_s2 , \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.sum_s1  };
assign \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.u2.a  = \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.ain_s1 ;
assign \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.u2.b  = \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.bin_s1 ;
assign \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.u2.cin  = \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.carry_s1 ;
assign \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.facout_s2  = \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.u2.cout ;
assign \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.fas_s2  = \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.u2.s ;
assign \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.u1.a  = \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.a [26:0];
assign \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.u1.b  = \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.b [26:0];
assign \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.u1.cin  = 1'h0;
assign \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.facout_s1  = \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.u1.cout ;
assign \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.fas_s1  = \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.u1.s ;
assign \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.a  = \add_54s_54s_54_2_1_U14.din0 ;
assign \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.b  = \add_54s_54s_54_2_1_U14.din1 ;
assign \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.ce  = \add_54s_54s_54_2_1_U14.ce ;
assign \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.clk  = \add_54s_54s_54_2_1_U14.clk ;
assign \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.reset  = \add_54s_54s_54_2_1_U14.reset ;
assign \add_54s_54s_54_2_1_U14.dout  = \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_9_U.s ;
assign \add_54s_54s_54_2_1_U14.ce  = 1'h1;
assign \add_54s_54s_54_2_1_U14.clk  = ap_clk;
assign \add_54s_54s_54_2_1_U14.din0  = { op_28_V_reg_970[31], op_28_V_reg_970, 21'h000000 };
assign \add_54s_54s_54_2_1_U14.din1  = { op_17[31], op_17[31], op_17[31], op_17[31], op_17[31], op_17[31], op_17[31], op_17[31], op_17[31], op_17[31], op_17[31], op_17[31], op_17[31], op_17[31], op_17[31], op_17[31], op_17[31], op_17[31], op_17[31], op_17[31], op_17[31], op_17[31], op_17 };
assign grp_fu_685_p2 = \add_54s_54s_54_2_1_U14.dout ;
assign \add_54s_54s_54_2_1_U14.reset  = ap_rst;
assign \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.ain_s0  = \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.a ;
assign \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.bin_s0  = \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.b ;
assign \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.s  = { \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.fas_s2 , \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.sum_s1  };
assign \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.u2.a  = \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.ain_s1 ;
assign \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.u2.b  = \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.bin_s1 ;
assign \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.u2.cin  = \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.carry_s1 ;
assign \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.facout_s2  = \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.u2.cout ;
assign \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.fas_s2  = \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.u2.s ;
assign \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.u1.a  = \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.a [19:0];
assign \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.u1.b  = \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.b [19:0];
assign \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.u1.cin  = 1'h0;
assign \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.facout_s1  = \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.u1.cout ;
assign \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.fas_s1  = \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.u1.s ;
assign \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.a  = \add_40s_40s_40_2_1_U9.din0 ;
assign \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.b  = \add_40s_40s_40_2_1_U9.din1 ;
assign \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.ce  = \add_40s_40s_40_2_1_U9.ce ;
assign \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.clk  = \add_40s_40s_40_2_1_U9.clk ;
assign \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.reset  = \add_40s_40s_40_2_1_U9.reset ;
assign \add_40s_40s_40_2_1_U9.dout  = \add_40s_40s_40_2_1_U9.top_add_40s_40s_40_2_1_Adder_7_U.s ;
assign \add_40s_40s_40_2_1_U9.ce  = 1'h1;
assign \add_40s_40s_40_2_1_U9.clk  = ap_clk;
assign \add_40s_40s_40_2_1_U9.din0  = { select_ln353_1_reg_886[31], select_ln353_1_reg_886, 7'h00 };
assign \add_40s_40s_40_2_1_U9.din1  = { op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14 };
assign grp_fu_540_p2 = \add_40s_40s_40_2_1_U9.dout ;
assign \add_40s_40s_40_2_1_U9.reset  = ap_rst;
assign \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.ain_s0  = \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.a ;
assign \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.bin_s0  = \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.b ;
assign \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.s  = { \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.fas_s2 , \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.sum_s1  };
assign \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.u2.a  = \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.ain_s1 ;
assign \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.u2.b  = \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.bin_s1 ;
assign \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.u2.cin  = \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.carry_s1 ;
assign \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.facout_s2  = \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.u2.cout ;
assign \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.fas_s2  = \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.u2.s ;
assign \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.u1.a  = \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.a [16:0];
assign \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.u1.b  = \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.b [16:0];
assign \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.u1.cin  = 1'h0;
assign \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.facout_s1  = \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.u1.cout ;
assign \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.fas_s1  = \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.u1.s ;
assign \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.a  = \add_35s_35s_35_2_1_U7.din0 ;
assign \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.b  = \add_35s_35s_35_2_1_U7.din1 ;
assign \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.ce  = \add_35s_35s_35_2_1_U7.ce ;
assign \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.clk  = \add_35s_35s_35_2_1_U7.clk ;
assign \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.reset  = \add_35s_35s_35_2_1_U7.reset ;
assign \add_35s_35s_35_2_1_U7.dout  = \add_35s_35s_35_2_1_U7.top_add_35s_35s_35_2_1_Adder_5_U.s ;
assign \add_35s_35s_35_2_1_U7.ce  = 1'h1;
assign \add_35s_35s_35_2_1_U7.clk  = ap_clk;
assign \add_35s_35s_35_2_1_U7.din0  = { select_ln353_reg_849[23], select_ln353_reg_849[23], select_ln353_reg_849[23], select_ln353_reg_849[23], select_ln353_reg_849[23], select_ln353_reg_849[23], select_ln353_reg_849[23], select_ln353_reg_849[23], select_ln353_reg_849[23], select_ln353_reg_849, 2'h0 };
assign \add_35s_35s_35_2_1_U7.din1  = { op_13[31], op_13[31], op_13[31], op_13 };
assign grp_fu_475_p2 = \add_35s_35s_35_2_1_U7.dout ;
assign \add_35s_35s_35_2_1_U7.reset  = ap_rst;
assign \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.ain_s0  = \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.a ;
assign \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.bin_s0  = \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.b ;
assign \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.s  = { \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.fas_s2 , \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.sum_s1  };
assign \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.u2.a  = \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.ain_s1 ;
assign \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.u2.b  = \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.bin_s1 ;
assign \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.u2.cin  = \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.carry_s1 ;
assign \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.facout_s2  = \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.u2.cout ;
assign \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.fas_s2  = \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.u2.s ;
assign \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.u1.a  = \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.a [16:0];
assign \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.u1.b  = \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.b [16:0];
assign \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.u1.cin  = 1'h0;
assign \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.facout_s1  = \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.u1.cout ;
assign \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.fas_s1  = \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.u1.s ;
assign \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.a  = \add_34s_34s_34_2_1_U11.din0 ;
assign \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.b  = \add_34s_34s_34_2_1_U11.din1 ;
assign \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.ce  = \add_34s_34s_34_2_1_U11.ce ;
assign \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.clk  = \add_34s_34s_34_2_1_U11.clk ;
assign \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.reset  = \add_34s_34s_34_2_1_U11.reset ;
assign \add_34s_34s_34_2_1_U11.dout  = \add_34s_34s_34_2_1_U11.top_add_34s_34s_34_2_1_Adder_8_U.s ;
assign \add_34s_34s_34_2_1_U11.ce  = 1'h1;
assign \add_34s_34s_34_2_1_U11.clk  = ap_clk;
assign \add_34s_34s_34_2_1_U11.din0  = { select_ln353_2_reg_923[31], select_ln353_2_reg_923, 1'h0 };
assign \add_34s_34s_34_2_1_U11.din1  = { op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15 };
assign grp_fu_605_p2 = \add_34s_34s_34_2_1_U11.dout ;
assign \add_34s_34s_34_2_1_U11.reset  = ap_rst;
assign \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.ain_s0  = \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.a ;
assign \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.bin_s0  = \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.b ;
assign \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.s  = { \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.fas_s2 , \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.sum_s1  };
assign \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.u2.a  = \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.ain_s1 ;
assign \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.u2.b  = \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.bin_s1 ;
assign \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.u2.cin  = \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.carry_s1 ;
assign \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.facout_s2  = \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.u2.cout ;
assign \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.fas_s2  = \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.u2.s ;
assign \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.u1.a  = \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.a [15:0];
assign \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.u1.b  = \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.b [15:0];
assign \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.u1.cin  = 1'h0;
assign \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.facout_s1  = \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.u1.cout ;
assign \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.fas_s1  = \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.u1.s ;
assign \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.a  = \add_33s_33s_33_2_1_U5.din0 ;
assign \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.b  = \add_33s_33s_33_2_1_U5.din1 ;
assign \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.ce  = \add_33s_33s_33_2_1_U5.ce ;
assign \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.clk  = \add_33s_33s_33_2_1_U5.clk ;
assign \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.reset  = \add_33s_33s_33_2_1_U5.reset ;
assign \add_33s_33s_33_2_1_U5.dout  = \add_33s_33s_33_2_1_U5.top_add_33s_33s_33_2_1_Adder_3_U.s ;
assign \add_33s_33s_33_2_1_U5.ce  = 1'h1;
assign \add_33s_33s_33_2_1_U5.clk  = ap_clk;
assign \add_33s_33s_33_2_1_U5.din0  = { op_23_V_reg_807[5], op_23_V_reg_807[5], op_23_V_reg_807[5], op_23_V_reg_807[5], op_23_V_reg_807[5], op_23_V_reg_807[5], op_23_V_reg_807[5], op_23_V_reg_807[5], op_23_V_reg_807[5], op_23_V_reg_807[5], op_23_V_reg_807[5], op_23_V_reg_807[5], op_23_V_reg_807[5], op_23_V_reg_807[5], op_23_V_reg_807[5], op_23_V_reg_807[5], op_23_V_reg_807[5], op_23_V_reg_807, 10'h000 };
assign \add_33s_33s_33_2_1_U5.din1  = { op_12[31], op_12 };
assign grp_fu_406_p2 = \add_33s_33s_33_2_1_U5.dout ;
assign \add_33s_33s_33_2_1_U5.reset  = ap_rst;
assign \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s0  = \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.a ;
assign \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s0  = \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.b ;
assign \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.s  = { \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s2 , \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.sum_s1  };
assign \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.a  = \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s1 ;
assign \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.b  = \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s1 ;
assign \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cin  = \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.carry_s1 ;
assign \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s2  = \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cout ;
assign \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s2  = \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.s ;
assign \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.a  = \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.a [15:0];
assign \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.b  = \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.b [15:0];
assign \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cin  = 1'h0;
assign \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s1  = \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cout ;
assign \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s1  = \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.s ;
assign \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.a  = \add_32ns_32ns_32_2_1_U8.din0 ;
assign \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.b  = \add_32ns_32ns_32_2_1_U8.din1 ;
assign \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  = \add_32ns_32ns_32_2_1_U8.ce ;
assign \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.clk  = \add_32ns_32ns_32_2_1_U8.clk ;
assign \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.reset  = \add_32ns_32ns_32_2_1_U8.reset ;
assign \add_32ns_32ns_32_2_1_U8.dout  = \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.s ;
assign \add_32ns_32ns_32_2_1_U8.ce  = 1'h1;
assign \add_32ns_32ns_32_2_1_U8.clk  = ap_clk;
assign \add_32ns_32ns_32_2_1_U8.din0  = ret_V_7_cast_reg_874;
assign \add_32ns_32ns_32_2_1_U8.din1  = 32'd1;
assign grp_fu_501_p2 = \add_32ns_32ns_32_2_1_U8.dout ;
assign \add_32ns_32ns_32_2_1_U8.reset  = ap_rst;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s0  = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.a ;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s0  = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.b ;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.s  = { \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s2 , \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.sum_s1  };
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.a  = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s1 ;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.b  = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s1 ;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cin  = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.carry_s1 ;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s2  = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cout ;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s2  = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.s ;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.a  = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.a [15:0];
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.b  = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.b [15:0];
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cin  = 1'h0;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s1  = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cout ;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s1  = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.s ;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.a  = \add_32ns_32ns_32_2_1_U17.din0 ;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.b  = \add_32ns_32ns_32_2_1_U17.din1 ;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  = \add_32ns_32ns_32_2_1_U17.ce ;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.clk  = \add_32ns_32ns_32_2_1_U17.clk ;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.reset  = \add_32ns_32ns_32_2_1_U17.reset ;
assign \add_32ns_32ns_32_2_1_U17.dout  = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.s ;
assign \add_32ns_32ns_32_2_1_U17.ce  = 1'h1;
assign \add_32ns_32ns_32_2_1_U17.clk  = ap_clk;
assign \add_32ns_32ns_32_2_1_U17.din0  = ret_V_21_reg_1017;
assign \add_32ns_32ns_32_2_1_U17.din1  = select_ln1192_1_reg_1022;
assign grp_fu_755_p2 = \add_32ns_32ns_32_2_1_U17.dout ;
assign \add_32ns_32ns_32_2_1_U17.reset  = ap_rst;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s0  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.a ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s0  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.b ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.s  = { \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s2 , \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.sum_s1  };
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.a  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s1 ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.b  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s1 ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cin  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.carry_s1 ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s2  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cout ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s2  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.s ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.a  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.a [15:0];
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.b  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.b [15:0];
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cin  = 1'h0;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s1  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cout ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s1  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.s ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.a  = \add_32ns_32ns_32_2_1_U16.din0 ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.b  = \add_32ns_32ns_32_2_1_U16.din1 ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  = \add_32ns_32ns_32_2_1_U16.ce ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.clk  = \add_32ns_32ns_32_2_1_U16.clk ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.reset  = \add_32ns_32ns_32_2_1_U16.reset ;
assign \add_32ns_32ns_32_2_1_U16.dout  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.s ;
assign \add_32ns_32ns_32_2_1_U16.ce  = 1'h1;
assign \add_32ns_32ns_32_2_1_U16.clk  = ap_clk;
assign \add_32ns_32ns_32_2_1_U16.din0  = ret_V_20_reg_1007;
assign \add_32ns_32ns_32_2_1_U16.din1  = select_ln1192_reg_1012;
assign grp_fu_743_p2 = \add_32ns_32ns_32_2_1_U16.dout ;
assign \add_32ns_32ns_32_2_1_U16.reset  = ap_rst;
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s0  = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.a ;
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s0  = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.b ;
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.s  = { \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s2 , \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.sum_s1  };
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.a  = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s1 ;
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.b  = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s1 ;
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cin  = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.carry_s1 ;
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s2  = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cout ;
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s2  = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.s ;
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.a  = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.a [15:0];
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.b  = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.b [15:0];
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cin  = 1'h0;
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s1  = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cout ;
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s1  = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.s ;
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.a  = \add_32ns_32ns_32_2_1_U15.din0 ;
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.b  = \add_32ns_32ns_32_2_1_U15.din1 ;
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  = \add_32ns_32ns_32_2_1_U15.ce ;
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.clk  = \add_32ns_32ns_32_2_1_U15.clk ;
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.reset  = \add_32ns_32ns_32_2_1_U15.reset ;
assign \add_32ns_32ns_32_2_1_U15.dout  = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_6_U.s ;
assign \add_32ns_32ns_32_2_1_U15.ce  = 1'h1;
assign \add_32ns_32ns_32_2_1_U15.clk  = ap_clk;
assign \add_32ns_32ns_32_2_1_U15.din0  = ret_V_22_cast_reg_995;
assign \add_32ns_32ns_32_2_1_U15.din1  = 32'd1;
assign grp_fu_711_p2 = \add_32ns_32ns_32_2_1_U15.dout ;
assign \add_32ns_32ns_32_2_1_U15.reset  = ap_rst;
assign \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s0  = \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.a ;
assign \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s0  = \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.b ;
assign \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.s  = { \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s2 , \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.sum_s1  };
assign \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.a  = \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s1 ;
assign \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.b  = \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s1 ;
assign \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cin  = \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.carry_s1 ;
assign \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s2  = \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cout ;
assign \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s2  = \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.s ;
assign \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.a  = \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.a [15:0];
assign \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.b  = \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.b [15:0];
assign \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cin  = 1'h0;
assign \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s1  = \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cout ;
assign \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s1  = \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.s ;
assign \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.a  = \add_32ns_32ns_32_2_1_U13.din0 ;
assign \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.b  = \add_32ns_32ns_32_2_1_U13.din1 ;
assign \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  = \add_32ns_32ns_32_2_1_U13.ce ;
assign \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.clk  = \add_32ns_32ns_32_2_1_U13.clk ;
assign \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.reset  = \add_32ns_32ns_32_2_1_U13.reset ;
assign \add_32ns_32ns_32_2_1_U13.dout  = \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.s ;
assign \add_32ns_32ns_32_2_1_U13.ce  = 1'h1;
assign \add_32ns_32ns_32_2_1_U13.clk  = ap_clk;
assign \add_32ns_32ns_32_2_1_U13.din0  = ret_V_18_reg_960;
assign \add_32ns_32ns_32_2_1_U13.din1  = select_ln69_1_reg_965;
assign grp_fu_666_p2 = \add_32ns_32ns_32_2_1_U13.dout ;
assign \add_32ns_32ns_32_2_1_U13.reset  = ap_rst;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s0  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.a ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s0  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.b ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.s  = { \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s2 , \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.sum_s1  };
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.a  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s1 ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.b  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s1 ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cin  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.carry_s1 ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s2  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cout ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s2  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.s ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.a  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.a [15:0];
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.b  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.b [15:0];
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cin  = 1'h0;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s1  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cout ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s1  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.s ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.a  = \add_32ns_32ns_32_2_1_U12.din0 ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.b  = \add_32ns_32ns_32_2_1_U12.din1 ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  = \add_32ns_32ns_32_2_1_U12.ce ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.clk  = \add_32ns_32ns_32_2_1_U12.clk ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.reset  = \add_32ns_32ns_32_2_1_U12.reset ;
assign \add_32ns_32ns_32_2_1_U12.dout  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_6_U.s ;
assign \add_32ns_32ns_32_2_1_U12.ce  = 1'h1;
assign \add_32ns_32ns_32_2_1_U12.clk  = ap_clk;
assign \add_32ns_32ns_32_2_1_U12.din0  = ret_V_20_cast_reg_948;
assign \add_32ns_32ns_32_2_1_U12.din1  = 32'd1;
assign grp_fu_621_p2 = \add_32ns_32ns_32_2_1_U12.dout ;
assign \add_32ns_32ns_32_2_1_U12.reset  = ap_rst;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s0  = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.a ;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s0  = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.b ;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.s  = { \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s2 , \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.sum_s1  };
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.a  = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s1 ;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.b  = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s1 ;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cin  = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.carry_s1 ;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s2  = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cout ;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s2  = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.s ;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.a  = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.a [15:0];
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.b  = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.b [15:0];
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cin  = 1'h0;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s1  = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cout ;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s1  = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.s ;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.a  = \add_32ns_32ns_32_2_1_U10.din0 ;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.b  = \add_32ns_32ns_32_2_1_U10.din1 ;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  = \add_32ns_32ns_32_2_1_U10.ce ;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.clk  = \add_32ns_32ns_32_2_1_U10.clk ;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.reset  = \add_32ns_32ns_32_2_1_U10.reset ;
assign \add_32ns_32ns_32_2_1_U10.dout  = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.s ;
assign \add_32ns_32ns_32_2_1_U10.ce  = 1'h1;
assign \add_32ns_32ns_32_2_1_U10.clk  = ap_clk;
assign \add_32ns_32ns_32_2_1_U10.din0  = ret_V_18_cast_reg_911;
assign \add_32ns_32ns_32_2_1_U10.din1  = 32'd1;
assign grp_fu_566_p2 = \add_32ns_32ns_32_2_1_U10.dout ;
assign \add_32ns_32ns_32_2_1_U10.reset  = ap_rst;
assign \add_2ns_2ns_2_1_1_U3.top_add_2ns_2ns_2_1_1_Adder_0_U.a  = \add_2ns_2ns_2_1_1_U3.din0 ;
assign \add_2ns_2ns_2_1_1_U3.top_add_2ns_2ns_2_1_1_Adder_0_U.b  = \add_2ns_2ns_2_1_1_U3.din1 ;
assign \add_2ns_2ns_2_1_1_U3.dout  = \add_2ns_2ns_2_1_1_U3.top_add_2ns_2ns_2_1_1_Adder_0_U.s ;
assign \add_2ns_2ns_2_1_1_U3.din0  = { 1'h0, icmp_ln1494_reg_782 };
assign \add_2ns_2ns_2_1_1_U3.din1  = add_ln69_1_fu_377_p1;
assign add_ln69_1_fu_377_p2 = \add_2ns_2ns_2_1_1_U3.dout ;
assign \add_2ns_2ns_2_1_1_U1.top_add_2ns_2ns_2_1_1_Adder_0_U.a  = \add_2ns_2ns_2_1_1_U1.din0 ;
assign \add_2ns_2ns_2_1_1_U1.top_add_2ns_2ns_2_1_1_Adder_0_U.b  = \add_2ns_2ns_2_1_1_U1.din1 ;
assign \add_2ns_2ns_2_1_1_U1.dout  = \add_2ns_2ns_2_1_1_U1.top_add_2ns_2ns_2_1_1_Adder_0_U.s ;
assign \add_2ns_2ns_2_1_1_U1.din0  = ret_V_cast_reg_770;
assign \add_2ns_2ns_2_1_1_U1.din1  = 2'h1;
assign ret_V_fu_321_p2 = \add_2ns_2ns_2_1_1_U1.dout ;
assign \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.ain_s0  = \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.a ;
assign \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.bin_s0  = \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.b ;
assign \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.s  = { \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.fas_s2 , \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.sum_s1  };
assign \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.u2.a  = \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.ain_s1 ;
assign \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.u2.b  = \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.bin_s1 ;
assign \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.u2.cin  = \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.carry_s1 ;
assign \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.facout_s2  = \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.u2.cout ;
assign \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.fas_s2  = \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.u2.s ;
assign \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.u1.a  = \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.a [11:0];
assign \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.u1.b  = \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.b [11:0];
assign \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.u1.cin  = 1'h0;
assign \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.facout_s1  = \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.u1.cout ;
assign \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.fas_s1  = \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.u1.s ;
assign \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.a  = \add_24s_24ns_24_2_1_U6.din0 ;
assign \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.b  = \add_24s_24ns_24_2_1_U6.din1 ;
assign \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.ce  = \add_24s_24ns_24_2_1_U6.ce ;
assign \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.clk  = \add_24s_24ns_24_2_1_U6.clk ;
assign \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.reset  = \add_24s_24ns_24_2_1_U6.reset ;
assign \add_24s_24ns_24_2_1_U6.dout  = \add_24s_24ns_24_2_1_U6.top_add_24s_24ns_24_2_1_Adder_4_U.s ;
assign \add_24s_24ns_24_2_1_U6.ce  = 1'h1;
assign \add_24s_24ns_24_2_1_U6.clk  = ap_clk;
assign \add_24s_24ns_24_2_1_U6.din0  = { tmp_reg_832[22], tmp_reg_832 };
assign \add_24s_24ns_24_2_1_U6.din1  = 24'h000001;
assign grp_fu_435_p2 = \add_24s_24ns_24_2_1_U6.dout ;
assign \add_24s_24ns_24_2_1_U6.reset  = ap_rst;
endmodule


// Product machine:
module top_A_times_top_B (ap_start, op_0, op_10, op_11, op_12, op_13, op_14, op_15, op_17, op_18, op_19, op_2, op_3, op_5, ap_clk, unsafe_signal);
input ap_start;
input [3:0] op_0;
input [1:0] op_10;
input op_11;
input [31:0] op_12;
input [31:0] op_13;
input [7:0] op_14;
input [3:0] op_15;
input [31:0] op_17;
input op_18;
input op_19;
input [1:0] op_2;
input [3:0] op_3;
input [3:0] op_5;
input ap_clk;
output unsafe_signal;
reg _setup;
initial _setup = 1'b0;
always @ (posedge ap_clk) _setup <= 1'b1;
reg ap_start_internal;
always @ (posedge ap_clk) if (!_setup) ap_start_internal <= ap_start;
reg [3:0] op_0_internal;
always @ (posedge ap_clk) if (!_setup) op_0_internal <= op_0;
reg [1:0] op_10_internal;
always @ (posedge ap_clk) if (!_setup) op_10_internal <= op_10;
reg op_11_internal;
always @ (posedge ap_clk) if (!_setup) op_11_internal <= op_11;
reg [31:0] op_12_internal;
always @ (posedge ap_clk) if (!_setup) op_12_internal <= op_12;
reg [31:0] op_13_internal;
always @ (posedge ap_clk) if (!_setup) op_13_internal <= op_13;
reg [7:0] op_14_internal;
always @ (posedge ap_clk) if (!_setup) op_14_internal <= op_14;
reg [3:0] op_15_internal;
always @ (posedge ap_clk) if (!_setup) op_15_internal <= op_15;
reg [31:0] op_17_internal;
always @ (posedge ap_clk) if (!_setup) op_17_internal <= op_17;
reg op_18_internal;
always @ (posedge ap_clk) if (!_setup) op_18_internal <= op_18;
reg op_19_internal;
always @ (posedge ap_clk) if (!_setup) op_19_internal <= op_19;
reg [1:0] op_2_internal;
always @ (posedge ap_clk) if (!_setup) op_2_internal <= op_2;
reg [3:0] op_3_internal;
always @ (posedge ap_clk) if (!_setup) op_3_internal <= op_3;
reg [3:0] op_5_internal;
always @ (posedge ap_clk) if (!_setup) op_5_internal <= op_5;
wire ap_done_A;
wire ap_done_B;
wire ap_done_eq;
assign ap_done_eq = ap_done_A == ap_done_B;
wire ap_idle_A;
wire ap_idle_B;
wire ap_idle_eq;
assign ap_idle_eq = ap_idle_A == ap_idle_B;
wire ap_ready_A;
wire ap_ready_B;
wire ap_ready_eq;
assign ap_ready_eq = ap_ready_A == ap_ready_B;
wire [31:0] op_31_A;
wire [31:0] op_31_B;
wire op_31_eq;
assign op_31_eq = op_31_A == op_31_B;
wire op_31_ap_vld_A;
wire op_31_ap_vld_B;
wire clk_enable_A;
wire clk_enable_B;
assign clk_enable_A = _setup & (~op_31_ap_vld_A | op_31_ap_vld_B);
assign clk_enable_B = _setup;
wire divergent;
assign divergent = ~(ap_done_eq & ap_idle_eq & ap_ready_eq & op_31_eq);
assign unsafe_signal = op_31_ap_vld_A & op_31_ap_vld_B & divergent;
top_A instance_A (
    .ap_clk(ap_clk),
    .clk_enable(clk_enable_A),
    .ap_start(ap_start_internal),
    .op_0(op_0_internal),
    .op_10(op_10_internal),
    .op_11(op_11_internal),
    .op_12(op_12_internal),
    .op_13(op_13_internal),
    .op_14(op_14_internal),
    .op_15(op_15_internal),
    .op_17(op_17_internal),
    .op_18(op_18_internal),
    .op_19(op_19_internal),
    .op_2(op_2_internal),
    .op_3(op_3_internal),
    .op_5(op_5_internal),
    .ap_done(ap_done_A),
    .ap_idle(ap_idle_A),
    .ap_ready(ap_ready_A),
    .op_31(op_31_A),
    .op_31_ap_vld(op_31_ap_vld_A)
);
top_B instance_B (
    .ap_clk(ap_clk),
    .clk_enable(clk_enable_B),
    .ap_start(ap_start_internal),
    .op_0(op_0_internal),
    .op_10(op_10_internal),
    .op_11(op_11_internal),
    .op_12(op_12_internal),
    .op_13(op_13_internal),
    .op_14(op_14_internal),
    .op_15(op_15_internal),
    .op_17(op_17_internal),
    .op_18(op_18_internal),
    .op_19(op_19_internal),
    .op_2(op_2_internal),
    .op_3(op_3_internal),
    .op_5(op_5_internal),
    .ap_done(ap_done_B),
    .ap_idle(ap_idle_B),
    .ap_ready(ap_ready_B),
    .op_31(op_31_B),
    .op_31_ap_vld(op_31_ap_vld_B)
);
endmodule
