// Processed by function `construct_kairos` in `verilog_tricks.py`.
// Machine A:
// Processed by function `add_clk_enable_signal` in `verilog_tricks.py`.
// Processed by function `remove_reset_signal` in `verilog_tricks.py`.
module top_A (
  ap_clk,
  ap_start,
  ap_done,
  ap_idle,
  ap_ready,
  op_0,
  op_2,
  op_3,
  op_4,
  op_5,
  op_6,
  op_7,
  op_8,
  op_10,
  op_12,
  op_13,
  op_14,
  op_15,
  op_19,
  op_31,
  op_31_ap_vld,
clk_enable
);
input clk_enable;


input ap_clk;
wire ap_rst;
assign ap_rst = op_31_ap_vld;
input ap_start;
input [3:0] op_0;
input [3:0] op_10;
input [15:0] op_12;
input [15:0] op_13;
input [3:0] op_14;
input [7:0] op_15;
input [31:0] op_19;
input [7:0] op_2;
input [7:0] op_3;
input [15:0] op_4;
input [7:0] op_5;
input [3:0] op_6;
input [7:0] op_7;
input [3:0] op_8;
output ap_done;
output ap_idle;
output ap_ready;
output [31:0] op_31;
output op_31_ap_vld;


reg [4:0] \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.ain_s1 ;
reg [4:0] \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.bin_s1 ;
reg \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.carry_s1 ;
reg [4:0] \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.sum_s1 ;
reg [4:0] \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.ain_s1 ;
reg [4:0] \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.bin_s1 ;
reg \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.carry_s1 ;
reg [4:0] \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.sum_s1 ;
reg [5:0] \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.ain_s1 ;
reg [5:0] \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.bin_s1 ;
reg \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.carry_s1 ;
reg [5:0] \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.sum_s1 ;
reg [8:0] \add_17s_17s_17_2_1_U22.top_add_17s_17s_17_2_1_Adder_13_U.ain_s1 ;
reg [8:0] \add_17s_17s_17_2_1_U22.top_add_17s_17s_17_2_1_Adder_13_U.bin_s1 ;
reg \add_17s_17s_17_2_1_U22.top_add_17s_17s_17_2_1_Adder_13_U.carry_s1 ;
reg [7:0] \add_17s_17s_17_2_1_U22.top_add_17s_17s_17_2_1_Adder_13_U.sum_s1 ;
reg \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_10_U.ain_s1 ;
reg \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_10_U.bin_s1 ;
reg \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_10_U.carry_s1 ;
reg \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_10_U.sum_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.ain_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.bin_s1 ;
reg \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.carry_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.sum_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_5_U.ain_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_5_U.bin_s1 ;
reg \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_5_U.carry_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_5_U.sum_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_5_U.ain_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_5_U.bin_s1 ;
reg \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_5_U.carry_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_5_U.sum_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_5_U.ain_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_5_U.bin_s1 ;
reg \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_5_U.carry_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_5_U.sum_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.ain_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.bin_s1 ;
reg \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.carry_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.sum_s1 ;
reg [15:0] \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_14_U.ain_s1 ;
reg [15:0] \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_14_U.bin_s1 ;
reg \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_14_U.carry_s1 ;
reg [15:0] \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_14_U.sum_s1 ;
reg [16:0] \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.ain_s1 ;
reg [16:0] \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.bin_s1 ;
reg \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.carry_s1 ;
reg [16:0] \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.sum_s1 ;
reg [17:0] \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.ain_s1 ;
reg [17:0] \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.bin_s1 ;
reg \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.carry_s1 ;
reg [16:0] \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.sum_s1 ;
reg [1:0] \add_3s_3ns_3_2_1_U20.top_add_3s_3ns_3_2_1_Adder_12_U.ain_s1 ;
reg [1:0] \add_3s_3ns_3_2_1_U20.top_add_3s_3ns_3_2_1_Adder_12_U.bin_s1 ;
reg \add_3s_3ns_3_2_1_U20.top_add_3s_3ns_3_2_1_Adder_12_U.carry_s1 ;
reg \add_3s_3ns_3_2_1_U20.top_add_3s_3ns_3_2_1_Adder_12_U.sum_s1 ;
reg [22:0] \add_45s_45s_45_2_1_U8.top_add_45s_45s_45_2_1_Adder_7_U.ain_s1 ;
reg [22:0] \add_45s_45s_45_2_1_U8.top_add_45s_45s_45_2_1_Adder_7_U.bin_s1 ;
reg \add_45s_45s_45_2_1_U8.top_add_45s_45s_45_2_1_Adder_7_U.carry_s1 ;
reg [21:0] \add_45s_45s_45_2_1_U8.top_add_45s_45s_45_2_1_Adder_7_U.sum_s1 ;
reg [22:0] \add_46s_46s_46_2_1_U5.top_add_46s_46s_46_2_1_Adder_4_U.ain_s1 ;
reg [22:0] \add_46s_46s_46_2_1_U5.top_add_46s_46s_46_2_1_Adder_4_U.bin_s1 ;
reg \add_46s_46s_46_2_1_U5.top_add_46s_46s_46_2_1_Adder_4_U.carry_s1 ;
reg [22:0] \add_46s_46s_46_2_1_U5.top_add_46s_46s_46_2_1_Adder_4_U.sum_s1 ;
reg [4:0] \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.ain_s1 ;
reg [4:0] \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.bin_s1 ;
reg \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.carry_s1 ;
reg [3:0] \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.sum_s1 ;
reg [31:0] add_ln691_1_reg_930;
reg [31:0] add_ln691_2_reg_1027;
reg [31:0] add_ln691_3_reg_1089;
reg [31:0] add_ln691_4_reg_1173;
reg [9:0] add_ln691_reg_861;
reg [2:0] add_ln69_1_reg_1188;
reg [16:0] add_ln69_2_reg_1213;
reg [31:0] add_ln69_reg_1208;
reg [32:0] ap_CS_fsm = 33'h000000001;
reg [3:0] \ashr_16ns_4ns_16_7_1_U14.din1_cast_array[0] ;
reg [3:0] \ashr_16ns_4ns_16_7_1_U14.din1_cast_array[1] ;
reg [3:0] \ashr_16ns_4ns_16_7_1_U14.din1_cast_array[2] ;
reg [3:0] \ashr_16ns_4ns_16_7_1_U14.din1_cast_array[3] ;
reg [3:0] \ashr_16ns_4ns_16_7_1_U14.din1_cast_array[4] ;
reg [3:0] \ashr_16ns_4ns_16_7_1_U14.din1_cast_array[5] ;
reg [15:0] \ashr_16ns_4ns_16_7_1_U14.dout_array[0] ;
reg [15:0] \ashr_16ns_4ns_16_7_1_U14.dout_array[1] ;
reg [15:0] \ashr_16ns_4ns_16_7_1_U14.dout_array[2] ;
reg [15:0] \ashr_16ns_4ns_16_7_1_U14.dout_array[3] ;
reg [15:0] \ashr_16ns_4ns_16_7_1_U14.dout_array[4] ;
reg [15:0] \ashr_16ns_4ns_16_7_1_U14.dout_array[5] ;
reg [31:0] \ashr_32s_32s_32_7_1_U10.din1_cast_array[0] ;
reg [31:0] \ashr_32s_32s_32_7_1_U10.din1_cast_array[1] ;
reg [31:0] \ashr_32s_32s_32_7_1_U10.din1_cast_array[2] ;
reg [31:0] \ashr_32s_32s_32_7_1_U10.din1_cast_array[3] ;
reg [31:0] \ashr_32s_32s_32_7_1_U10.din1_cast_array[4] ;
reg [31:0] \ashr_32s_32s_32_7_1_U10.din1_cast_array[5] ;
reg [31:0] \ashr_32s_32s_32_7_1_U10.dout_array[0] ;
reg [31:0] \ashr_32s_32s_32_7_1_U10.dout_array[1] ;
reg [31:0] \ashr_32s_32s_32_7_1_U10.dout_array[2] ;
reg [31:0] \ashr_32s_32s_32_7_1_U10.dout_array[3] ;
reg [31:0] \ashr_32s_32s_32_7_1_U10.dout_array[4] ;
reg [31:0] \ashr_32s_32s_32_7_1_U10.dout_array[5] ;
reg [31:0] ashr_ln1333_reg_1079;
reg [15:0] ashr_ln799_reg_1126;
reg icmp_ln850_reg_1022;
reg icmp_ln851_1_reg_839;
reg icmp_ln851_2_reg_902;
reg icmp_ln851_3_reg_961;
reg icmp_ln851_4_reg_1062;
reg icmp_ln851_reg_1131;
reg [3:0] op_11_V_reg_872;
reg [8:0] op_21_V_reg_824;
reg [9:0] op_23_V_reg_887;
reg p_Result_7_reg_989;
reg [15:0] r_1_reg_1146;
reg [7:0] r_reg_919;
reg [11:0] ret_V_14_reg_844;
reg [9:0] ret_V_15_reg_877;
reg [45:0] ret_V_16_reg_907;
reg [44:0] ret_V_17_reg_971;
reg [34:0] ret_V_18_reg_1067;
reg [33:0] ret_V_19_reg_1156;
reg [31:0] ret_V_20_reg_1183;
reg [31:0] ret_V_21_cast_reg_912;
reg [31:0] ret_V_23_cast_reg_976;
reg [31:0] ret_V_25_cast_reg_1072;
reg [31:0] ret_V_27_cast_reg_1161;
reg [1:0] ret_V_3_reg_1151;
reg [1:0] ret_V_4_reg_1168;
reg [1:0] ret_V_reg_1099;
reg [31:0] select_ln1358_reg_1094;
reg [31:0] select_ln353_1_reg_1042;
reg [31:0] select_ln353_2_reg_1111;
reg [31:0] select_ln353_reg_941;
reg [2:0] select_ln69_reg_1047;
reg [8:0] sext_ln15_reg_935;
reg [9:0] sext_ln850_reg_854;
reg [3:0] sh_reg_1017;
reg [3:0] \shl_16ns_4ns_16_7_1_U13.din1_cast_array[0] ;
reg [3:0] \shl_16ns_4ns_16_7_1_U13.din1_cast_array[1] ;
reg [3:0] \shl_16ns_4ns_16_7_1_U13.din1_cast_array[2] ;
reg [3:0] \shl_16ns_4ns_16_7_1_U13.din1_cast_array[3] ;
reg [3:0] \shl_16ns_4ns_16_7_1_U13.din1_cast_array[4] ;
reg [3:0] \shl_16ns_4ns_16_7_1_U13.din1_cast_array[5] ;
reg [15:0] \shl_16ns_4ns_16_7_1_U13.dout_array[0] ;
reg [15:0] \shl_16ns_4ns_16_7_1_U13.dout_array[1] ;
reg [15:0] \shl_16ns_4ns_16_7_1_U13.dout_array[2] ;
reg [15:0] \shl_16ns_4ns_16_7_1_U13.dout_array[3] ;
reg [15:0] \shl_16ns_4ns_16_7_1_U13.dout_array[4] ;
reg [15:0] \shl_16ns_4ns_16_7_1_U13.dout_array[5] ;
reg [31:0] \shl_32s_32s_32_7_1_U11.din1_cast_array[0] ;
reg [31:0] \shl_32s_32s_32_7_1_U11.din1_cast_array[1] ;
reg [31:0] \shl_32s_32s_32_7_1_U11.din1_cast_array[2] ;
reg [31:0] \shl_32s_32s_32_7_1_U11.din1_cast_array[3] ;
reg [31:0] \shl_32s_32s_32_7_1_U11.din1_cast_array[4] ;
reg [31:0] \shl_32s_32s_32_7_1_U11.din1_cast_array[5] ;
reg [31:0] \shl_32s_32s_32_7_1_U11.dout_array[0] ;
reg [31:0] \shl_32s_32s_32_7_1_U11.dout_array[1] ;
reg [31:0] \shl_32s_32s_32_7_1_U11.dout_array[2] ;
reg [31:0] \shl_32s_32s_32_7_1_U11.dout_array[3] ;
reg [31:0] \shl_32s_32s_32_7_1_U11.dout_array[4] ;
reg [31:0] \shl_32s_32s_32_7_1_U11.dout_array[5] ;
reg [31:0] shl_ln1299_reg_1084;
reg [15:0] shl_ln781_reg_1121;
reg [1:0] \sub_4ns_4ns_4_2_1_U9.top_sub_4ns_4ns_4_2_1_Adder_8_U.ain_s1 ;
reg [1:0] \sub_4ns_4ns_4_2_1_U9.top_sub_4ns_4ns_4_2_1_Adder_8_U.bin_s1 ;
reg \sub_4ns_4ns_4_2_1_U9.top_sub_4ns_4ns_4_2_1_Adder_8_U.carry_s1 ;
reg [1:0] \sub_4ns_4ns_4_2_1_U9.top_sub_4ns_4ns_4_2_1_Adder_8_U.sum_s1 ;
reg [4:0] \sub_9ns_9s_9_2_1_U7.top_sub_9ns_9s_9_2_1_Adder_6_U.ain_s1 ;
reg [4:0] \sub_9ns_9s_9_2_1_U7.top_sub_9ns_9s_9_2_1_Adder_6_U.bin_s1 ;
reg \sub_9ns_9s_9_2_1_U7.top_sub_9ns_9s_9_2_1_Adder_6_U.carry_s1 ;
reg [3:0] \sub_9ns_9s_9_2_1_U7.top_sub_9ns_9s_9_2_1_Adder_6_U.sum_s1 ;
reg [8:0] sub_ln1357_reg_946;
reg [8:0] tmp_1_reg_849;
reg tmp_3_reg_924;
reg [5:0] trunc_ln851_1_reg_1106;
reg [5:0] trunc_ln851_reg_1000;
reg [8:0] ush_reg_966;
reg [3:0] _784_;
wire [31:0] _000_;
wire [31:0] _001_;
wire [31:0] _002_;
wire [31:0] _003_;
wire [9:0] _004_;
wire [2:0] _005_;
wire [16:0] _006_;
wire [31:0] _007_;
wire [32:0] _008_;
wire [31:0] _009_;
wire [15:0] _010_;
wire _011_;
wire _012_;
wire _013_;
wire _014_;
wire _015_;
wire _016_;
wire [3:0] _017_;
wire [8:0] _018_;
wire [9:0] _019_;
wire _020_;
wire [15:0] _021_;
wire [7:0] _022_;
wire [3:0] _023_;
wire [11:0] _024_;
wire [9:0] _025_;
wire [45:0] _026_;
wire [44:0] _027_;
wire [34:0] _028_;
wire [33:0] _029_;
wire [31:0] _030_;
wire [31:0] _031_;
wire [31:0] _032_;
wire [31:0] _033_;
wire [31:0] _034_;
wire [1:0] _035_;
wire [1:0] _036_;
wire [1:0] _037_;
wire [31:0] _038_;
wire [31:0] _039_;
wire [31:0] _040_;
wire [31:0] _041_;
wire [2:0] _042_;
wire [8:0] _043_;
wire [9:0] _044_;
wire [3:0] _045_;
wire [31:0] _046_;
wire [15:0] _047_;
wire [8:0] _048_;
wire [8:0] _049_;
wire _050_;
wire [5:0] _051_;
wire [8:0] _052_;
wire [1:0] _053_;
wire _054_;
wire _055_;
wire _056_;
wire _057_;
wire _058_;
wire _059_;
wire _060_;
wire _061_;
wire _062_;
wire _063_;
wire _064_;
wire _065_;
wire _066_;
wire _067_;
wire _068_;
wire [4:0] _069_;
wire [4:0] _070_;
wire _071_;
wire [4:0] _072_;
wire [5:0] _073_;
wire [5:0] _074_;
wire [4:0] _075_;
wire [4:0] _076_;
wire _077_;
wire [4:0] _078_;
wire [5:0] _079_;
wire [5:0] _080_;
wire [5:0] _081_;
wire [5:0] _082_;
wire _083_;
wire [5:0] _084_;
wire [6:0] _085_;
wire [6:0] _086_;
wire [8:0] _087_;
wire [8:0] _088_;
wire _089_;
wire [7:0] _090_;
wire [8:0] _091_;
wire [9:0] _092_;
wire _093_;
wire _094_;
wire _095_;
wire _096_;
wire [1:0] _097_;
wire [1:0] _098_;
wire [15:0] _099_;
wire [15:0] _100_;
wire _101_;
wire [15:0] _102_;
wire [16:0] _103_;
wire [16:0] _104_;
wire [15:0] _105_;
wire [15:0] _106_;
wire _107_;
wire [15:0] _108_;
wire [16:0] _109_;
wire [16:0] _110_;
wire [15:0] _111_;
wire [15:0] _112_;
wire _113_;
wire [15:0] _114_;
wire [16:0] _115_;
wire [16:0] _116_;
wire [15:0] _117_;
wire [15:0] _118_;
wire _119_;
wire [15:0] _120_;
wire [16:0] _121_;
wire [16:0] _122_;
wire [15:0] _123_;
wire [15:0] _124_;
wire _125_;
wire [15:0] _126_;
wire [16:0] _127_;
wire [16:0] _128_;
wire [15:0] _129_;
wire [15:0] _130_;
wire _131_;
wire [15:0] _132_;
wire [16:0] _133_;
wire [16:0] _134_;
wire [16:0] _135_;
wire [16:0] _136_;
wire _137_;
wire [16:0] _138_;
wire [17:0] _139_;
wire [17:0] _140_;
wire [17:0] _141_;
wire [17:0] _142_;
wire _143_;
wire [16:0] _144_;
wire [17:0] _145_;
wire [18:0] _146_;
wire [1:0] _147_;
wire [1:0] _148_;
wire _149_;
wire _150_;
wire [1:0] _151_;
wire [2:0] _152_;
wire [22:0] _153_;
wire [22:0] _154_;
wire _155_;
wire [21:0] _156_;
wire [22:0] _157_;
wire [23:0] _158_;
wire [22:0] _159_;
wire [22:0] _160_;
wire _161_;
wire [22:0] _162_;
wire [23:0] _163_;
wire [23:0] _164_;
wire [4:0] _165_;
wire [4:0] _166_;
wire _167_;
wire [3:0] _168_;
wire [4:0] _169_;
wire [5:0] _170_;
wire [3:0] _171_;
wire [3:0] _172_;
wire [3:0] _173_;
wire [3:0] _174_;
wire [3:0] _175_;
wire [3:0] _176_;
wire [15:0] _177_;
wire [15:0] _178_;
wire [15:0] _179_;
wire [15:0] _180_;
wire [15:0] _181_;
wire [15:0] _182_;
wire [3:0] _183_;
wire [15:0] _184_;
wire [3:0] _185_;
wire [15:0] _186_;
wire [3:0] _187_;
wire [15:0] _188_;
wire [3:0] _189_;
wire [15:0] _190_;
wire [3:0] _191_;
wire [15:0] _192_;
wire [3:0] _193_;
wire [15:0] _194_;
wire [15:0] _195_;
wire [15:0] _196_;
wire [15:0] _197_;
wire [31:0] _198_;
wire [31:0] _199_;
wire [31:0] _200_;
wire [31:0] _201_;
wire [31:0] _202_;
wire [31:0] _203_;
wire [31:0] _204_;
wire [31:0] _205_;
wire [31:0] _206_;
wire [31:0] _207_;
wire [31:0] _208_;
wire [31:0] _209_;
wire [31:0] _210_;
wire [31:0] _211_;
wire [31:0] _212_;
wire [31:0] _213_;
wire [31:0] _214_;
wire [31:0] _215_;
wire [31:0] _216_;
wire [31:0] _217_;
wire [31:0] _218_;
wire [31:0] _219_;
wire [31:0] _220_;
wire [31:0] _221_;
wire [31:0] _222_;
wire [31:0] _223_;
wire [31:0] _224_;
wire [31:0] _225_;
wire [31:0] _226_;
wire [31:0] _227_;
wire [3:0] _228_;
wire [3:0] _229_;
wire [3:0] _230_;
wire [3:0] _231_;
wire [3:0] _232_;
wire [3:0] _233_;
wire [15:0] _234_;
wire [15:0] _235_;
wire [15:0] _236_;
wire [15:0] _237_;
wire [15:0] _238_;
wire [15:0] _239_;
wire [3:0] _240_;
wire [15:0] _241_;
wire [3:0] _242_;
wire [15:0] _243_;
wire [3:0] _244_;
wire [15:0] _245_;
wire [3:0] _246_;
wire [15:0] _247_;
wire [3:0] _248_;
wire [15:0] _249_;
wire [3:0] _250_;
wire [15:0] _251_;
wire [15:0] _252_;
wire [15:0] _253_;
wire [15:0] _254_;
wire [31:0] _255_;
wire [31:0] _256_;
wire [31:0] _257_;
wire [31:0] _258_;
wire [31:0] _259_;
wire [31:0] _260_;
wire [31:0] _261_;
wire [31:0] _262_;
wire [31:0] _263_;
wire [31:0] _264_;
wire [31:0] _265_;
wire [31:0] _266_;
wire [31:0] _267_;
wire [31:0] _268_;
wire [31:0] _269_;
wire [31:0] _270_;
wire [31:0] _271_;
wire [31:0] _272_;
wire [31:0] _273_;
wire [31:0] _274_;
wire [31:0] _275_;
wire [31:0] _276_;
wire [31:0] _277_;
wire [31:0] _278_;
wire [31:0] _279_;
wire [31:0] _280_;
wire [31:0] _281_;
wire [31:0] _282_;
wire [31:0] _283_;
wire [31:0] _284_;
wire [1:0] _285_;
wire [1:0] _286_;
wire _287_;
wire [1:0] _288_;
wire [2:0] _289_;
wire [2:0] _290_;
wire [4:0] _291_;
wire [4:0] _292_;
wire _293_;
wire [3:0] _294_;
wire [4:0] _295_;
wire [5:0] _296_;
wire _297_;
wire _298_;
wire _299_;
wire _300_;
wire _301_;
wire _302_;
wire _303_;
wire _304_;
wire _305_;
wire _306_;
wire _307_;
wire _308_;
wire _309_;
wire _310_;
wire _311_;
wire _312_;
wire _313_;
wire _314_;
wire _315_;
wire _316_;
wire _317_;
wire _318_;
wire _319_;
wire _320_;
wire _321_;
wire _322_;
wire _323_;
wire _324_;
wire _325_;
wire _326_;
wire _327_;
wire _328_;
wire _329_;
wire _330_;
wire _331_;
wire _332_;
wire _333_;
wire _334_;
wire \add_10ns_10s_10_2_1_U4.ce ;
wire \add_10ns_10s_10_2_1_U4.clk ;
wire [9:0] \add_10ns_10s_10_2_1_U4.din0 ;
wire [9:0] \add_10ns_10s_10_2_1_U4.din1 ;
wire [9:0] \add_10ns_10s_10_2_1_U4.dout ;
wire \add_10ns_10s_10_2_1_U4.reset ;
wire [9:0] \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.a ;
wire [9:0] \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.ain_s0 ;
wire [9:0] \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.b ;
wire [9:0] \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.bin_s0 ;
wire \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.ce ;
wire \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.clk ;
wire \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.facout_s1 ;
wire \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.facout_s2 ;
wire [4:0] \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.fas_s1 ;
wire [4:0] \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.fas_s2 ;
wire \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.reset ;
wire [9:0] \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.s ;
wire [4:0] \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.u1.a ;
wire [4:0] \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.u1.b ;
wire \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.u1.cin ;
wire \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.u1.cout ;
wire [4:0] \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.u1.s ;
wire [4:0] \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.u2.a ;
wire [4:0] \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.u2.b ;
wire \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.u2.cin ;
wire \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.u2.cout ;
wire [4:0] \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.u2.s ;
wire \add_10s_10ns_10_2_1_U3.ce ;
wire \add_10s_10ns_10_2_1_U3.clk ;
wire [9:0] \add_10s_10ns_10_2_1_U3.din0 ;
wire [9:0] \add_10s_10ns_10_2_1_U3.din1 ;
wire [9:0] \add_10s_10ns_10_2_1_U3.dout ;
wire \add_10s_10ns_10_2_1_U3.reset ;
wire [9:0] \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.a ;
wire [9:0] \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.ain_s0 ;
wire [9:0] \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.b ;
wire [9:0] \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.bin_s0 ;
wire \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.ce ;
wire \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.clk ;
wire \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.facout_s1 ;
wire \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.facout_s2 ;
wire [4:0] \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.fas_s1 ;
wire [4:0] \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.fas_s2 ;
wire \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.reset ;
wire [9:0] \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.s ;
wire [4:0] \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.u1.a ;
wire [4:0] \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.u1.b ;
wire \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.u1.cin ;
wire \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.u1.cout ;
wire [4:0] \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.u1.s ;
wire [4:0] \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.u2.a ;
wire [4:0] \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.u2.b ;
wire \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.u2.cin ;
wire \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.u2.cout ;
wire [4:0] \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.u2.s ;
wire \add_12ns_12s_12_2_1_U2.ce ;
wire \add_12ns_12s_12_2_1_U2.clk ;
wire [11:0] \add_12ns_12s_12_2_1_U2.din0 ;
wire [11:0] \add_12ns_12s_12_2_1_U2.din1 ;
wire [11:0] \add_12ns_12s_12_2_1_U2.dout ;
wire \add_12ns_12s_12_2_1_U2.reset ;
wire [11:0] \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.a ;
wire [11:0] \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.ain_s0 ;
wire [11:0] \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.b ;
wire [11:0] \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.bin_s0 ;
wire \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.ce ;
wire \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.clk ;
wire \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.facout_s1 ;
wire \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.facout_s2 ;
wire [5:0] \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.fas_s1 ;
wire [5:0] \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.fas_s2 ;
wire \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.reset ;
wire [11:0] \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.s ;
wire [5:0] \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.u1.a ;
wire [5:0] \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.u1.b ;
wire \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.u1.cin ;
wire \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.u1.cout ;
wire [5:0] \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.u1.s ;
wire [5:0] \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.u2.a ;
wire [5:0] \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.u2.b ;
wire \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.u2.cin ;
wire \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.u2.cout ;
wire [5:0] \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.u2.s ;
wire \add_17s_17s_17_2_1_U22.ce ;
wire \add_17s_17s_17_2_1_U22.clk ;
wire [16:0] \add_17s_17s_17_2_1_U22.din0 ;
wire [16:0] \add_17s_17s_17_2_1_U22.din1 ;
wire [16:0] \add_17s_17s_17_2_1_U22.dout ;
wire \add_17s_17s_17_2_1_U22.reset ;
wire [16:0] \add_17s_17s_17_2_1_U22.top_add_17s_17s_17_2_1_Adder_13_U.a ;
wire [16:0] \add_17s_17s_17_2_1_U22.top_add_17s_17s_17_2_1_Adder_13_U.ain_s0 ;
wire [16:0] \add_17s_17s_17_2_1_U22.top_add_17s_17s_17_2_1_Adder_13_U.b ;
wire [16:0] \add_17s_17s_17_2_1_U22.top_add_17s_17s_17_2_1_Adder_13_U.bin_s0 ;
wire \add_17s_17s_17_2_1_U22.top_add_17s_17s_17_2_1_Adder_13_U.ce ;
wire \add_17s_17s_17_2_1_U22.top_add_17s_17s_17_2_1_Adder_13_U.clk ;
wire \add_17s_17s_17_2_1_U22.top_add_17s_17s_17_2_1_Adder_13_U.facout_s1 ;
wire \add_17s_17s_17_2_1_U22.top_add_17s_17s_17_2_1_Adder_13_U.facout_s2 ;
wire [7:0] \add_17s_17s_17_2_1_U22.top_add_17s_17s_17_2_1_Adder_13_U.fas_s1 ;
wire [8:0] \add_17s_17s_17_2_1_U22.top_add_17s_17s_17_2_1_Adder_13_U.fas_s2 ;
wire \add_17s_17s_17_2_1_U22.top_add_17s_17s_17_2_1_Adder_13_U.reset ;
wire [16:0] \add_17s_17s_17_2_1_U22.top_add_17s_17s_17_2_1_Adder_13_U.s ;
wire [7:0] \add_17s_17s_17_2_1_U22.top_add_17s_17s_17_2_1_Adder_13_U.u1.a ;
wire [7:0] \add_17s_17s_17_2_1_U22.top_add_17s_17s_17_2_1_Adder_13_U.u1.b ;
wire \add_17s_17s_17_2_1_U22.top_add_17s_17s_17_2_1_Adder_13_U.u1.cin ;
wire \add_17s_17s_17_2_1_U22.top_add_17s_17s_17_2_1_Adder_13_U.u1.cout ;
wire [7:0] \add_17s_17s_17_2_1_U22.top_add_17s_17s_17_2_1_Adder_13_U.u1.s ;
wire [8:0] \add_17s_17s_17_2_1_U22.top_add_17s_17s_17_2_1_Adder_13_U.u2.a ;
wire [8:0] \add_17s_17s_17_2_1_U22.top_add_17s_17s_17_2_1_Adder_13_U.u2.b ;
wire \add_17s_17s_17_2_1_U22.top_add_17s_17s_17_2_1_Adder_13_U.u2.cin ;
wire \add_17s_17s_17_2_1_U22.top_add_17s_17s_17_2_1_Adder_13_U.u2.cout ;
wire [8:0] \add_17s_17s_17_2_1_U22.top_add_17s_17s_17_2_1_Adder_13_U.u2.s ;
wire \add_2ns_2ns_2_2_1_U17.ce ;
wire \add_2ns_2ns_2_2_1_U17.clk ;
wire [1:0] \add_2ns_2ns_2_2_1_U17.din0 ;
wire [1:0] \add_2ns_2ns_2_2_1_U17.din1 ;
wire [1:0] \add_2ns_2ns_2_2_1_U17.dout ;
wire \add_2ns_2ns_2_2_1_U17.reset ;
wire [1:0] \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_10_U.a ;
wire [1:0] \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_10_U.ain_s0 ;
wire [1:0] \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_10_U.b ;
wire [1:0] \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_10_U.bin_s0 ;
wire \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_10_U.ce ;
wire \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_10_U.clk ;
wire \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_10_U.facout_s1 ;
wire \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_10_U.facout_s2 ;
wire \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_10_U.fas_s1 ;
wire \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_10_U.fas_s2 ;
wire \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_10_U.reset ;
wire [1:0] \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_10_U.s ;
wire \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_10_U.u1.a ;
wire \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_10_U.u1.b ;
wire \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_10_U.u1.cin ;
wire \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_10_U.u1.cout ;
wire \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_10_U.u1.s ;
wire \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_10_U.u2.a ;
wire \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_10_U.u2.b ;
wire \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_10_U.u2.cin ;
wire \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_10_U.u2.cout ;
wire \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_10_U.u2.s ;
wire \add_32ns_32ns_32_2_1_U12.ce ;
wire \add_32ns_32ns_32_2_1_U12.clk ;
wire [31:0] \add_32ns_32ns_32_2_1_U12.din0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U12.din1 ;
wire [31:0] \add_32ns_32ns_32_2_1_U12.dout ;
wire \add_32ns_32ns_32_2_1_U12.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.a ;
wire [31:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.ain_s0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.b ;
wire [31:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.bin_s0 ;
wire \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.ce ;
wire \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.clk ;
wire \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.facout_s1 ;
wire \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.facout_s2 ;
wire [15:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.fas_s1 ;
wire [15:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.fas_s2 ;
wire \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.b ;
wire \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.cin ;
wire \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.b ;
wire \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.cin ;
wire \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.s ;
wire \add_32ns_32ns_32_2_1_U16.ce ;
wire \add_32ns_32ns_32_2_1_U16.clk ;
wire [31:0] \add_32ns_32ns_32_2_1_U16.din0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U16.din1 ;
wire [31:0] \add_32ns_32ns_32_2_1_U16.dout ;
wire \add_32ns_32ns_32_2_1_U16.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_5_U.a ;
wire [31:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_5_U.ain_s0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_5_U.b ;
wire [31:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_5_U.bin_s0 ;
wire \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_5_U.ce ;
wire \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_5_U.clk ;
wire \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_5_U.facout_s1 ;
wire \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_5_U.facout_s2 ;
wire [15:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_5_U.fas_s1 ;
wire [15:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_5_U.fas_s2 ;
wire \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_5_U.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_5_U.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.b ;
wire \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.cin ;
wire \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.b ;
wire \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.cin ;
wire \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.s ;
wire \add_32ns_32ns_32_2_1_U19.ce ;
wire \add_32ns_32ns_32_2_1_U19.clk ;
wire [31:0] \add_32ns_32ns_32_2_1_U19.din0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U19.din1 ;
wire [31:0] \add_32ns_32ns_32_2_1_U19.dout ;
wire \add_32ns_32ns_32_2_1_U19.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_5_U.a ;
wire [31:0] \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_5_U.ain_s0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_5_U.b ;
wire [31:0] \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_5_U.bin_s0 ;
wire \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_5_U.ce ;
wire \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_5_U.clk ;
wire \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_5_U.facout_s1 ;
wire \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_5_U.facout_s2 ;
wire [15:0] \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_5_U.fas_s1 ;
wire [15:0] \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_5_U.fas_s2 ;
wire \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_5_U.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_5_U.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.b ;
wire \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.cin ;
wire \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.b ;
wire \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.cin ;
wire \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.s ;
wire \add_32ns_32ns_32_2_1_U21.ce ;
wire \add_32ns_32ns_32_2_1_U21.clk ;
wire [31:0] \add_32ns_32ns_32_2_1_U21.din0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U21.din1 ;
wire [31:0] \add_32ns_32ns_32_2_1_U21.dout ;
wire \add_32ns_32ns_32_2_1_U21.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_5_U.a ;
wire [31:0] \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_5_U.ain_s0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_5_U.b ;
wire [31:0] \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_5_U.bin_s0 ;
wire \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_5_U.ce ;
wire \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_5_U.clk ;
wire \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_5_U.facout_s1 ;
wire \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_5_U.facout_s2 ;
wire [15:0] \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_5_U.fas_s1 ;
wire [15:0] \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_5_U.fas_s2 ;
wire \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_5_U.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_5_U.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.b ;
wire \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.cin ;
wire \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.b ;
wire \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.cin ;
wire \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.s ;
wire \add_32ns_32ns_32_2_1_U6.ce ;
wire \add_32ns_32ns_32_2_1_U6.clk ;
wire [31:0] \add_32ns_32ns_32_2_1_U6.din0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U6.din1 ;
wire [31:0] \add_32ns_32ns_32_2_1_U6.dout ;
wire \add_32ns_32ns_32_2_1_U6.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.a ;
wire [31:0] \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.ain_s0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.b ;
wire [31:0] \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.bin_s0 ;
wire \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.ce ;
wire \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.clk ;
wire \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.facout_s1 ;
wire \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.facout_s2 ;
wire [15:0] \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.fas_s1 ;
wire [15:0] \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.fas_s2 ;
wire \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.b ;
wire \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.cin ;
wire \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.b ;
wire \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.cin ;
wire \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.s ;
wire \add_32s_32ns_32_2_1_U23.ce ;
wire \add_32s_32ns_32_2_1_U23.clk ;
wire [31:0] \add_32s_32ns_32_2_1_U23.din0 ;
wire [31:0] \add_32s_32ns_32_2_1_U23.din1 ;
wire [31:0] \add_32s_32ns_32_2_1_U23.dout ;
wire \add_32s_32ns_32_2_1_U23.reset ;
wire [31:0] \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_14_U.a ;
wire [31:0] \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_14_U.ain_s0 ;
wire [31:0] \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_14_U.b ;
wire [31:0] \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_14_U.bin_s0 ;
wire \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_14_U.ce ;
wire \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_14_U.clk ;
wire \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_14_U.facout_s1 ;
wire \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_14_U.facout_s2 ;
wire [15:0] \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_14_U.fas_s1 ;
wire [15:0] \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_14_U.fas_s2 ;
wire \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_14_U.reset ;
wire [31:0] \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_14_U.s ;
wire [15:0] \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_14_U.u1.a ;
wire [15:0] \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_14_U.u1.b ;
wire \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_14_U.u1.cin ;
wire \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_14_U.u1.cout ;
wire [15:0] \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_14_U.u1.s ;
wire [15:0] \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_14_U.u2.a ;
wire [15:0] \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_14_U.u2.b ;
wire \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_14_U.u2.cin ;
wire \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_14_U.u2.cout ;
wire [15:0] \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_14_U.u2.s ;
wire \add_34s_34s_34_2_1_U18.ce ;
wire \add_34s_34s_34_2_1_U18.clk ;
wire [33:0] \add_34s_34s_34_2_1_U18.din0 ;
wire [33:0] \add_34s_34s_34_2_1_U18.din1 ;
wire [33:0] \add_34s_34s_34_2_1_U18.dout ;
wire \add_34s_34s_34_2_1_U18.reset ;
wire [33:0] \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.a ;
wire [33:0] \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.ain_s0 ;
wire [33:0] \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.b ;
wire [33:0] \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.bin_s0 ;
wire \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.ce ;
wire \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.clk ;
wire \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.facout_s1 ;
wire \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.facout_s2 ;
wire [16:0] \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.fas_s1 ;
wire [16:0] \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.fas_s2 ;
wire \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.reset ;
wire [33:0] \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.s ;
wire [16:0] \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.u1.a ;
wire [16:0] \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.u1.b ;
wire \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.u1.cin ;
wire \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.u1.cout ;
wire [16:0] \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.u1.s ;
wire [16:0] \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.u2.a ;
wire [16:0] \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.u2.b ;
wire \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.u2.cin ;
wire \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.u2.cout ;
wire [16:0] \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.u2.s ;
wire \add_35s_35s_35_2_1_U15.ce ;
wire \add_35s_35s_35_2_1_U15.clk ;
wire [34:0] \add_35s_35s_35_2_1_U15.din0 ;
wire [34:0] \add_35s_35s_35_2_1_U15.din1 ;
wire [34:0] \add_35s_35s_35_2_1_U15.dout ;
wire \add_35s_35s_35_2_1_U15.reset ;
wire [34:0] \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.a ;
wire [34:0] \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.ain_s0 ;
wire [34:0] \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.b ;
wire [34:0] \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.bin_s0 ;
wire \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.ce ;
wire \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.clk ;
wire \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.facout_s1 ;
wire \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.facout_s2 ;
wire [16:0] \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.fas_s1 ;
wire [17:0] \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.fas_s2 ;
wire \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.reset ;
wire [34:0] \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.s ;
wire [16:0] \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.u1.a ;
wire [16:0] \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.u1.b ;
wire \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.u1.cin ;
wire \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.u1.cout ;
wire [16:0] \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.u1.s ;
wire [17:0] \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.u2.a ;
wire [17:0] \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.u2.b ;
wire \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.u2.cin ;
wire \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.u2.cout ;
wire [17:0] \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.u2.s ;
wire \add_3s_3ns_3_2_1_U20.ce ;
wire \add_3s_3ns_3_2_1_U20.clk ;
wire [2:0] \add_3s_3ns_3_2_1_U20.din0 ;
wire [2:0] \add_3s_3ns_3_2_1_U20.din1 ;
wire [2:0] \add_3s_3ns_3_2_1_U20.dout ;
wire \add_3s_3ns_3_2_1_U20.reset ;
wire [2:0] \add_3s_3ns_3_2_1_U20.top_add_3s_3ns_3_2_1_Adder_12_U.a ;
wire [2:0] \add_3s_3ns_3_2_1_U20.top_add_3s_3ns_3_2_1_Adder_12_U.ain_s0 ;
wire [2:0] \add_3s_3ns_3_2_1_U20.top_add_3s_3ns_3_2_1_Adder_12_U.b ;
wire [2:0] \add_3s_3ns_3_2_1_U20.top_add_3s_3ns_3_2_1_Adder_12_U.bin_s0 ;
wire \add_3s_3ns_3_2_1_U20.top_add_3s_3ns_3_2_1_Adder_12_U.ce ;
wire \add_3s_3ns_3_2_1_U20.top_add_3s_3ns_3_2_1_Adder_12_U.clk ;
wire \add_3s_3ns_3_2_1_U20.top_add_3s_3ns_3_2_1_Adder_12_U.facout_s1 ;
wire \add_3s_3ns_3_2_1_U20.top_add_3s_3ns_3_2_1_Adder_12_U.facout_s2 ;
wire \add_3s_3ns_3_2_1_U20.top_add_3s_3ns_3_2_1_Adder_12_U.fas_s1 ;
wire [1:0] \add_3s_3ns_3_2_1_U20.top_add_3s_3ns_3_2_1_Adder_12_U.fas_s2 ;
wire \add_3s_3ns_3_2_1_U20.top_add_3s_3ns_3_2_1_Adder_12_U.reset ;
wire [2:0] \add_3s_3ns_3_2_1_U20.top_add_3s_3ns_3_2_1_Adder_12_U.s ;
wire \add_3s_3ns_3_2_1_U20.top_add_3s_3ns_3_2_1_Adder_12_U.u1.a ;
wire \add_3s_3ns_3_2_1_U20.top_add_3s_3ns_3_2_1_Adder_12_U.u1.b ;
wire \add_3s_3ns_3_2_1_U20.top_add_3s_3ns_3_2_1_Adder_12_U.u1.cin ;
wire \add_3s_3ns_3_2_1_U20.top_add_3s_3ns_3_2_1_Adder_12_U.u1.cout ;
wire \add_3s_3ns_3_2_1_U20.top_add_3s_3ns_3_2_1_Adder_12_U.u1.s ;
wire [1:0] \add_3s_3ns_3_2_1_U20.top_add_3s_3ns_3_2_1_Adder_12_U.u2.a ;
wire [1:0] \add_3s_3ns_3_2_1_U20.top_add_3s_3ns_3_2_1_Adder_12_U.u2.b ;
wire \add_3s_3ns_3_2_1_U20.top_add_3s_3ns_3_2_1_Adder_12_U.u2.cin ;
wire \add_3s_3ns_3_2_1_U20.top_add_3s_3ns_3_2_1_Adder_12_U.u2.cout ;
wire [1:0] \add_3s_3ns_3_2_1_U20.top_add_3s_3ns_3_2_1_Adder_12_U.u2.s ;
wire \add_45s_45s_45_2_1_U8.ce ;
wire \add_45s_45s_45_2_1_U8.clk ;
wire [44:0] \add_45s_45s_45_2_1_U8.din0 ;
wire [44:0] \add_45s_45s_45_2_1_U8.din1 ;
wire [44:0] \add_45s_45s_45_2_1_U8.dout ;
wire \add_45s_45s_45_2_1_U8.reset ;
wire [44:0] \add_45s_45s_45_2_1_U8.top_add_45s_45s_45_2_1_Adder_7_U.a ;
wire [44:0] \add_45s_45s_45_2_1_U8.top_add_45s_45s_45_2_1_Adder_7_U.ain_s0 ;
wire [44:0] \add_45s_45s_45_2_1_U8.top_add_45s_45s_45_2_1_Adder_7_U.b ;
wire [44:0] \add_45s_45s_45_2_1_U8.top_add_45s_45s_45_2_1_Adder_7_U.bin_s0 ;
wire \add_45s_45s_45_2_1_U8.top_add_45s_45s_45_2_1_Adder_7_U.ce ;
wire \add_45s_45s_45_2_1_U8.top_add_45s_45s_45_2_1_Adder_7_U.clk ;
wire \add_45s_45s_45_2_1_U8.top_add_45s_45s_45_2_1_Adder_7_U.facout_s1 ;
wire \add_45s_45s_45_2_1_U8.top_add_45s_45s_45_2_1_Adder_7_U.facout_s2 ;
wire [21:0] \add_45s_45s_45_2_1_U8.top_add_45s_45s_45_2_1_Adder_7_U.fas_s1 ;
wire [22:0] \add_45s_45s_45_2_1_U8.top_add_45s_45s_45_2_1_Adder_7_U.fas_s2 ;
wire \add_45s_45s_45_2_1_U8.top_add_45s_45s_45_2_1_Adder_7_U.reset ;
wire [44:0] \add_45s_45s_45_2_1_U8.top_add_45s_45s_45_2_1_Adder_7_U.s ;
wire [21:0] \add_45s_45s_45_2_1_U8.top_add_45s_45s_45_2_1_Adder_7_U.u1.a ;
wire [21:0] \add_45s_45s_45_2_1_U8.top_add_45s_45s_45_2_1_Adder_7_U.u1.b ;
wire \add_45s_45s_45_2_1_U8.top_add_45s_45s_45_2_1_Adder_7_U.u1.cin ;
wire \add_45s_45s_45_2_1_U8.top_add_45s_45s_45_2_1_Adder_7_U.u1.cout ;
wire [21:0] \add_45s_45s_45_2_1_U8.top_add_45s_45s_45_2_1_Adder_7_U.u1.s ;
wire [22:0] \add_45s_45s_45_2_1_U8.top_add_45s_45s_45_2_1_Adder_7_U.u2.a ;
wire [22:0] \add_45s_45s_45_2_1_U8.top_add_45s_45s_45_2_1_Adder_7_U.u2.b ;
wire \add_45s_45s_45_2_1_U8.top_add_45s_45s_45_2_1_Adder_7_U.u2.cin ;
wire \add_45s_45s_45_2_1_U8.top_add_45s_45s_45_2_1_Adder_7_U.u2.cout ;
wire [22:0] \add_45s_45s_45_2_1_U8.top_add_45s_45s_45_2_1_Adder_7_U.u2.s ;
wire \add_46s_46s_46_2_1_U5.ce ;
wire \add_46s_46s_46_2_1_U5.clk ;
wire [45:0] \add_46s_46s_46_2_1_U5.din0 ;
wire [45:0] \add_46s_46s_46_2_1_U5.din1 ;
wire [45:0] \add_46s_46s_46_2_1_U5.dout ;
wire \add_46s_46s_46_2_1_U5.reset ;
wire [45:0] \add_46s_46s_46_2_1_U5.top_add_46s_46s_46_2_1_Adder_4_U.a ;
wire [45:0] \add_46s_46s_46_2_1_U5.top_add_46s_46s_46_2_1_Adder_4_U.ain_s0 ;
wire [45:0] \add_46s_46s_46_2_1_U5.top_add_46s_46s_46_2_1_Adder_4_U.b ;
wire [45:0] \add_46s_46s_46_2_1_U5.top_add_46s_46s_46_2_1_Adder_4_U.bin_s0 ;
wire \add_46s_46s_46_2_1_U5.top_add_46s_46s_46_2_1_Adder_4_U.ce ;
wire \add_46s_46s_46_2_1_U5.top_add_46s_46s_46_2_1_Adder_4_U.clk ;
wire \add_46s_46s_46_2_1_U5.top_add_46s_46s_46_2_1_Adder_4_U.facout_s1 ;
wire \add_46s_46s_46_2_1_U5.top_add_46s_46s_46_2_1_Adder_4_U.facout_s2 ;
wire [22:0] \add_46s_46s_46_2_1_U5.top_add_46s_46s_46_2_1_Adder_4_U.fas_s1 ;
wire [22:0] \add_46s_46s_46_2_1_U5.top_add_46s_46s_46_2_1_Adder_4_U.fas_s2 ;
wire \add_46s_46s_46_2_1_U5.top_add_46s_46s_46_2_1_Adder_4_U.reset ;
wire [45:0] \add_46s_46s_46_2_1_U5.top_add_46s_46s_46_2_1_Adder_4_U.s ;
wire [22:0] \add_46s_46s_46_2_1_U5.top_add_46s_46s_46_2_1_Adder_4_U.u1.a ;
wire [22:0] \add_46s_46s_46_2_1_U5.top_add_46s_46s_46_2_1_Adder_4_U.u1.b ;
wire \add_46s_46s_46_2_1_U5.top_add_46s_46s_46_2_1_Adder_4_U.u1.cin ;
wire \add_46s_46s_46_2_1_U5.top_add_46s_46s_46_2_1_Adder_4_U.u1.cout ;
wire [22:0] \add_46s_46s_46_2_1_U5.top_add_46s_46s_46_2_1_Adder_4_U.u1.s ;
wire [22:0] \add_46s_46s_46_2_1_U5.top_add_46s_46s_46_2_1_Adder_4_U.u2.a ;
wire [22:0] \add_46s_46s_46_2_1_U5.top_add_46s_46s_46_2_1_Adder_4_U.u2.b ;
wire \add_46s_46s_46_2_1_U5.top_add_46s_46s_46_2_1_Adder_4_U.u2.cin ;
wire \add_46s_46s_46_2_1_U5.top_add_46s_46s_46_2_1_Adder_4_U.u2.cout ;
wire [22:0] \add_46s_46s_46_2_1_U5.top_add_46s_46s_46_2_1_Adder_4_U.u2.s ;
wire \add_9s_9s_9_2_1_U1.ce ;
wire \add_9s_9s_9_2_1_U1.clk ;
wire [8:0] \add_9s_9s_9_2_1_U1.din0 ;
wire [8:0] \add_9s_9s_9_2_1_U1.din1 ;
wire [8:0] \add_9s_9s_9_2_1_U1.dout ;
wire \add_9s_9s_9_2_1_U1.reset ;
wire [8:0] \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.a ;
wire [8:0] \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.ain_s0 ;
wire [8:0] \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.b ;
wire [8:0] \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.bin_s0 ;
wire \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.ce ;
wire \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.clk ;
wire \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.facout_s1 ;
wire \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.facout_s2 ;
wire [3:0] \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.fas_s1 ;
wire [4:0] \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.fas_s2 ;
wire \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.reset ;
wire [8:0] \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.s ;
wire [3:0] \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.u1.a ;
wire [3:0] \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.u1.b ;
wire \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.u1.cin ;
wire \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.u1.cout ;
wire [3:0] \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.u1.s ;
wire [4:0] \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.u2.a ;
wire [4:0] \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.u2.b ;
wire \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.u2.cin ;
wire \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.u2.cout ;
wire [4:0] \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.u2.s ;
wire and_ln353_fu_565_p2;
wire ap_CS_fsm_state1;
wire ap_CS_fsm_state10;
wire ap_CS_fsm_state11;
wire ap_CS_fsm_state12;
wire ap_CS_fsm_state13;
wire ap_CS_fsm_state14;
wire ap_CS_fsm_state15;
wire ap_CS_fsm_state16;
wire ap_CS_fsm_state17;
wire ap_CS_fsm_state18;
wire ap_CS_fsm_state19;
wire ap_CS_fsm_state2;
wire ap_CS_fsm_state20;
wire ap_CS_fsm_state21;
wire ap_CS_fsm_state22;
wire ap_CS_fsm_state23;
wire ap_CS_fsm_state24;
wire ap_CS_fsm_state25;
wire ap_CS_fsm_state26;
wire ap_CS_fsm_state27;
wire ap_CS_fsm_state28;
wire ap_CS_fsm_state29;
wire ap_CS_fsm_state3;
wire ap_CS_fsm_state30;
wire ap_CS_fsm_state31;
wire ap_CS_fsm_state32;
wire ap_CS_fsm_state33;
wire ap_CS_fsm_state4;
wire ap_CS_fsm_state5;
wire ap_CS_fsm_state6;
wire ap_CS_fsm_state7;
wire ap_CS_fsm_state8;
wire ap_CS_fsm_state9;
wire [32:0] ap_NS_fsm;
wire ap_clk;
wire ap_done;
wire ap_idle;
wire ap_ready;
wire ap_rst;
wire ap_start;
wire \ashr_16ns_4ns_16_7_1_U14.ce ;
wire \ashr_16ns_4ns_16_7_1_U14.clk ;
wire [15:0] \ashr_16ns_4ns_16_7_1_U14.din0 ;
wire [15:0] \ashr_16ns_4ns_16_7_1_U14.din1 ;
wire [3:0] \ashr_16ns_4ns_16_7_1_U14.din1_cast ;
wire [3:0] \ashr_16ns_4ns_16_7_1_U14.din1_mask ;
wire [15:0] \ashr_16ns_4ns_16_7_1_U14.dout ;
wire \ashr_16ns_4ns_16_7_1_U14.reset ;
wire \ashr_32s_32s_32_7_1_U10.ce ;
wire \ashr_32s_32s_32_7_1_U10.clk ;
wire [31:0] \ashr_32s_32s_32_7_1_U10.din0 ;
wire [31:0] \ashr_32s_32s_32_7_1_U10.din1 ;
wire [31:0] \ashr_32s_32s_32_7_1_U10.din1_cast ;
wire [31:0] \ashr_32s_32s_32_7_1_U10.din1_mask ;
wire [31:0] \ashr_32s_32s_32_7_1_U10.dout ;
wire \ashr_32s_32s_32_7_1_U10.reset ;
wire [7:0] conv_i_i_i357_fu_509_p0;
wire [31:0] conv_i_i_i357_fu_509_p1;
wire [8:0] grp_fu_243_p0;
wire [8:0] grp_fu_243_p1;
wire [8:0] grp_fu_243_p2;
wire [11:0] grp_fu_260_p0;
wire [11:0] grp_fu_260_p1;
wire [11:0] grp_fu_260_p2;
wire [9:0] grp_fu_289_p0;
wire [9:0] grp_fu_289_p2;
wire [9:0] grp_fu_331_p1;
wire [9:0] grp_fu_331_p2;
wire [45:0] grp_fu_351_p0;
wire [45:0] grp_fu_351_p1;
wire [45:0] grp_fu_351_p2;
wire [31:0] grp_fu_377_p2;
wire [8:0] grp_fu_399_p1;
wire [8:0] grp_fu_399_p2;
wire [44:0] grp_fu_439_p0;
wire [44:0] grp_fu_439_p1;
wire [44:0] grp_fu_439_p2;
wire [3:0] grp_fu_478_p2;
wire [31:0] grp_fu_513_p2;
wire [31:0] grp_fu_519_p2;
wire [31:0] grp_fu_525_p2;
wire [15:0] grp_fu_538_p1;
wire [15:0] grp_fu_538_p2;
wire [15:0] grp_fu_546_p1;
wire [15:0] grp_fu_546_p2;
wire [34:0] grp_fu_618_p0;
wire [34:0] grp_fu_618_p1;
wire [34:0] grp_fu_618_p2;
wire [31:0] grp_fu_644_p2;
wire [1:0] grp_fu_692_p2;
wire [33:0] grp_fu_712_p0;
wire [33:0] grp_fu_712_p1;
wire [33:0] grp_fu_712_p2;
wire [31:0] grp_fu_752_p2;
wire [2:0] grp_fu_760_p0;
wire [2:0] grp_fu_760_p2;
wire [31:0] grp_fu_791_p2;
wire [16:0] grp_fu_799_p0;
wire [16:0] grp_fu_799_p1;
wire [16:0] grp_fu_799_p2;
wire [31:0] grp_fu_808_p0;
wire [31:0] grp_fu_808_p2;
wire icmp_ln850_fu_530_p2;
wire icmp_ln851_1_fu_270_p2;
wire icmp_ln851_2_fu_361_p2;
wire icmp_ln851_3_fu_449_p2;
wire icmp_ln851_4_fu_628_p2;
wire icmp_ln851_fu_687_p2;
wire [9:0] lhs_fu_484_p3;
wire [3:0] op_0;
wire [3:0] op_10;
wire [3:0] op_11_V_fu_303_p2;
wire [15:0] op_12;
wire [15:0] op_13;
wire [3:0] op_14;
wire [7:0] op_15;
wire [31:0] op_19;
wire [7:0] op_2;
wire [7:0] op_3;
wire [31:0] op_31;
wire op_31_ap_vld;
wire [15:0] op_4;
wire [7:0] op_5;
wire [3:0] op_6;
wire [7:0] op_7;
wire [3:0] op_8;
wire p_Result_1_fu_733_p3;
wire p_Result_2_fu_309_p3;
wire p_Result_3_fu_405_p3;
wire p_Result_4_fu_576_p3;
wire p_Result_5_fu_668_p3;
wire p_Result_6_fu_765_p3;
wire p_Result_s_fu_558_p3;
wire [15:0] r_1_fu_718_p3;
wire [7:0] r_fu_382_p2;
wire [9:0] ret_V_12_fu_496_p2;
wire [9:0] ret_V_12_reg_994;
wire ret_V_13_fu_570_p2;
wire [9:0] ret_V_15_fu_321_p3;
wire [31:0] ret_V_20_fu_781_p3;
wire [1:0] ret_V_4_fu_745_p3;
wire [43:0] rhs_3_fu_428_p3;
wire [33:0] rhs_4_fu_607_p3;
wire [32:0] rhs_5_fu_701_p3;
wire [31:0] select_ln1358_fu_649_p3;
wire [31:0] select_ln353_1_fu_588_p3;
wire [31:0] select_ln353_2_fu_680_p3;
wire [31:0] select_ln353_fu_417_p3;
wire [2:0] select_ln69_fu_595_p3;
wire [9:0] select_ln850_2_fu_316_p3;
wire [31:0] select_ln850_3_fu_412_p3;
wire [31:0] select_ln850_4_fu_583_p3;
wire [31:0] select_ln850_5_fu_675_p3;
wire [31:0] select_ln850_6_fu_775_p3;
wire [1:0] select_ln850_fu_740_p3;
wire [3:0] sext_ln1192_fu_249_p0;
wire [31:0] sext_ln1357_fu_506_p1;
wire [8:0] sext_ln15_fu_396_p1;
wire [15:0] sext_ln703_1_fu_336_p0;
wire [15:0] sext_ln703_2_fu_424_p0;
wire [3:0] sext_ln703_3_fu_603_p0;
wire [7:0] sext_ln703_4_fu_697_p0;
wire [7:0] sext_ln703_fu_492_p0;
wire [9:0] sext_ln703_fu_492_p1;
wire [9:0] sext_ln850_fu_286_p1;
wire \shl_16ns_4ns_16_7_1_U13.ce ;
wire \shl_16ns_4ns_16_7_1_U13.clk ;
wire [15:0] \shl_16ns_4ns_16_7_1_U13.din0 ;
wire [15:0] \shl_16ns_4ns_16_7_1_U13.din1 ;
wire [3:0] \shl_16ns_4ns_16_7_1_U13.din1_cast ;
wire [3:0] \shl_16ns_4ns_16_7_1_U13.din1_mask ;
wire [15:0] \shl_16ns_4ns_16_7_1_U13.dout ;
wire \shl_16ns_4ns_16_7_1_U13.reset ;
wire \shl_32s_32s_32_7_1_U11.ce ;
wire \shl_32s_32s_32_7_1_U11.clk ;
wire [31:0] \shl_32s_32s_32_7_1_U11.din0 ;
wire [31:0] \shl_32s_32s_32_7_1_U11.din1 ;
wire [31:0] \shl_32s_32s_32_7_1_U11.din1_cast ;
wire [31:0] \shl_32s_32s_32_7_1_U11.din1_mask ;
wire [31:0] \shl_32s_32s_32_7_1_U11.dout ;
wire \shl_32s_32s_32_7_1_U11.reset ;
wire \sub_4ns_4ns_4_2_1_U9.ce ;
wire \sub_4ns_4ns_4_2_1_U9.clk ;
wire [3:0] \sub_4ns_4ns_4_2_1_U9.din0 ;
wire [3:0] \sub_4ns_4ns_4_2_1_U9.din1 ;
wire [3:0] \sub_4ns_4ns_4_2_1_U9.dout ;
wire \sub_4ns_4ns_4_2_1_U9.reset ;
wire [3:0] \sub_4ns_4ns_4_2_1_U9.top_sub_4ns_4ns_4_2_1_Adder_8_U.a ;
wire [3:0] \sub_4ns_4ns_4_2_1_U9.top_sub_4ns_4ns_4_2_1_Adder_8_U.ain_s0 ;
wire [3:0] \sub_4ns_4ns_4_2_1_U9.top_sub_4ns_4ns_4_2_1_Adder_8_U.b ;
wire [3:0] \sub_4ns_4ns_4_2_1_U9.top_sub_4ns_4ns_4_2_1_Adder_8_U.bin_s0 ;
wire \sub_4ns_4ns_4_2_1_U9.top_sub_4ns_4ns_4_2_1_Adder_8_U.ce ;
wire \sub_4ns_4ns_4_2_1_U9.top_sub_4ns_4ns_4_2_1_Adder_8_U.clk ;
wire \sub_4ns_4ns_4_2_1_U9.top_sub_4ns_4ns_4_2_1_Adder_8_U.facout_s1 ;
wire \sub_4ns_4ns_4_2_1_U9.top_sub_4ns_4ns_4_2_1_Adder_8_U.facout_s2 ;
wire [1:0] \sub_4ns_4ns_4_2_1_U9.top_sub_4ns_4ns_4_2_1_Adder_8_U.fas_s1 ;
wire [1:0] \sub_4ns_4ns_4_2_1_U9.top_sub_4ns_4ns_4_2_1_Adder_8_U.fas_s2 ;
wire \sub_4ns_4ns_4_2_1_U9.top_sub_4ns_4ns_4_2_1_Adder_8_U.reset ;
wire [3:0] \sub_4ns_4ns_4_2_1_U9.top_sub_4ns_4ns_4_2_1_Adder_8_U.s ;
wire [1:0] \sub_4ns_4ns_4_2_1_U9.top_sub_4ns_4ns_4_2_1_Adder_8_U.u1.a ;
wire [1:0] \sub_4ns_4ns_4_2_1_U9.top_sub_4ns_4ns_4_2_1_Adder_8_U.u1.b ;
wire \sub_4ns_4ns_4_2_1_U9.top_sub_4ns_4ns_4_2_1_Adder_8_U.u1.cin ;
wire \sub_4ns_4ns_4_2_1_U9.top_sub_4ns_4ns_4_2_1_Adder_8_U.u1.cout ;
wire [1:0] \sub_4ns_4ns_4_2_1_U9.top_sub_4ns_4ns_4_2_1_Adder_8_U.u1.s ;
wire [1:0] \sub_4ns_4ns_4_2_1_U9.top_sub_4ns_4ns_4_2_1_Adder_8_U.u2.a ;
wire [1:0] \sub_4ns_4ns_4_2_1_U9.top_sub_4ns_4ns_4_2_1_Adder_8_U.u2.b ;
wire \sub_4ns_4ns_4_2_1_U9.top_sub_4ns_4ns_4_2_1_Adder_8_U.u2.cin ;
wire \sub_4ns_4ns_4_2_1_U9.top_sub_4ns_4ns_4_2_1_Adder_8_U.u2.cout ;
wire [1:0] \sub_4ns_4ns_4_2_1_U9.top_sub_4ns_4ns_4_2_1_Adder_8_U.u2.s ;
wire \sub_9ns_9s_9_2_1_U7.ce ;
wire \sub_9ns_9s_9_2_1_U7.clk ;
wire [8:0] \sub_9ns_9s_9_2_1_U7.din0 ;
wire [8:0] \sub_9ns_9s_9_2_1_U7.din1 ;
wire [8:0] \sub_9ns_9s_9_2_1_U7.dout ;
wire \sub_9ns_9s_9_2_1_U7.reset ;
wire [8:0] \sub_9ns_9s_9_2_1_U7.top_sub_9ns_9s_9_2_1_Adder_6_U.a ;
wire [8:0] \sub_9ns_9s_9_2_1_U7.top_sub_9ns_9s_9_2_1_Adder_6_U.ain_s0 ;
wire [8:0] \sub_9ns_9s_9_2_1_U7.top_sub_9ns_9s_9_2_1_Adder_6_U.b ;
wire [8:0] \sub_9ns_9s_9_2_1_U7.top_sub_9ns_9s_9_2_1_Adder_6_U.bin_s0 ;
wire \sub_9ns_9s_9_2_1_U7.top_sub_9ns_9s_9_2_1_Adder_6_U.ce ;
wire \sub_9ns_9s_9_2_1_U7.top_sub_9ns_9s_9_2_1_Adder_6_U.clk ;
wire \sub_9ns_9s_9_2_1_U7.top_sub_9ns_9s_9_2_1_Adder_6_U.facout_s1 ;
wire \sub_9ns_9s_9_2_1_U7.top_sub_9ns_9s_9_2_1_Adder_6_U.facout_s2 ;
wire [3:0] \sub_9ns_9s_9_2_1_U7.top_sub_9ns_9s_9_2_1_Adder_6_U.fas_s1 ;
wire [4:0] \sub_9ns_9s_9_2_1_U7.top_sub_9ns_9s_9_2_1_Adder_6_U.fas_s2 ;
wire \sub_9ns_9s_9_2_1_U7.top_sub_9ns_9s_9_2_1_Adder_6_U.reset ;
wire [8:0] \sub_9ns_9s_9_2_1_U7.top_sub_9ns_9s_9_2_1_Adder_6_U.s ;
wire [3:0] \sub_9ns_9s_9_2_1_U7.top_sub_9ns_9s_9_2_1_Adder_6_U.u1.a ;
wire [3:0] \sub_9ns_9s_9_2_1_U7.top_sub_9ns_9s_9_2_1_Adder_6_U.u1.b ;
wire \sub_9ns_9s_9_2_1_U7.top_sub_9ns_9s_9_2_1_Adder_6_U.u1.cin ;
wire \sub_9ns_9s_9_2_1_U7.top_sub_9ns_9s_9_2_1_Adder_6_U.u1.cout ;
wire [3:0] \sub_9ns_9s_9_2_1_U7.top_sub_9ns_9s_9_2_1_Adder_6_U.u1.s ;
wire [4:0] \sub_9ns_9s_9_2_1_U7.top_sub_9ns_9s_9_2_1_Adder_6_U.u2.a ;
wire [4:0] \sub_9ns_9s_9_2_1_U7.top_sub_9ns_9s_9_2_1_Adder_6_U.u2.b ;
wire \sub_9ns_9s_9_2_1_U7.top_sub_9ns_9s_9_2_1_Adder_6_U.u2.cin ;
wire \sub_9ns_9s_9_2_1_U7.top_sub_9ns_9s_9_2_1_Adder_6_U.u2.cout ;
wire [4:0] \sub_9ns_9s_9_2_1_U7.top_sub_9ns_9s_9_2_1_Adder_6_U.u2.s ;
wire [22:0] tmp_6_fu_340_p3;
wire tmp_fu_551_p3;
wire [3:0] trunc_ln1350_1_fu_299_p1;
wire [3:0] trunc_ln1350_fu_295_p1;
wire [5:0] trunc_ln851_1_fu_664_p1;
wire [3:0] trunc_ln851_2_fu_266_p0;
wire [2:0] trunc_ln851_2_fu_266_p1;
wire [15:0] trunc_ln851_3_fu_357_p0;
wire [12:0] trunc_ln851_3_fu_357_p1;
wire [15:0] trunc_ln851_4_fu_445_p0;
wire [11:0] trunc_ln851_4_fu_445_p1;
wire [3:0] trunc_ln851_5_fu_624_p0;
wire [1:0] trunc_ln851_5_fu_624_p1;
wire [7:0] trunc_ln851_6_fu_772_p0;
wire trunc_ln851_6_fu_772_p1;
wire [5:0] trunc_ln851_fu_502_p1;
wire [8:0] ush_fu_455_p3;


assign _054_ = ap_CS_fsm[12] & icmp_ln851_2_reg_902;
assign _055_ = ap_CS_fsm[17] & icmp_ln851_3_reg_961;
assign _056_ = icmp_ln851_4_reg_1062 & ap_CS_fsm[22];
assign _057_ = icmp_ln851_1_reg_839 & ap_CS_fsm[5];
assign _058_ = ap_CS_fsm[22] & _065_;
assign _059_ = _066_ & ap_CS_fsm[24];
assign _060_ = ap_CS_fsm[22] & tmp_3_reg_924;
assign _061_ = p_Result_7_reg_989 & ap_CS_fsm[24];
assign _062_ = ap_CS_fsm[14] & _065_;
assign _063_ = _067_ & ap_CS_fsm[0];
assign _064_ = ap_start & ap_CS_fsm[0];
assign and_ln353_fu_565_p2 = ret_V_12_reg_994[9] & icmp_ln850_reg_1022;
assign ret_V_12_fu_496_p2 = { op_7[7], op_7[7], op_7 } & { op_6, 6'h00 };
assign r_fu_382_p2 = ~ op_3;
assign _065_ = ~ tmp_3_reg_924;
assign _066_ = ~ p_Result_7_reg_989;
assign _067_ = ~ ap_start;
assign _068_ = ! trunc_ln851_1_reg_1106;
always @(posedge \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.clk )
\add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.bin_s1  <= _070_;
always @(posedge \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.clk )
\add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.ain_s1  <= _069_;
always @(posedge \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.clk )
\add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.sum_s1  <= _072_;
always @(posedge \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.clk )
\add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.carry_s1  <= _071_;
assign _070_ = \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.ce  ? \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.b [9:5] : \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.bin_s1 ;
assign _069_ = \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.ce  ? \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.a [9:5] : \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.ain_s1 ;
assign _071_ = \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.ce  ? \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.facout_s1  : \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.carry_s1 ;
assign _072_ = \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.ce  ? \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.fas_s1  : \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.sum_s1 ;
assign _073_ = \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.u1.a  + \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.u1.b ;
assign { \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.u1.cout , \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.u1.s  } = _073_ + \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.u1.cin ;
assign _074_ = \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.u2.a  + \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.u2.b ;
assign { \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.u2.cout , \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.u2.s  } = _074_ + \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.u2.cin ;
always @(posedge \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.clk )
\add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.bin_s1  <= _076_;
always @(posedge \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.clk )
\add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.ain_s1  <= _075_;
always @(posedge \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.clk )
\add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.sum_s1  <= _078_;
always @(posedge \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.clk )
\add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.carry_s1  <= _077_;
assign _076_ = \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.ce  ? \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.b [9:5] : \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.bin_s1 ;
assign _075_ = \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.ce  ? \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.a [9:5] : \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.ain_s1 ;
assign _077_ = \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.ce  ? \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.facout_s1  : \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.carry_s1 ;
assign _078_ = \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.ce  ? \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.fas_s1  : \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.sum_s1 ;
assign _079_ = \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.u1.a  + \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.u1.b ;
assign { \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.u1.cout , \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.u1.s  } = _079_ + \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.u1.cin ;
assign _080_ = \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.u2.a  + \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.u2.b ;
assign { \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.u2.cout , \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.u2.s  } = _080_ + \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.u2.cin ;
always @(posedge \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.clk )
\add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.bin_s1  <= _082_;
always @(posedge \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.clk )
\add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.ain_s1  <= _081_;
always @(posedge \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.clk )
\add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.sum_s1  <= _084_;
always @(posedge \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.clk )
\add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.carry_s1  <= _083_;
assign _082_ = \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.ce  ? \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.b [11:6] : \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.bin_s1 ;
assign _081_ = \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.ce  ? \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.a [11:6] : \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.ain_s1 ;
assign _083_ = \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.ce  ? \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.facout_s1  : \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.carry_s1 ;
assign _084_ = \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.ce  ? \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.fas_s1  : \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.sum_s1 ;
assign _085_ = \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.u1.a  + \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.u1.b ;
assign { \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.u1.cout , \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.u1.s  } = _085_ + \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.u1.cin ;
assign _086_ = \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.u2.a  + \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.u2.b ;
assign { \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.u2.cout , \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.u2.s  } = _086_ + \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.u2.cin ;
always @(posedge \add_17s_17s_17_2_1_U22.top_add_17s_17s_17_2_1_Adder_13_U.clk )
\add_17s_17s_17_2_1_U22.top_add_17s_17s_17_2_1_Adder_13_U.bin_s1  <= _088_;
always @(posedge \add_17s_17s_17_2_1_U22.top_add_17s_17s_17_2_1_Adder_13_U.clk )
\add_17s_17s_17_2_1_U22.top_add_17s_17s_17_2_1_Adder_13_U.ain_s1  <= _087_;
always @(posedge \add_17s_17s_17_2_1_U22.top_add_17s_17s_17_2_1_Adder_13_U.clk )
\add_17s_17s_17_2_1_U22.top_add_17s_17s_17_2_1_Adder_13_U.sum_s1  <= _090_;
always @(posedge \add_17s_17s_17_2_1_U22.top_add_17s_17s_17_2_1_Adder_13_U.clk )
\add_17s_17s_17_2_1_U22.top_add_17s_17s_17_2_1_Adder_13_U.carry_s1  <= _089_;
assign _088_ = \add_17s_17s_17_2_1_U22.top_add_17s_17s_17_2_1_Adder_13_U.ce  ? \add_17s_17s_17_2_1_U22.top_add_17s_17s_17_2_1_Adder_13_U.b [16:8] : \add_17s_17s_17_2_1_U22.top_add_17s_17s_17_2_1_Adder_13_U.bin_s1 ;
assign _087_ = \add_17s_17s_17_2_1_U22.top_add_17s_17s_17_2_1_Adder_13_U.ce  ? \add_17s_17s_17_2_1_U22.top_add_17s_17s_17_2_1_Adder_13_U.a [16:8] : \add_17s_17s_17_2_1_U22.top_add_17s_17s_17_2_1_Adder_13_U.ain_s1 ;
assign _089_ = \add_17s_17s_17_2_1_U22.top_add_17s_17s_17_2_1_Adder_13_U.ce  ? \add_17s_17s_17_2_1_U22.top_add_17s_17s_17_2_1_Adder_13_U.facout_s1  : \add_17s_17s_17_2_1_U22.top_add_17s_17s_17_2_1_Adder_13_U.carry_s1 ;
assign _090_ = \add_17s_17s_17_2_1_U22.top_add_17s_17s_17_2_1_Adder_13_U.ce  ? \add_17s_17s_17_2_1_U22.top_add_17s_17s_17_2_1_Adder_13_U.fas_s1  : \add_17s_17s_17_2_1_U22.top_add_17s_17s_17_2_1_Adder_13_U.sum_s1 ;
assign _091_ = \add_17s_17s_17_2_1_U22.top_add_17s_17s_17_2_1_Adder_13_U.u1.a  + \add_17s_17s_17_2_1_U22.top_add_17s_17s_17_2_1_Adder_13_U.u1.b ;
assign { \add_17s_17s_17_2_1_U22.top_add_17s_17s_17_2_1_Adder_13_U.u1.cout , \add_17s_17s_17_2_1_U22.top_add_17s_17s_17_2_1_Adder_13_U.u1.s  } = _091_ + \add_17s_17s_17_2_1_U22.top_add_17s_17s_17_2_1_Adder_13_U.u1.cin ;
assign _092_ = \add_17s_17s_17_2_1_U22.top_add_17s_17s_17_2_1_Adder_13_U.u2.a  + \add_17s_17s_17_2_1_U22.top_add_17s_17s_17_2_1_Adder_13_U.u2.b ;
assign { \add_17s_17s_17_2_1_U22.top_add_17s_17s_17_2_1_Adder_13_U.u2.cout , \add_17s_17s_17_2_1_U22.top_add_17s_17s_17_2_1_Adder_13_U.u2.s  } = _092_ + \add_17s_17s_17_2_1_U22.top_add_17s_17s_17_2_1_Adder_13_U.u2.cin ;
always @(posedge \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_10_U.clk )
\add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_10_U.bin_s1  <= _094_;
always @(posedge \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_10_U.clk )
\add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_10_U.ain_s1  <= _093_;
always @(posedge \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_10_U.clk )
\add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_10_U.sum_s1  <= _096_;
always @(posedge \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_10_U.clk )
\add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_10_U.carry_s1  <= _095_;
assign _094_ = \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_10_U.ce  ? \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_10_U.b [1] : \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_10_U.bin_s1 ;
assign _093_ = \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_10_U.ce  ? \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_10_U.a [1] : \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_10_U.ain_s1 ;
assign _095_ = \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_10_U.ce  ? \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_10_U.facout_s1  : \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_10_U.carry_s1 ;
assign _096_ = \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_10_U.ce  ? \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_10_U.fas_s1  : \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_10_U.sum_s1 ;
assign _097_ = \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_10_U.u1.a  + \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_10_U.u1.b ;
assign { \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_10_U.u1.cout , \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_10_U.u1.s  } = _097_ + \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_10_U.u1.cin ;
assign _098_ = \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_10_U.u2.a  + \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_10_U.u2.b ;
assign { \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_10_U.u2.cout , \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_10_U.u2.s  } = _098_ + \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_10_U.u2.cin ;
always @(posedge \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.clk )
\add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.bin_s1  <= _100_;
always @(posedge \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.clk )
\add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.ain_s1  <= _099_;
always @(posedge \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.clk )
\add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.sum_s1  <= _102_;
always @(posedge \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.clk )
\add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.carry_s1  <= _101_;
assign _100_ = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.ce  ? \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.b [31:16] : \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.bin_s1 ;
assign _099_ = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.ce  ? \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.a [31:16] : \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.ain_s1 ;
assign _101_ = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.ce  ? \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.facout_s1  : \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.carry_s1 ;
assign _102_ = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.ce  ? \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.fas_s1  : \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.sum_s1 ;
assign _103_ = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.a  + \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.b ;
assign { \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.cout , \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.s  } = _103_ + \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.cin ;
assign _104_ = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.a  + \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.b ;
assign { \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.cout , \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.s  } = _104_ + \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.cin ;
always @(posedge \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_5_U.clk )
\add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_5_U.bin_s1  <= _106_;
always @(posedge \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_5_U.clk )
\add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_5_U.ain_s1  <= _105_;
always @(posedge \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_5_U.clk )
\add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_5_U.sum_s1  <= _108_;
always @(posedge \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_5_U.clk )
\add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_5_U.carry_s1  <= _107_;
assign _106_ = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_5_U.ce  ? \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_5_U.b [31:16] : \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_5_U.bin_s1 ;
assign _105_ = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_5_U.ce  ? \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_5_U.a [31:16] : \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_5_U.ain_s1 ;
assign _107_ = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_5_U.ce  ? \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_5_U.facout_s1  : \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_5_U.carry_s1 ;
assign _108_ = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_5_U.ce  ? \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_5_U.fas_s1  : \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_5_U.sum_s1 ;
assign _109_ = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.a  + \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.b ;
assign { \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.cout , \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.s  } = _109_ + \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.cin ;
assign _110_ = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.a  + \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.b ;
assign { \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.cout , \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.s  } = _110_ + \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.cin ;
always @(posedge \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_5_U.clk )
\add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_5_U.bin_s1  <= _112_;
always @(posedge \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_5_U.clk )
\add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_5_U.ain_s1  <= _111_;
always @(posedge \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_5_U.clk )
\add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_5_U.sum_s1  <= _114_;
always @(posedge \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_5_U.clk )
\add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_5_U.carry_s1  <= _113_;
assign _112_ = \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_5_U.ce  ? \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_5_U.b [31:16] : \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_5_U.bin_s1 ;
assign _111_ = \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_5_U.ce  ? \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_5_U.a [31:16] : \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_5_U.ain_s1 ;
assign _113_ = \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_5_U.ce  ? \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_5_U.facout_s1  : \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_5_U.carry_s1 ;
assign _114_ = \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_5_U.ce  ? \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_5_U.fas_s1  : \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_5_U.sum_s1 ;
assign _115_ = \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.a  + \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.b ;
assign { \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.cout , \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.s  } = _115_ + \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.cin ;
assign _116_ = \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.a  + \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.b ;
assign { \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.cout , \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.s  } = _116_ + \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.cin ;
always @(posedge \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_5_U.clk )
\add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_5_U.bin_s1  <= _118_;
always @(posedge \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_5_U.clk )
\add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_5_U.ain_s1  <= _117_;
always @(posedge \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_5_U.clk )
\add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_5_U.sum_s1  <= _120_;
always @(posedge \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_5_U.clk )
\add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_5_U.carry_s1  <= _119_;
assign _118_ = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_5_U.ce  ? \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_5_U.b [31:16] : \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_5_U.bin_s1 ;
assign _117_ = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_5_U.ce  ? \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_5_U.a [31:16] : \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_5_U.ain_s1 ;
assign _119_ = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_5_U.ce  ? \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_5_U.facout_s1  : \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_5_U.carry_s1 ;
assign _120_ = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_5_U.ce  ? \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_5_U.fas_s1  : \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_5_U.sum_s1 ;
assign _121_ = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.a  + \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.b ;
assign { \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.cout , \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.s  } = _121_ + \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.cin ;
assign _122_ = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.a  + \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.b ;
assign { \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.cout , \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.s  } = _122_ + \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.cin ;
always @(posedge \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.clk )
\add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.bin_s1  <= _124_;
always @(posedge \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.clk )
\add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.ain_s1  <= _123_;
always @(posedge \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.clk )
\add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.sum_s1  <= _126_;
always @(posedge \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.clk )
\add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.carry_s1  <= _125_;
assign _124_ = \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.ce  ? \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.b [31:16] : \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.bin_s1 ;
assign _123_ = \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.ce  ? \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.a [31:16] : \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.ain_s1 ;
assign _125_ = \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.ce  ? \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.facout_s1  : \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.carry_s1 ;
assign _126_ = \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.ce  ? \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.fas_s1  : \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.sum_s1 ;
assign _127_ = \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.a  + \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.b ;
assign { \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.cout , \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.s  } = _127_ + \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.cin ;
assign _128_ = \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.a  + \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.b ;
assign { \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.cout , \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.s  } = _128_ + \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.cin ;
always @(posedge \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_14_U.clk )
\add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_14_U.bin_s1  <= _130_;
always @(posedge \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_14_U.clk )
\add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_14_U.ain_s1  <= _129_;
always @(posedge \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_14_U.clk )
\add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_14_U.sum_s1  <= _132_;
always @(posedge \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_14_U.clk )
\add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_14_U.carry_s1  <= _131_;
assign _130_ = \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_14_U.ce  ? \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_14_U.b [31:16] : \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_14_U.bin_s1 ;
assign _129_ = \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_14_U.ce  ? \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_14_U.a [31:16] : \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_14_U.ain_s1 ;
assign _131_ = \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_14_U.ce  ? \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_14_U.facout_s1  : \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_14_U.carry_s1 ;
assign _132_ = \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_14_U.ce  ? \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_14_U.fas_s1  : \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_14_U.sum_s1 ;
assign _133_ = \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_14_U.u1.a  + \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_14_U.u1.b ;
assign { \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_14_U.u1.cout , \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_14_U.u1.s  } = _133_ + \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_14_U.u1.cin ;
assign _134_ = \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_14_U.u2.a  + \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_14_U.u2.b ;
assign { \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_14_U.u2.cout , \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_14_U.u2.s  } = _134_ + \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_14_U.u2.cin ;
always @(posedge \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.clk )
\add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.bin_s1  <= _136_;
always @(posedge \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.clk )
\add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.ain_s1  <= _135_;
always @(posedge \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.clk )
\add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.sum_s1  <= _138_;
always @(posedge \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.clk )
\add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.carry_s1  <= _137_;
assign _136_ = \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.ce  ? \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.b [33:17] : \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.bin_s1 ;
assign _135_ = \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.ce  ? \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.a [33:17] : \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.ain_s1 ;
assign _137_ = \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.ce  ? \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.facout_s1  : \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.carry_s1 ;
assign _138_ = \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.ce  ? \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.fas_s1  : \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.sum_s1 ;
assign _139_ = \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.u1.a  + \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.u1.b ;
assign { \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.u1.cout , \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.u1.s  } = _139_ + \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.u1.cin ;
assign _140_ = \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.u2.a  + \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.u2.b ;
assign { \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.u2.cout , \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.u2.s  } = _140_ + \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.u2.cin ;
always @(posedge \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.clk )
\add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.bin_s1  <= _142_;
always @(posedge \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.clk )
\add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.ain_s1  <= _141_;
always @(posedge \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.clk )
\add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.sum_s1  <= _144_;
always @(posedge \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.clk )
\add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.carry_s1  <= _143_;
assign _142_ = \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.ce  ? \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.b [34:17] : \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.bin_s1 ;
assign _141_ = \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.ce  ? \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.a [34:17] : \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.ain_s1 ;
assign _143_ = \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.ce  ? \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.facout_s1  : \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.carry_s1 ;
assign _144_ = \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.ce  ? \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.fas_s1  : \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.sum_s1 ;
assign _145_ = \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.u1.a  + \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.u1.b ;
assign { \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.u1.cout , \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.u1.s  } = _145_ + \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.u1.cin ;
assign _146_ = \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.u2.a  + \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.u2.b ;
assign { \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.u2.cout , \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.u2.s  } = _146_ + \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.u2.cin ;
always @(posedge \add_3s_3ns_3_2_1_U20.top_add_3s_3ns_3_2_1_Adder_12_U.clk )
\add_3s_3ns_3_2_1_U20.top_add_3s_3ns_3_2_1_Adder_12_U.bin_s1  <= _148_;
always @(posedge \add_3s_3ns_3_2_1_U20.top_add_3s_3ns_3_2_1_Adder_12_U.clk )
\add_3s_3ns_3_2_1_U20.top_add_3s_3ns_3_2_1_Adder_12_U.ain_s1  <= _147_;
always @(posedge \add_3s_3ns_3_2_1_U20.top_add_3s_3ns_3_2_1_Adder_12_U.clk )
\add_3s_3ns_3_2_1_U20.top_add_3s_3ns_3_2_1_Adder_12_U.sum_s1  <= _150_;
always @(posedge \add_3s_3ns_3_2_1_U20.top_add_3s_3ns_3_2_1_Adder_12_U.clk )
\add_3s_3ns_3_2_1_U20.top_add_3s_3ns_3_2_1_Adder_12_U.carry_s1  <= _149_;
assign _148_ = \add_3s_3ns_3_2_1_U20.top_add_3s_3ns_3_2_1_Adder_12_U.ce  ? \add_3s_3ns_3_2_1_U20.top_add_3s_3ns_3_2_1_Adder_12_U.b [2:1] : \add_3s_3ns_3_2_1_U20.top_add_3s_3ns_3_2_1_Adder_12_U.bin_s1 ;
assign _147_ = \add_3s_3ns_3_2_1_U20.top_add_3s_3ns_3_2_1_Adder_12_U.ce  ? \add_3s_3ns_3_2_1_U20.top_add_3s_3ns_3_2_1_Adder_12_U.a [2:1] : \add_3s_3ns_3_2_1_U20.top_add_3s_3ns_3_2_1_Adder_12_U.ain_s1 ;
assign _149_ = \add_3s_3ns_3_2_1_U20.top_add_3s_3ns_3_2_1_Adder_12_U.ce  ? \add_3s_3ns_3_2_1_U20.top_add_3s_3ns_3_2_1_Adder_12_U.facout_s1  : \add_3s_3ns_3_2_1_U20.top_add_3s_3ns_3_2_1_Adder_12_U.carry_s1 ;
assign _150_ = \add_3s_3ns_3_2_1_U20.top_add_3s_3ns_3_2_1_Adder_12_U.ce  ? \add_3s_3ns_3_2_1_U20.top_add_3s_3ns_3_2_1_Adder_12_U.fas_s1  : \add_3s_3ns_3_2_1_U20.top_add_3s_3ns_3_2_1_Adder_12_U.sum_s1 ;
assign _151_ = \add_3s_3ns_3_2_1_U20.top_add_3s_3ns_3_2_1_Adder_12_U.u1.a  + \add_3s_3ns_3_2_1_U20.top_add_3s_3ns_3_2_1_Adder_12_U.u1.b ;
assign { \add_3s_3ns_3_2_1_U20.top_add_3s_3ns_3_2_1_Adder_12_U.u1.cout , \add_3s_3ns_3_2_1_U20.top_add_3s_3ns_3_2_1_Adder_12_U.u1.s  } = _151_ + \add_3s_3ns_3_2_1_U20.top_add_3s_3ns_3_2_1_Adder_12_U.u1.cin ;
assign _152_ = \add_3s_3ns_3_2_1_U20.top_add_3s_3ns_3_2_1_Adder_12_U.u2.a  + \add_3s_3ns_3_2_1_U20.top_add_3s_3ns_3_2_1_Adder_12_U.u2.b ;
assign { \add_3s_3ns_3_2_1_U20.top_add_3s_3ns_3_2_1_Adder_12_U.u2.cout , \add_3s_3ns_3_2_1_U20.top_add_3s_3ns_3_2_1_Adder_12_U.u2.s  } = _152_ + \add_3s_3ns_3_2_1_U20.top_add_3s_3ns_3_2_1_Adder_12_U.u2.cin ;
always @(posedge \add_45s_45s_45_2_1_U8.top_add_45s_45s_45_2_1_Adder_7_U.clk )
\add_45s_45s_45_2_1_U8.top_add_45s_45s_45_2_1_Adder_7_U.bin_s1  <= _154_;
always @(posedge \add_45s_45s_45_2_1_U8.top_add_45s_45s_45_2_1_Adder_7_U.clk )
\add_45s_45s_45_2_1_U8.top_add_45s_45s_45_2_1_Adder_7_U.ain_s1  <= _153_;
always @(posedge \add_45s_45s_45_2_1_U8.top_add_45s_45s_45_2_1_Adder_7_U.clk )
\add_45s_45s_45_2_1_U8.top_add_45s_45s_45_2_1_Adder_7_U.sum_s1  <= _156_;
always @(posedge \add_45s_45s_45_2_1_U8.top_add_45s_45s_45_2_1_Adder_7_U.clk )
\add_45s_45s_45_2_1_U8.top_add_45s_45s_45_2_1_Adder_7_U.carry_s1  <= _155_;
assign _154_ = \add_45s_45s_45_2_1_U8.top_add_45s_45s_45_2_1_Adder_7_U.ce  ? \add_45s_45s_45_2_1_U8.top_add_45s_45s_45_2_1_Adder_7_U.b [44:22] : \add_45s_45s_45_2_1_U8.top_add_45s_45s_45_2_1_Adder_7_U.bin_s1 ;
assign _153_ = \add_45s_45s_45_2_1_U8.top_add_45s_45s_45_2_1_Adder_7_U.ce  ? \add_45s_45s_45_2_1_U8.top_add_45s_45s_45_2_1_Adder_7_U.a [44:22] : \add_45s_45s_45_2_1_U8.top_add_45s_45s_45_2_1_Adder_7_U.ain_s1 ;
assign _155_ = \add_45s_45s_45_2_1_U8.top_add_45s_45s_45_2_1_Adder_7_U.ce  ? \add_45s_45s_45_2_1_U8.top_add_45s_45s_45_2_1_Adder_7_U.facout_s1  : \add_45s_45s_45_2_1_U8.top_add_45s_45s_45_2_1_Adder_7_U.carry_s1 ;
assign _156_ = \add_45s_45s_45_2_1_U8.top_add_45s_45s_45_2_1_Adder_7_U.ce  ? \add_45s_45s_45_2_1_U8.top_add_45s_45s_45_2_1_Adder_7_U.fas_s1  : \add_45s_45s_45_2_1_U8.top_add_45s_45s_45_2_1_Adder_7_U.sum_s1 ;
assign _157_ = \add_45s_45s_45_2_1_U8.top_add_45s_45s_45_2_1_Adder_7_U.u1.a  + \add_45s_45s_45_2_1_U8.top_add_45s_45s_45_2_1_Adder_7_U.u1.b ;
assign { \add_45s_45s_45_2_1_U8.top_add_45s_45s_45_2_1_Adder_7_U.u1.cout , \add_45s_45s_45_2_1_U8.top_add_45s_45s_45_2_1_Adder_7_U.u1.s  } = _157_ + \add_45s_45s_45_2_1_U8.top_add_45s_45s_45_2_1_Adder_7_U.u1.cin ;
assign _158_ = \add_45s_45s_45_2_1_U8.top_add_45s_45s_45_2_1_Adder_7_U.u2.a  + \add_45s_45s_45_2_1_U8.top_add_45s_45s_45_2_1_Adder_7_U.u2.b ;
assign { \add_45s_45s_45_2_1_U8.top_add_45s_45s_45_2_1_Adder_7_U.u2.cout , \add_45s_45s_45_2_1_U8.top_add_45s_45s_45_2_1_Adder_7_U.u2.s  } = _158_ + \add_45s_45s_45_2_1_U8.top_add_45s_45s_45_2_1_Adder_7_U.u2.cin ;
always @(posedge \add_46s_46s_46_2_1_U5.top_add_46s_46s_46_2_1_Adder_4_U.clk )
\add_46s_46s_46_2_1_U5.top_add_46s_46s_46_2_1_Adder_4_U.bin_s1  <= _160_;
always @(posedge \add_46s_46s_46_2_1_U5.top_add_46s_46s_46_2_1_Adder_4_U.clk )
\add_46s_46s_46_2_1_U5.top_add_46s_46s_46_2_1_Adder_4_U.ain_s1  <= _159_;
always @(posedge \add_46s_46s_46_2_1_U5.top_add_46s_46s_46_2_1_Adder_4_U.clk )
\add_46s_46s_46_2_1_U5.top_add_46s_46s_46_2_1_Adder_4_U.sum_s1  <= _162_;
always @(posedge \add_46s_46s_46_2_1_U5.top_add_46s_46s_46_2_1_Adder_4_U.clk )
\add_46s_46s_46_2_1_U5.top_add_46s_46s_46_2_1_Adder_4_U.carry_s1  <= _161_;
assign _160_ = \add_46s_46s_46_2_1_U5.top_add_46s_46s_46_2_1_Adder_4_U.ce  ? \add_46s_46s_46_2_1_U5.top_add_46s_46s_46_2_1_Adder_4_U.b [45:23] : \add_46s_46s_46_2_1_U5.top_add_46s_46s_46_2_1_Adder_4_U.bin_s1 ;
assign _159_ = \add_46s_46s_46_2_1_U5.top_add_46s_46s_46_2_1_Adder_4_U.ce  ? \add_46s_46s_46_2_1_U5.top_add_46s_46s_46_2_1_Adder_4_U.a [45:23] : \add_46s_46s_46_2_1_U5.top_add_46s_46s_46_2_1_Adder_4_U.ain_s1 ;
assign _161_ = \add_46s_46s_46_2_1_U5.top_add_46s_46s_46_2_1_Adder_4_U.ce  ? \add_46s_46s_46_2_1_U5.top_add_46s_46s_46_2_1_Adder_4_U.facout_s1  : \add_46s_46s_46_2_1_U5.top_add_46s_46s_46_2_1_Adder_4_U.carry_s1 ;
assign _162_ = \add_46s_46s_46_2_1_U5.top_add_46s_46s_46_2_1_Adder_4_U.ce  ? \add_46s_46s_46_2_1_U5.top_add_46s_46s_46_2_1_Adder_4_U.fas_s1  : \add_46s_46s_46_2_1_U5.top_add_46s_46s_46_2_1_Adder_4_U.sum_s1 ;
assign _163_ = \add_46s_46s_46_2_1_U5.top_add_46s_46s_46_2_1_Adder_4_U.u1.a  + \add_46s_46s_46_2_1_U5.top_add_46s_46s_46_2_1_Adder_4_U.u1.b ;
assign { \add_46s_46s_46_2_1_U5.top_add_46s_46s_46_2_1_Adder_4_U.u1.cout , \add_46s_46s_46_2_1_U5.top_add_46s_46s_46_2_1_Adder_4_U.u1.s  } = _163_ + \add_46s_46s_46_2_1_U5.top_add_46s_46s_46_2_1_Adder_4_U.u1.cin ;
assign _164_ = \add_46s_46s_46_2_1_U5.top_add_46s_46s_46_2_1_Adder_4_U.u2.a  + \add_46s_46s_46_2_1_U5.top_add_46s_46s_46_2_1_Adder_4_U.u2.b ;
assign { \add_46s_46s_46_2_1_U5.top_add_46s_46s_46_2_1_Adder_4_U.u2.cout , \add_46s_46s_46_2_1_U5.top_add_46s_46s_46_2_1_Adder_4_U.u2.s  } = _164_ + \add_46s_46s_46_2_1_U5.top_add_46s_46s_46_2_1_Adder_4_U.u2.cin ;
always @(posedge \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.clk )
\add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.bin_s1  <= _166_;
always @(posedge \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.clk )
\add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.ain_s1  <= _165_;
always @(posedge \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.clk )
\add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.sum_s1  <= _168_;
always @(posedge \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.clk )
\add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.carry_s1  <= _167_;
assign _166_ = \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.ce  ? \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.b [8:4] : \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.bin_s1 ;
assign _165_ = \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.ce  ? \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.a [8:4] : \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.ain_s1 ;
assign _167_ = \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.ce  ? \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.facout_s1  : \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.carry_s1 ;
assign _168_ = \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.ce  ? \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.fas_s1  : \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.sum_s1 ;
assign _169_ = \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.u1.a  + \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.u1.b ;
assign { \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.u1.cout , \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.u1.s  } = _169_ + \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.u1.cin ;
assign _170_ = \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.u2.a  + \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.u2.b ;
assign { \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.u2.cout , \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.u2.s  } = _170_ + \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.u2.cin ;
always @(posedge \ashr_16ns_4ns_16_7_1_U14.clk )
\ashr_16ns_4ns_16_7_1_U14.dout_array[5]  <= _182_;
always @(posedge \ashr_16ns_4ns_16_7_1_U14.clk )
\ashr_16ns_4ns_16_7_1_U14.din1_cast_array[5]  <= _176_;
always @(posedge \ashr_16ns_4ns_16_7_1_U14.clk )
\ashr_16ns_4ns_16_7_1_U14.dout_array[4]  <= _181_;
always @(posedge \ashr_16ns_4ns_16_7_1_U14.clk )
\ashr_16ns_4ns_16_7_1_U14.din1_cast_array[4]  <= _175_;
always @(posedge \ashr_16ns_4ns_16_7_1_U14.clk )
\ashr_16ns_4ns_16_7_1_U14.dout_array[3]  <= _180_;
always @(posedge \ashr_16ns_4ns_16_7_1_U14.clk )
\ashr_16ns_4ns_16_7_1_U14.din1_cast_array[3]  <= _174_;
always @(posedge \ashr_16ns_4ns_16_7_1_U14.clk )
\ashr_16ns_4ns_16_7_1_U14.dout_array[2]  <= _179_;
always @(posedge \ashr_16ns_4ns_16_7_1_U14.clk )
\ashr_16ns_4ns_16_7_1_U14.din1_cast_array[2]  <= _173_;
always @(posedge \ashr_16ns_4ns_16_7_1_U14.clk )
\ashr_16ns_4ns_16_7_1_U14.dout_array[1]  <= _178_;
always @(posedge \ashr_16ns_4ns_16_7_1_U14.clk )
\ashr_16ns_4ns_16_7_1_U14.din1_cast_array[1]  <= _172_;
always @(posedge \ashr_16ns_4ns_16_7_1_U14.clk )
\ashr_16ns_4ns_16_7_1_U14.dout_array[0]  <= _177_;
always @(posedge \ashr_16ns_4ns_16_7_1_U14.clk )
\ashr_16ns_4ns_16_7_1_U14.din1_cast_array[0]  <= _171_;
assign _183_ = \ashr_16ns_4ns_16_7_1_U14.ce  ? \ashr_16ns_4ns_16_7_1_U14.din1_cast_array[4]  : \ashr_16ns_4ns_16_7_1_U14.din1_cast_array[5] ;
assign _176_ = \ashr_16ns_4ns_16_7_1_U14.reset  ? 4'h0 : _183_;
assign _184_ = \ashr_16ns_4ns_16_7_1_U14.ce  ? _197_ : \ashr_16ns_4ns_16_7_1_U14.dout_array[5] ;
assign _182_ = \ashr_16ns_4ns_16_7_1_U14.reset  ? 16'h0000 : _184_;
assign _185_ = \ashr_16ns_4ns_16_7_1_U14.ce  ? \ashr_16ns_4ns_16_7_1_U14.din1_cast_array[3]  : \ashr_16ns_4ns_16_7_1_U14.din1_cast_array[4] ;
assign _175_ = \ashr_16ns_4ns_16_7_1_U14.reset  ? 4'h0 : _185_;
assign _186_ = \ashr_16ns_4ns_16_7_1_U14.ce  ? _196_ : \ashr_16ns_4ns_16_7_1_U14.dout_array[4] ;
assign _181_ = \ashr_16ns_4ns_16_7_1_U14.reset  ? 16'h0000 : _186_;
assign _187_ = \ashr_16ns_4ns_16_7_1_U14.ce  ? \ashr_16ns_4ns_16_7_1_U14.din1_cast_array[2]  : \ashr_16ns_4ns_16_7_1_U14.din1_cast_array[3] ;
assign _174_ = \ashr_16ns_4ns_16_7_1_U14.reset  ? 4'h0 : _187_;
assign _188_ = \ashr_16ns_4ns_16_7_1_U14.ce  ? _195_ : \ashr_16ns_4ns_16_7_1_U14.dout_array[3] ;
assign _180_ = \ashr_16ns_4ns_16_7_1_U14.reset  ? 16'h0000 : _188_;
assign _189_ = \ashr_16ns_4ns_16_7_1_U14.ce  ? \ashr_16ns_4ns_16_7_1_U14.din1_cast_array[1]  : \ashr_16ns_4ns_16_7_1_U14.din1_cast_array[2] ;
assign _173_ = \ashr_16ns_4ns_16_7_1_U14.reset  ? 4'h0 : _189_;
assign _190_ = \ashr_16ns_4ns_16_7_1_U14.ce  ? \ashr_16ns_4ns_16_7_1_U14.dout_array[1]  : \ashr_16ns_4ns_16_7_1_U14.dout_array[2] ;
assign _179_ = \ashr_16ns_4ns_16_7_1_U14.reset  ? 16'h0000 : _190_;
assign _191_ = \ashr_16ns_4ns_16_7_1_U14.ce  ? \ashr_16ns_4ns_16_7_1_U14.din1_cast_array[0]  : \ashr_16ns_4ns_16_7_1_U14.din1_cast_array[1] ;
assign _172_ = \ashr_16ns_4ns_16_7_1_U14.reset  ? 4'h0 : _191_;
assign _192_ = \ashr_16ns_4ns_16_7_1_U14.ce  ? \ashr_16ns_4ns_16_7_1_U14.dout_array[0]  : \ashr_16ns_4ns_16_7_1_U14.dout_array[1] ;
assign _178_ = \ashr_16ns_4ns_16_7_1_U14.reset  ? 16'h0000 : _192_;
assign _193_ = \ashr_16ns_4ns_16_7_1_U14.ce  ? \ashr_16ns_4ns_16_7_1_U14.din1 [3:0] : \ashr_16ns_4ns_16_7_1_U14.din1_cast_array[0] ;
assign _171_ = \ashr_16ns_4ns_16_7_1_U14.reset  ? 4'h0 : _193_;
assign _194_ = \ashr_16ns_4ns_16_7_1_U14.ce  ? \ashr_16ns_4ns_16_7_1_U14.din0  : \ashr_16ns_4ns_16_7_1_U14.dout_array[0] ;
assign _177_ = \ashr_16ns_4ns_16_7_1_U14.reset  ? 16'h0000 : _194_;
assign _195_ = $signed(\ashr_16ns_4ns_16_7_1_U14.dout_array[2] ) >>> { \ashr_16ns_4ns_16_7_1_U14.din1_cast_array[2] [3], 3'h0 };
assign _196_ = $signed(\ashr_16ns_4ns_16_7_1_U14.dout_array[3] ) >>> { \ashr_16ns_4ns_16_7_1_U14.din1_cast_array[3] [2], 2'h0 };
assign _197_ = $signed(\ashr_16ns_4ns_16_7_1_U14.dout_array[4] ) >>> { \ashr_16ns_4ns_16_7_1_U14.din1_cast_array[4] [1], 1'h0 };
assign \ashr_16ns_4ns_16_7_1_U14.dout  = $signed(\ashr_16ns_4ns_16_7_1_U14.dout_array[5] ) >>> \ashr_16ns_4ns_16_7_1_U14.din1_cast_array[5] [0];
always @(posedge \ashr_32s_32s_32_7_1_U10.clk )
\ashr_32s_32s_32_7_1_U10.dout_array[5]  <= _209_;
always @(posedge \ashr_32s_32s_32_7_1_U10.clk )
\ashr_32s_32s_32_7_1_U10.din1_cast_array[5]  <= _203_;
always @(posedge \ashr_32s_32s_32_7_1_U10.clk )
\ashr_32s_32s_32_7_1_U10.dout_array[4]  <= _208_;
always @(posedge \ashr_32s_32s_32_7_1_U10.clk )
\ashr_32s_32s_32_7_1_U10.din1_cast_array[4]  <= _202_;
always @(posedge \ashr_32s_32s_32_7_1_U10.clk )
\ashr_32s_32s_32_7_1_U10.dout_array[3]  <= _207_;
always @(posedge \ashr_32s_32s_32_7_1_U10.clk )
\ashr_32s_32s_32_7_1_U10.din1_cast_array[3]  <= _201_;
always @(posedge \ashr_32s_32s_32_7_1_U10.clk )
\ashr_32s_32s_32_7_1_U10.dout_array[2]  <= _206_;
always @(posedge \ashr_32s_32s_32_7_1_U10.clk )
\ashr_32s_32s_32_7_1_U10.din1_cast_array[2]  <= _200_;
always @(posedge \ashr_32s_32s_32_7_1_U10.clk )
\ashr_32s_32s_32_7_1_U10.dout_array[1]  <= _205_;
always @(posedge \ashr_32s_32s_32_7_1_U10.clk )
\ashr_32s_32s_32_7_1_U10.din1_cast_array[1]  <= _199_;
always @(posedge \ashr_32s_32s_32_7_1_U10.clk )
\ashr_32s_32s_32_7_1_U10.dout_array[0]  <= _204_;
always @(posedge \ashr_32s_32s_32_7_1_U10.clk )
\ashr_32s_32s_32_7_1_U10.din1_cast_array[0]  <= _198_;
assign _210_ = \ashr_32s_32s_32_7_1_U10.ce  ? \ashr_32s_32s_32_7_1_U10.din1_cast_array[4]  : \ashr_32s_32s_32_7_1_U10.din1_cast_array[5] ;
assign _203_ = \ashr_32s_32s_32_7_1_U10.reset  ? 32'd0 : _210_;
assign _211_ = \ashr_32s_32s_32_7_1_U10.ce  ? _227_ : \ashr_32s_32s_32_7_1_U10.dout_array[5] ;
assign _209_ = \ashr_32s_32s_32_7_1_U10.reset  ? 32'd0 : _211_;
assign _212_ = \ashr_32s_32s_32_7_1_U10.ce  ? \ashr_32s_32s_32_7_1_U10.din1_cast_array[3]  : \ashr_32s_32s_32_7_1_U10.din1_cast_array[4] ;
assign _202_ = \ashr_32s_32s_32_7_1_U10.reset  ? 32'd0 : _212_;
assign _213_ = \ashr_32s_32s_32_7_1_U10.ce  ? _226_ : \ashr_32s_32s_32_7_1_U10.dout_array[4] ;
assign _208_ = \ashr_32s_32s_32_7_1_U10.reset  ? 32'd0 : _213_;
assign _214_ = \ashr_32s_32s_32_7_1_U10.ce  ? \ashr_32s_32s_32_7_1_U10.din1_cast_array[2]  : \ashr_32s_32s_32_7_1_U10.din1_cast_array[3] ;
assign _201_ = \ashr_32s_32s_32_7_1_U10.reset  ? 32'd0 : _214_;
assign _215_ = \ashr_32s_32s_32_7_1_U10.ce  ? _225_ : \ashr_32s_32s_32_7_1_U10.dout_array[3] ;
assign _207_ = \ashr_32s_32s_32_7_1_U10.reset  ? 32'd0 : _215_;
assign _216_ = \ashr_32s_32s_32_7_1_U10.ce  ? \ashr_32s_32s_32_7_1_U10.din1_cast_array[1]  : \ashr_32s_32s_32_7_1_U10.din1_cast_array[2] ;
assign _200_ = \ashr_32s_32s_32_7_1_U10.reset  ? 32'd0 : _216_;
assign _217_ = \ashr_32s_32s_32_7_1_U10.ce  ? _224_ : \ashr_32s_32s_32_7_1_U10.dout_array[2] ;
assign _206_ = \ashr_32s_32s_32_7_1_U10.reset  ? 32'd0 : _217_;
assign _218_ = \ashr_32s_32s_32_7_1_U10.ce  ? \ashr_32s_32s_32_7_1_U10.din1_cast_array[0]  : \ashr_32s_32s_32_7_1_U10.din1_cast_array[1] ;
assign _199_ = \ashr_32s_32s_32_7_1_U10.reset  ? 32'd0 : _218_;
assign _219_ = \ashr_32s_32s_32_7_1_U10.ce  ? _223_ : \ashr_32s_32s_32_7_1_U10.dout_array[1] ;
assign _205_ = \ashr_32s_32s_32_7_1_U10.reset  ? 32'd0 : _219_;
assign _220_ = \ashr_32s_32s_32_7_1_U10.ce  ? \ashr_32s_32s_32_7_1_U10.din1  : \ashr_32s_32s_32_7_1_U10.din1_cast_array[0] ;
assign _198_ = \ashr_32s_32s_32_7_1_U10.reset  ? 32'd0 : _220_;
assign _221_ = \ashr_32s_32s_32_7_1_U10.ce  ? _222_ : \ashr_32s_32s_32_7_1_U10.dout_array[0] ;
assign _204_ = \ashr_32s_32s_32_7_1_U10.reset  ? 32'd0 : _221_;
assign _222_ = $signed(\ashr_32s_32s_32_7_1_U10.din0 ) >>> { \ashr_32s_32s_32_7_1_U10.din1 [31:30], 30'h00000000 };
assign _223_ = $signed(\ashr_32s_32s_32_7_1_U10.dout_array[0] ) >>> { \ashr_32s_32s_32_7_1_U10.din1_cast_array[0] [29:25], 25'h0000000 };
assign _224_ = $signed(\ashr_32s_32s_32_7_1_U10.dout_array[1] ) >>> { \ashr_32s_32s_32_7_1_U10.din1_cast_array[1] [24:20], 20'h00000 };
assign _225_ = $signed(\ashr_32s_32s_32_7_1_U10.dout_array[2] ) >>> { \ashr_32s_32s_32_7_1_U10.din1_cast_array[2] [19:15], 15'h0000 };
assign _226_ = $signed(\ashr_32s_32s_32_7_1_U10.dout_array[3] ) >>> { \ashr_32s_32s_32_7_1_U10.din1_cast_array[3] [14:10], 10'h000 };
assign _227_ = $signed(\ashr_32s_32s_32_7_1_U10.dout_array[4] ) >>> { \ashr_32s_32s_32_7_1_U10.din1_cast_array[4] [9:5], 5'h00 };
assign \ashr_32s_32s_32_7_1_U10.dout  = $signed(\ashr_32s_32s_32_7_1_U10.dout_array[5] ) >>> \ashr_32s_32s_32_7_1_U10.din1_cast_array[5] [4:0];
always @(posedge \shl_16ns_4ns_16_7_1_U13.clk )
\shl_16ns_4ns_16_7_1_U13.dout_array[5]  <= _239_;
always @(posedge \shl_16ns_4ns_16_7_1_U13.clk )
\shl_16ns_4ns_16_7_1_U13.din1_cast_array[5]  <= _233_;
always @(posedge \shl_16ns_4ns_16_7_1_U13.clk )
\shl_16ns_4ns_16_7_1_U13.dout_array[4]  <= _238_;
always @(posedge \shl_16ns_4ns_16_7_1_U13.clk )
\shl_16ns_4ns_16_7_1_U13.din1_cast_array[4]  <= _232_;
always @(posedge \shl_16ns_4ns_16_7_1_U13.clk )
\shl_16ns_4ns_16_7_1_U13.dout_array[3]  <= _237_;
always @(posedge \shl_16ns_4ns_16_7_1_U13.clk )
\shl_16ns_4ns_16_7_1_U13.din1_cast_array[3]  <= _231_;
always @(posedge \shl_16ns_4ns_16_7_1_U13.clk )
\shl_16ns_4ns_16_7_1_U13.dout_array[2]  <= _236_;
always @(posedge \shl_16ns_4ns_16_7_1_U13.clk )
\shl_16ns_4ns_16_7_1_U13.din1_cast_array[2]  <= _230_;
always @(posedge \shl_16ns_4ns_16_7_1_U13.clk )
\shl_16ns_4ns_16_7_1_U13.dout_array[1]  <= _235_;
always @(posedge \shl_16ns_4ns_16_7_1_U13.clk )
\shl_16ns_4ns_16_7_1_U13.din1_cast_array[1]  <= _229_;
always @(posedge \shl_16ns_4ns_16_7_1_U13.clk )
\shl_16ns_4ns_16_7_1_U13.dout_array[0]  <= _234_;
always @(posedge \shl_16ns_4ns_16_7_1_U13.clk )
\shl_16ns_4ns_16_7_1_U13.din1_cast_array[0]  <= _228_;
assign _240_ = \shl_16ns_4ns_16_7_1_U13.ce  ? \shl_16ns_4ns_16_7_1_U13.din1_cast_array[4]  : \shl_16ns_4ns_16_7_1_U13.din1_cast_array[5] ;
assign _233_ = \shl_16ns_4ns_16_7_1_U13.reset  ? 4'h0 : _240_;
assign _241_ = \shl_16ns_4ns_16_7_1_U13.ce  ? _254_ : \shl_16ns_4ns_16_7_1_U13.dout_array[5] ;
assign _239_ = \shl_16ns_4ns_16_7_1_U13.reset  ? 16'h0000 : _241_;
assign _242_ = \shl_16ns_4ns_16_7_1_U13.ce  ? \shl_16ns_4ns_16_7_1_U13.din1_cast_array[3]  : \shl_16ns_4ns_16_7_1_U13.din1_cast_array[4] ;
assign _232_ = \shl_16ns_4ns_16_7_1_U13.reset  ? 4'h0 : _242_;
assign _243_ = \shl_16ns_4ns_16_7_1_U13.ce  ? _253_ : \shl_16ns_4ns_16_7_1_U13.dout_array[4] ;
assign _238_ = \shl_16ns_4ns_16_7_1_U13.reset  ? 16'h0000 : _243_;
assign _244_ = \shl_16ns_4ns_16_7_1_U13.ce  ? \shl_16ns_4ns_16_7_1_U13.din1_cast_array[2]  : \shl_16ns_4ns_16_7_1_U13.din1_cast_array[3] ;
assign _231_ = \shl_16ns_4ns_16_7_1_U13.reset  ? 4'h0 : _244_;
assign _245_ = \shl_16ns_4ns_16_7_1_U13.ce  ? _252_ : \shl_16ns_4ns_16_7_1_U13.dout_array[3] ;
assign _237_ = \shl_16ns_4ns_16_7_1_U13.reset  ? 16'h0000 : _245_;
assign _246_ = \shl_16ns_4ns_16_7_1_U13.ce  ? \shl_16ns_4ns_16_7_1_U13.din1_cast_array[1]  : \shl_16ns_4ns_16_7_1_U13.din1_cast_array[2] ;
assign _230_ = \shl_16ns_4ns_16_7_1_U13.reset  ? 4'h0 : _246_;
assign _247_ = \shl_16ns_4ns_16_7_1_U13.ce  ? \shl_16ns_4ns_16_7_1_U13.dout_array[1]  : \shl_16ns_4ns_16_7_1_U13.dout_array[2] ;
assign _236_ = \shl_16ns_4ns_16_7_1_U13.reset  ? 16'h0000 : _247_;
assign _248_ = \shl_16ns_4ns_16_7_1_U13.ce  ? \shl_16ns_4ns_16_7_1_U13.din1_cast_array[0]  : \shl_16ns_4ns_16_7_1_U13.din1_cast_array[1] ;
assign _229_ = \shl_16ns_4ns_16_7_1_U13.reset  ? 4'h0 : _248_;
assign _249_ = \shl_16ns_4ns_16_7_1_U13.ce  ? \shl_16ns_4ns_16_7_1_U13.dout_array[0]  : \shl_16ns_4ns_16_7_1_U13.dout_array[1] ;
assign _235_ = \shl_16ns_4ns_16_7_1_U13.reset  ? 16'h0000 : _249_;
assign _250_ = \shl_16ns_4ns_16_7_1_U13.ce  ? \shl_16ns_4ns_16_7_1_U13.din1 [3:0] : \shl_16ns_4ns_16_7_1_U13.din1_cast_array[0] ;
assign _228_ = \shl_16ns_4ns_16_7_1_U13.reset  ? 4'h0 : _250_;
assign _251_ = \shl_16ns_4ns_16_7_1_U13.ce  ? \shl_16ns_4ns_16_7_1_U13.din0  : \shl_16ns_4ns_16_7_1_U13.dout_array[0] ;
assign _234_ = \shl_16ns_4ns_16_7_1_U13.reset  ? 16'h0000 : _251_;
assign _252_ = \shl_16ns_4ns_16_7_1_U13.dout_array[2]  << { \shl_16ns_4ns_16_7_1_U13.din1_cast_array[2] [3], 3'h0 };
assign _253_ = \shl_16ns_4ns_16_7_1_U13.dout_array[3]  << { \shl_16ns_4ns_16_7_1_U13.din1_cast_array[3] [2], 2'h0 };
assign _254_ = \shl_16ns_4ns_16_7_1_U13.dout_array[4]  << { \shl_16ns_4ns_16_7_1_U13.din1_cast_array[4] [1], 1'h0 };
assign \shl_16ns_4ns_16_7_1_U13.dout  = \shl_16ns_4ns_16_7_1_U13.dout_array[5]  << \shl_16ns_4ns_16_7_1_U13.din1_cast_array[5] [0];
always @(posedge \shl_32s_32s_32_7_1_U11.clk )
\shl_32s_32s_32_7_1_U11.dout_array[5]  <= _266_;
always @(posedge \shl_32s_32s_32_7_1_U11.clk )
\shl_32s_32s_32_7_1_U11.din1_cast_array[5]  <= _260_;
always @(posedge \shl_32s_32s_32_7_1_U11.clk )
\shl_32s_32s_32_7_1_U11.dout_array[4]  <= _265_;
always @(posedge \shl_32s_32s_32_7_1_U11.clk )
\shl_32s_32s_32_7_1_U11.din1_cast_array[4]  <= _259_;
always @(posedge \shl_32s_32s_32_7_1_U11.clk )
\shl_32s_32s_32_7_1_U11.dout_array[3]  <= _264_;
always @(posedge \shl_32s_32s_32_7_1_U11.clk )
\shl_32s_32s_32_7_1_U11.din1_cast_array[3]  <= _258_;
always @(posedge \shl_32s_32s_32_7_1_U11.clk )
\shl_32s_32s_32_7_1_U11.dout_array[2]  <= _263_;
always @(posedge \shl_32s_32s_32_7_1_U11.clk )
\shl_32s_32s_32_7_1_U11.din1_cast_array[2]  <= _257_;
always @(posedge \shl_32s_32s_32_7_1_U11.clk )
\shl_32s_32s_32_7_1_U11.dout_array[1]  <= _262_;
always @(posedge \shl_32s_32s_32_7_1_U11.clk )
\shl_32s_32s_32_7_1_U11.din1_cast_array[1]  <= _256_;
always @(posedge \shl_32s_32s_32_7_1_U11.clk )
\shl_32s_32s_32_7_1_U11.dout_array[0]  <= _261_;
always @(posedge \shl_32s_32s_32_7_1_U11.clk )
\shl_32s_32s_32_7_1_U11.din1_cast_array[0]  <= _255_;
assign _267_ = \shl_32s_32s_32_7_1_U11.ce  ? \shl_32s_32s_32_7_1_U11.din1_cast_array[4]  : \shl_32s_32s_32_7_1_U11.din1_cast_array[5] ;
assign _260_ = \shl_32s_32s_32_7_1_U11.reset  ? 32'd0 : _267_;
assign _268_ = \shl_32s_32s_32_7_1_U11.ce  ? _284_ : \shl_32s_32s_32_7_1_U11.dout_array[5] ;
assign _266_ = \shl_32s_32s_32_7_1_U11.reset  ? 32'd0 : _268_;
assign _269_ = \shl_32s_32s_32_7_1_U11.ce  ? \shl_32s_32s_32_7_1_U11.din1_cast_array[3]  : \shl_32s_32s_32_7_1_U11.din1_cast_array[4] ;
assign _259_ = \shl_32s_32s_32_7_1_U11.reset  ? 32'd0 : _269_;
assign _270_ = \shl_32s_32s_32_7_1_U11.ce  ? _283_ : \shl_32s_32s_32_7_1_U11.dout_array[4] ;
assign _265_ = \shl_32s_32s_32_7_1_U11.reset  ? 32'd0 : _270_;
assign _271_ = \shl_32s_32s_32_7_1_U11.ce  ? \shl_32s_32s_32_7_1_U11.din1_cast_array[2]  : \shl_32s_32s_32_7_1_U11.din1_cast_array[3] ;
assign _258_ = \shl_32s_32s_32_7_1_U11.reset  ? 32'd0 : _271_;
assign _272_ = \shl_32s_32s_32_7_1_U11.ce  ? _282_ : \shl_32s_32s_32_7_1_U11.dout_array[3] ;
assign _264_ = \shl_32s_32s_32_7_1_U11.reset  ? 32'd0 : _272_;
assign _273_ = \shl_32s_32s_32_7_1_U11.ce  ? \shl_32s_32s_32_7_1_U11.din1_cast_array[1]  : \shl_32s_32s_32_7_1_U11.din1_cast_array[2] ;
assign _257_ = \shl_32s_32s_32_7_1_U11.reset  ? 32'd0 : _273_;
assign _274_ = \shl_32s_32s_32_7_1_U11.ce  ? _281_ : \shl_32s_32s_32_7_1_U11.dout_array[2] ;
assign _263_ = \shl_32s_32s_32_7_1_U11.reset  ? 32'd0 : _274_;
assign _275_ = \shl_32s_32s_32_7_1_U11.ce  ? \shl_32s_32s_32_7_1_U11.din1_cast_array[0]  : \shl_32s_32s_32_7_1_U11.din1_cast_array[1] ;
assign _256_ = \shl_32s_32s_32_7_1_U11.reset  ? 32'd0 : _275_;
assign _276_ = \shl_32s_32s_32_7_1_U11.ce  ? _280_ : \shl_32s_32s_32_7_1_U11.dout_array[1] ;
assign _262_ = \shl_32s_32s_32_7_1_U11.reset  ? 32'd0 : _276_;
assign _277_ = \shl_32s_32s_32_7_1_U11.ce  ? \shl_32s_32s_32_7_1_U11.din1  : \shl_32s_32s_32_7_1_U11.din1_cast_array[0] ;
assign _255_ = \shl_32s_32s_32_7_1_U11.reset  ? 32'd0 : _277_;
assign _278_ = \shl_32s_32s_32_7_1_U11.ce  ? _279_ : \shl_32s_32s_32_7_1_U11.dout_array[0] ;
assign _261_ = \shl_32s_32s_32_7_1_U11.reset  ? 32'd0 : _278_;
assign _279_ = \shl_32s_32s_32_7_1_U11.din0  << { \shl_32s_32s_32_7_1_U11.din1 [31:30], 30'h00000000 };
assign _280_ = \shl_32s_32s_32_7_1_U11.dout_array[0]  << { \shl_32s_32s_32_7_1_U11.din1_cast_array[0] [29:25], 25'h0000000 };
assign _281_ = \shl_32s_32s_32_7_1_U11.dout_array[1]  << { \shl_32s_32s_32_7_1_U11.din1_cast_array[1] [24:20], 20'h00000 };
assign _282_ = \shl_32s_32s_32_7_1_U11.dout_array[2]  << { \shl_32s_32s_32_7_1_U11.din1_cast_array[2] [19:15], 15'h0000 };
assign _283_ = \shl_32s_32s_32_7_1_U11.dout_array[3]  << { \shl_32s_32s_32_7_1_U11.din1_cast_array[3] [14:10], 10'h000 };
assign _284_ = \shl_32s_32s_32_7_1_U11.dout_array[4]  << { \shl_32s_32s_32_7_1_U11.din1_cast_array[4] [9:5], 5'h00 };
assign \shl_32s_32s_32_7_1_U11.dout  = \shl_32s_32s_32_7_1_U11.dout_array[5]  << \shl_32s_32s_32_7_1_U11.din1_cast_array[5] [4:0];
assign \sub_4ns_4ns_4_2_1_U9.top_sub_4ns_4ns_4_2_1_Adder_8_U.bin_s0  = ~ \sub_4ns_4ns_4_2_1_U9.top_sub_4ns_4ns_4_2_1_Adder_8_U.b ;
always @(posedge \sub_4ns_4ns_4_2_1_U9.top_sub_4ns_4ns_4_2_1_Adder_8_U.clk )
\sub_4ns_4ns_4_2_1_U9.top_sub_4ns_4ns_4_2_1_Adder_8_U.bin_s1  <= _286_;
always @(posedge \sub_4ns_4ns_4_2_1_U9.top_sub_4ns_4ns_4_2_1_Adder_8_U.clk )
\sub_4ns_4ns_4_2_1_U9.top_sub_4ns_4ns_4_2_1_Adder_8_U.ain_s1  <= _285_;
always @(posedge \sub_4ns_4ns_4_2_1_U9.top_sub_4ns_4ns_4_2_1_Adder_8_U.clk )
\sub_4ns_4ns_4_2_1_U9.top_sub_4ns_4ns_4_2_1_Adder_8_U.sum_s1  <= _288_;
always @(posedge \sub_4ns_4ns_4_2_1_U9.top_sub_4ns_4ns_4_2_1_Adder_8_U.clk )
\sub_4ns_4ns_4_2_1_U9.top_sub_4ns_4ns_4_2_1_Adder_8_U.carry_s1  <= _287_;
assign _286_ = \sub_4ns_4ns_4_2_1_U9.top_sub_4ns_4ns_4_2_1_Adder_8_U.ce  ? \sub_4ns_4ns_4_2_1_U9.top_sub_4ns_4ns_4_2_1_Adder_8_U.bin_s0 [3:2] : \sub_4ns_4ns_4_2_1_U9.top_sub_4ns_4ns_4_2_1_Adder_8_U.bin_s1 ;
assign _285_ = \sub_4ns_4ns_4_2_1_U9.top_sub_4ns_4ns_4_2_1_Adder_8_U.ce  ? \sub_4ns_4ns_4_2_1_U9.top_sub_4ns_4ns_4_2_1_Adder_8_U.a [3:2] : \sub_4ns_4ns_4_2_1_U9.top_sub_4ns_4ns_4_2_1_Adder_8_U.ain_s1 ;
assign _287_ = \sub_4ns_4ns_4_2_1_U9.top_sub_4ns_4ns_4_2_1_Adder_8_U.ce  ? \sub_4ns_4ns_4_2_1_U9.top_sub_4ns_4ns_4_2_1_Adder_8_U.facout_s1  : \sub_4ns_4ns_4_2_1_U9.top_sub_4ns_4ns_4_2_1_Adder_8_U.carry_s1 ;
assign _288_ = \sub_4ns_4ns_4_2_1_U9.top_sub_4ns_4ns_4_2_1_Adder_8_U.ce  ? \sub_4ns_4ns_4_2_1_U9.top_sub_4ns_4ns_4_2_1_Adder_8_U.fas_s1  : \sub_4ns_4ns_4_2_1_U9.top_sub_4ns_4ns_4_2_1_Adder_8_U.sum_s1 ;
assign _289_ = \sub_4ns_4ns_4_2_1_U9.top_sub_4ns_4ns_4_2_1_Adder_8_U.u1.a  + \sub_4ns_4ns_4_2_1_U9.top_sub_4ns_4ns_4_2_1_Adder_8_U.u1.b ;
assign { \sub_4ns_4ns_4_2_1_U9.top_sub_4ns_4ns_4_2_1_Adder_8_U.u1.cout , \sub_4ns_4ns_4_2_1_U9.top_sub_4ns_4ns_4_2_1_Adder_8_U.u1.s  } = _289_ + \sub_4ns_4ns_4_2_1_U9.top_sub_4ns_4ns_4_2_1_Adder_8_U.u1.cin ;
assign _290_ = \sub_4ns_4ns_4_2_1_U9.top_sub_4ns_4ns_4_2_1_Adder_8_U.u2.a  + \sub_4ns_4ns_4_2_1_U9.top_sub_4ns_4ns_4_2_1_Adder_8_U.u2.b ;
assign { \sub_4ns_4ns_4_2_1_U9.top_sub_4ns_4ns_4_2_1_Adder_8_U.u2.cout , \sub_4ns_4ns_4_2_1_U9.top_sub_4ns_4ns_4_2_1_Adder_8_U.u2.s  } = _290_ + \sub_4ns_4ns_4_2_1_U9.top_sub_4ns_4ns_4_2_1_Adder_8_U.u2.cin ;
assign \sub_9ns_9s_9_2_1_U7.top_sub_9ns_9s_9_2_1_Adder_6_U.bin_s0  = ~ \sub_9ns_9s_9_2_1_U7.top_sub_9ns_9s_9_2_1_Adder_6_U.b ;
always @(posedge \sub_9ns_9s_9_2_1_U7.top_sub_9ns_9s_9_2_1_Adder_6_U.clk )
\sub_9ns_9s_9_2_1_U7.top_sub_9ns_9s_9_2_1_Adder_6_U.bin_s1  <= _292_;
always @(posedge \sub_9ns_9s_9_2_1_U7.top_sub_9ns_9s_9_2_1_Adder_6_U.clk )
\sub_9ns_9s_9_2_1_U7.top_sub_9ns_9s_9_2_1_Adder_6_U.ain_s1  <= _291_;
always @(posedge \sub_9ns_9s_9_2_1_U7.top_sub_9ns_9s_9_2_1_Adder_6_U.clk )
\sub_9ns_9s_9_2_1_U7.top_sub_9ns_9s_9_2_1_Adder_6_U.sum_s1  <= _294_;
always @(posedge \sub_9ns_9s_9_2_1_U7.top_sub_9ns_9s_9_2_1_Adder_6_U.clk )
\sub_9ns_9s_9_2_1_U7.top_sub_9ns_9s_9_2_1_Adder_6_U.carry_s1  <= _293_;
assign _292_ = \sub_9ns_9s_9_2_1_U7.top_sub_9ns_9s_9_2_1_Adder_6_U.ce  ? \sub_9ns_9s_9_2_1_U7.top_sub_9ns_9s_9_2_1_Adder_6_U.bin_s0 [8:4] : \sub_9ns_9s_9_2_1_U7.top_sub_9ns_9s_9_2_1_Adder_6_U.bin_s1 ;
assign _291_ = \sub_9ns_9s_9_2_1_U7.top_sub_9ns_9s_9_2_1_Adder_6_U.ce  ? \sub_9ns_9s_9_2_1_U7.top_sub_9ns_9s_9_2_1_Adder_6_U.a [8:4] : \sub_9ns_9s_9_2_1_U7.top_sub_9ns_9s_9_2_1_Adder_6_U.ain_s1 ;
assign _293_ = \sub_9ns_9s_9_2_1_U7.top_sub_9ns_9s_9_2_1_Adder_6_U.ce  ? \sub_9ns_9s_9_2_1_U7.top_sub_9ns_9s_9_2_1_Adder_6_U.facout_s1  : \sub_9ns_9s_9_2_1_U7.top_sub_9ns_9s_9_2_1_Adder_6_U.carry_s1 ;
assign _294_ = \sub_9ns_9s_9_2_1_U7.top_sub_9ns_9s_9_2_1_Adder_6_U.ce  ? \sub_9ns_9s_9_2_1_U7.top_sub_9ns_9s_9_2_1_Adder_6_U.fas_s1  : \sub_9ns_9s_9_2_1_U7.top_sub_9ns_9s_9_2_1_Adder_6_U.sum_s1 ;
assign _295_ = \sub_9ns_9s_9_2_1_U7.top_sub_9ns_9s_9_2_1_Adder_6_U.u1.a  + \sub_9ns_9s_9_2_1_U7.top_sub_9ns_9s_9_2_1_Adder_6_U.u1.b ;
assign { \sub_9ns_9s_9_2_1_U7.top_sub_9ns_9s_9_2_1_Adder_6_U.u1.cout , \sub_9ns_9s_9_2_1_U7.top_sub_9ns_9s_9_2_1_Adder_6_U.u1.s  } = _295_ + \sub_9ns_9s_9_2_1_U7.top_sub_9ns_9s_9_2_1_Adder_6_U.u1.cin ;
assign _296_ = \sub_9ns_9s_9_2_1_U7.top_sub_9ns_9s_9_2_1_Adder_6_U.u2.a  + \sub_9ns_9s_9_2_1_U7.top_sub_9ns_9s_9_2_1_Adder_6_U.u2.b ;
assign { \sub_9ns_9s_9_2_1_U7.top_sub_9ns_9s_9_2_1_Adder_6_U.u2.cout , \sub_9ns_9s_9_2_1_U7.top_sub_9ns_9s_9_2_1_Adder_6_U.u2.s  } = _296_ + \sub_9ns_9s_9_2_1_U7.top_sub_9ns_9s_9_2_1_Adder_6_U.u2.cin ;
assign _297_ = | trunc_ln851_reg_1000;
assign _298_ = | op_10[2:0];
assign _299_ = | op_12[12:0];
assign _300_ = | op_13[11:0];
assign _301_ = | op_14[1:0];
always @(posedge ap_clk)
trunc_ln851_reg_1000 <= 6'h00;
always @(posedge ap_clk)
sub_ln1357_reg_946 <= _048_;
always @(posedge ap_clk)
shl_ln781_reg_1121 <= _047_;
always @(posedge ap_clk)
shl_ln1299_reg_1084 <= _046_;
always @(posedge ap_clk)
sext_ln850_reg_854 <= _044_;
always @(posedge ap_clk)
sext_ln15_reg_935 <= _043_;
always @(posedge ap_clk)
select_ln353_reg_941 <= _041_;
always @(posedge ap_clk)
select_ln353_1_reg_1042 <= _039_;
always @(posedge ap_clk)
select_ln69_reg_1047 <= _042_;
always @(posedge ap_clk)
select_ln1358_reg_1094 <= _038_;
always @(posedge ap_clk)
ret_V_reg_1099 <= _037_;
always @(posedge ap_clk)
trunc_ln851_1_reg_1106 <= _051_;
always @(posedge ap_clk)
select_ln353_2_reg_1111 <= _040_;
always @(posedge ap_clk)
ret_V_4_reg_1168 <= _036_;
always @(posedge ap_clk)
ret_V_18_reg_1067 <= _028_;
always @(posedge ap_clk)
ret_V_25_cast_reg_1072 <= _033_;
always @(posedge ap_clk)
ush_reg_966 <= _052_;
always @(posedge ap_clk)
ret_V_17_reg_971 <= _027_;
always @(posedge ap_clk)
ret_V_23_cast_reg_976 <= _032_;
always @(posedge ap_clk)
ret_V_16_reg_907 <= _026_;
always @(posedge ap_clk)
ret_V_21_cast_reg_912 <= _031_;
always @(posedge ap_clk)
ret_V_14_reg_844 <= _024_;
always @(posedge ap_clk)
tmp_1_reg_849 <= _049_;
always @(posedge ap_clk)
r_reg_919 <= _022_;
always @(posedge ap_clk)
tmp_3_reg_924 <= _050_;
always @(posedge ap_clk)
r_1_reg_1146 <= _021_;
always @(posedge ap_clk)
ret_V_3_reg_1151 <= _035_;
always @(posedge ap_clk)
ret_V_19_reg_1156 <= _029_;
always @(posedge ap_clk)
ret_V_27_cast_reg_1161 <= _034_;
always @(posedge ap_clk)
p_Result_7_reg_989 <= _020_;
always @(posedge ap_clk)
_784_ <= _023_;
assign ret_V_12_reg_994[9:6] = _784_;
always @(posedge ap_clk)
op_23_V_reg_887 <= _019_;
always @(posedge ap_clk)
op_21_V_reg_824 <= _018_;
always @(posedge ap_clk)
op_11_V_reg_872 <= _017_;
always @(posedge ap_clk)
ret_V_15_reg_877 <= _025_;
always @(posedge ap_clk)
icmp_ln851_reg_1131 <= _016_;
always @(posedge ap_clk)
icmp_ln851_4_reg_1062 <= _015_;
always @(posedge ap_clk)
icmp_ln851_3_reg_961 <= _014_;
always @(posedge ap_clk)
icmp_ln851_2_reg_902 <= _013_;
always @(posedge ap_clk)
icmp_ln851_1_reg_839 <= _012_;
always @(posedge ap_clk)
sh_reg_1017 <= _045_;
always @(posedge ap_clk)
icmp_ln850_reg_1022 <= _011_;
always @(posedge ap_clk)
ashr_ln799_reg_1126 <= _010_;
always @(posedge ap_clk)
ashr_ln1333_reg_1079 <= _009_;
always @(posedge ap_clk)
add_ln69_reg_1208 <= _007_;
always @(posedge ap_clk)
add_ln69_2_reg_1213 <= _006_;
always @(posedge ap_clk)
ret_V_20_reg_1183 <= _030_;
always @(posedge ap_clk)
add_ln69_1_reg_1188 <= _005_;
always @(posedge ap_clk)
add_ln691_reg_861 <= _004_;
always @(posedge ap_clk)
add_ln691_4_reg_1173 <= _003_;
always @(posedge ap_clk)
add_ln691_3_reg_1089 <= _002_;
always @(posedge ap_clk)
add_ln691_2_reg_1027 <= _001_;
always @(posedge ap_clk)
add_ln691_1_reg_930 <= _000_;
always @(posedge ap_clk)
ap_CS_fsm <= _008_;
assign _053_ = _064_ ? 2'h2 : 2'h1;
assign _302_ = ap_CS_fsm == 1'h1;
function [32:0] _810_;
input [32:0] a;
input [1088:0] b;
input [32:0] s;
case (s)
33'b000000000000000000000000000000001:
_810_ = b[32:0];
33'b000000000000000000000000000000010:
_810_ = b[65:33];
33'b000000000000000000000000000000100:
_810_ = b[98:66];
33'b000000000000000000000000000001000:
_810_ = b[131:99];
33'b000000000000000000000000000010000:
_810_ = b[164:132];
33'b000000000000000000000000000100000:
_810_ = b[197:165];
33'b000000000000000000000000001000000:
_810_ = b[230:198];
33'b000000000000000000000000010000000:
_810_ = b[263:231];
33'b000000000000000000000000100000000:
_810_ = b[296:264];
33'b000000000000000000000001000000000:
_810_ = b[329:297];
33'b000000000000000000000010000000000:
_810_ = b[362:330];
33'b000000000000000000000100000000000:
_810_ = b[395:363];
33'b000000000000000000001000000000000:
_810_ = b[428:396];
33'b000000000000000000010000000000000:
_810_ = b[461:429];
33'b000000000000000000100000000000000:
_810_ = b[494:462];
33'b000000000000000001000000000000000:
_810_ = b[527:495];
33'b000000000000000010000000000000000:
_810_ = b[560:528];
33'b000000000000000100000000000000000:
_810_ = b[593:561];
33'b000000000000001000000000000000000:
_810_ = b[626:594];
33'b000000000000010000000000000000000:
_810_ = b[659:627];
33'b000000000000100000000000000000000:
_810_ = b[692:660];
33'b000000000001000000000000000000000:
_810_ = b[725:693];
33'b000000000010000000000000000000000:
_810_ = b[758:726];
33'b000000000100000000000000000000000:
_810_ = b[791:759];
33'b000000001000000000000000000000000:
_810_ = b[824:792];
33'b000000010000000000000000000000000:
_810_ = b[857:825];
33'b000000100000000000000000000000000:
_810_ = b[890:858];
33'b000001000000000000000000000000000:
_810_ = b[923:891];
33'b000010000000000000000000000000000:
_810_ = b[956:924];
33'b000100000000000000000000000000000:
_810_ = b[989:957];
33'b001000000000000000000000000000000:
_810_ = b[1022:990];
33'b010000000000000000000000000000000:
_810_ = b[1055:1023];
33'b100000000000000000000000000000000:
_810_ = b[1088:1056];
33'b000000000000000000000000000000000:
_810_ = a;
default:
_810_ = 33'bx;
endcase
endfunction
assign ap_NS_fsm = _810_(33'hxxxxxxxxx, { 31'h00000000, _053_, 1056'h000000020000000200000002000000020000000200000002000000020000000200000002000000020000000200000002000000020000000200000002000000020000000200000002000000020000000200000002000000020000000200000002000000020000000200000002000000020000000200000002000000020000000000000001 }, { _302_, _334_, _333_, _332_, _331_, _330_, _329_, _328_, _327_, _326_, _325_, _324_, _323_, _322_, _321_, _320_, _319_, _318_, _317_, _316_, _315_, _314_, _313_, _312_, _311_, _310_, _309_, _308_, _307_, _306_, _305_, _304_, _303_ });
assign _303_ = ap_CS_fsm == 33'h100000000;
assign _304_ = ap_CS_fsm == 32'd2147483648;
assign _305_ = ap_CS_fsm == 31'h40000000;
assign _306_ = ap_CS_fsm == 30'h20000000;
assign _307_ = ap_CS_fsm == 29'h10000000;
assign _308_ = ap_CS_fsm == 28'h8000000;
assign _309_ = ap_CS_fsm == 27'h4000000;
assign _310_ = ap_CS_fsm == 26'h2000000;
assign _311_ = ap_CS_fsm == 25'h1000000;
assign _312_ = ap_CS_fsm == 24'h800000;
assign _313_ = ap_CS_fsm == 23'h400000;
assign _314_ = ap_CS_fsm == 22'h200000;
assign _315_ = ap_CS_fsm == 21'h100000;
assign _316_ = ap_CS_fsm == 20'h80000;
assign _317_ = ap_CS_fsm == 19'h40000;
assign _318_ = ap_CS_fsm == 18'h20000;
assign _319_ = ap_CS_fsm == 17'h10000;
assign _320_ = ap_CS_fsm == 16'h8000;
assign _321_ = ap_CS_fsm == 15'h4000;
assign _322_ = ap_CS_fsm == 14'h2000;
assign _323_ = ap_CS_fsm == 13'h1000;
assign _324_ = ap_CS_fsm == 12'h800;
assign _325_ = ap_CS_fsm == 11'h400;
assign _326_ = ap_CS_fsm == 10'h200;
assign _327_ = ap_CS_fsm == 9'h100;
assign _328_ = ap_CS_fsm == 8'h80;
assign _329_ = ap_CS_fsm == 7'h40;
assign _330_ = ap_CS_fsm == 6'h20;
assign _331_ = ap_CS_fsm == 5'h10;
assign _332_ = ap_CS_fsm == 4'h8;
assign _333_ = ap_CS_fsm == 3'h4;
assign _334_ = ap_CS_fsm == 2'h2;
assign op_31_ap_vld = ap_CS_fsm[32] ? 1'h1 : 1'h0;
assign ap_idle = _063_ ? 1'h1 : 1'h0;
assign _048_ = _062_ ? grp_fu_399_p2 : sub_ln1357_reg_946;
assign _047_ = _061_ ? grp_fu_538_p2 : shl_ln781_reg_1121;
assign _046_ = _060_ ? grp_fu_519_p2 : shl_ln1299_reg_1084;
assign _044_ = ap_CS_fsm[4] ? { tmp_1_reg_849[8], tmp_1_reg_849 } : sext_ln850_reg_854;
assign _041_ = ap_CS_fsm[13] ? select_ln353_fu_417_p3 : select_ln353_reg_941;
assign _043_ = ap_CS_fsm[13] ? { r_reg_919[7], r_reg_919 } : sext_ln15_reg_935;
assign _042_ = ap_CS_fsm[18] ? select_ln69_fu_595_p3 : select_ln69_reg_1047;
assign _039_ = ap_CS_fsm[18] ? select_ln353_1_fu_588_p3 : select_ln353_1_reg_1042;
assign _040_ = ap_CS_fsm[23] ? select_ln353_2_fu_680_p3 : select_ln353_2_reg_1111;
assign _051_ = ap_CS_fsm[23] ? select_ln1358_fu_649_p3[5:0] : trunc_ln851_1_reg_1106;
assign _037_ = ap_CS_fsm[23] ? select_ln1358_fu_649_p3[7:6] : ret_V_reg_1099;
assign _038_ = ap_CS_fsm[23] ? select_ln1358_fu_649_p3 : select_ln1358_reg_1094;
assign _036_ = ap_CS_fsm[26] ? ret_V_4_fu_745_p3 : ret_V_4_reg_1168;
assign _033_ = ap_CS_fsm[20] ? grp_fu_618_p2[33:2] : ret_V_25_cast_reg_1072;
assign _028_ = ap_CS_fsm[20] ? grp_fu_618_p2 : ret_V_18_reg_1067;
assign _032_ = ap_CS_fsm[15] ? grp_fu_439_p2[43:12] : ret_V_23_cast_reg_976;
assign _027_ = ap_CS_fsm[15] ? grp_fu_439_p2 : ret_V_17_reg_971;
assign _052_ = ap_CS_fsm[15] ? ush_fu_455_p3 : ush_reg_966;
assign _031_ = ap_CS_fsm[10] ? grp_fu_351_p2[44:13] : ret_V_21_cast_reg_912;
assign _026_ = ap_CS_fsm[10] ? grp_fu_351_p2 : ret_V_16_reg_907;
assign _049_ = ap_CS_fsm[3] ? grp_fu_260_p2[11:3] : tmp_1_reg_849;
assign _024_ = ap_CS_fsm[3] ? grp_fu_260_p2 : ret_V_14_reg_844;
assign _050_ = ap_CS_fsm[12] ? op_3[7] : tmp_3_reg_924;
assign _022_ = ap_CS_fsm[12] ? r_fu_382_p2 : r_reg_919;
assign _034_ = ap_CS_fsm[25] ? grp_fu_712_p2[32:1] : ret_V_27_cast_reg_1161;
assign _029_ = ap_CS_fsm[25] ? grp_fu_712_p2 : ret_V_19_reg_1156;
assign _035_ = ap_CS_fsm[25] ? grp_fu_692_p2 : ret_V_3_reg_1151;
assign _021_ = ap_CS_fsm[25] ? r_1_fu_718_p3 : r_1_reg_1146;
assign _023_ = ap_CS_fsm[16] ? ret_V_12_fu_496_p2[9:6] : ret_V_12_reg_994[9:6];
assign _020_ = ap_CS_fsm[16] ? op_6[3] : p_Result_7_reg_989;
assign _019_ = ap_CS_fsm[8] ? grp_fu_331_p2 : op_23_V_reg_887;
assign _018_ = ap_CS_fsm[1] ? grp_fu_243_p2 : op_21_V_reg_824;
assign _025_ = ap_CS_fsm[6] ? ret_V_15_fu_321_p3 : ret_V_15_reg_877;
assign _017_ = ap_CS_fsm[6] ? op_11_V_fu_303_p2 : op_11_V_reg_872;
assign _016_ = ap_CS_fsm[24] ? icmp_ln851_fu_687_p2 : icmp_ln851_reg_1131;
assign _015_ = ap_CS_fsm[19] ? icmp_ln851_4_fu_628_p2 : icmp_ln851_4_reg_1062;
assign _014_ = ap_CS_fsm[14] ? icmp_ln851_3_fu_449_p2 : icmp_ln851_3_reg_961;
assign _013_ = ap_CS_fsm[9] ? icmp_ln851_2_fu_361_p2 : icmp_ln851_2_reg_902;
assign _012_ = ap_CS_fsm[2] ? icmp_ln851_1_fu_270_p2 : icmp_ln851_1_reg_839;
assign _011_ = ap_CS_fsm[17] ? icmp_ln850_fu_530_p2 : icmp_ln850_reg_1022;
assign _045_ = ap_CS_fsm[17] ? grp_fu_478_p2 : sh_reg_1017;
assign _010_ = _059_ ? grp_fu_546_p2 : ashr_ln799_reg_1126;
assign _009_ = _058_ ? grp_fu_513_p2 : ashr_ln1333_reg_1079;
assign _006_ = ap_CS_fsm[30] ? grp_fu_799_p2 : add_ln69_2_reg_1213;
assign _007_ = ap_CS_fsm[30] ? grp_fu_791_p2 : add_ln69_reg_1208;
assign _005_ = ap_CS_fsm[28] ? grp_fu_760_p2 : add_ln69_1_reg_1188;
assign _030_ = ap_CS_fsm[28] ? ret_V_20_fu_781_p3 : ret_V_20_reg_1183;
assign _004_ = _057_ ? grp_fu_289_p2 : add_ln691_reg_861;
assign _003_ = ap_CS_fsm[27] ? grp_fu_752_p2 : add_ln691_4_reg_1173;
assign _002_ = _056_ ? grp_fu_644_p2 : add_ln691_3_reg_1089;
assign _001_ = _055_ ? grp_fu_525_p2 : add_ln691_2_reg_1027;
assign _000_ = _054_ ? grp_fu_377_p2 : add_ln691_1_reg_930;
assign _008_ = ap_rst ? 33'h000000001 : ap_NS_fsm;
assign icmp_ln850_fu_530_p2 = _297_ ? 1'h1 : 1'h0;
assign icmp_ln851_1_fu_270_p2 = _298_ ? 1'h1 : 1'h0;
assign icmp_ln851_2_fu_361_p2 = _299_ ? 1'h1 : 1'h0;
assign icmp_ln851_3_fu_449_p2 = _300_ ? 1'h1 : 1'h0;
assign icmp_ln851_4_fu_628_p2 = _301_ ? 1'h1 : 1'h0;
assign icmp_ln851_fu_687_p2 = _068_ ? 1'h1 : 1'h0;
assign r_1_fu_718_p3 = p_Result_7_reg_989 ? shl_ln781_reg_1121 : ashr_ln799_reg_1126;
assign ret_V_15_fu_321_p3 = ret_V_14_reg_844[11] ? select_ln850_2_fu_316_p3 : sext_ln850_reg_854;
assign ret_V_20_fu_781_p3 = ret_V_19_reg_1156[33] ? select_ln850_6_fu_775_p3 : ret_V_27_cast_reg_1161;
assign ret_V_4_fu_745_p3 = select_ln1358_reg_1094[7] ? select_ln850_fu_740_p3 : ret_V_reg_1099;
assign select_ln1358_fu_649_p3 = tmp_3_reg_924 ? shl_ln1299_reg_1084 : ashr_ln1333_reg_1079;
assign select_ln353_1_fu_588_p3 = ret_V_17_reg_971[44] ? select_ln850_4_fu_583_p3 : ret_V_23_cast_reg_976;
assign select_ln353_2_fu_680_p3 = ret_V_18_reg_1067[34] ? select_ln850_5_fu_675_p3 : ret_V_25_cast_reg_1072;
assign select_ln353_fu_417_p3 = ret_V_16_reg_907[45] ? select_ln850_3_fu_412_p3 : ret_V_21_cast_reg_912;
assign select_ln69_fu_595_p3 = ret_V_13_fu_570_p2 ? 3'h7 : 3'h0;
assign select_ln850_2_fu_316_p3 = icmp_ln851_1_reg_839 ? add_ln691_reg_861 : sext_ln850_reg_854;
assign select_ln850_3_fu_412_p3 = icmp_ln851_2_reg_902 ? add_ln691_1_reg_930 : ret_V_21_cast_reg_912;
assign select_ln850_4_fu_583_p3 = icmp_ln851_3_reg_961 ? add_ln691_2_reg_1027 : ret_V_23_cast_reg_976;
assign select_ln850_5_fu_675_p3 = icmp_ln851_4_reg_1062 ? add_ln691_3_reg_1089 : ret_V_25_cast_reg_1072;
assign select_ln850_6_fu_775_p3 = op_15[0] ? add_ln691_4_reg_1173 : ret_V_27_cast_reg_1161;
assign select_ln850_fu_740_p3 = icmp_ln851_reg_1131 ? ret_V_reg_1099 : ret_V_3_reg_1151;
assign ush_fu_455_p3 = tmp_3_reg_924 ? sext_ln15_reg_935 : sub_ln1357_reg_946;
assign op_11_V_fu_303_p2 = op_2[3:0] ^ op_4[3:0];
assign ret_V_13_fu_570_p2 = ret_V_12_reg_994[6] ^ and_ln353_fu_565_p2;
assign ap_CS_fsm_state1 = ap_CS_fsm[0];
assign ap_CS_fsm_state10 = ap_CS_fsm[9];
assign ap_CS_fsm_state11 = ap_CS_fsm[10];
assign ap_CS_fsm_state12 = ap_CS_fsm[11];
assign ap_CS_fsm_state13 = ap_CS_fsm[12];
assign ap_CS_fsm_state14 = ap_CS_fsm[13];
assign ap_CS_fsm_state15 = ap_CS_fsm[14];
assign ap_CS_fsm_state16 = ap_CS_fsm[15];
assign ap_CS_fsm_state17 = ap_CS_fsm[16];
assign ap_CS_fsm_state18 = ap_CS_fsm[17];
assign ap_CS_fsm_state19 = ap_CS_fsm[18];
assign ap_CS_fsm_state2 = ap_CS_fsm[1];
assign ap_CS_fsm_state20 = ap_CS_fsm[19];
assign ap_CS_fsm_state21 = ap_CS_fsm[20];
assign ap_CS_fsm_state22 = ap_CS_fsm[21];
assign ap_CS_fsm_state23 = ap_CS_fsm[22];
assign ap_CS_fsm_state24 = ap_CS_fsm[23];
assign ap_CS_fsm_state25 = ap_CS_fsm[24];
assign ap_CS_fsm_state26 = ap_CS_fsm[25];
assign ap_CS_fsm_state27 = ap_CS_fsm[26];
assign ap_CS_fsm_state28 = ap_CS_fsm[27];
assign ap_CS_fsm_state29 = ap_CS_fsm[28];
assign ap_CS_fsm_state3 = ap_CS_fsm[2];
assign ap_CS_fsm_state30 = ap_CS_fsm[29];
assign ap_CS_fsm_state31 = ap_CS_fsm[30];
assign ap_CS_fsm_state32 = ap_CS_fsm[31];
assign ap_CS_fsm_state33 = ap_CS_fsm[32];
assign ap_CS_fsm_state4 = ap_CS_fsm[3];
assign ap_CS_fsm_state5 = ap_CS_fsm[4];
assign ap_CS_fsm_state6 = ap_CS_fsm[5];
assign ap_CS_fsm_state7 = ap_CS_fsm[6];
assign ap_CS_fsm_state8 = ap_CS_fsm[7];
assign ap_CS_fsm_state9 = ap_CS_fsm[8];
assign ap_done = op_31_ap_vld;
assign ap_ready = op_31_ap_vld;
assign conv_i_i_i357_fu_509_p0 = op_7;
assign conv_i_i_i357_fu_509_p1 = { op_7[7], op_7[7], op_7[7], op_7[7], op_7[7], op_7[7], op_7[7], op_7[7], op_7[7], op_7[7], op_7[7], op_7[7], op_7[7], op_7[7], op_7[7], op_7[7], op_7[7], op_7[7], op_7[7], op_7[7], op_7[7], op_7[7], op_7[7], op_7[7], op_7 };
assign grp_fu_243_p0 = { op_5[7], op_5 };
assign grp_fu_243_p1 = { op_8[3], op_8[3], op_8[3], op_8[3], op_8[3], op_8 };
assign grp_fu_260_p0 = { op_21_V_reg_824, 3'h0 };
assign grp_fu_260_p1 = { op_10[3], op_10[3], op_10[3], op_10[3], op_10[3], op_10[3], op_10[3], op_10[3], op_10 };
assign grp_fu_289_p0 = { tmp_1_reg_849[8], tmp_1_reg_849 };
assign grp_fu_331_p1 = { op_11_V_reg_872[3], op_11_V_reg_872[3], op_11_V_reg_872[3], op_11_V_reg_872[3], op_11_V_reg_872[3], op_11_V_reg_872[3], op_11_V_reg_872 };
assign grp_fu_351_p0 = { op_23_V_reg_887[9], op_23_V_reg_887[9], op_23_V_reg_887[9], op_23_V_reg_887[9], op_23_V_reg_887[9], op_23_V_reg_887[9], op_23_V_reg_887[9], op_23_V_reg_887[9], op_23_V_reg_887[9], op_23_V_reg_887[9], op_23_V_reg_887[9], op_23_V_reg_887[9], op_23_V_reg_887[9], op_23_V_reg_887[9], op_23_V_reg_887[9], op_23_V_reg_887[9], op_23_V_reg_887[9], op_23_V_reg_887[9], op_23_V_reg_887[9], op_23_V_reg_887[9], op_23_V_reg_887[9], op_23_V_reg_887[9], op_23_V_reg_887[9], op_23_V_reg_887, 13'h0000 };
assign grp_fu_351_p1 = { op_12[15], op_12[15], op_12[15], op_12[15], op_12[15], op_12[15], op_12[15], op_12[15], op_12[15], op_12[15], op_12[15], op_12[15], op_12[15], op_12[15], op_12[15], op_12[15], op_12[15], op_12[15], op_12[15], op_12[15], op_12[15], op_12[15], op_12[15], op_12[15], op_12[15], op_12[15], op_12[15], op_12[15], op_12[15], op_12[15], op_12 };
assign grp_fu_399_p1 = { r_reg_919[7], r_reg_919 };
assign grp_fu_439_p0 = { select_ln353_reg_941[31], select_ln353_reg_941, 12'h000 };
assign grp_fu_439_p1 = { op_13[15], op_13[15], op_13[15], op_13[15], op_13[15], op_13[15], op_13[15], op_13[15], op_13[15], op_13[15], op_13[15], op_13[15], op_13[15], op_13[15], op_13[15], op_13[15], op_13[15], op_13[15], op_13[15], op_13[15], op_13[15], op_13[15], op_13[15], op_13[15], op_13[15], op_13[15], op_13[15], op_13[15], op_13[15], op_13 };
assign grp_fu_538_p1 = { 12'h000, sh_reg_1017 };
assign grp_fu_546_p1 = { 12'h000, op_6 };
assign grp_fu_618_p0 = { select_ln353_1_reg_1042[31], select_ln353_1_reg_1042, 2'h0 };
assign grp_fu_618_p1 = { op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14 };
assign grp_fu_712_p0 = { select_ln353_2_reg_1111[31], select_ln353_2_reg_1111, 1'h0 };
assign grp_fu_712_p1 = { op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15 };
assign grp_fu_760_p0 = { ret_V_4_reg_1168[1], ret_V_4_reg_1168 };
assign grp_fu_799_p0 = { add_ln69_1_reg_1188[2], add_ln69_1_reg_1188[2], add_ln69_1_reg_1188[2], add_ln69_1_reg_1188[2], add_ln69_1_reg_1188[2], add_ln69_1_reg_1188[2], add_ln69_1_reg_1188[2], add_ln69_1_reg_1188[2], add_ln69_1_reg_1188[2], add_ln69_1_reg_1188[2], add_ln69_1_reg_1188[2], add_ln69_1_reg_1188[2], add_ln69_1_reg_1188[2], add_ln69_1_reg_1188[2], add_ln69_1_reg_1188 };
assign grp_fu_799_p1 = { r_1_reg_1146[15], r_1_reg_1146 };
assign grp_fu_808_p0 = { add_ln69_2_reg_1213[16], add_ln69_2_reg_1213[16], add_ln69_2_reg_1213[16], add_ln69_2_reg_1213[16], add_ln69_2_reg_1213[16], add_ln69_2_reg_1213[16], add_ln69_2_reg_1213[16], add_ln69_2_reg_1213[16], add_ln69_2_reg_1213[16], add_ln69_2_reg_1213[16], add_ln69_2_reg_1213[16], add_ln69_2_reg_1213[16], add_ln69_2_reg_1213[16], add_ln69_2_reg_1213[16], add_ln69_2_reg_1213[16], add_ln69_2_reg_1213 };
assign lhs_fu_484_p3 = { op_6, 6'h00 };
assign op_31 = grp_fu_808_p2;
assign p_Result_1_fu_733_p3 = select_ln1358_reg_1094[7];
assign p_Result_2_fu_309_p3 = ret_V_14_reg_844[11];
assign p_Result_3_fu_405_p3 = ret_V_16_reg_907[45];
assign p_Result_4_fu_576_p3 = ret_V_17_reg_971[44];
assign p_Result_5_fu_668_p3 = ret_V_18_reg_1067[34];
assign p_Result_6_fu_765_p3 = ret_V_19_reg_1156[33];
assign p_Result_s_fu_558_p3 = ret_V_12_reg_994[9];
assign rhs_3_fu_428_p3 = { select_ln353_reg_941, 12'h000 };
assign rhs_4_fu_607_p3 = { select_ln353_1_reg_1042, 2'h0 };
assign rhs_5_fu_701_p3 = { select_ln353_2_reg_1111, 1'h0 };
assign sext_ln1192_fu_249_p0 = op_10;
assign sext_ln1357_fu_506_p1 = { ush_reg_966[8], ush_reg_966[8], ush_reg_966[8], ush_reg_966[8], ush_reg_966[8], ush_reg_966[8], ush_reg_966[8], ush_reg_966[8], ush_reg_966[8], ush_reg_966[8], ush_reg_966[8], ush_reg_966[8], ush_reg_966[8], ush_reg_966[8], ush_reg_966[8], ush_reg_966[8], ush_reg_966[8], ush_reg_966[8], ush_reg_966[8], ush_reg_966[8], ush_reg_966[8], ush_reg_966[8], ush_reg_966[8], ush_reg_966 };
assign sext_ln15_fu_396_p1 = { r_reg_919[7], r_reg_919 };
assign sext_ln703_1_fu_336_p0 = op_12;
assign sext_ln703_2_fu_424_p0 = op_13;
assign sext_ln703_3_fu_603_p0 = op_14;
assign sext_ln703_4_fu_697_p0 = op_15;
assign sext_ln703_fu_492_p0 = op_7;
assign sext_ln703_fu_492_p1 = { op_7[7], op_7[7], op_7 };
assign sext_ln850_fu_286_p1 = { tmp_1_reg_849[8], tmp_1_reg_849 };
assign tmp_6_fu_340_p3 = { op_23_V_reg_887, 13'h0000 };
assign tmp_fu_551_p3 = ret_V_12_reg_994[6];
assign trunc_ln1350_1_fu_299_p1 = op_4[3:0];
assign trunc_ln1350_fu_295_p1 = op_2[3:0];
assign trunc_ln851_1_fu_664_p1 = select_ln1358_fu_649_p3[5:0];
assign trunc_ln851_2_fu_266_p0 = op_10;
assign trunc_ln851_2_fu_266_p1 = op_10[2:0];
assign trunc_ln851_3_fu_357_p0 = op_12;
assign trunc_ln851_3_fu_357_p1 = op_12[12:0];
assign trunc_ln851_4_fu_445_p0 = op_13;
assign trunc_ln851_4_fu_445_p1 = op_13[11:0];
assign trunc_ln851_5_fu_624_p0 = op_14;
assign trunc_ln851_5_fu_624_p1 = op_14[1:0];
assign trunc_ln851_6_fu_772_p0 = op_15;
assign trunc_ln851_6_fu_772_p1 = op_15[0];
assign trunc_ln851_fu_502_p1 = ret_V_12_fu_496_p2[5:0];
assign \sub_9ns_9s_9_2_1_U7.top_sub_9ns_9s_9_2_1_Adder_6_U.ain_s0  = \sub_9ns_9s_9_2_1_U7.top_sub_9ns_9s_9_2_1_Adder_6_U.a ;
assign \sub_9ns_9s_9_2_1_U7.top_sub_9ns_9s_9_2_1_Adder_6_U.s  = { \sub_9ns_9s_9_2_1_U7.top_sub_9ns_9s_9_2_1_Adder_6_U.fas_s2 , \sub_9ns_9s_9_2_1_U7.top_sub_9ns_9s_9_2_1_Adder_6_U.sum_s1  };
assign \sub_9ns_9s_9_2_1_U7.top_sub_9ns_9s_9_2_1_Adder_6_U.u2.a  = \sub_9ns_9s_9_2_1_U7.top_sub_9ns_9s_9_2_1_Adder_6_U.ain_s1 ;
assign \sub_9ns_9s_9_2_1_U7.top_sub_9ns_9s_9_2_1_Adder_6_U.u2.b  = \sub_9ns_9s_9_2_1_U7.top_sub_9ns_9s_9_2_1_Adder_6_U.bin_s1 ;
assign \sub_9ns_9s_9_2_1_U7.top_sub_9ns_9s_9_2_1_Adder_6_U.u2.cin  = \sub_9ns_9s_9_2_1_U7.top_sub_9ns_9s_9_2_1_Adder_6_U.carry_s1 ;
assign \sub_9ns_9s_9_2_1_U7.top_sub_9ns_9s_9_2_1_Adder_6_U.facout_s2  = \sub_9ns_9s_9_2_1_U7.top_sub_9ns_9s_9_2_1_Adder_6_U.u2.cout ;
assign \sub_9ns_9s_9_2_1_U7.top_sub_9ns_9s_9_2_1_Adder_6_U.fas_s2  = \sub_9ns_9s_9_2_1_U7.top_sub_9ns_9s_9_2_1_Adder_6_U.u2.s ;
assign \sub_9ns_9s_9_2_1_U7.top_sub_9ns_9s_9_2_1_Adder_6_U.u1.a  = \sub_9ns_9s_9_2_1_U7.top_sub_9ns_9s_9_2_1_Adder_6_U.a [3:0];
assign \sub_9ns_9s_9_2_1_U7.top_sub_9ns_9s_9_2_1_Adder_6_U.u1.b  = \sub_9ns_9s_9_2_1_U7.top_sub_9ns_9s_9_2_1_Adder_6_U.bin_s0 [3:0];
assign \sub_9ns_9s_9_2_1_U7.top_sub_9ns_9s_9_2_1_Adder_6_U.u1.cin  = 1'h1;
assign \sub_9ns_9s_9_2_1_U7.top_sub_9ns_9s_9_2_1_Adder_6_U.facout_s1  = \sub_9ns_9s_9_2_1_U7.top_sub_9ns_9s_9_2_1_Adder_6_U.u1.cout ;
assign \sub_9ns_9s_9_2_1_U7.top_sub_9ns_9s_9_2_1_Adder_6_U.fas_s1  = \sub_9ns_9s_9_2_1_U7.top_sub_9ns_9s_9_2_1_Adder_6_U.u1.s ;
assign \sub_9ns_9s_9_2_1_U7.top_sub_9ns_9s_9_2_1_Adder_6_U.a  = \sub_9ns_9s_9_2_1_U7.din0 ;
assign \sub_9ns_9s_9_2_1_U7.top_sub_9ns_9s_9_2_1_Adder_6_U.b  = \sub_9ns_9s_9_2_1_U7.din1 ;
assign \sub_9ns_9s_9_2_1_U7.top_sub_9ns_9s_9_2_1_Adder_6_U.ce  = \sub_9ns_9s_9_2_1_U7.ce ;
assign \sub_9ns_9s_9_2_1_U7.top_sub_9ns_9s_9_2_1_Adder_6_U.clk  = \sub_9ns_9s_9_2_1_U7.clk ;
assign \sub_9ns_9s_9_2_1_U7.top_sub_9ns_9s_9_2_1_Adder_6_U.reset  = \sub_9ns_9s_9_2_1_U7.reset ;
assign \sub_9ns_9s_9_2_1_U7.dout  = \sub_9ns_9s_9_2_1_U7.top_sub_9ns_9s_9_2_1_Adder_6_U.s ;
assign \sub_9ns_9s_9_2_1_U7.ce  = 1'h1;
assign \sub_9ns_9s_9_2_1_U7.clk  = ap_clk;
assign \sub_9ns_9s_9_2_1_U7.din0  = 9'h000;
assign \sub_9ns_9s_9_2_1_U7.din1  = { r_reg_919[7], r_reg_919 };
assign grp_fu_399_p2 = \sub_9ns_9s_9_2_1_U7.dout ;
assign \sub_9ns_9s_9_2_1_U7.reset  = ap_rst;
assign \sub_4ns_4ns_4_2_1_U9.top_sub_4ns_4ns_4_2_1_Adder_8_U.ain_s0  = \sub_4ns_4ns_4_2_1_U9.top_sub_4ns_4ns_4_2_1_Adder_8_U.a ;
assign \sub_4ns_4ns_4_2_1_U9.top_sub_4ns_4ns_4_2_1_Adder_8_U.s  = { \sub_4ns_4ns_4_2_1_U9.top_sub_4ns_4ns_4_2_1_Adder_8_U.fas_s2 , \sub_4ns_4ns_4_2_1_U9.top_sub_4ns_4ns_4_2_1_Adder_8_U.sum_s1  };
assign \sub_4ns_4ns_4_2_1_U9.top_sub_4ns_4ns_4_2_1_Adder_8_U.u2.a  = \sub_4ns_4ns_4_2_1_U9.top_sub_4ns_4ns_4_2_1_Adder_8_U.ain_s1 ;
assign \sub_4ns_4ns_4_2_1_U9.top_sub_4ns_4ns_4_2_1_Adder_8_U.u2.b  = \sub_4ns_4ns_4_2_1_U9.top_sub_4ns_4ns_4_2_1_Adder_8_U.bin_s1 ;
assign \sub_4ns_4ns_4_2_1_U9.top_sub_4ns_4ns_4_2_1_Adder_8_U.u2.cin  = \sub_4ns_4ns_4_2_1_U9.top_sub_4ns_4ns_4_2_1_Adder_8_U.carry_s1 ;
assign \sub_4ns_4ns_4_2_1_U9.top_sub_4ns_4ns_4_2_1_Adder_8_U.facout_s2  = \sub_4ns_4ns_4_2_1_U9.top_sub_4ns_4ns_4_2_1_Adder_8_U.u2.cout ;
assign \sub_4ns_4ns_4_2_1_U9.top_sub_4ns_4ns_4_2_1_Adder_8_U.fas_s2  = \sub_4ns_4ns_4_2_1_U9.top_sub_4ns_4ns_4_2_1_Adder_8_U.u2.s ;
assign \sub_4ns_4ns_4_2_1_U9.top_sub_4ns_4ns_4_2_1_Adder_8_U.u1.a  = \sub_4ns_4ns_4_2_1_U9.top_sub_4ns_4ns_4_2_1_Adder_8_U.a [1:0];
assign \sub_4ns_4ns_4_2_1_U9.top_sub_4ns_4ns_4_2_1_Adder_8_U.u1.b  = \sub_4ns_4ns_4_2_1_U9.top_sub_4ns_4ns_4_2_1_Adder_8_U.bin_s0 [1:0];
assign \sub_4ns_4ns_4_2_1_U9.top_sub_4ns_4ns_4_2_1_Adder_8_U.u1.cin  = 1'h1;
assign \sub_4ns_4ns_4_2_1_U9.top_sub_4ns_4ns_4_2_1_Adder_8_U.facout_s1  = \sub_4ns_4ns_4_2_1_U9.top_sub_4ns_4ns_4_2_1_Adder_8_U.u1.cout ;
assign \sub_4ns_4ns_4_2_1_U9.top_sub_4ns_4ns_4_2_1_Adder_8_U.fas_s1  = \sub_4ns_4ns_4_2_1_U9.top_sub_4ns_4ns_4_2_1_Adder_8_U.u1.s ;
assign \sub_4ns_4ns_4_2_1_U9.top_sub_4ns_4ns_4_2_1_Adder_8_U.a  = \sub_4ns_4ns_4_2_1_U9.din0 ;
assign \sub_4ns_4ns_4_2_1_U9.top_sub_4ns_4ns_4_2_1_Adder_8_U.b  = \sub_4ns_4ns_4_2_1_U9.din1 ;
assign \sub_4ns_4ns_4_2_1_U9.top_sub_4ns_4ns_4_2_1_Adder_8_U.ce  = \sub_4ns_4ns_4_2_1_U9.ce ;
assign \sub_4ns_4ns_4_2_1_U9.top_sub_4ns_4ns_4_2_1_Adder_8_U.clk  = \sub_4ns_4ns_4_2_1_U9.clk ;
assign \sub_4ns_4ns_4_2_1_U9.top_sub_4ns_4ns_4_2_1_Adder_8_U.reset  = \sub_4ns_4ns_4_2_1_U9.reset ;
assign \sub_4ns_4ns_4_2_1_U9.dout  = \sub_4ns_4ns_4_2_1_U9.top_sub_4ns_4ns_4_2_1_Adder_8_U.s ;
assign \sub_4ns_4ns_4_2_1_U9.ce  = 1'h1;
assign \sub_4ns_4ns_4_2_1_U9.clk  = ap_clk;
assign \sub_4ns_4ns_4_2_1_U9.din0  = 4'h0;
assign \sub_4ns_4ns_4_2_1_U9.din1  = op_6;
assign grp_fu_478_p2 = \sub_4ns_4ns_4_2_1_U9.dout ;
assign \sub_4ns_4ns_4_2_1_U9.reset  = ap_rst;
assign \shl_32s_32s_32_7_1_U11.din1_cast  = \shl_32s_32s_32_7_1_U11.din1 ;
assign \shl_32s_32s_32_7_1_U11.din1_mask  = 32'd31;
assign \shl_32s_32s_32_7_1_U11.ce  = 1'h1;
assign \shl_32s_32s_32_7_1_U11.clk  = ap_clk;
assign \shl_32s_32s_32_7_1_U11.din0  = { op_7[7], op_7[7], op_7[7], op_7[7], op_7[7], op_7[7], op_7[7], op_7[7], op_7[7], op_7[7], op_7[7], op_7[7], op_7[7], op_7[7], op_7[7], op_7[7], op_7[7], op_7[7], op_7[7], op_7[7], op_7[7], op_7[7], op_7[7], op_7[7], op_7 };
assign \shl_32s_32s_32_7_1_U11.din1  = { ush_reg_966[8], ush_reg_966[8], ush_reg_966[8], ush_reg_966[8], ush_reg_966[8], ush_reg_966[8], ush_reg_966[8], ush_reg_966[8], ush_reg_966[8], ush_reg_966[8], ush_reg_966[8], ush_reg_966[8], ush_reg_966[8], ush_reg_966[8], ush_reg_966[8], ush_reg_966[8], ush_reg_966[8], ush_reg_966[8], ush_reg_966[8], ush_reg_966[8], ush_reg_966[8], ush_reg_966[8], ush_reg_966[8], ush_reg_966 };
assign grp_fu_519_p2 = \shl_32s_32s_32_7_1_U11.dout ;
assign \shl_32s_32s_32_7_1_U11.reset  = ap_rst;
assign \shl_16ns_4ns_16_7_1_U13.din1_cast  = \shl_16ns_4ns_16_7_1_U13.din1 [3:0];
assign \shl_16ns_4ns_16_7_1_U13.din1_mask  = 4'h1;
assign \shl_16ns_4ns_16_7_1_U13.ce  = 1'h1;
assign \shl_16ns_4ns_16_7_1_U13.clk  = ap_clk;
assign \shl_16ns_4ns_16_7_1_U13.din0  = op_4;
assign \shl_16ns_4ns_16_7_1_U13.din1  = { 12'h000, sh_reg_1017 };
assign grp_fu_538_p2 = \shl_16ns_4ns_16_7_1_U13.dout ;
assign \shl_16ns_4ns_16_7_1_U13.reset  = ap_rst;
assign \ashr_32s_32s_32_7_1_U10.din1_cast  = \ashr_32s_32s_32_7_1_U10.din1 ;
assign \ashr_32s_32s_32_7_1_U10.din1_mask  = 32'd31;
assign \ashr_32s_32s_32_7_1_U10.ce  = 1'h1;
assign \ashr_32s_32s_32_7_1_U10.clk  = ap_clk;
assign \ashr_32s_32s_32_7_1_U10.din0  = { op_7[7], op_7[7], op_7[7], op_7[7], op_7[7], op_7[7], op_7[7], op_7[7], op_7[7], op_7[7], op_7[7], op_7[7], op_7[7], op_7[7], op_7[7], op_7[7], op_7[7], op_7[7], op_7[7], op_7[7], op_7[7], op_7[7], op_7[7], op_7[7], op_7 };
assign \ashr_32s_32s_32_7_1_U10.din1  = { ush_reg_966[8], ush_reg_966[8], ush_reg_966[8], ush_reg_966[8], ush_reg_966[8], ush_reg_966[8], ush_reg_966[8], ush_reg_966[8], ush_reg_966[8], ush_reg_966[8], ush_reg_966[8], ush_reg_966[8], ush_reg_966[8], ush_reg_966[8], ush_reg_966[8], ush_reg_966[8], ush_reg_966[8], ush_reg_966[8], ush_reg_966[8], ush_reg_966[8], ush_reg_966[8], ush_reg_966[8], ush_reg_966[8], ush_reg_966 };
assign grp_fu_513_p2 = \ashr_32s_32s_32_7_1_U10.dout ;
assign \ashr_32s_32s_32_7_1_U10.reset  = ap_rst;
assign \ashr_16ns_4ns_16_7_1_U14.din1_cast  = \ashr_16ns_4ns_16_7_1_U14.din1 [3:0];
assign \ashr_16ns_4ns_16_7_1_U14.din1_mask  = 4'h1;
assign \ashr_16ns_4ns_16_7_1_U14.ce  = 1'h1;
assign \ashr_16ns_4ns_16_7_1_U14.clk  = ap_clk;
assign \ashr_16ns_4ns_16_7_1_U14.din0  = op_4;
assign \ashr_16ns_4ns_16_7_1_U14.din1  = { 12'h000, op_6 };
assign grp_fu_546_p2 = \ashr_16ns_4ns_16_7_1_U14.dout ;
assign \ashr_16ns_4ns_16_7_1_U14.reset  = ap_rst;
assign \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.ain_s0  = \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.a ;
assign \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.bin_s0  = \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.b ;
assign \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.s  = { \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.fas_s2 , \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.sum_s1  };
assign \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.u2.a  = \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.ain_s1 ;
assign \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.u2.b  = \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.bin_s1 ;
assign \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.u2.cin  = \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.carry_s1 ;
assign \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.facout_s2  = \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.u2.cout ;
assign \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.fas_s2  = \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.u2.s ;
assign \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.u1.a  = \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.a [3:0];
assign \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.u1.b  = \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.b [3:0];
assign \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.u1.cin  = 1'h0;
assign \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.facout_s1  = \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.u1.cout ;
assign \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.fas_s1  = \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.u1.s ;
assign \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.a  = \add_9s_9s_9_2_1_U1.din0 ;
assign \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.b  = \add_9s_9s_9_2_1_U1.din1 ;
assign \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.ce  = \add_9s_9s_9_2_1_U1.ce ;
assign \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.clk  = \add_9s_9s_9_2_1_U1.clk ;
assign \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.reset  = \add_9s_9s_9_2_1_U1.reset ;
assign \add_9s_9s_9_2_1_U1.dout  = \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.s ;
assign \add_9s_9s_9_2_1_U1.ce  = 1'h1;
assign \add_9s_9s_9_2_1_U1.clk  = ap_clk;
assign \add_9s_9s_9_2_1_U1.din0  = { op_5[7], op_5 };
assign \add_9s_9s_9_2_1_U1.din1  = { op_8[3], op_8[3], op_8[3], op_8[3], op_8[3], op_8 };
assign grp_fu_243_p2 = \add_9s_9s_9_2_1_U1.dout ;
assign \add_9s_9s_9_2_1_U1.reset  = ap_rst;
assign \add_46s_46s_46_2_1_U5.top_add_46s_46s_46_2_1_Adder_4_U.ain_s0  = \add_46s_46s_46_2_1_U5.top_add_46s_46s_46_2_1_Adder_4_U.a ;
assign \add_46s_46s_46_2_1_U5.top_add_46s_46s_46_2_1_Adder_4_U.bin_s0  = \add_46s_46s_46_2_1_U5.top_add_46s_46s_46_2_1_Adder_4_U.b ;
assign \add_46s_46s_46_2_1_U5.top_add_46s_46s_46_2_1_Adder_4_U.s  = { \add_46s_46s_46_2_1_U5.top_add_46s_46s_46_2_1_Adder_4_U.fas_s2 , \add_46s_46s_46_2_1_U5.top_add_46s_46s_46_2_1_Adder_4_U.sum_s1  };
assign \add_46s_46s_46_2_1_U5.top_add_46s_46s_46_2_1_Adder_4_U.u2.a  = \add_46s_46s_46_2_1_U5.top_add_46s_46s_46_2_1_Adder_4_U.ain_s1 ;
assign \add_46s_46s_46_2_1_U5.top_add_46s_46s_46_2_1_Adder_4_U.u2.b  = \add_46s_46s_46_2_1_U5.top_add_46s_46s_46_2_1_Adder_4_U.bin_s1 ;
assign \add_46s_46s_46_2_1_U5.top_add_46s_46s_46_2_1_Adder_4_U.u2.cin  = \add_46s_46s_46_2_1_U5.top_add_46s_46s_46_2_1_Adder_4_U.carry_s1 ;
assign \add_46s_46s_46_2_1_U5.top_add_46s_46s_46_2_1_Adder_4_U.facout_s2  = \add_46s_46s_46_2_1_U5.top_add_46s_46s_46_2_1_Adder_4_U.u2.cout ;
assign \add_46s_46s_46_2_1_U5.top_add_46s_46s_46_2_1_Adder_4_U.fas_s2  = \add_46s_46s_46_2_1_U5.top_add_46s_46s_46_2_1_Adder_4_U.u2.s ;
assign \add_46s_46s_46_2_1_U5.top_add_46s_46s_46_2_1_Adder_4_U.u1.a  = \add_46s_46s_46_2_1_U5.top_add_46s_46s_46_2_1_Adder_4_U.a [22:0];
assign \add_46s_46s_46_2_1_U5.top_add_46s_46s_46_2_1_Adder_4_U.u1.b  = \add_46s_46s_46_2_1_U5.top_add_46s_46s_46_2_1_Adder_4_U.b [22:0];
assign \add_46s_46s_46_2_1_U5.top_add_46s_46s_46_2_1_Adder_4_U.u1.cin  = 1'h0;
assign \add_46s_46s_46_2_1_U5.top_add_46s_46s_46_2_1_Adder_4_U.facout_s1  = \add_46s_46s_46_2_1_U5.top_add_46s_46s_46_2_1_Adder_4_U.u1.cout ;
assign \add_46s_46s_46_2_1_U5.top_add_46s_46s_46_2_1_Adder_4_U.fas_s1  = \add_46s_46s_46_2_1_U5.top_add_46s_46s_46_2_1_Adder_4_U.u1.s ;
assign \add_46s_46s_46_2_1_U5.top_add_46s_46s_46_2_1_Adder_4_U.a  = \add_46s_46s_46_2_1_U5.din0 ;
assign \add_46s_46s_46_2_1_U5.top_add_46s_46s_46_2_1_Adder_4_U.b  = \add_46s_46s_46_2_1_U5.din1 ;
assign \add_46s_46s_46_2_1_U5.top_add_46s_46s_46_2_1_Adder_4_U.ce  = \add_46s_46s_46_2_1_U5.ce ;
assign \add_46s_46s_46_2_1_U5.top_add_46s_46s_46_2_1_Adder_4_U.clk  = \add_46s_46s_46_2_1_U5.clk ;
assign \add_46s_46s_46_2_1_U5.top_add_46s_46s_46_2_1_Adder_4_U.reset  = \add_46s_46s_46_2_1_U5.reset ;
assign \add_46s_46s_46_2_1_U5.dout  = \add_46s_46s_46_2_1_U5.top_add_46s_46s_46_2_1_Adder_4_U.s ;
assign \add_46s_46s_46_2_1_U5.ce  = 1'h1;
assign \add_46s_46s_46_2_1_U5.clk  = ap_clk;
assign \add_46s_46s_46_2_1_U5.din0  = { op_23_V_reg_887[9], op_23_V_reg_887[9], op_23_V_reg_887[9], op_23_V_reg_887[9], op_23_V_reg_887[9], op_23_V_reg_887[9], op_23_V_reg_887[9], op_23_V_reg_887[9], op_23_V_reg_887[9], op_23_V_reg_887[9], op_23_V_reg_887[9], op_23_V_reg_887[9], op_23_V_reg_887[9], op_23_V_reg_887[9], op_23_V_reg_887[9], op_23_V_reg_887[9], op_23_V_reg_887[9], op_23_V_reg_887[9], op_23_V_reg_887[9], op_23_V_reg_887[9], op_23_V_reg_887[9], op_23_V_reg_887[9], op_23_V_reg_887[9], op_23_V_reg_887, 13'h0000 };
assign \add_46s_46s_46_2_1_U5.din1  = { op_12[15], op_12[15], op_12[15], op_12[15], op_12[15], op_12[15], op_12[15], op_12[15], op_12[15], op_12[15], op_12[15], op_12[15], op_12[15], op_12[15], op_12[15], op_12[15], op_12[15], op_12[15], op_12[15], op_12[15], op_12[15], op_12[15], op_12[15], op_12[15], op_12[15], op_12[15], op_12[15], op_12[15], op_12[15], op_12[15], op_12 };
assign grp_fu_351_p2 = \add_46s_46s_46_2_1_U5.dout ;
assign \add_46s_46s_46_2_1_U5.reset  = ap_rst;
assign \add_45s_45s_45_2_1_U8.top_add_45s_45s_45_2_1_Adder_7_U.ain_s0  = \add_45s_45s_45_2_1_U8.top_add_45s_45s_45_2_1_Adder_7_U.a ;
assign \add_45s_45s_45_2_1_U8.top_add_45s_45s_45_2_1_Adder_7_U.bin_s0  = \add_45s_45s_45_2_1_U8.top_add_45s_45s_45_2_1_Adder_7_U.b ;
assign \add_45s_45s_45_2_1_U8.top_add_45s_45s_45_2_1_Adder_7_U.s  = { \add_45s_45s_45_2_1_U8.top_add_45s_45s_45_2_1_Adder_7_U.fas_s2 , \add_45s_45s_45_2_1_U8.top_add_45s_45s_45_2_1_Adder_7_U.sum_s1  };
assign \add_45s_45s_45_2_1_U8.top_add_45s_45s_45_2_1_Adder_7_U.u2.a  = \add_45s_45s_45_2_1_U8.top_add_45s_45s_45_2_1_Adder_7_U.ain_s1 ;
assign \add_45s_45s_45_2_1_U8.top_add_45s_45s_45_2_1_Adder_7_U.u2.b  = \add_45s_45s_45_2_1_U8.top_add_45s_45s_45_2_1_Adder_7_U.bin_s1 ;
assign \add_45s_45s_45_2_1_U8.top_add_45s_45s_45_2_1_Adder_7_U.u2.cin  = \add_45s_45s_45_2_1_U8.top_add_45s_45s_45_2_1_Adder_7_U.carry_s1 ;
assign \add_45s_45s_45_2_1_U8.top_add_45s_45s_45_2_1_Adder_7_U.facout_s2  = \add_45s_45s_45_2_1_U8.top_add_45s_45s_45_2_1_Adder_7_U.u2.cout ;
assign \add_45s_45s_45_2_1_U8.top_add_45s_45s_45_2_1_Adder_7_U.fas_s2  = \add_45s_45s_45_2_1_U8.top_add_45s_45s_45_2_1_Adder_7_U.u2.s ;
assign \add_45s_45s_45_2_1_U8.top_add_45s_45s_45_2_1_Adder_7_U.u1.a  = \add_45s_45s_45_2_1_U8.top_add_45s_45s_45_2_1_Adder_7_U.a [21:0];
assign \add_45s_45s_45_2_1_U8.top_add_45s_45s_45_2_1_Adder_7_U.u1.b  = \add_45s_45s_45_2_1_U8.top_add_45s_45s_45_2_1_Adder_7_U.b [21:0];
assign \add_45s_45s_45_2_1_U8.top_add_45s_45s_45_2_1_Adder_7_U.u1.cin  = 1'h0;
assign \add_45s_45s_45_2_1_U8.top_add_45s_45s_45_2_1_Adder_7_U.facout_s1  = \add_45s_45s_45_2_1_U8.top_add_45s_45s_45_2_1_Adder_7_U.u1.cout ;
assign \add_45s_45s_45_2_1_U8.top_add_45s_45s_45_2_1_Adder_7_U.fas_s1  = \add_45s_45s_45_2_1_U8.top_add_45s_45s_45_2_1_Adder_7_U.u1.s ;
assign \add_45s_45s_45_2_1_U8.top_add_45s_45s_45_2_1_Adder_7_U.a  = \add_45s_45s_45_2_1_U8.din0 ;
assign \add_45s_45s_45_2_1_U8.top_add_45s_45s_45_2_1_Adder_7_U.b  = \add_45s_45s_45_2_1_U8.din1 ;
assign \add_45s_45s_45_2_1_U8.top_add_45s_45s_45_2_1_Adder_7_U.ce  = \add_45s_45s_45_2_1_U8.ce ;
assign \add_45s_45s_45_2_1_U8.top_add_45s_45s_45_2_1_Adder_7_U.clk  = \add_45s_45s_45_2_1_U8.clk ;
assign \add_45s_45s_45_2_1_U8.top_add_45s_45s_45_2_1_Adder_7_U.reset  = \add_45s_45s_45_2_1_U8.reset ;
assign \add_45s_45s_45_2_1_U8.dout  = \add_45s_45s_45_2_1_U8.top_add_45s_45s_45_2_1_Adder_7_U.s ;
assign \add_45s_45s_45_2_1_U8.ce  = 1'h1;
assign \add_45s_45s_45_2_1_U8.clk  = ap_clk;
assign \add_45s_45s_45_2_1_U8.din0  = { select_ln353_reg_941[31], select_ln353_reg_941, 12'h000 };
assign \add_45s_45s_45_2_1_U8.din1  = { op_13[15], op_13[15], op_13[15], op_13[15], op_13[15], op_13[15], op_13[15], op_13[15], op_13[15], op_13[15], op_13[15], op_13[15], op_13[15], op_13[15], op_13[15], op_13[15], op_13[15], op_13[15], op_13[15], op_13[15], op_13[15], op_13[15], op_13[15], op_13[15], op_13[15], op_13[15], op_13[15], op_13[15], op_13[15], op_13 };
assign grp_fu_439_p2 = \add_45s_45s_45_2_1_U8.dout ;
assign \add_45s_45s_45_2_1_U8.reset  = ap_rst;
assign \add_3s_3ns_3_2_1_U20.top_add_3s_3ns_3_2_1_Adder_12_U.ain_s0  = \add_3s_3ns_3_2_1_U20.top_add_3s_3ns_3_2_1_Adder_12_U.a ;
assign \add_3s_3ns_3_2_1_U20.top_add_3s_3ns_3_2_1_Adder_12_U.bin_s0  = \add_3s_3ns_3_2_1_U20.top_add_3s_3ns_3_2_1_Adder_12_U.b ;
assign \add_3s_3ns_3_2_1_U20.top_add_3s_3ns_3_2_1_Adder_12_U.s  = { \add_3s_3ns_3_2_1_U20.top_add_3s_3ns_3_2_1_Adder_12_U.fas_s2 , \add_3s_3ns_3_2_1_U20.top_add_3s_3ns_3_2_1_Adder_12_U.sum_s1  };
assign \add_3s_3ns_3_2_1_U20.top_add_3s_3ns_3_2_1_Adder_12_U.u2.a  = \add_3s_3ns_3_2_1_U20.top_add_3s_3ns_3_2_1_Adder_12_U.ain_s1 ;
assign \add_3s_3ns_3_2_1_U20.top_add_3s_3ns_3_2_1_Adder_12_U.u2.b  = \add_3s_3ns_3_2_1_U20.top_add_3s_3ns_3_2_1_Adder_12_U.bin_s1 ;
assign \add_3s_3ns_3_2_1_U20.top_add_3s_3ns_3_2_1_Adder_12_U.u2.cin  = \add_3s_3ns_3_2_1_U20.top_add_3s_3ns_3_2_1_Adder_12_U.carry_s1 ;
assign \add_3s_3ns_3_2_1_U20.top_add_3s_3ns_3_2_1_Adder_12_U.facout_s2  = \add_3s_3ns_3_2_1_U20.top_add_3s_3ns_3_2_1_Adder_12_U.u2.cout ;
assign \add_3s_3ns_3_2_1_U20.top_add_3s_3ns_3_2_1_Adder_12_U.fas_s2  = \add_3s_3ns_3_2_1_U20.top_add_3s_3ns_3_2_1_Adder_12_U.u2.s ;
assign \add_3s_3ns_3_2_1_U20.top_add_3s_3ns_3_2_1_Adder_12_U.u1.a  = \add_3s_3ns_3_2_1_U20.top_add_3s_3ns_3_2_1_Adder_12_U.a [0];
assign \add_3s_3ns_3_2_1_U20.top_add_3s_3ns_3_2_1_Adder_12_U.u1.b  = \add_3s_3ns_3_2_1_U20.top_add_3s_3ns_3_2_1_Adder_12_U.b [0];
assign \add_3s_3ns_3_2_1_U20.top_add_3s_3ns_3_2_1_Adder_12_U.u1.cin  = 1'h0;
assign \add_3s_3ns_3_2_1_U20.top_add_3s_3ns_3_2_1_Adder_12_U.facout_s1  = \add_3s_3ns_3_2_1_U20.top_add_3s_3ns_3_2_1_Adder_12_U.u1.cout ;
assign \add_3s_3ns_3_2_1_U20.top_add_3s_3ns_3_2_1_Adder_12_U.fas_s1  = \add_3s_3ns_3_2_1_U20.top_add_3s_3ns_3_2_1_Adder_12_U.u1.s ;
assign \add_3s_3ns_3_2_1_U20.top_add_3s_3ns_3_2_1_Adder_12_U.a  = \add_3s_3ns_3_2_1_U20.din0 ;
assign \add_3s_3ns_3_2_1_U20.top_add_3s_3ns_3_2_1_Adder_12_U.b  = \add_3s_3ns_3_2_1_U20.din1 ;
assign \add_3s_3ns_3_2_1_U20.top_add_3s_3ns_3_2_1_Adder_12_U.ce  = \add_3s_3ns_3_2_1_U20.ce ;
assign \add_3s_3ns_3_2_1_U20.top_add_3s_3ns_3_2_1_Adder_12_U.clk  = \add_3s_3ns_3_2_1_U20.clk ;
assign \add_3s_3ns_3_2_1_U20.top_add_3s_3ns_3_2_1_Adder_12_U.reset  = \add_3s_3ns_3_2_1_U20.reset ;
assign \add_3s_3ns_3_2_1_U20.dout  = \add_3s_3ns_3_2_1_U20.top_add_3s_3ns_3_2_1_Adder_12_U.s ;
assign \add_3s_3ns_3_2_1_U20.ce  = 1'h1;
assign \add_3s_3ns_3_2_1_U20.clk  = ap_clk;
assign \add_3s_3ns_3_2_1_U20.din0  = { ret_V_4_reg_1168[1], ret_V_4_reg_1168 };
assign \add_3s_3ns_3_2_1_U20.din1  = select_ln69_reg_1047;
assign grp_fu_760_p2 = \add_3s_3ns_3_2_1_U20.dout ;
assign \add_3s_3ns_3_2_1_U20.reset  = ap_rst;
assign \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.ain_s0  = \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.a ;
assign \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.bin_s0  = \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.b ;
assign \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.s  = { \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.fas_s2 , \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.sum_s1  };
assign \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.u2.a  = \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.ain_s1 ;
assign \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.u2.b  = \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.bin_s1 ;
assign \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.u2.cin  = \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.carry_s1 ;
assign \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.facout_s2  = \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.u2.cout ;
assign \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.fas_s2  = \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.u2.s ;
assign \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.u1.a  = \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.a [16:0];
assign \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.u1.b  = \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.b [16:0];
assign \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.u1.cin  = 1'h0;
assign \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.facout_s1  = \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.u1.cout ;
assign \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.fas_s1  = \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.u1.s ;
assign \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.a  = \add_35s_35s_35_2_1_U15.din0 ;
assign \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.b  = \add_35s_35s_35_2_1_U15.din1 ;
assign \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.ce  = \add_35s_35s_35_2_1_U15.ce ;
assign \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.clk  = \add_35s_35s_35_2_1_U15.clk ;
assign \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.reset  = \add_35s_35s_35_2_1_U15.reset ;
assign \add_35s_35s_35_2_1_U15.dout  = \add_35s_35s_35_2_1_U15.top_add_35s_35s_35_2_1_Adder_9_U.s ;
assign \add_35s_35s_35_2_1_U15.ce  = 1'h1;
assign \add_35s_35s_35_2_1_U15.clk  = ap_clk;
assign \add_35s_35s_35_2_1_U15.din0  = { select_ln353_1_reg_1042[31], select_ln353_1_reg_1042, 2'h0 };
assign \add_35s_35s_35_2_1_U15.din1  = { op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14 };
assign grp_fu_618_p2 = \add_35s_35s_35_2_1_U15.dout ;
assign \add_35s_35s_35_2_1_U15.reset  = ap_rst;
assign \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.ain_s0  = \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.a ;
assign \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.bin_s0  = \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.b ;
assign \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.s  = { \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.fas_s2 , \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.sum_s1  };
assign \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.u2.a  = \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.ain_s1 ;
assign \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.u2.b  = \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.bin_s1 ;
assign \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.u2.cin  = \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.carry_s1 ;
assign \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.facout_s2  = \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.u2.cout ;
assign \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.fas_s2  = \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.u2.s ;
assign \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.u1.a  = \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.a [16:0];
assign \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.u1.b  = \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.b [16:0];
assign \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.u1.cin  = 1'h0;
assign \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.facout_s1  = \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.u1.cout ;
assign \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.fas_s1  = \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.u1.s ;
assign \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.a  = \add_34s_34s_34_2_1_U18.din0 ;
assign \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.b  = \add_34s_34s_34_2_1_U18.din1 ;
assign \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.ce  = \add_34s_34s_34_2_1_U18.ce ;
assign \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.clk  = \add_34s_34s_34_2_1_U18.clk ;
assign \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.reset  = \add_34s_34s_34_2_1_U18.reset ;
assign \add_34s_34s_34_2_1_U18.dout  = \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.s ;
assign \add_34s_34s_34_2_1_U18.ce  = 1'h1;
assign \add_34s_34s_34_2_1_U18.clk  = ap_clk;
assign \add_34s_34s_34_2_1_U18.din0  = { select_ln353_2_reg_1111[31], select_ln353_2_reg_1111, 1'h0 };
assign \add_34s_34s_34_2_1_U18.din1  = { op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15 };
assign grp_fu_712_p2 = \add_34s_34s_34_2_1_U18.dout ;
assign \add_34s_34s_34_2_1_U18.reset  = ap_rst;
assign \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_14_U.ain_s0  = \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_14_U.a ;
assign \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_14_U.bin_s0  = \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_14_U.b ;
assign \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_14_U.s  = { \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_14_U.fas_s2 , \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_14_U.sum_s1  };
assign \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_14_U.u2.a  = \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_14_U.ain_s1 ;
assign \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_14_U.u2.b  = \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_14_U.bin_s1 ;
assign \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_14_U.u2.cin  = \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_14_U.carry_s1 ;
assign \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_14_U.facout_s2  = \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_14_U.u2.cout ;
assign \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_14_U.fas_s2  = \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_14_U.u2.s ;
assign \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_14_U.u1.a  = \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_14_U.a [15:0];
assign \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_14_U.u1.b  = \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_14_U.b [15:0];
assign \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_14_U.u1.cin  = 1'h0;
assign \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_14_U.facout_s1  = \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_14_U.u1.cout ;
assign \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_14_U.fas_s1  = \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_14_U.u1.s ;
assign \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_14_U.a  = \add_32s_32ns_32_2_1_U23.din0 ;
assign \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_14_U.b  = \add_32s_32ns_32_2_1_U23.din1 ;
assign \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_14_U.ce  = \add_32s_32ns_32_2_1_U23.ce ;
assign \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_14_U.clk  = \add_32s_32ns_32_2_1_U23.clk ;
assign \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_14_U.reset  = \add_32s_32ns_32_2_1_U23.reset ;
assign \add_32s_32ns_32_2_1_U23.dout  = \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_14_U.s ;
assign \add_32s_32ns_32_2_1_U23.ce  = 1'h1;
assign \add_32s_32ns_32_2_1_U23.clk  = ap_clk;
assign \add_32s_32ns_32_2_1_U23.din0  = { add_ln69_2_reg_1213[16], add_ln69_2_reg_1213[16], add_ln69_2_reg_1213[16], add_ln69_2_reg_1213[16], add_ln69_2_reg_1213[16], add_ln69_2_reg_1213[16], add_ln69_2_reg_1213[16], add_ln69_2_reg_1213[16], add_ln69_2_reg_1213[16], add_ln69_2_reg_1213[16], add_ln69_2_reg_1213[16], add_ln69_2_reg_1213[16], add_ln69_2_reg_1213[16], add_ln69_2_reg_1213[16], add_ln69_2_reg_1213[16], add_ln69_2_reg_1213 };
assign \add_32s_32ns_32_2_1_U23.din1  = add_ln69_reg_1208;
assign grp_fu_808_p2 = \add_32s_32ns_32_2_1_U23.dout ;
assign \add_32s_32ns_32_2_1_U23.reset  = ap_rst;
assign \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.ain_s0  = \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.a ;
assign \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.bin_s0  = \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.b ;
assign \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.s  = { \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.fas_s2 , \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.sum_s1  };
assign \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.a  = \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.ain_s1 ;
assign \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.b  = \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.bin_s1 ;
assign \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.cin  = \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.carry_s1 ;
assign \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.facout_s2  = \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.cout ;
assign \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.fas_s2  = \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.s ;
assign \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.a  = \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.a [15:0];
assign \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.b  = \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.b [15:0];
assign \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.cin  = 1'h0;
assign \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.facout_s1  = \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.cout ;
assign \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.fas_s1  = \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.s ;
assign \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.a  = \add_32ns_32ns_32_2_1_U6.din0 ;
assign \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.b  = \add_32ns_32ns_32_2_1_U6.din1 ;
assign \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.ce  = \add_32ns_32ns_32_2_1_U6.ce ;
assign \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.clk  = \add_32ns_32ns_32_2_1_U6.clk ;
assign \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.reset  = \add_32ns_32ns_32_2_1_U6.reset ;
assign \add_32ns_32ns_32_2_1_U6.dout  = \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.s ;
assign \add_32ns_32ns_32_2_1_U6.ce  = 1'h1;
assign \add_32ns_32ns_32_2_1_U6.clk  = ap_clk;
assign \add_32ns_32ns_32_2_1_U6.din0  = ret_V_21_cast_reg_912;
assign \add_32ns_32ns_32_2_1_U6.din1  = 32'd1;
assign grp_fu_377_p2 = \add_32ns_32ns_32_2_1_U6.dout ;
assign \add_32ns_32ns_32_2_1_U6.reset  = ap_rst;
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_5_U.ain_s0  = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_5_U.a ;
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_5_U.bin_s0  = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_5_U.b ;
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_5_U.s  = { \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_5_U.fas_s2 , \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_5_U.sum_s1  };
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.a  = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_5_U.ain_s1 ;
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.b  = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_5_U.bin_s1 ;
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.cin  = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_5_U.carry_s1 ;
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_5_U.facout_s2  = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.cout ;
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_5_U.fas_s2  = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.s ;
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.a  = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_5_U.a [15:0];
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.b  = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_5_U.b [15:0];
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.cin  = 1'h0;
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_5_U.facout_s1  = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.cout ;
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_5_U.fas_s1  = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.s ;
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_5_U.a  = \add_32ns_32ns_32_2_1_U21.din0 ;
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_5_U.b  = \add_32ns_32ns_32_2_1_U21.din1 ;
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_5_U.ce  = \add_32ns_32ns_32_2_1_U21.ce ;
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_5_U.clk  = \add_32ns_32ns_32_2_1_U21.clk ;
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_5_U.reset  = \add_32ns_32ns_32_2_1_U21.reset ;
assign \add_32ns_32ns_32_2_1_U21.dout  = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_5_U.s ;
assign \add_32ns_32ns_32_2_1_U21.ce  = 1'h1;
assign \add_32ns_32ns_32_2_1_U21.clk  = ap_clk;
assign \add_32ns_32ns_32_2_1_U21.din0  = ret_V_20_reg_1183;
assign \add_32ns_32ns_32_2_1_U21.din1  = op_19;
assign grp_fu_791_p2 = \add_32ns_32ns_32_2_1_U21.dout ;
assign \add_32ns_32ns_32_2_1_U21.reset  = ap_rst;
assign \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_5_U.ain_s0  = \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_5_U.a ;
assign \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_5_U.bin_s0  = \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_5_U.b ;
assign \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_5_U.s  = { \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_5_U.fas_s2 , \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_5_U.sum_s1  };
assign \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.a  = \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_5_U.ain_s1 ;
assign \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.b  = \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_5_U.bin_s1 ;
assign \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.cin  = \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_5_U.carry_s1 ;
assign \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_5_U.facout_s2  = \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.cout ;
assign \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_5_U.fas_s2  = \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.s ;
assign \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.a  = \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_5_U.a [15:0];
assign \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.b  = \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_5_U.b [15:0];
assign \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.cin  = 1'h0;
assign \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_5_U.facout_s1  = \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.cout ;
assign \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_5_U.fas_s1  = \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.s ;
assign \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_5_U.a  = \add_32ns_32ns_32_2_1_U19.din0 ;
assign \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_5_U.b  = \add_32ns_32ns_32_2_1_U19.din1 ;
assign \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_5_U.ce  = \add_32ns_32ns_32_2_1_U19.ce ;
assign \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_5_U.clk  = \add_32ns_32ns_32_2_1_U19.clk ;
assign \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_5_U.reset  = \add_32ns_32ns_32_2_1_U19.reset ;
assign \add_32ns_32ns_32_2_1_U19.dout  = \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_5_U.s ;
assign \add_32ns_32ns_32_2_1_U19.ce  = 1'h1;
assign \add_32ns_32ns_32_2_1_U19.clk  = ap_clk;
assign \add_32ns_32ns_32_2_1_U19.din0  = ret_V_27_cast_reg_1161;
assign \add_32ns_32ns_32_2_1_U19.din1  = 32'd1;
assign grp_fu_752_p2 = \add_32ns_32ns_32_2_1_U19.dout ;
assign \add_32ns_32ns_32_2_1_U19.reset  = ap_rst;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_5_U.ain_s0  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_5_U.a ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_5_U.bin_s0  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_5_U.b ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_5_U.s  = { \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_5_U.fas_s2 , \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_5_U.sum_s1  };
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.a  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_5_U.ain_s1 ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.b  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_5_U.bin_s1 ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.cin  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_5_U.carry_s1 ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_5_U.facout_s2  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.cout ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_5_U.fas_s2  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.s ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.a  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_5_U.a [15:0];
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.b  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_5_U.b [15:0];
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.cin  = 1'h0;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_5_U.facout_s1  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.cout ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_5_U.fas_s1  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.s ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_5_U.a  = \add_32ns_32ns_32_2_1_U16.din0 ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_5_U.b  = \add_32ns_32ns_32_2_1_U16.din1 ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_5_U.ce  = \add_32ns_32ns_32_2_1_U16.ce ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_5_U.clk  = \add_32ns_32ns_32_2_1_U16.clk ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_5_U.reset  = \add_32ns_32ns_32_2_1_U16.reset ;
assign \add_32ns_32ns_32_2_1_U16.dout  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_5_U.s ;
assign \add_32ns_32ns_32_2_1_U16.ce  = 1'h1;
assign \add_32ns_32ns_32_2_1_U16.clk  = ap_clk;
assign \add_32ns_32ns_32_2_1_U16.din0  = ret_V_25_cast_reg_1072;
assign \add_32ns_32ns_32_2_1_U16.din1  = 32'd1;
assign grp_fu_644_p2 = \add_32ns_32ns_32_2_1_U16.dout ;
assign \add_32ns_32ns_32_2_1_U16.reset  = ap_rst;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.ain_s0  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.a ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.bin_s0  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.b ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.s  = { \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.fas_s2 , \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.sum_s1  };
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.a  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.ain_s1 ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.b  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.bin_s1 ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.cin  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.carry_s1 ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.facout_s2  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.cout ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.fas_s2  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.s ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.a  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.a [15:0];
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.b  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.b [15:0];
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.cin  = 1'h0;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.facout_s1  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.cout ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.fas_s1  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.s ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.a  = \add_32ns_32ns_32_2_1_U12.din0 ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.b  = \add_32ns_32ns_32_2_1_U12.din1 ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.ce  = \add_32ns_32ns_32_2_1_U12.ce ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.clk  = \add_32ns_32ns_32_2_1_U12.clk ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.reset  = \add_32ns_32ns_32_2_1_U12.reset ;
assign \add_32ns_32ns_32_2_1_U12.dout  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.s ;
assign \add_32ns_32ns_32_2_1_U12.ce  = 1'h1;
assign \add_32ns_32ns_32_2_1_U12.clk  = ap_clk;
assign \add_32ns_32ns_32_2_1_U12.din0  = ret_V_23_cast_reg_976;
assign \add_32ns_32ns_32_2_1_U12.din1  = 32'd1;
assign grp_fu_525_p2 = \add_32ns_32ns_32_2_1_U12.dout ;
assign \add_32ns_32ns_32_2_1_U12.reset  = ap_rst;
assign \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_10_U.ain_s0  = \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_10_U.a ;
assign \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_10_U.bin_s0  = \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_10_U.b ;
assign \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_10_U.s  = { \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_10_U.fas_s2 , \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_10_U.sum_s1  };
assign \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_10_U.u2.a  = \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_10_U.ain_s1 ;
assign \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_10_U.u2.b  = \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_10_U.bin_s1 ;
assign \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_10_U.u2.cin  = \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_10_U.carry_s1 ;
assign \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_10_U.facout_s2  = \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_10_U.u2.cout ;
assign \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_10_U.fas_s2  = \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_10_U.u2.s ;
assign \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_10_U.u1.a  = \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_10_U.a [0];
assign \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_10_U.u1.b  = \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_10_U.b [0];
assign \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_10_U.u1.cin  = 1'h0;
assign \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_10_U.facout_s1  = \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_10_U.u1.cout ;
assign \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_10_U.fas_s1  = \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_10_U.u1.s ;
assign \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_10_U.a  = \add_2ns_2ns_2_2_1_U17.din0 ;
assign \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_10_U.b  = \add_2ns_2ns_2_2_1_U17.din1 ;
assign \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_10_U.ce  = \add_2ns_2ns_2_2_1_U17.ce ;
assign \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_10_U.clk  = \add_2ns_2ns_2_2_1_U17.clk ;
assign \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_10_U.reset  = \add_2ns_2ns_2_2_1_U17.reset ;
assign \add_2ns_2ns_2_2_1_U17.dout  = \add_2ns_2ns_2_2_1_U17.top_add_2ns_2ns_2_2_1_Adder_10_U.s ;
assign \add_2ns_2ns_2_2_1_U17.ce  = 1'h1;
assign \add_2ns_2ns_2_2_1_U17.clk  = ap_clk;
assign \add_2ns_2ns_2_2_1_U17.din0  = ret_V_reg_1099;
assign \add_2ns_2ns_2_2_1_U17.din1  = 2'h1;
assign grp_fu_692_p2 = \add_2ns_2ns_2_2_1_U17.dout ;
assign \add_2ns_2ns_2_2_1_U17.reset  = ap_rst;
assign \add_17s_17s_17_2_1_U22.top_add_17s_17s_17_2_1_Adder_13_U.ain_s0  = \add_17s_17s_17_2_1_U22.top_add_17s_17s_17_2_1_Adder_13_U.a ;
assign \add_17s_17s_17_2_1_U22.top_add_17s_17s_17_2_1_Adder_13_U.bin_s0  = \add_17s_17s_17_2_1_U22.top_add_17s_17s_17_2_1_Adder_13_U.b ;
assign \add_17s_17s_17_2_1_U22.top_add_17s_17s_17_2_1_Adder_13_U.s  = { \add_17s_17s_17_2_1_U22.top_add_17s_17s_17_2_1_Adder_13_U.fas_s2 , \add_17s_17s_17_2_1_U22.top_add_17s_17s_17_2_1_Adder_13_U.sum_s1  };
assign \add_17s_17s_17_2_1_U22.top_add_17s_17s_17_2_1_Adder_13_U.u2.a  = \add_17s_17s_17_2_1_U22.top_add_17s_17s_17_2_1_Adder_13_U.ain_s1 ;
assign \add_17s_17s_17_2_1_U22.top_add_17s_17s_17_2_1_Adder_13_U.u2.b  = \add_17s_17s_17_2_1_U22.top_add_17s_17s_17_2_1_Adder_13_U.bin_s1 ;
assign \add_17s_17s_17_2_1_U22.top_add_17s_17s_17_2_1_Adder_13_U.u2.cin  = \add_17s_17s_17_2_1_U22.top_add_17s_17s_17_2_1_Adder_13_U.carry_s1 ;
assign \add_17s_17s_17_2_1_U22.top_add_17s_17s_17_2_1_Adder_13_U.facout_s2  = \add_17s_17s_17_2_1_U22.top_add_17s_17s_17_2_1_Adder_13_U.u2.cout ;
assign \add_17s_17s_17_2_1_U22.top_add_17s_17s_17_2_1_Adder_13_U.fas_s2  = \add_17s_17s_17_2_1_U22.top_add_17s_17s_17_2_1_Adder_13_U.u2.s ;
assign \add_17s_17s_17_2_1_U22.top_add_17s_17s_17_2_1_Adder_13_U.u1.a  = \add_17s_17s_17_2_1_U22.top_add_17s_17s_17_2_1_Adder_13_U.a [7:0];
assign \add_17s_17s_17_2_1_U22.top_add_17s_17s_17_2_1_Adder_13_U.u1.b  = \add_17s_17s_17_2_1_U22.top_add_17s_17s_17_2_1_Adder_13_U.b [7:0];
assign \add_17s_17s_17_2_1_U22.top_add_17s_17s_17_2_1_Adder_13_U.u1.cin  = 1'h0;
assign \add_17s_17s_17_2_1_U22.top_add_17s_17s_17_2_1_Adder_13_U.facout_s1  = \add_17s_17s_17_2_1_U22.top_add_17s_17s_17_2_1_Adder_13_U.u1.cout ;
assign \add_17s_17s_17_2_1_U22.top_add_17s_17s_17_2_1_Adder_13_U.fas_s1  = \add_17s_17s_17_2_1_U22.top_add_17s_17s_17_2_1_Adder_13_U.u1.s ;
assign \add_17s_17s_17_2_1_U22.top_add_17s_17s_17_2_1_Adder_13_U.a  = \add_17s_17s_17_2_1_U22.din0 ;
assign \add_17s_17s_17_2_1_U22.top_add_17s_17s_17_2_1_Adder_13_U.b  = \add_17s_17s_17_2_1_U22.din1 ;
assign \add_17s_17s_17_2_1_U22.top_add_17s_17s_17_2_1_Adder_13_U.ce  = \add_17s_17s_17_2_1_U22.ce ;
assign \add_17s_17s_17_2_1_U22.top_add_17s_17s_17_2_1_Adder_13_U.clk  = \add_17s_17s_17_2_1_U22.clk ;
assign \add_17s_17s_17_2_1_U22.top_add_17s_17s_17_2_1_Adder_13_U.reset  = \add_17s_17s_17_2_1_U22.reset ;
assign \add_17s_17s_17_2_1_U22.dout  = \add_17s_17s_17_2_1_U22.top_add_17s_17s_17_2_1_Adder_13_U.s ;
assign \add_17s_17s_17_2_1_U22.ce  = 1'h1;
assign \add_17s_17s_17_2_1_U22.clk  = ap_clk;
assign \add_17s_17s_17_2_1_U22.din0  = { add_ln69_1_reg_1188[2], add_ln69_1_reg_1188[2], add_ln69_1_reg_1188[2], add_ln69_1_reg_1188[2], add_ln69_1_reg_1188[2], add_ln69_1_reg_1188[2], add_ln69_1_reg_1188[2], add_ln69_1_reg_1188[2], add_ln69_1_reg_1188[2], add_ln69_1_reg_1188[2], add_ln69_1_reg_1188[2], add_ln69_1_reg_1188[2], add_ln69_1_reg_1188[2], add_ln69_1_reg_1188[2], add_ln69_1_reg_1188 };
assign \add_17s_17s_17_2_1_U22.din1  = { r_1_reg_1146[15], r_1_reg_1146 };
assign grp_fu_799_p2 = \add_17s_17s_17_2_1_U22.dout ;
assign \add_17s_17s_17_2_1_U22.reset  = ap_rst;
assign \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.ain_s0  = \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.a ;
assign \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.bin_s0  = \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.b ;
assign \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.s  = { \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.fas_s2 , \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.sum_s1  };
assign \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.u2.a  = \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.ain_s1 ;
assign \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.u2.b  = \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.bin_s1 ;
assign \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.u2.cin  = \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.carry_s1 ;
assign \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.facout_s2  = \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.u2.cout ;
assign \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.fas_s2  = \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.u2.s ;
assign \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.u1.a  = \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.a [5:0];
assign \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.u1.b  = \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.b [5:0];
assign \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.u1.cin  = 1'h0;
assign \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.facout_s1  = \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.u1.cout ;
assign \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.fas_s1  = \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.u1.s ;
assign \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.a  = \add_12ns_12s_12_2_1_U2.din0 ;
assign \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.b  = \add_12ns_12s_12_2_1_U2.din1 ;
assign \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.ce  = \add_12ns_12s_12_2_1_U2.ce ;
assign \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.clk  = \add_12ns_12s_12_2_1_U2.clk ;
assign \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.reset  = \add_12ns_12s_12_2_1_U2.reset ;
assign \add_12ns_12s_12_2_1_U2.dout  = \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.s ;
assign \add_12ns_12s_12_2_1_U2.ce  = 1'h1;
assign \add_12ns_12s_12_2_1_U2.clk  = ap_clk;
assign \add_12ns_12s_12_2_1_U2.din0  = { op_21_V_reg_824, 3'h0 };
assign \add_12ns_12s_12_2_1_U2.din1  = { op_10[3], op_10[3], op_10[3], op_10[3], op_10[3], op_10[3], op_10[3], op_10[3], op_10 };
assign grp_fu_260_p2 = \add_12ns_12s_12_2_1_U2.dout ;
assign \add_12ns_12s_12_2_1_U2.reset  = ap_rst;
assign \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.ain_s0  = \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.a ;
assign \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.bin_s0  = \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.b ;
assign \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.s  = { \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.fas_s2 , \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.sum_s1  };
assign \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.u2.a  = \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.ain_s1 ;
assign \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.u2.b  = \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.bin_s1 ;
assign \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.u2.cin  = \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.carry_s1 ;
assign \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.facout_s2  = \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.u2.cout ;
assign \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.fas_s2  = \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.u2.s ;
assign \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.u1.a  = \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.a [4:0];
assign \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.u1.b  = \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.b [4:0];
assign \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.u1.cin  = 1'h0;
assign \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.facout_s1  = \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.u1.cout ;
assign \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.fas_s1  = \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.u1.s ;
assign \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.a  = \add_10s_10ns_10_2_1_U3.din0 ;
assign \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.b  = \add_10s_10ns_10_2_1_U3.din1 ;
assign \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.ce  = \add_10s_10ns_10_2_1_U3.ce ;
assign \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.clk  = \add_10s_10ns_10_2_1_U3.clk ;
assign \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.reset  = \add_10s_10ns_10_2_1_U3.reset ;
assign \add_10s_10ns_10_2_1_U3.dout  = \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.s ;
assign \add_10s_10ns_10_2_1_U3.ce  = 1'h1;
assign \add_10s_10ns_10_2_1_U3.clk  = ap_clk;
assign \add_10s_10ns_10_2_1_U3.din0  = { tmp_1_reg_849[8], tmp_1_reg_849 };
assign \add_10s_10ns_10_2_1_U3.din1  = 10'h001;
assign grp_fu_289_p2 = \add_10s_10ns_10_2_1_U3.dout ;
assign \add_10s_10ns_10_2_1_U3.reset  = ap_rst;
assign \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.ain_s0  = \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.a ;
assign \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.bin_s0  = \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.b ;
assign \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.s  = { \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.fas_s2 , \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.sum_s1  };
assign \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.u2.a  = \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.ain_s1 ;
assign \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.u2.b  = \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.bin_s1 ;
assign \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.u2.cin  = \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.carry_s1 ;
assign \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.facout_s2  = \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.u2.cout ;
assign \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.fas_s2  = \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.u2.s ;
assign \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.u1.a  = \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.a [4:0];
assign \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.u1.b  = \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.b [4:0];
assign \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.u1.cin  = 1'h0;
assign \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.facout_s1  = \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.u1.cout ;
assign \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.fas_s1  = \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.u1.s ;
assign \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.a  = \add_10ns_10s_10_2_1_U4.din0 ;
assign \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.b  = \add_10ns_10s_10_2_1_U4.din1 ;
assign \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.ce  = \add_10ns_10s_10_2_1_U4.ce ;
assign \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.clk  = \add_10ns_10s_10_2_1_U4.clk ;
assign \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.reset  = \add_10ns_10s_10_2_1_U4.reset ;
assign \add_10ns_10s_10_2_1_U4.dout  = \add_10ns_10s_10_2_1_U4.top_add_10ns_10s_10_2_1_Adder_3_U.s ;
assign \add_10ns_10s_10_2_1_U4.ce  = 1'h1;
assign \add_10ns_10s_10_2_1_U4.clk  = ap_clk;
assign \add_10ns_10s_10_2_1_U4.din0  = ret_V_15_reg_877;
assign \add_10ns_10s_10_2_1_U4.din1  = { op_11_V_reg_872[3], op_11_V_reg_872[3], op_11_V_reg_872[3], op_11_V_reg_872[3], op_11_V_reg_872[3], op_11_V_reg_872[3], op_11_V_reg_872 };
assign grp_fu_331_p2 = \add_10ns_10s_10_2_1_U4.dout ;
assign \add_10ns_10s_10_2_1_U4.reset  = ap_rst;
endmodule


// Machine B:
// Processed by function `add_clk_enable_signal` in `verilog_tricks.py`.
// Processed by function `remove_reset_signal` in `verilog_tricks.py`.
module top_B (
  ap_clk,
  ap_start,
  ap_done,
  ap_idle,
  ap_ready,
  op_0,
  op_2,
  op_3,
  op_4,
  op_5,
  op_6,
  op_7,
  op_8,
  op_10,
  op_12,
  op_13,
  op_14,
  op_15,
  op_19,
  op_31,
  op_31_ap_vld,
clk_enable
);
input clk_enable;


input ap_clk;
wire ap_rst;
assign ap_rst = op_31_ap_vld;
input ap_start;
input [3:0] op_0;
input [3:0] op_10;
input [15:0] op_12;
input [15:0] op_13;
input [3:0] op_14;
input [7:0] op_15;
input [31:0] op_19;
input [7:0] op_2;
input [7:0] op_3;
input [15:0] op_4;
input [7:0] op_5;
input [3:0] op_6;
input [7:0] op_7;
input [3:0] op_8;
output ap_done;
output ap_idle;
output ap_ready;
output [31:0] op_31;
output op_31_ap_vld;


reg [31:0] add_ln691_1_reg_880;
reg [31:0] add_ln691_2_reg_911;
reg [31:0] add_ln691_3_reg_960;
reg [31:0] add_ln691_4_reg_986;
reg [16:0] add_ln69_2_reg_991;
reg [6:0] ap_CS_fsm = 7'h01;
reg icmp_ln851_2_reg_875;
reg icmp_ln851_3_reg_906;
reg icmp_ln851_4_reg_955;
reg icmp_ln851_reg_934;
reg [8:0] op_21_V_reg_848;
reg [9:0] op_23_V_reg_859;
reg [45:0] ret_V_16_reg_864;
reg [44:0] ret_V_17_reg_895;
reg [34:0] ret_V_18_reg_944;
reg [33:0] ret_V_19_reg_975;
reg [31:0] ret_V_21_cast_reg_869;
reg [31:0] ret_V_23_cast_reg_900;
reg [31:0] ret_V_25_cast_reg_949;
reg [31:0] ret_V_27_cast_reg_980;
reg [1:0] ret_V_3_reg_939;
reg [1:0] ret_V_reg_928;
reg [31:0] select_ln1358_reg_923;
reg [2:0] select_ln69_reg_965;
reg tmp_3_reg_885;
reg [8:0] ush_reg_890;
wire [31:0] _000_;
wire [31:0] _001_;
wire [31:0] _002_;
wire [31:0] _003_;
wire [16:0] _004_;
wire [6:0] _005_;
wire _006_;
wire _007_;
wire _008_;
wire _009_;
wire [8:0] _010_;
wire [9:0] _011_;
wire [45:0] _012_;
wire [44:0] _013_;
wire [34:0] _014_;
wire [33:0] _015_;
wire [31:0] _016_;
wire [31:0] _017_;
wire [31:0] _018_;
wire [31:0] _019_;
wire [1:0] _020_;
wire [1:0] _021_;
wire [31:0] _022_;
wire [2:0] _023_;
wire _024_;
wire [8:0] _025_;
wire [1:0] _026_;
wire _027_;
wire _028_;
wire _029_;
wire _030_;
wire _031_;
wire _032_;
wire _033_;
wire _034_;
wire _035_;
wire _036_;
wire _037_;
wire _038_;
wire _039_;
wire _040_;
wire _041_;
wire _042_;
wire [31:0] add_ln691_1_fu_385_p2;
wire [31:0] add_ln691_2_fu_484_p2;
wire [31:0] add_ln691_3_fu_659_p2;
wire [31:0] add_ln691_4_fu_780_p2;
wire [9:0] add_ln691_fu_312_p2;
wire [2:0] add_ln69_1_fu_794_p2;
wire [16:0] add_ln69_2_fu_803_p2;
wire [31:0] add_ln69_fu_832_p2;
wire and_ln353_fu_534_p2;
wire ap_CS_fsm_state1;
wire ap_CS_fsm_state2;
wire ap_CS_fsm_state3;
wire ap_CS_fsm_state4;
wire ap_CS_fsm_state5;
wire ap_CS_fsm_state6;
wire ap_CS_fsm_state7;
wire [6:0] ap_NS_fsm;
wire ap_clk;
wire ap_done;
wire ap_idle;
wire ap_ready;
wire ap_rst;
wire ap_start;
wire [31:0] ashr_ln1333_fu_553_p2;
wire [15:0] ashr_ln799_fu_697_p2;
wire [7:0] conv_i_i_i357_fu_549_p0;
wire [31:0] conv_i_i_i357_fu_549_p1;
wire icmp_ln850_fu_528_p2;
wire icmp_ln851_1_fu_306_p2;
wire icmp_ln851_2_fu_379_p2;
wire icmp_ln851_3_fu_478_p2;
wire icmp_ln851_4_fu_653_p2;
wire icmp_ln851_fu_586_p2;
wire [9:0] lhs_fu_490_p3;
wire [3:0] op_0;
wire [3:0] op_10;
wire [3:0] op_11_V_fu_257_p2;
wire [15:0] op_12;
wire [15:0] op_13;
wire [3:0] op_14;
wire [7:0] op_15;
wire [31:0] op_19;
wire [7:0] op_2;
wire [8:0] op_21_V_fu_243_p2;
wire [9:0] op_23_V_fu_338_p2;
wire [7:0] op_3;
wire [31:0] op_31;
wire op_31_ap_vld;
wire [15:0] op_4;
wire [7:0] op_5;
wire [3:0] op_6;
wire [7:0] op_7;
wire [3:0] op_8;
wire p_Result_1_fu_710_p3;
wire p_Result_2_fu_294_p3;
wire p_Result_3_fu_423_p3;
wire p_Result_4_fu_598_p3;
wire p_Result_5_fu_729_p3;
wire p_Result_6_fu_809_p3;
wire p_Result_7_fu_673_p3;
wire p_Result_s_fu_516_p3;
wire [15:0] r_1_fu_702_p3;
wire [7:0] r_fu_391_p2;
wire [9:0] ret_V_12_fu_502_p2;
wire ret_V_13_fu_540_p2;
wire [11:0] ret_V_14_fu_274_p2;
wire [9:0] ret_V_15_fu_326_p3;
wire [45:0] ret_V_16_fu_359_p2;
wire [44:0] ret_V_17_fu_458_p2;
wire [34:0] ret_V_18_fu_633_p2;
wire [33:0] ret_V_19_fu_764_p2;
wire [31:0] ret_V_20_fu_825_p3;
wire [31:0] ret_V_21_cast_fu_365_p4;
wire [31:0] ret_V_23_cast_fu_464_p4;
wire [31:0] ret_V_25_cast_fu_639_p4;
wire [31:0] ret_V_27_cast_fu_770_p4;
wire [1:0] ret_V_3_fu_592_p2;
wire [1:0] ret_V_4_fu_722_p3;
wire [1:0] ret_V_fu_572_p4;
wire [11:0] rhs_1_fu_267_p3;
wire [43:0] rhs_3_fu_446_p3;
wire [33:0] rhs_4_fu_621_p3;
wire [32:0] rhs_5_fu_752_p3;
wire [31:0] select_ln1358_fu_565_p3;
wire [31:0] select_ln353_1_fu_614_p3;
wire [31:0] select_ln353_2_fu_745_p3;
wire [31:0] select_ln353_fu_439_p3;
wire [2:0] select_ln69_fu_665_p3;
wire [9:0] select_ln850_2_fu_318_p3;
wire [31:0] select_ln850_3_fu_434_p3;
wire [31:0] select_ln850_4_fu_609_p3;
wire [31:0] select_ln850_5_fu_740_p3;
wire [31:0] select_ln850_6_fu_819_p3;
wire [1:0] select_ln850_fu_717_p3;
wire [45:0] sext_ln1192_1_fu_355_p1;
wire [44:0] sext_ln1192_2_fu_454_p1;
wire [34:0] sext_ln1192_3_fu_629_p1;
wire [33:0] sext_ln1192_4_fu_760_p1;
wire [3:0] sext_ln1192_fu_263_p0;
wire [11:0] sext_ln1192_fu_263_p1;
wire [31:0] sext_ln1357_fu_546_p1;
wire [8:0] sext_ln15_fu_397_p1;
wire [8:0] sext_ln20_fu_235_p1;
wire [9:0] sext_ln69_1_fu_334_p1;
wire [16:0] sext_ln69_2_fu_786_p1;
wire [2:0] sext_ln69_3_fu_790_p1;
wire [16:0] sext_ln69_4_fu_799_p1;
wire [31:0] sext_ln69_5_fu_838_p1;
wire [8:0] sext_ln69_fu_239_p1;
wire [15:0] sext_ln703_1_fu_344_p0;
wire [45:0] sext_ln703_1_fu_344_p1;
wire [15:0] sext_ln703_2_fu_430_p0;
wire [44:0] sext_ln703_2_fu_430_p1;
wire [3:0] sext_ln703_3_fu_605_p0;
wire [34:0] sext_ln703_3_fu_605_p1;
wire [7:0] sext_ln703_4_fu_736_p0;
wire [33:0] sext_ln703_4_fu_736_p1;
wire [7:0] sext_ln703_fu_498_p0;
wire [9:0] sext_ln703_fu_498_p1;
wire [9:0] sext_ln850_fu_290_p1;
wire [3:0] sh_fu_680_p2;
wire [31:0] shl_ln1299_fu_559_p2;
wire [15:0] shl_ln781_fu_689_p2;
wire [8:0] sub_ln1357_fu_409_p2;
wire [8:0] tmp_1_fu_280_p4;
wire tmp_3_fu_401_p3;
wire [22:0] tmp_6_fu_348_p3;
wire tmp_fu_508_p3;
wire [3:0] trunc_ln1350_1_fu_253_p1;
wire [3:0] trunc_ln1350_fu_249_p1;
wire [5:0] trunc_ln851_1_fu_582_p1;
wire [3:0] trunc_ln851_2_fu_302_p0;
wire [2:0] trunc_ln851_2_fu_302_p1;
wire [15:0] trunc_ln851_3_fu_375_p0;
wire [12:0] trunc_ln851_3_fu_375_p1;
wire [15:0] trunc_ln851_4_fu_474_p0;
wire [11:0] trunc_ln851_4_fu_474_p1;
wire [3:0] trunc_ln851_5_fu_649_p0;
wire [1:0] trunc_ln851_5_fu_649_p1;
wire [7:0] trunc_ln851_6_fu_816_p0;
wire trunc_ln851_6_fu_816_p1;
wire [5:0] trunc_ln851_fu_524_p1;
wire [8:0] ush_fu_415_p3;
wire [15:0] zext_ln781_fu_685_p1;
wire [15:0] zext_ln799_fu_694_p1;


assign add_ln691_1_fu_385_p2 = { ret_V_16_fu_359_p2[45], ret_V_16_fu_359_p2[45], ret_V_16_fu_359_p2[45], ret_V_16_fu_359_p2[45], ret_V_16_fu_359_p2[45], ret_V_16_fu_359_p2[45], ret_V_16_fu_359_p2[45], ret_V_16_fu_359_p2[45], ret_V_16_fu_359_p2[45], ret_V_16_fu_359_p2[45], ret_V_16_fu_359_p2[45], ret_V_16_fu_359_p2[45], ret_V_16_fu_359_p2[45], ret_V_16_fu_359_p2[45], ret_V_16_fu_359_p2[45], ret_V_16_fu_359_p2[45], ret_V_16_fu_359_p2[45], ret_V_16_fu_359_p2[45], ret_V_16_fu_359_p2[45], ret_V_16_fu_359_p2[45], ret_V_16_fu_359_p2[45], ret_V_16_fu_359_p2[45], ret_V_16_fu_359_p2[22:13] } + 1'h1;
assign add_ln691_2_fu_484_p2 = ret_V_17_fu_458_p2[43:12] + 1'h1;
assign add_ln691_3_fu_659_p2 = ret_V_18_fu_633_p2[33:2] + 1'h1;
assign add_ln691_4_fu_780_p2 = ret_V_19_fu_764_p2[32:1] + 1'h1;
assign add_ln691_fu_312_p2 = $signed(ret_V_14_fu_274_p2[11:3]) + $signed(2'h1);
assign add_ln69_1_fu_794_p2 = $signed(ret_V_4_fu_722_p3) + $signed(select_ln69_reg_965);
assign add_ln69_2_fu_803_p2 = $signed(add_ln69_1_fu_794_p2) + $signed(r_1_fu_702_p3);
assign add_ln69_fu_832_p2 = ret_V_20_fu_825_p3 + op_19;
assign op_21_V_fu_243_p2 = $signed(op_5) + $signed(op_8);
assign op_23_V_fu_338_p2 = $signed(ret_V_15_fu_326_p3) + $signed(op_11_V_fu_257_p2);
assign op_31 = $signed(add_ln69_2_reg_991) + $signed(add_ln69_fu_832_p2);
assign ret_V_14_fu_274_p2 = $signed({ op_21_V_reg_848, 3'h0 }) + $signed(op_10);
assign { ret_V_16_fu_359_p2[45], ret_V_16_fu_359_p2[22:0] } = $signed({ op_23_V_reg_859, 13'h0000 }) + $signed(op_12);
assign ret_V_17_fu_458_p2 = $signed({ select_ln353_fu_439_p3, 12'h000 }) + $signed(op_13);
assign ret_V_18_fu_633_p2 = $signed({ select_ln353_1_fu_614_p3, 2'h0 }) + $signed(op_14);
assign ret_V_19_fu_764_p2 = $signed({ select_ln353_2_fu_745_p3, 1'h0 }) + $signed(op_15);
assign ret_V_3_fu_592_p2 = select_ln1358_fu_565_p3[7:6] + 1'h1;
assign _027_ = ap_CS_fsm[0] & _029_;
assign _028_ = ap_CS_fsm[0] & ap_start;
assign and_ln353_fu_534_p2 = ret_V_12_fu_502_p2[9] & icmp_ln850_fu_528_p2;
assign ret_V_12_fu_502_p2 = { op_7[7], op_7[7], op_7 } & { op_6, 6'h00 };
assign r_fu_391_p2 = ~ op_3;
assign _029_ = ~ ap_start;
assign _030_ = ! select_ln1358_fu_565_p3[5:0];
assign _031_ = | ret_V_12_fu_502_p2[5:0];
assign _032_ = | op_10[2:0];
assign _033_ = | op_12[12:0];
assign _034_ = | op_13[11:0];
assign _035_ = | op_14[1:0];
always @(posedge ap_clk)
op_23_V_reg_859 <= _011_;
always @(posedge ap_clk)
op_21_V_reg_848 <= _010_;
always @(posedge ap_clk)
ret_V_19_reg_975 <= _015_;
always @(posedge ap_clk)
ret_V_27_cast_reg_980 <= _019_;
always @(posedge ap_clk)
add_ln691_4_reg_986 <= _003_;
always @(posedge ap_clk)
add_ln69_2_reg_991 <= _004_;
always @(posedge ap_clk)
select_ln1358_reg_923 <= _022_;
always @(posedge ap_clk)
ret_V_reg_928 <= _021_;
always @(posedge ap_clk)
icmp_ln851_reg_934 <= _009_;
always @(posedge ap_clk)
ret_V_3_reg_939 <= _020_;
always @(posedge ap_clk)
ret_V_18_reg_944 <= _014_;
always @(posedge ap_clk)
ret_V_25_cast_reg_949 <= _018_;
always @(posedge ap_clk)
icmp_ln851_4_reg_955 <= _008_;
always @(posedge ap_clk)
add_ln691_3_reg_960 <= _002_;
always @(posedge ap_clk)
select_ln69_reg_965 <= _023_;
always @(posedge ap_clk)
tmp_3_reg_885 <= _024_;
always @(posedge ap_clk)
ush_reg_890 <= _025_;
always @(posedge ap_clk)
ret_V_17_reg_895 <= _013_;
always @(posedge ap_clk)
ret_V_23_cast_reg_900 <= _017_;
always @(posedge ap_clk)
icmp_ln851_3_reg_906 <= _007_;
always @(posedge ap_clk)
add_ln691_2_reg_911 <= _001_;
always @(posedge ap_clk)
ret_V_16_reg_864 <= _012_;
always @(posedge ap_clk)
ret_V_21_cast_reg_869 <= _016_;
always @(posedge ap_clk)
icmp_ln851_2_reg_875 <= _006_;
always @(posedge ap_clk)
add_ln691_1_reg_880 <= _000_;
always @(posedge ap_clk)
ap_CS_fsm <= _005_;
assign _026_ = _028_ ? 2'h2 : 2'h1;
assign _036_ = ap_CS_fsm == 1'h1;
function [6:0] _100_;
input [6:0] a;
input [48:0] b;
input [6:0] s;
case (s)
7'b0000001:
_100_ = b[6:0];
7'b0000010:
_100_ = b[13:7];
7'b0000100:
_100_ = b[20:14];
7'b0001000:
_100_ = b[27:21];
7'b0010000:
_100_ = b[34:28];
7'b0100000:
_100_ = b[41:35];
7'b1000000:
_100_ = b[48:42];
7'b0000000:
_100_ = a;
default:
_100_ = 7'bx;
endcase
endfunction
assign ap_NS_fsm = _100_(7'hxx, { 5'h00, _026_, 42'h02082082001 }, { _036_, _042_, _041_, _040_, _039_, _038_, _037_ });
assign _037_ = ap_CS_fsm == 7'h40;
assign _038_ = ap_CS_fsm == 6'h20;
assign _039_ = ap_CS_fsm == 5'h10;
assign _040_ = ap_CS_fsm == 4'h8;
assign _041_ = ap_CS_fsm == 3'h4;
assign _042_ = ap_CS_fsm == 2'h2;
assign op_31_ap_vld = ap_CS_fsm[6] ? 1'h1 : 1'h0;
assign ap_idle = _027_ ? 1'h1 : 1'h0;
assign _011_ = ap_CS_fsm[1] ? op_23_V_fu_338_p2 : op_23_V_reg_859;
assign _010_ = ap_CS_fsm[0] ? op_21_V_fu_243_p2 : op_21_V_reg_848;
assign _004_ = ap_CS_fsm[5] ? add_ln69_2_fu_803_p2 : add_ln69_2_reg_991;
assign _003_ = ap_CS_fsm[5] ? add_ln691_4_fu_780_p2 : add_ln691_4_reg_986;
assign _019_ = ap_CS_fsm[5] ? ret_V_19_fu_764_p2[32:1] : ret_V_27_cast_reg_980;
assign _015_ = ap_CS_fsm[5] ? ret_V_19_fu_764_p2 : ret_V_19_reg_975;
assign _023_ = ap_CS_fsm[4] ? select_ln69_fu_665_p3 : select_ln69_reg_965;
assign _002_ = ap_CS_fsm[4] ? add_ln691_3_fu_659_p2 : add_ln691_3_reg_960;
assign _008_ = ap_CS_fsm[4] ? icmp_ln851_4_fu_653_p2 : icmp_ln851_4_reg_955;
assign _018_ = ap_CS_fsm[4] ? ret_V_18_fu_633_p2[33:2] : ret_V_25_cast_reg_949;
assign _014_ = ap_CS_fsm[4] ? ret_V_18_fu_633_p2 : ret_V_18_reg_944;
assign _020_ = ap_CS_fsm[4] ? ret_V_3_fu_592_p2 : ret_V_3_reg_939;
assign _009_ = ap_CS_fsm[4] ? icmp_ln851_fu_586_p2 : icmp_ln851_reg_934;
assign _021_ = ap_CS_fsm[4] ? select_ln1358_fu_565_p3[7:6] : ret_V_reg_928;
assign _022_ = ap_CS_fsm[4] ? select_ln1358_fu_565_p3 : select_ln1358_reg_923;
assign _001_ = ap_CS_fsm[3] ? add_ln691_2_fu_484_p2 : add_ln691_2_reg_911;
assign _007_ = ap_CS_fsm[3] ? icmp_ln851_3_fu_478_p2 : icmp_ln851_3_reg_906;
assign _017_ = ap_CS_fsm[3] ? ret_V_17_fu_458_p2[43:12] : ret_V_23_cast_reg_900;
assign _013_ = ap_CS_fsm[3] ? ret_V_17_fu_458_p2 : ret_V_17_reg_895;
assign _025_ = ap_CS_fsm[3] ? ush_fu_415_p3 : ush_reg_890;
assign _024_ = ap_CS_fsm[3] ? op_3[7] : tmp_3_reg_885;
assign _000_ = ap_CS_fsm[2] ? add_ln691_1_fu_385_p2 : add_ln691_1_reg_880;
assign _006_ = ap_CS_fsm[2] ? icmp_ln851_2_fu_379_p2 : icmp_ln851_2_reg_875;
assign _016_ = ap_CS_fsm[2] ? { ret_V_16_fu_359_p2[45], ret_V_16_fu_359_p2[45], ret_V_16_fu_359_p2[45], ret_V_16_fu_359_p2[45], ret_V_16_fu_359_p2[45], ret_V_16_fu_359_p2[45], ret_V_16_fu_359_p2[45], ret_V_16_fu_359_p2[45], ret_V_16_fu_359_p2[45], ret_V_16_fu_359_p2[45], ret_V_16_fu_359_p2[45], ret_V_16_fu_359_p2[45], ret_V_16_fu_359_p2[45], ret_V_16_fu_359_p2[45], ret_V_16_fu_359_p2[45], ret_V_16_fu_359_p2[45], ret_V_16_fu_359_p2[45], ret_V_16_fu_359_p2[45], ret_V_16_fu_359_p2[45], ret_V_16_fu_359_p2[45], ret_V_16_fu_359_p2[45], ret_V_16_fu_359_p2[45], ret_V_16_fu_359_p2[22:13] } : ret_V_21_cast_reg_869;
assign _012_ = ap_CS_fsm[2] ? { ret_V_16_fu_359_p2[45], ret_V_16_fu_359_p2[45], ret_V_16_fu_359_p2[45], ret_V_16_fu_359_p2[45], ret_V_16_fu_359_p2[45], ret_V_16_fu_359_p2[45], ret_V_16_fu_359_p2[45], ret_V_16_fu_359_p2[45], ret_V_16_fu_359_p2[45], ret_V_16_fu_359_p2[45], ret_V_16_fu_359_p2[45], ret_V_16_fu_359_p2[45], ret_V_16_fu_359_p2[45], ret_V_16_fu_359_p2[45], ret_V_16_fu_359_p2[45], ret_V_16_fu_359_p2[45], ret_V_16_fu_359_p2[45], ret_V_16_fu_359_p2[45], ret_V_16_fu_359_p2[45], ret_V_16_fu_359_p2[45], ret_V_16_fu_359_p2[45], ret_V_16_fu_359_p2[45], ret_V_16_fu_359_p2[45], ret_V_16_fu_359_p2[22:0] } : ret_V_16_reg_864;
assign _005_ = ap_rst ? 7'h01 : ap_NS_fsm;
assign shl_ln1299_fu_559_p2 = $signed(op_7) << { ush_reg_890[8], ush_reg_890[8], ush_reg_890[8], ush_reg_890[8], ush_reg_890[8], ush_reg_890[8], ush_reg_890[8], ush_reg_890[8], ush_reg_890[8], ush_reg_890[8], ush_reg_890[8], ush_reg_890[8], ush_reg_890[8], ush_reg_890[8], ush_reg_890[8], ush_reg_890[8], ush_reg_890[8], ush_reg_890[8], ush_reg_890[8], ush_reg_890[8], ush_reg_890[8], ush_reg_890[8], ush_reg_890[8], ush_reg_890 };
assign shl_ln781_fu_689_p2 = op_4 << sh_fu_680_p2;
assign ashr_ln1333_fu_553_p2 = $signed(op_7) >>> { ush_reg_890[8], ush_reg_890[8], ush_reg_890[8], ush_reg_890[8], ush_reg_890[8], ush_reg_890[8], ush_reg_890[8], ush_reg_890[8], ush_reg_890[8], ush_reg_890[8], ush_reg_890[8], ush_reg_890[8], ush_reg_890[8], ush_reg_890[8], ush_reg_890[8], ush_reg_890[8], ush_reg_890[8], ush_reg_890[8], ush_reg_890[8], ush_reg_890[8], ush_reg_890[8], ush_reg_890[8], ush_reg_890[8], ush_reg_890 };
assign ashr_ln799_fu_697_p2 = $signed(op_4) >>> op_6;
assign sh_fu_680_p2 = 1'h0 - op_6;
assign sub_ln1357_fu_409_p2 = $signed(1'h0) - $signed(r_fu_391_p2);
assign icmp_ln850_fu_528_p2 = _031_ ? 1'h1 : 1'h0;
assign icmp_ln851_1_fu_306_p2 = _032_ ? 1'h1 : 1'h0;
assign icmp_ln851_2_fu_379_p2 = _033_ ? 1'h1 : 1'h0;
assign icmp_ln851_3_fu_478_p2 = _034_ ? 1'h1 : 1'h0;
assign icmp_ln851_4_fu_653_p2 = _035_ ? 1'h1 : 1'h0;
assign icmp_ln851_fu_586_p2 = _030_ ? 1'h1 : 1'h0;
assign r_1_fu_702_p3 = op_6[3] ? shl_ln781_fu_689_p2 : ashr_ln799_fu_697_p2;
assign ret_V_15_fu_326_p3 = ret_V_14_fu_274_p2[11] ? select_ln850_2_fu_318_p3 : { 2'h0, ret_V_14_fu_274_p2[10:3] };
assign ret_V_20_fu_825_p3 = ret_V_19_reg_975[33] ? select_ln850_6_fu_819_p3 : ret_V_27_cast_reg_980;
assign ret_V_4_fu_722_p3 = select_ln1358_reg_923[7] ? select_ln850_fu_717_p3 : ret_V_reg_928;
assign select_ln1358_fu_565_p3 = tmp_3_reg_885 ? shl_ln1299_fu_559_p2 : ashr_ln1333_fu_553_p2;
assign select_ln353_1_fu_614_p3 = ret_V_17_reg_895[44] ? select_ln850_4_fu_609_p3 : ret_V_23_cast_reg_900;
assign select_ln353_2_fu_745_p3 = ret_V_18_reg_944[34] ? select_ln850_5_fu_740_p3 : ret_V_25_cast_reg_949;
assign select_ln353_fu_439_p3 = ret_V_16_reg_864[45] ? select_ln850_3_fu_434_p3 : ret_V_21_cast_reg_869;
assign select_ln69_fu_665_p3 = ret_V_13_fu_540_p2 ? 3'h7 : 3'h0;
assign select_ln850_2_fu_318_p3 = icmp_ln851_1_fu_306_p2 ? add_ln691_fu_312_p2 : { 2'h3, ret_V_14_fu_274_p2[10:3] };
assign select_ln850_3_fu_434_p3 = icmp_ln851_2_reg_875 ? add_ln691_1_reg_880 : ret_V_21_cast_reg_869;
assign select_ln850_4_fu_609_p3 = icmp_ln851_3_reg_906 ? add_ln691_2_reg_911 : ret_V_23_cast_reg_900;
assign select_ln850_5_fu_740_p3 = icmp_ln851_4_reg_955 ? add_ln691_3_reg_960 : ret_V_25_cast_reg_949;
assign select_ln850_6_fu_819_p3 = op_15[0] ? add_ln691_4_reg_986 : ret_V_27_cast_reg_980;
assign select_ln850_fu_717_p3 = icmp_ln851_reg_934 ? ret_V_reg_928 : ret_V_3_reg_939;
assign ush_fu_415_p3 = op_3[7] ? { r_fu_391_p2[7], r_fu_391_p2 } : sub_ln1357_fu_409_p2;
assign op_11_V_fu_257_p2 = op_2[3:0] ^ op_4[3:0];
assign ret_V_13_fu_540_p2 = ret_V_12_fu_502_p2[6] ^ and_ln353_fu_534_p2;
assign ap_CS_fsm_state1 = ap_CS_fsm[0];
assign ap_CS_fsm_state2 = ap_CS_fsm[1];
assign ap_CS_fsm_state3 = ap_CS_fsm[2];
assign ap_CS_fsm_state4 = ap_CS_fsm[3];
assign ap_CS_fsm_state5 = ap_CS_fsm[4];
assign ap_CS_fsm_state6 = ap_CS_fsm[5];
assign ap_CS_fsm_state7 = ap_CS_fsm[6];
assign ap_done = op_31_ap_vld;
assign ap_ready = op_31_ap_vld;
assign conv_i_i_i357_fu_549_p0 = op_7;
assign conv_i_i_i357_fu_549_p1 = { op_7[7], op_7[7], op_7[7], op_7[7], op_7[7], op_7[7], op_7[7], op_7[7], op_7[7], op_7[7], op_7[7], op_7[7], op_7[7], op_7[7], op_7[7], op_7[7], op_7[7], op_7[7], op_7[7], op_7[7], op_7[7], op_7[7], op_7[7], op_7[7], op_7 };
assign lhs_fu_490_p3 = { op_6, 6'h00 };
assign p_Result_1_fu_710_p3 = select_ln1358_reg_923[7];
assign p_Result_2_fu_294_p3 = ret_V_14_fu_274_p2[11];
assign p_Result_3_fu_423_p3 = ret_V_16_reg_864[45];
assign p_Result_4_fu_598_p3 = ret_V_17_reg_895[44];
assign p_Result_5_fu_729_p3 = ret_V_18_reg_944[34];
assign p_Result_6_fu_809_p3 = ret_V_19_reg_975[33];
assign p_Result_7_fu_673_p3 = op_6[3];
assign p_Result_s_fu_516_p3 = ret_V_12_fu_502_p2[9];
assign ret_V_16_fu_359_p2[44:23] = { ret_V_16_fu_359_p2[45], ret_V_16_fu_359_p2[45], ret_V_16_fu_359_p2[45], ret_V_16_fu_359_p2[45], ret_V_16_fu_359_p2[45], ret_V_16_fu_359_p2[45], ret_V_16_fu_359_p2[45], ret_V_16_fu_359_p2[45], ret_V_16_fu_359_p2[45], ret_V_16_fu_359_p2[45], ret_V_16_fu_359_p2[45], ret_V_16_fu_359_p2[45], ret_V_16_fu_359_p2[45], ret_V_16_fu_359_p2[45], ret_V_16_fu_359_p2[45], ret_V_16_fu_359_p2[45], ret_V_16_fu_359_p2[45], ret_V_16_fu_359_p2[45], ret_V_16_fu_359_p2[45], ret_V_16_fu_359_p2[45], ret_V_16_fu_359_p2[45], ret_V_16_fu_359_p2[45] };
assign ret_V_21_cast_fu_365_p4 = { ret_V_16_fu_359_p2[45], ret_V_16_fu_359_p2[45], ret_V_16_fu_359_p2[45], ret_V_16_fu_359_p2[45], ret_V_16_fu_359_p2[45], ret_V_16_fu_359_p2[45], ret_V_16_fu_359_p2[45], ret_V_16_fu_359_p2[45], ret_V_16_fu_359_p2[45], ret_V_16_fu_359_p2[45], ret_V_16_fu_359_p2[45], ret_V_16_fu_359_p2[45], ret_V_16_fu_359_p2[45], ret_V_16_fu_359_p2[45], ret_V_16_fu_359_p2[45], ret_V_16_fu_359_p2[45], ret_V_16_fu_359_p2[45], ret_V_16_fu_359_p2[45], ret_V_16_fu_359_p2[45], ret_V_16_fu_359_p2[45], ret_V_16_fu_359_p2[45], ret_V_16_fu_359_p2[45], ret_V_16_fu_359_p2[22:13] };
assign ret_V_23_cast_fu_464_p4 = ret_V_17_fu_458_p2[43:12];
assign ret_V_25_cast_fu_639_p4 = ret_V_18_fu_633_p2[33:2];
assign ret_V_27_cast_fu_770_p4 = ret_V_19_fu_764_p2[32:1];
assign ret_V_fu_572_p4 = select_ln1358_fu_565_p3[7:6];
assign rhs_1_fu_267_p3 = { op_21_V_reg_848, 3'h0 };
assign rhs_3_fu_446_p3 = { select_ln353_fu_439_p3, 12'h000 };
assign rhs_4_fu_621_p3 = { select_ln353_1_fu_614_p3, 2'h0 };
assign rhs_5_fu_752_p3 = { select_ln353_2_fu_745_p3, 1'h0 };
assign sext_ln1192_1_fu_355_p1 = { op_23_V_reg_859[9], op_23_V_reg_859[9], op_23_V_reg_859[9], op_23_V_reg_859[9], op_23_V_reg_859[9], op_23_V_reg_859[9], op_23_V_reg_859[9], op_23_V_reg_859[9], op_23_V_reg_859[9], op_23_V_reg_859[9], op_23_V_reg_859[9], op_23_V_reg_859[9], op_23_V_reg_859[9], op_23_V_reg_859[9], op_23_V_reg_859[9], op_23_V_reg_859[9], op_23_V_reg_859[9], op_23_V_reg_859[9], op_23_V_reg_859[9], op_23_V_reg_859[9], op_23_V_reg_859[9], op_23_V_reg_859[9], op_23_V_reg_859[9], op_23_V_reg_859, 13'h0000 };
assign sext_ln1192_2_fu_454_p1 = { select_ln353_fu_439_p3[31], select_ln353_fu_439_p3, 12'h000 };
assign sext_ln1192_3_fu_629_p1 = { select_ln353_1_fu_614_p3[31], select_ln353_1_fu_614_p3, 2'h0 };
assign sext_ln1192_4_fu_760_p1 = { select_ln353_2_fu_745_p3[31], select_ln353_2_fu_745_p3, 1'h0 };
assign sext_ln1192_fu_263_p0 = op_10;
assign sext_ln1192_fu_263_p1 = { op_10[3], op_10[3], op_10[3], op_10[3], op_10[3], op_10[3], op_10[3], op_10[3], op_10 };
assign sext_ln1357_fu_546_p1 = { ush_reg_890[8], ush_reg_890[8], ush_reg_890[8], ush_reg_890[8], ush_reg_890[8], ush_reg_890[8], ush_reg_890[8], ush_reg_890[8], ush_reg_890[8], ush_reg_890[8], ush_reg_890[8], ush_reg_890[8], ush_reg_890[8], ush_reg_890[8], ush_reg_890[8], ush_reg_890[8], ush_reg_890[8], ush_reg_890[8], ush_reg_890[8], ush_reg_890[8], ush_reg_890[8], ush_reg_890[8], ush_reg_890[8], ush_reg_890 };
assign sext_ln15_fu_397_p1 = { r_fu_391_p2[7], r_fu_391_p2 };
assign sext_ln20_fu_235_p1 = { op_5[7], op_5 };
assign sext_ln69_1_fu_334_p1 = { op_11_V_fu_257_p2[3], op_11_V_fu_257_p2[3], op_11_V_fu_257_p2[3], op_11_V_fu_257_p2[3], op_11_V_fu_257_p2[3], op_11_V_fu_257_p2[3], op_11_V_fu_257_p2 };
assign sext_ln69_2_fu_786_p1 = { r_1_fu_702_p3[15], r_1_fu_702_p3 };
assign sext_ln69_3_fu_790_p1 = { ret_V_4_fu_722_p3[1], ret_V_4_fu_722_p3 };
assign sext_ln69_4_fu_799_p1 = { add_ln69_1_fu_794_p2[2], add_ln69_1_fu_794_p2[2], add_ln69_1_fu_794_p2[2], add_ln69_1_fu_794_p2[2], add_ln69_1_fu_794_p2[2], add_ln69_1_fu_794_p2[2], add_ln69_1_fu_794_p2[2], add_ln69_1_fu_794_p2[2], add_ln69_1_fu_794_p2[2], add_ln69_1_fu_794_p2[2], add_ln69_1_fu_794_p2[2], add_ln69_1_fu_794_p2[2], add_ln69_1_fu_794_p2[2], add_ln69_1_fu_794_p2[2], add_ln69_1_fu_794_p2 };
assign sext_ln69_5_fu_838_p1 = { add_ln69_2_reg_991[16], add_ln69_2_reg_991[16], add_ln69_2_reg_991[16], add_ln69_2_reg_991[16], add_ln69_2_reg_991[16], add_ln69_2_reg_991[16], add_ln69_2_reg_991[16], add_ln69_2_reg_991[16], add_ln69_2_reg_991[16], add_ln69_2_reg_991[16], add_ln69_2_reg_991[16], add_ln69_2_reg_991[16], add_ln69_2_reg_991[16], add_ln69_2_reg_991[16], add_ln69_2_reg_991[16], add_ln69_2_reg_991 };
assign sext_ln69_fu_239_p1 = { op_8[3], op_8[3], op_8[3], op_8[3], op_8[3], op_8 };
assign sext_ln703_1_fu_344_p0 = op_12;
assign sext_ln703_1_fu_344_p1 = { op_12[15], op_12[15], op_12[15], op_12[15], op_12[15], op_12[15], op_12[15], op_12[15], op_12[15], op_12[15], op_12[15], op_12[15], op_12[15], op_12[15], op_12[15], op_12[15], op_12[15], op_12[15], op_12[15], op_12[15], op_12[15], op_12[15], op_12[15], op_12[15], op_12[15], op_12[15], op_12[15], op_12[15], op_12[15], op_12[15], op_12 };
assign sext_ln703_2_fu_430_p0 = op_13;
assign sext_ln703_2_fu_430_p1 = { op_13[15], op_13[15], op_13[15], op_13[15], op_13[15], op_13[15], op_13[15], op_13[15], op_13[15], op_13[15], op_13[15], op_13[15], op_13[15], op_13[15], op_13[15], op_13[15], op_13[15], op_13[15], op_13[15], op_13[15], op_13[15], op_13[15], op_13[15], op_13[15], op_13[15], op_13[15], op_13[15], op_13[15], op_13[15], op_13 };
assign sext_ln703_3_fu_605_p0 = op_14;
assign sext_ln703_3_fu_605_p1 = { op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14 };
assign sext_ln703_4_fu_736_p0 = op_15;
assign sext_ln703_4_fu_736_p1 = { op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15 };
assign sext_ln703_fu_498_p0 = op_7;
assign sext_ln703_fu_498_p1 = { op_7[7], op_7[7], op_7 };
assign sext_ln850_fu_290_p1 = { ret_V_14_fu_274_p2[11], ret_V_14_fu_274_p2[11:3] };
assign tmp_1_fu_280_p4 = ret_V_14_fu_274_p2[11:3];
assign tmp_3_fu_401_p3 = op_3[7];
assign tmp_6_fu_348_p3 = { op_23_V_reg_859, 13'h0000 };
assign tmp_fu_508_p3 = ret_V_12_fu_502_p2[6];
assign trunc_ln1350_1_fu_253_p1 = op_4[3:0];
assign trunc_ln1350_fu_249_p1 = op_2[3:0];
assign trunc_ln851_1_fu_582_p1 = select_ln1358_fu_565_p3[5:0];
assign trunc_ln851_2_fu_302_p0 = op_10;
assign trunc_ln851_2_fu_302_p1 = op_10[2:0];
assign trunc_ln851_3_fu_375_p0 = op_12;
assign trunc_ln851_3_fu_375_p1 = op_12[12:0];
assign trunc_ln851_4_fu_474_p0 = op_13;
assign trunc_ln851_4_fu_474_p1 = op_13[11:0];
assign trunc_ln851_5_fu_649_p0 = op_14;
assign trunc_ln851_5_fu_649_p1 = op_14[1:0];
assign trunc_ln851_6_fu_816_p0 = op_15;
assign trunc_ln851_6_fu_816_p1 = op_15[0];
assign trunc_ln851_fu_524_p1 = ret_V_12_fu_502_p2[5:0];
assign zext_ln781_fu_685_p1 = { 12'h000, sh_fu_680_p2 };
assign zext_ln799_fu_694_p1 = { 12'h000, op_6 };
endmodule


// Product machine:
module top_A_times_top_B (ap_start, op_0, op_10, op_12, op_13, op_14, op_15, op_19, op_2, op_3, op_4, op_5, op_6, op_7, op_8, ap_clk, unsafe_signal);
input ap_start;
input [3:0] op_0;
input [3:0] op_10;
input [15:0] op_12;
input [15:0] op_13;
input [3:0] op_14;
input [7:0] op_15;
input [31:0] op_19;
input [7:0] op_2;
input [7:0] op_3;
input [15:0] op_4;
input [7:0] op_5;
input [3:0] op_6;
input [7:0] op_7;
input [3:0] op_8;
input ap_clk;
output unsafe_signal;
reg _setup;
initial _setup = 1'b0;
always @ (posedge ap_clk) _setup <= 1'b1;
reg ap_start_internal;
always @ (posedge ap_clk) if (!_setup) ap_start_internal <= ap_start;
reg [3:0] op_0_internal;
always @ (posedge ap_clk) if (!_setup) op_0_internal <= op_0;
reg [3:0] op_10_internal;
always @ (posedge ap_clk) if (!_setup) op_10_internal <= op_10;
reg [15:0] op_12_internal;
always @ (posedge ap_clk) if (!_setup) op_12_internal <= op_12;
reg [15:0] op_13_internal;
always @ (posedge ap_clk) if (!_setup) op_13_internal <= op_13;
reg [3:0] op_14_internal;
always @ (posedge ap_clk) if (!_setup) op_14_internal <= op_14;
reg [7:0] op_15_internal;
always @ (posedge ap_clk) if (!_setup) op_15_internal <= op_15;
reg [31:0] op_19_internal;
always @ (posedge ap_clk) if (!_setup) op_19_internal <= op_19;
reg [7:0] op_2_internal;
always @ (posedge ap_clk) if (!_setup) op_2_internal <= op_2;
reg [7:0] op_3_internal;
always @ (posedge ap_clk) if (!_setup) op_3_internal <= op_3;
reg [15:0] op_4_internal;
always @ (posedge ap_clk) if (!_setup) op_4_internal <= op_4;
reg [7:0] op_5_internal;
always @ (posedge ap_clk) if (!_setup) op_5_internal <= op_5;
reg [3:0] op_6_internal;
always @ (posedge ap_clk) if (!_setup) op_6_internal <= op_6;
reg [7:0] op_7_internal;
always @ (posedge ap_clk) if (!_setup) op_7_internal <= op_7;
reg [3:0] op_8_internal;
always @ (posedge ap_clk) if (!_setup) op_8_internal <= op_8;
wire ap_done_A;
wire ap_done_B;
wire ap_done_eq;
assign ap_done_eq = ap_done_A == ap_done_B;
wire ap_idle_A;
wire ap_idle_B;
wire ap_idle_eq;
assign ap_idle_eq = ap_idle_A == ap_idle_B;
wire ap_ready_A;
wire ap_ready_B;
wire ap_ready_eq;
assign ap_ready_eq = ap_ready_A == ap_ready_B;
wire [31:0] op_31_A;
wire [31:0] op_31_B;
wire op_31_eq;
assign op_31_eq = op_31_A == op_31_B;
wire op_31_ap_vld_A;
wire op_31_ap_vld_B;
wire clk_enable_A;
wire clk_enable_B;
assign clk_enable_A = _setup & (~op_31_ap_vld_A | op_31_ap_vld_B);
assign clk_enable_B = _setup;
wire divergent;
assign divergent = ~(ap_done_eq & ap_idle_eq & ap_ready_eq & op_31_eq);
assign unsafe_signal = op_31_ap_vld_A & op_31_ap_vld_B & divergent;
top_A instance_A (
    .ap_clk(ap_clk),
    .clk_enable(clk_enable_A),
    .ap_start(ap_start_internal),
    .op_0(op_0_internal),
    .op_10(op_10_internal),
    .op_12(op_12_internal),
    .op_13(op_13_internal),
    .op_14(op_14_internal),
    .op_15(op_15_internal),
    .op_19(op_19_internal),
    .op_2(op_2_internal),
    .op_3(op_3_internal),
    .op_4(op_4_internal),
    .op_5(op_5_internal),
    .op_6(op_6_internal),
    .op_7(op_7_internal),
    .op_8(op_8_internal),
    .ap_done(ap_done_A),
    .ap_idle(ap_idle_A),
    .ap_ready(ap_ready_A),
    .op_31(op_31_A),
    .op_31_ap_vld(op_31_ap_vld_A)
);
top_B instance_B (
    .ap_clk(ap_clk),
    .clk_enable(clk_enable_B),
    .ap_start(ap_start_internal),
    .op_0(op_0_internal),
    .op_10(op_10_internal),
    .op_12(op_12_internal),
    .op_13(op_13_internal),
    .op_14(op_14_internal),
    .op_15(op_15_internal),
    .op_19(op_19_internal),
    .op_2(op_2_internal),
    .op_3(op_3_internal),
    .op_4(op_4_internal),
    .op_5(op_5_internal),
    .op_6(op_6_internal),
    .op_7(op_7_internal),
    .op_8(op_8_internal),
    .ap_done(ap_done_B),
    .ap_idle(ap_idle_B),
    .ap_ready(ap_ready_B),
    .op_31(op_31_B),
    .op_31_ap_vld(op_31_ap_vld_B)
);
endmodule
