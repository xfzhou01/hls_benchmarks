// Processed by function `construct_kairos` in `verilog_tricks.py`.
// Machine A:
// Processed by function `add_clk_enable_signal` in `verilog_tricks.py`.
// Processed by function `remove_reset_signal` in `verilog_tricks.py`.
module top_A (
  ap_clk,
  ap_start,
  ap_done,
  ap_idle,
  ap_ready,
  op_0,
  op_6,
  op_7,
  op_8,
  op_11,
  op_16,
  op_17,
  op_18,
  op_29,
  op_29_ap_vld,
clk_enable
);
input clk_enable;


input ap_clk;
wire ap_rst;
assign ap_rst = op_29_ap_vld;
input ap_start;
input [3:0] op_0;
input [15:0] op_11;
input [15:0] op_16;
input [31:0] op_17;
input [3:0] op_18;
input [7:0] op_6;
input [15:0] op_7;
input [3:0] op_8;
output ap_done;
output ap_idle;
output ap_ready;
output [31:0] op_29;
output op_29_ap_vld;


reg Range1_all_ones_reg_2030;
reg Range1_all_zeros_reg_2037;
reg Range2_all_ones_reg_2025;
reg [4:0] \add_10ns_10ns_10_2_1_U13.top_add_10ns_10ns_10_2_1_Adder_9_U.ain_s1 ;
reg [4:0] \add_10ns_10ns_10_2_1_U13.top_add_10ns_10ns_10_2_1_Adder_9_U.bin_s1 ;
reg \add_10ns_10ns_10_2_1_U13.top_add_10ns_10ns_10_2_1_Adder_9_U.carry_s1 ;
reg [4:0] \add_10ns_10ns_10_2_1_U13.top_add_10ns_10ns_10_2_1_Adder_9_U.sum_s1 ;
reg [5:0] \add_12s_12ns_12_2_1_U17.top_add_12s_12ns_12_2_1_Adder_13_U.ain_s1 ;
reg [5:0] \add_12s_12ns_12_2_1_U17.top_add_12s_12ns_12_2_1_Adder_13_U.bin_s1 ;
reg \add_12s_12ns_12_2_1_U17.top_add_12s_12ns_12_2_1_Adder_13_U.carry_s1 ;
reg [5:0] \add_12s_12ns_12_2_1_U17.top_add_12s_12ns_12_2_1_Adder_13_U.sum_s1 ;
reg [6:0] \add_13ns_13s_13_2_1_U10.top_add_13ns_13s_13_2_1_Adder_7_U.ain_s1 ;
reg [6:0] \add_13ns_13s_13_2_1_U10.top_add_13ns_13s_13_2_1_Adder_7_U.bin_s1 ;
reg \add_13ns_13s_13_2_1_U10.top_add_13ns_13s_13_2_1_Adder_7_U.carry_s1 ;
reg [5:0] \add_13ns_13s_13_2_1_U10.top_add_13ns_13s_13_2_1_Adder_7_U.sum_s1 ;
reg [8:0] \add_17s_17s_17_2_1_U28.top_add_17s_17s_17_2_1_Adder_18_U.ain_s1 ;
reg [8:0] \add_17s_17s_17_2_1_U28.top_add_17s_17s_17_2_1_Adder_18_U.bin_s1 ;
reg \add_17s_17s_17_2_1_U28.top_add_17s_17s_17_2_1_Adder_18_U.carry_s1 ;
reg [7:0] \add_17s_17s_17_2_1_U28.top_add_17s_17s_17_2_1_Adder_18_U.sum_s1 ;
reg [11:0] \add_24s_24s_24_2_1_U16.top_add_24s_24s_24_2_1_Adder_12_U.ain_s1 ;
reg [11:0] \add_24s_24s_24_2_1_U16.top_add_24s_24s_24_2_1_Adder_12_U.bin_s1 ;
reg \add_24s_24s_24_2_1_U16.top_add_24s_24s_24_2_1_Adder_12_U.carry_s1 ;
reg [11:0] \add_24s_24s_24_2_1_U16.top_add_24s_24s_24_2_1_Adder_12_U.sum_s1 ;
reg \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.ain_s1 ;
reg \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.bin_s1 ;
reg \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.carry_s1 ;
reg \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.sum_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_15_U.ain_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_15_U.bin_s1 ;
reg \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_15_U.carry_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_15_U.sum_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_15_U.ain_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_15_U.bin_s1 ;
reg \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_15_U.carry_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_15_U.sum_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.ain_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.bin_s1 ;
reg \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.carry_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.sum_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.ain_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.bin_s1 ;
reg \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.carry_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.sum_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U27.top_add_32ns_32ns_32_2_1_Adder_15_U.ain_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U27.top_add_32ns_32ns_32_2_1_Adder_15_U.bin_s1 ;
reg \add_32ns_32ns_32_2_1_U27.top_add_32ns_32ns_32_2_1_Adder_15_U.carry_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U27.top_add_32ns_32ns_32_2_1_Adder_15_U.sum_s1 ;
reg [15:0] \add_32s_32ns_32_2_1_U29.top_add_32s_32ns_32_2_1_Adder_19_U.ain_s1 ;
reg [15:0] \add_32s_32ns_32_2_1_U29.top_add_32s_32ns_32_2_1_Adder_19_U.bin_s1 ;
reg \add_32s_32ns_32_2_1_U29.top_add_32s_32ns_32_2_1_Adder_19_U.carry_s1 ;
reg [15:0] \add_32s_32ns_32_2_1_U29.top_add_32s_32ns_32_2_1_Adder_19_U.sum_s1 ;
reg [16:0] \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_16_U.ain_s1 ;
reg [16:0] \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_16_U.bin_s1 ;
reg \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_16_U.carry_s1 ;
reg [16:0] \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_16_U.sum_s1 ;
reg [17:0] \add_35s_35s_35_2_1_U19.top_add_35s_35s_35_2_1_Adder_14_U.ain_s1 ;
reg [17:0] \add_35s_35s_35_2_1_U19.top_add_35s_35s_35_2_1_Adder_14_U.bin_s1 ;
reg \add_35s_35s_35_2_1_U19.top_add_35s_35s_35_2_1_Adder_14_U.carry_s1 ;
reg [16:0] \add_35s_35s_35_2_1_U19.top_add_35s_35s_35_2_1_Adder_14_U.sum_s1 ;
reg [17:0] \add_35s_35s_35_2_1_U21.top_add_35s_35s_35_2_1_Adder_14_U.ain_s1 ;
reg [17:0] \add_35s_35s_35_2_1_U21.top_add_35s_35s_35_2_1_Adder_14_U.bin_s1 ;
reg \add_35s_35s_35_2_1_U21.top_add_35s_35s_35_2_1_Adder_14_U.carry_s1 ;
reg [16:0] \add_35s_35s_35_2_1_U21.top_add_35s_35s_35_2_1_Adder_14_U.sum_s1 ;
reg [1:0] \add_3ns_3ns_3_2_1_U1.top_add_3ns_3ns_3_2_1_Adder_0_U.ain_s1 ;
reg [1:0] \add_3ns_3ns_3_2_1_U1.top_add_3ns_3ns_3_2_1_Adder_0_U.bin_s1 ;
reg \add_3ns_3ns_3_2_1_U1.top_add_3ns_3ns_3_2_1_Adder_0_U.carry_s1 ;
reg \add_3ns_3ns_3_2_1_U1.top_add_3ns_3ns_3_2_1_Adder_0_U.sum_s1 ;
reg [1:0] \add_4ns_4ns_4_2_1_U18.top_add_4ns_4ns_4_2_1_Adder_5_U.ain_s1 ;
reg [1:0] \add_4ns_4ns_4_2_1_U18.top_add_4ns_4ns_4_2_1_Adder_5_U.bin_s1 ;
reg \add_4ns_4ns_4_2_1_U18.top_add_4ns_4ns_4_2_1_Adder_5_U.carry_s1 ;
reg [1:0] \add_4ns_4ns_4_2_1_U18.top_add_4ns_4ns_4_2_1_Adder_5_U.sum_s1 ;
reg [1:0] \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_5_U.ain_s1 ;
reg [1:0] \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_5_U.bin_s1 ;
reg \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_5_U.carry_s1 ;
reg [1:0] \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_5_U.sum_s1 ;
reg [1:0] \add_4s_4ns_4_2_1_U4.top_add_4s_4ns_4_2_1_Adder_3_U.ain_s1 ;
reg [1:0] \add_4s_4ns_4_2_1_U4.top_add_4s_4ns_4_2_1_Adder_3_U.bin_s1 ;
reg \add_4s_4ns_4_2_1_U4.top_add_4s_4ns_4_2_1_Adder_3_U.carry_s1 ;
reg [1:0] \add_4s_4ns_4_2_1_U4.top_add_4s_4ns_4_2_1_Adder_3_U.sum_s1 ;
reg [2:0] \add_5ns_5s_5_2_1_U3.top_add_5ns_5s_5_2_1_Adder_2_U.ain_s1 ;
reg [2:0] \add_5ns_5s_5_2_1_U3.top_add_5ns_5s_5_2_1_Adder_2_U.bin_s1 ;
reg \add_5ns_5s_5_2_1_U3.top_add_5ns_5s_5_2_1_Adder_2_U.carry_s1 ;
reg [1:0] \add_5ns_5s_5_2_1_U3.top_add_5ns_5s_5_2_1_Adder_2_U.sum_s1 ;
reg [3:0] \add_7s_7s_7_2_1_U2.top_add_7s_7s_7_2_1_Adder_1_U.ain_s1 ;
reg [3:0] \add_7s_7s_7_2_1_U2.top_add_7s_7s_7_2_1_Adder_1_U.bin_s1 ;
reg \add_7s_7s_7_2_1_U2.top_add_7s_7s_7_2_1_Adder_1_U.carry_s1 ;
reg [2:0] \add_7s_7s_7_2_1_U2.top_add_7s_7s_7_2_1_Adder_1_U.sum_s1 ;
reg [4:0] \add_9s_9ns_9_2_1_U26.top_add_9s_9ns_9_2_1_Adder_17_U.ain_s1 ;
reg [4:0] \add_9s_9ns_9_2_1_U26.top_add_9s_9ns_9_2_1_Adder_17_U.bin_s1 ;
reg \add_9s_9ns_9_2_1_U26.top_add_9s_9ns_9_2_1_Adder_17_U.carry_s1 ;
reg [3:0] \add_9s_9ns_9_2_1_U26.top_add_9s_9ns_9_2_1_Adder_17_U.sum_s1 ;
reg [4:0] add_ln1192_1_reg_1826;
reg [11:0] add_ln691_3_reg_2407;
reg [31:0] add_ln691_4_reg_2469;
reg [31:0] add_ln691_5_reg_2501;
reg [31:0] add_ln691_6_reg_2543;
reg [3:0] add_ln691_reg_2057;
reg [8:0] add_ln69_1_reg_2563;
reg [16:0] add_ln69_2_reg_2588;
reg [31:0] add_ln69_reg_2583;
reg and_ln412_reg_2020;
reg and_ln786_1_reg_1896;
reg and_ln786_2_reg_2355;
reg and_ln786_reg_2194;
reg [51:0] ap_CS_fsm = 52'h0000000000001;
reg carry_1_reg_2141;
reg deleted_zeros_reg_2188;
reg icmp_ln768_1_reg_1861;
reg icmp_ln768_3_reg_2205;
reg icmp_ln768_4_reg_2269;
reg icmp_ln768_reg_1751;
reg icmp_ln786_1_reg_1866;
reg icmp_ln786_2_reg_2210;
reg icmp_ln786_3_reg_2274;
reg icmp_ln786_reg_1767;
reg icmp_ln851_1_reg_2092;
reg icmp_ln851_2_reg_2305;
reg icmp_ln851_3_reg_2452;
reg icmp_ln851_4_reg_2402;
reg icmp_ln851_reg_2042;
reg [31:0] \mul_32ns_4s_36_7_1_U5.top_mul_32ns_4s_36_7_1_Mul_DSP_0_U.a_reg0 ;
reg [3:0] \mul_32ns_4s_36_7_1_U5.top_mul_32ns_4s_36_7_1_Mul_DSP_0_U.b_reg0 ;
reg [35:0] \mul_32ns_4s_36_7_1_U5.top_mul_32ns_4s_36_7_1_Mul_DSP_0_U.buff0 ;
reg [35:0] \mul_32ns_4s_36_7_1_U5.top_mul_32ns_4s_36_7_1_Mul_DSP_0_U.buff1 ;
reg [35:0] \mul_32ns_4s_36_7_1_U5.top_mul_32ns_4s_36_7_1_Mul_DSP_0_U.buff2 ;
reg [35:0] \mul_32ns_4s_36_7_1_U5.top_mul_32ns_4s_36_7_1_Mul_DSP_0_U.buff3 ;
reg [35:0] \mul_32ns_4s_36_7_1_U5.top_mul_32ns_4s_36_7_1_Mul_DSP_0_U.buff4 ;
reg [31:0] \mul_32ns_4s_36_7_1_U6.top_mul_32ns_4s_36_7_1_Mul_DSP_0_U.a_reg0 ;
reg [3:0] \mul_32ns_4s_36_7_1_U6.top_mul_32ns_4s_36_7_1_Mul_DSP_0_U.b_reg0 ;
reg [35:0] \mul_32ns_4s_36_7_1_U6.top_mul_32ns_4s_36_7_1_Mul_DSP_0_U.buff0 ;
reg [35:0] \mul_32ns_4s_36_7_1_U6.top_mul_32ns_4s_36_7_1_Mul_DSP_0_U.buff1 ;
reg [35:0] \mul_32ns_4s_36_7_1_U6.top_mul_32ns_4s_36_7_1_Mul_DSP_0_U.buff2 ;
reg [35:0] \mul_32ns_4s_36_7_1_U6.top_mul_32ns_4s_36_7_1_Mul_DSP_0_U.buff3 ;
reg [35:0] \mul_32ns_4s_36_7_1_U6.top_mul_32ns_4s_36_7_1_Mul_DSP_0_U.buff4 ;
reg [3:0] \mul_4ns_3s_7_7_1_U12.top_mul_4ns_3s_7_7_1_Mul_DSP_1_U.a_reg0 ;
reg [2:0] \mul_4ns_3s_7_7_1_U12.top_mul_4ns_3s_7_7_1_Mul_DSP_1_U.b_reg0 ;
reg [6:0] \mul_4ns_3s_7_7_1_U12.top_mul_4ns_3s_7_7_1_Mul_DSP_1_U.buff0 ;
reg [6:0] \mul_4ns_3s_7_7_1_U12.top_mul_4ns_3s_7_7_1_Mul_DSP_1_U.buff1 ;
reg [6:0] \mul_4ns_3s_7_7_1_U12.top_mul_4ns_3s_7_7_1_Mul_DSP_1_U.buff2 ;
reg [6:0] \mul_4ns_3s_7_7_1_U12.top_mul_4ns_3s_7_7_1_Mul_DSP_1_U.buff3 ;
reg [6:0] \mul_4ns_3s_7_7_1_U12.top_mul_4ns_3s_7_7_1_Mul_DSP_1_U.buff4 ;
reg [7:0] op_10_V_reg_2047;
reg [7:0] op_12_V_reg_2422;
reg [15:0] op_13_V_reg_2328;
reg [1:0] op_15_V_reg_2322;
reg [7:0] op_19_V_reg_2248;
reg [3:0] op_1_V_reg_1789;
reg [31:0] op_24_V_reg_2516;
reg [3:0] op_3_V_reg_1917;
reg or_ln340_1_reg_1890;
reg or_ln340_2_reg_2253;
reg or_ln340_4_reg_2349;
reg or_ln785_1_reg_1872;
reg or_ln785_3_reg_2258;
reg or_ln785_4_reg_2310;
reg or_ln785_reg_1761;
reg or_ln786_1_reg_1884;
reg or_ln786_3_reg_2343;
reg p_Result_11_reg_1966;
reg [31:0] p_Result_1_reg_1976;
reg p_Result_26_reg_1736;
reg p_Result_27_reg_1832;
reg p_Result_28_reg_1848;
reg p_Result_30_reg_1954;
reg p_Result_31_reg_1949;
reg p_Result_32_reg_1971;
reg p_Result_33_reg_2068;
reg p_Result_34_reg_2148;
reg p_Result_35_reg_2160;
reg p_Result_36_reg_2223;
reg p_Result_37_reg_2235;
reg [32:0] p_Result_3_reg_1981;
reg [2:0] p_Result_4_reg_2167;
reg [2:0] p_Result_s_22_reg_1855;
reg p_Result_s_reg_1722;
reg [15:0] p_Val2_10_reg_2285;
reg [7:0] p_Val2_14_reg_2386;
reg [3:0] p_Val2_2_reg_1839;
reg [1:0] p_Val2_5_reg_1961;
reg [1:0] p_Val2_6_reg_2062;
reg [3:0] p_Val2_s_reg_1730;
reg [35:0] r_V_5_reg_1944;
reg [35:0] r_V_6_reg_1987;
reg [6:0] r_V_7_reg_2366;
reg [2:0] r_V_reg_1796;
reg [32:0] ret_1_reg_2216;
reg [3:0] ret_V_10_cast_reg_2372;
reg [2:0] ret_V_16_reg_1783;
reg [31:0] ret_V_17_cast_reg_2462;
reg [3:0] ret_V_18_reg_2075;
reg [12:0] ret_V_19_reg_2103;
reg [2:0] ret_V_1_reg_1773;
reg [31:0] ret_V_20_cast_reg_2494;
reg [3:0] ret_V_20_reg_2437;
reg [23:0] ret_V_21_reg_2333;
reg [34:0] ret_V_22_reg_2457;
reg [31:0] ret_V_23_cast_reg_2536;
reg [34:0] ret_V_23_reg_2489;
reg [31:0] ret_V_24_reg_2506;
reg [33:0] ret_V_25_reg_2531;
reg [31:0] ret_V_26_reg_2558;
reg [3:0] ret_V_4_cast_reg_1992;
reg [9:0] ret_V_6_reg_2108;
reg [9:0] ret_V_7_reg_2200;
reg [3:0] ret_V_8_reg_2417;
reg [2:0] ret_V_reg_1743;
reg rhs_4_reg_2120;
reg sel_tmp19_reg_1907;
reg sel_tmp51_reg_2397;
reg [3:0] select_ln340_1_reg_1902;
reg [1:0] select_ln340_2_reg_2280;
reg [15:0] select_ln340_3_reg_2290;
reg [7:0] select_ln340_4_reg_2392;
reg [3:0] select_ln340_reg_1778;
reg [31:0] select_ln353_1_reg_2474;
reg [11:0] select_ln353_reg_2427;
reg [7:0] select_ln785_3_reg_2412;
reg [3:0] select_ln785_reg_1912;
reg [9:0] select_ln850_4_reg_2264;
reg [31:0] sext_ln1116_reg_1923;
reg [11:0] sext_ln850_reg_2379;
reg [8:0] \sub_17ns_17ns_17_2_1_U11.top_sub_17ns_17ns_17_2_1_Adder_8_U.ain_s1 ;
reg [8:0] \sub_17ns_17ns_17_2_1_U11.top_sub_17ns_17ns_17_2_1_Adder_8_U.bin_s1 ;
reg \sub_17ns_17ns_17_2_1_U11.top_sub_17ns_17ns_17_2_1_Adder_8_U.carry_s1 ;
reg [7:0] \sub_17ns_17ns_17_2_1_U11.top_sub_17ns_17ns_17_2_1_Adder_8_U.sum_s1 ;
reg [16:0] \sub_33ns_33ns_33_2_1_U14.top_sub_33ns_33ns_33_2_1_Adder_10_U.ain_s1 ;
reg [16:0] \sub_33ns_33ns_33_2_1_U14.top_sub_33ns_33ns_33_2_1_Adder_10_U.bin_s1 ;
reg \sub_33ns_33ns_33_2_1_U14.top_sub_33ns_33ns_33_2_1_Adder_10_U.carry_s1 ;
reg [15:0] \sub_33ns_33ns_33_2_1_U14.top_sub_33ns_33ns_33_2_1_Adder_10_U.sum_s1 ;
reg [3:0] \sub_8ns_8ns_8_2_1_U15.top_sub_8ns_8ns_8_2_1_Adder_11_U.ain_s1 ;
reg [3:0] \sub_8ns_8ns_8_2_1_U15.top_sub_8ns_8ns_8_2_1_Adder_11_U.bin_s1 ;
reg \sub_8ns_8ns_8_2_1_U15.top_sub_8ns_8ns_8_2_1_Adder_11_U.carry_s1 ;
reg [3:0] \sub_8ns_8ns_8_2_1_U15.top_sub_8ns_8ns_8_2_1_Adder_11_U.sum_s1 ;
reg [3:0] \sub_8s_8ns_8_2_1_U7.top_sub_8s_8ns_8_2_1_Adder_4_U.ain_s1 ;
reg [3:0] \sub_8s_8ns_8_2_1_U7.top_sub_8s_8ns_8_2_1_Adder_4_U.bin_s1 ;
reg \sub_8s_8ns_8_2_1_U7.top_sub_8s_8ns_8_2_1_Adder_4_U.carry_s1 ;
reg [3:0] \sub_8s_8ns_8_2_1_U7.top_sub_8s_8ns_8_2_1_Adder_4_U.sum_s1 ;
reg [26:0] tmp_1_reg_2242;
reg [10:0] tmp_reg_2338;
reg [2:0] trunc_ln1192_reg_1756;
reg [7:0] trunc_ln213_reg_2014;
reg [13:0] trunc_ln731_1_reg_2155;
reg [5:0] trunc_ln731_2_reg_2230;
reg [1:0] trunc_ln851_4_reg_2432;
reg [1:0] trunc_ln851_5_reg_2361;
reg [2:0] trunc_ln851_reg_1999;
reg xor_ln416_reg_2097;
reg xor_ln785_1_reg_1878;
reg xor_ln785_5_reg_2316;
wire _0000_;
wire _0001_;
wire _0002_;
wire [4:0] _0003_;
wire [11:0] _0004_;
wire [31:0] _0005_;
wire [31:0] _0006_;
wire [31:0] _0007_;
wire [3:0] _0008_;
wire [8:0] _0009_;
wire [16:0] _0010_;
wire [31:0] _0011_;
wire _0012_;
wire _0013_;
wire _0014_;
wire _0015_;
wire [51:0] _0016_;
wire _0017_;
wire _0018_;
wire _0019_;
wire _0020_;
wire _0021_;
wire _0022_;
wire _0023_;
wire _0024_;
wire _0025_;
wire _0026_;
wire _0027_;
wire _0028_;
wire _0029_;
wire _0030_;
wire _0031_;
wire [7:0] _0032_;
wire [7:0] _0033_;
wire [13:0] _0034_;
wire [1:0] _0035_;
wire [7:0] _0036_;
wire _0037_;
wire [31:0] _0038_;
wire [3:0] _0039_;
wire _0040_;
wire _0041_;
wire _0042_;
wire _0043_;
wire _0044_;
wire _0045_;
wire _0046_;
wire _0047_;
wire _0048_;
wire _0049_;
wire [31:0] _0050_;
wire _0051_;
wire _0052_;
wire _0053_;
wire _0054_;
wire _0055_;
wire _0056_;
wire _0057_;
wire _0058_;
wire _0059_;
wire _0060_;
wire _0061_;
wire [32:0] _0062_;
wire [2:0] _0063_;
wire [2:0] _0064_;
wire _0065_;
wire [13:0] _0066_;
wire [5:0] _0067_;
wire [3:0] _0068_;
wire [1:0] _0069_;
wire [1:0] _0070_;
wire _0071_;
wire [35:0] _0072_;
wire [35:0] _0073_;
wire [6:0] _0074_;
wire [2:0] _0075_;
wire [32:0] _0076_;
wire [3:0] _0077_;
wire [2:0] _0078_;
wire [31:0] _0079_;
wire [3:0] _0080_;
wire [12:0] _0081_;
wire [2:0] _0082_;
wire [31:0] _0083_;
wire [3:0] _0084_;
wire [23:0] _0085_;
wire [34:0] _0086_;
wire [31:0] _0087_;
wire [34:0] _0088_;
wire [31:0] _0089_;
wire [33:0] _0090_;
wire [31:0] _0091_;
wire [3:0] _0092_;
wire [9:0] _0093_;
wire [9:0] _0094_;
wire [3:0] _0095_;
wire [2:0] _0096_;
wire _0097_;
wire _0098_;
wire _0099_;
wire [3:0] _0100_;
wire [1:0] _0101_;
wire [13:0] _0102_;
wire [7:0] _0103_;
wire _0104_;
wire [31:0] _0105_;
wire [11:0] _0106_;
wire [7:0] _0107_;
wire [3:0] _0108_;
wire [9:0] _0109_;
wire [31:0] _0110_;
wire [11:0] _0111_;
wire [26:0] _0112_;
wire [10:0] _0113_;
wire [2:0] _0114_;
wire [7:0] _0115_;
wire [13:0] _0116_;
wire [5:0] _0117_;
wire [1:0] _0118_;
wire [2:0] _0119_;
wire _0120_;
wire _0121_;
wire _0122_;
wire [1:0] _0123_;
wire _0124_;
wire _0125_;
wire _0126_;
wire _0127_;
wire _0128_;
wire _0129_;
wire _0130_;
wire _0131_;
wire _0132_;
wire _0133_;
wire _0134_;
wire _0135_;
wire _0136_;
wire _0137_;
wire _0138_;
wire _0139_;
wire [4:0] _0140_;
wire [4:0] _0141_;
wire _0142_;
wire [4:0] _0143_;
wire [5:0] _0144_;
wire [5:0] _0145_;
wire [5:0] _0146_;
wire [5:0] _0147_;
wire _0148_;
wire [5:0] _0149_;
wire [6:0] _0150_;
wire [6:0] _0151_;
wire [6:0] _0152_;
wire [6:0] _0153_;
wire _0154_;
wire [5:0] _0155_;
wire [6:0] _0156_;
wire [7:0] _0157_;
wire [8:0] _0158_;
wire [8:0] _0159_;
wire _0160_;
wire [7:0] _0161_;
wire [8:0] _0162_;
wire [9:0] _0163_;
wire [11:0] _0164_;
wire [11:0] _0165_;
wire _0166_;
wire [11:0] _0167_;
wire [12:0] _0168_;
wire [12:0] _0169_;
wire _0170_;
wire _0171_;
wire _0172_;
wire _0173_;
wire [1:0] _0174_;
wire [1:0] _0175_;
wire [15:0] _0176_;
wire [15:0] _0177_;
wire _0178_;
wire [15:0] _0179_;
wire [16:0] _0180_;
wire [16:0] _0181_;
wire [15:0] _0182_;
wire [15:0] _0183_;
wire _0184_;
wire [15:0] _0185_;
wire [16:0] _0186_;
wire [16:0] _0187_;
wire [15:0] _0188_;
wire [15:0] _0189_;
wire _0190_;
wire [15:0] _0191_;
wire [16:0] _0192_;
wire [16:0] _0193_;
wire [15:0] _0194_;
wire [15:0] _0195_;
wire _0196_;
wire [15:0] _0197_;
wire [16:0] _0198_;
wire [16:0] _0199_;
wire [15:0] _0200_;
wire [15:0] _0201_;
wire _0202_;
wire [15:0] _0203_;
wire [16:0] _0204_;
wire [16:0] _0205_;
wire [15:0] _0206_;
wire [15:0] _0207_;
wire _0208_;
wire [15:0] _0209_;
wire [16:0] _0210_;
wire [16:0] _0211_;
wire [16:0] _0212_;
wire [16:0] _0213_;
wire _0214_;
wire [16:0] _0215_;
wire [17:0] _0216_;
wire [17:0] _0217_;
wire [17:0] _0218_;
wire [17:0] _0219_;
wire _0220_;
wire [16:0] _0221_;
wire [17:0] _0222_;
wire [18:0] _0223_;
wire [17:0] _0224_;
wire [17:0] _0225_;
wire _0226_;
wire [16:0] _0227_;
wire [17:0] _0228_;
wire [18:0] _0229_;
wire [1:0] _0230_;
wire [1:0] _0231_;
wire _0232_;
wire _0233_;
wire [1:0] _0234_;
wire [2:0] _0235_;
wire [1:0] _0236_;
wire [1:0] _0237_;
wire _0238_;
wire [1:0] _0239_;
wire [2:0] _0240_;
wire [2:0] _0241_;
wire [1:0] _0242_;
wire [1:0] _0243_;
wire _0244_;
wire [1:0] _0245_;
wire [2:0] _0246_;
wire [2:0] _0247_;
wire [1:0] _0248_;
wire [1:0] _0249_;
wire _0250_;
wire [1:0] _0251_;
wire [2:0] _0252_;
wire [2:0] _0253_;
wire [2:0] _0254_;
wire [2:0] _0255_;
wire _0256_;
wire [1:0] _0257_;
wire [2:0] _0258_;
wire [3:0] _0259_;
wire [3:0] _0260_;
wire [3:0] _0261_;
wire _0262_;
wire [2:0] _0263_;
wire [3:0] _0264_;
wire [4:0] _0265_;
wire [4:0] _0266_;
wire [4:0] _0267_;
wire _0268_;
wire [3:0] _0269_;
wire [4:0] _0270_;
wire [5:0] _0271_;
wire [31:0] _0272_;
wire [3:0] _0273_;
wire [35:0] _0274_;
wire [35:0] _0275_;
wire [35:0] _0276_;
wire [35:0] _0277_;
wire [35:0] _0278_;
wire [31:0] _0279_;
wire [3:0] _0280_;
wire [35:0] _0281_;
wire [35:0] _0282_;
wire [35:0] _0283_;
wire [35:0] _0284_;
wire [35:0] _0285_;
wire [3:0] _0286_;
wire [2:0] _0287_;
wire [6:0] _0288_;
wire [6:0] _0289_;
wire [6:0] _0290_;
wire [6:0] _0291_;
wire [6:0] _0292_;
wire [8:0] _0293_;
wire [8:0] _0294_;
wire _0295_;
wire [7:0] _0296_;
wire [8:0] _0297_;
wire [9:0] _0298_;
wire [16:0] _0299_;
wire [16:0] _0300_;
wire _0301_;
wire [15:0] _0302_;
wire [16:0] _0303_;
wire [17:0] _0304_;
wire [3:0] _0305_;
wire [3:0] _0306_;
wire _0307_;
wire [3:0] _0308_;
wire [4:0] _0309_;
wire [4:0] _0310_;
wire [3:0] _0311_;
wire [3:0] _0312_;
wire _0313_;
wire [3:0] _0314_;
wire [4:0] _0315_;
wire [4:0] _0316_;
wire _0317_;
wire _0318_;
wire _0319_;
wire _0320_;
wire _0321_;
wire _0322_;
wire _0323_;
wire _0324_;
wire _0325_;
wire _0326_;
wire _0327_;
wire _0328_;
wire _0329_;
wire _0330_;
wire _0331_;
wire _0332_;
wire _0333_;
wire _0334_;
wire _0335_;
wire _0336_;
wire _0337_;
wire _0338_;
wire _0339_;
wire _0340_;
wire _0341_;
wire _0342_;
wire _0343_;
wire _0344_;
wire _0345_;
wire _0346_;
wire _0347_;
wire _0348_;
wire _0349_;
wire _0350_;
wire _0351_;
wire _0352_;
wire _0353_;
wire _0354_;
wire _0355_;
wire _0356_;
wire _0357_;
wire _0358_;
wire _0359_;
wire _0360_;
wire _0361_;
wire _0362_;
wire _0363_;
wire _0364_;
wire _0365_;
wire _0366_;
wire _0367_;
wire _0368_;
wire _0369_;
wire _0370_;
wire _0371_;
wire _0372_;
wire _0373_;
wire _0374_;
wire _0375_;
wire _0376_;
wire _0377_;
wire _0378_;
wire _0379_;
wire _0380_;
wire _0381_;
wire Range1_all_ones_fu_750_p2;
wire Range1_all_zeros_fu_755_p2;
wire Range2_all_ones_fu_745_p2;
wire \add_10ns_10ns_10_2_1_U13.ce ;
wire \add_10ns_10ns_10_2_1_U13.clk ;
wire [9:0] \add_10ns_10ns_10_2_1_U13.din0 ;
wire [9:0] \add_10ns_10ns_10_2_1_U13.din1 ;
wire [9:0] \add_10ns_10ns_10_2_1_U13.dout ;
wire \add_10ns_10ns_10_2_1_U13.reset ;
wire [9:0] \add_10ns_10ns_10_2_1_U13.top_add_10ns_10ns_10_2_1_Adder_9_U.a ;
wire [9:0] \add_10ns_10ns_10_2_1_U13.top_add_10ns_10ns_10_2_1_Adder_9_U.ain_s0 ;
wire [9:0] \add_10ns_10ns_10_2_1_U13.top_add_10ns_10ns_10_2_1_Adder_9_U.b ;
wire [9:0] \add_10ns_10ns_10_2_1_U13.top_add_10ns_10ns_10_2_1_Adder_9_U.bin_s0 ;
wire \add_10ns_10ns_10_2_1_U13.top_add_10ns_10ns_10_2_1_Adder_9_U.ce ;
wire \add_10ns_10ns_10_2_1_U13.top_add_10ns_10ns_10_2_1_Adder_9_U.clk ;
wire \add_10ns_10ns_10_2_1_U13.top_add_10ns_10ns_10_2_1_Adder_9_U.facout_s1 ;
wire \add_10ns_10ns_10_2_1_U13.top_add_10ns_10ns_10_2_1_Adder_9_U.facout_s2 ;
wire [4:0] \add_10ns_10ns_10_2_1_U13.top_add_10ns_10ns_10_2_1_Adder_9_U.fas_s1 ;
wire [4:0] \add_10ns_10ns_10_2_1_U13.top_add_10ns_10ns_10_2_1_Adder_9_U.fas_s2 ;
wire \add_10ns_10ns_10_2_1_U13.top_add_10ns_10ns_10_2_1_Adder_9_U.reset ;
wire [9:0] \add_10ns_10ns_10_2_1_U13.top_add_10ns_10ns_10_2_1_Adder_9_U.s ;
wire [4:0] \add_10ns_10ns_10_2_1_U13.top_add_10ns_10ns_10_2_1_Adder_9_U.u1.a ;
wire [4:0] \add_10ns_10ns_10_2_1_U13.top_add_10ns_10ns_10_2_1_Adder_9_U.u1.b ;
wire \add_10ns_10ns_10_2_1_U13.top_add_10ns_10ns_10_2_1_Adder_9_U.u1.cin ;
wire \add_10ns_10ns_10_2_1_U13.top_add_10ns_10ns_10_2_1_Adder_9_U.u1.cout ;
wire [4:0] \add_10ns_10ns_10_2_1_U13.top_add_10ns_10ns_10_2_1_Adder_9_U.u1.s ;
wire [4:0] \add_10ns_10ns_10_2_1_U13.top_add_10ns_10ns_10_2_1_Adder_9_U.u2.a ;
wire [4:0] \add_10ns_10ns_10_2_1_U13.top_add_10ns_10ns_10_2_1_Adder_9_U.u2.b ;
wire \add_10ns_10ns_10_2_1_U13.top_add_10ns_10ns_10_2_1_Adder_9_U.u2.cin ;
wire \add_10ns_10ns_10_2_1_U13.top_add_10ns_10ns_10_2_1_Adder_9_U.u2.cout ;
wire [4:0] \add_10ns_10ns_10_2_1_U13.top_add_10ns_10ns_10_2_1_Adder_9_U.u2.s ;
wire \add_12s_12ns_12_2_1_U17.ce ;
wire \add_12s_12ns_12_2_1_U17.clk ;
wire [11:0] \add_12s_12ns_12_2_1_U17.din0 ;
wire [11:0] \add_12s_12ns_12_2_1_U17.din1 ;
wire [11:0] \add_12s_12ns_12_2_1_U17.dout ;
wire \add_12s_12ns_12_2_1_U17.reset ;
wire [11:0] \add_12s_12ns_12_2_1_U17.top_add_12s_12ns_12_2_1_Adder_13_U.a ;
wire [11:0] \add_12s_12ns_12_2_1_U17.top_add_12s_12ns_12_2_1_Adder_13_U.ain_s0 ;
wire [11:0] \add_12s_12ns_12_2_1_U17.top_add_12s_12ns_12_2_1_Adder_13_U.b ;
wire [11:0] \add_12s_12ns_12_2_1_U17.top_add_12s_12ns_12_2_1_Adder_13_U.bin_s0 ;
wire \add_12s_12ns_12_2_1_U17.top_add_12s_12ns_12_2_1_Adder_13_U.ce ;
wire \add_12s_12ns_12_2_1_U17.top_add_12s_12ns_12_2_1_Adder_13_U.clk ;
wire \add_12s_12ns_12_2_1_U17.top_add_12s_12ns_12_2_1_Adder_13_U.facout_s1 ;
wire \add_12s_12ns_12_2_1_U17.top_add_12s_12ns_12_2_1_Adder_13_U.facout_s2 ;
wire [5:0] \add_12s_12ns_12_2_1_U17.top_add_12s_12ns_12_2_1_Adder_13_U.fas_s1 ;
wire [5:0] \add_12s_12ns_12_2_1_U17.top_add_12s_12ns_12_2_1_Adder_13_U.fas_s2 ;
wire \add_12s_12ns_12_2_1_U17.top_add_12s_12ns_12_2_1_Adder_13_U.reset ;
wire [11:0] \add_12s_12ns_12_2_1_U17.top_add_12s_12ns_12_2_1_Adder_13_U.s ;
wire [5:0] \add_12s_12ns_12_2_1_U17.top_add_12s_12ns_12_2_1_Adder_13_U.u1.a ;
wire [5:0] \add_12s_12ns_12_2_1_U17.top_add_12s_12ns_12_2_1_Adder_13_U.u1.b ;
wire \add_12s_12ns_12_2_1_U17.top_add_12s_12ns_12_2_1_Adder_13_U.u1.cin ;
wire \add_12s_12ns_12_2_1_U17.top_add_12s_12ns_12_2_1_Adder_13_U.u1.cout ;
wire [5:0] \add_12s_12ns_12_2_1_U17.top_add_12s_12ns_12_2_1_Adder_13_U.u1.s ;
wire [5:0] \add_12s_12ns_12_2_1_U17.top_add_12s_12ns_12_2_1_Adder_13_U.u2.a ;
wire [5:0] \add_12s_12ns_12_2_1_U17.top_add_12s_12ns_12_2_1_Adder_13_U.u2.b ;
wire \add_12s_12ns_12_2_1_U17.top_add_12s_12ns_12_2_1_Adder_13_U.u2.cin ;
wire \add_12s_12ns_12_2_1_U17.top_add_12s_12ns_12_2_1_Adder_13_U.u2.cout ;
wire [5:0] \add_12s_12ns_12_2_1_U17.top_add_12s_12ns_12_2_1_Adder_13_U.u2.s ;
wire \add_13ns_13s_13_2_1_U10.ce ;
wire \add_13ns_13s_13_2_1_U10.clk ;
wire [12:0] \add_13ns_13s_13_2_1_U10.din0 ;
wire [12:0] \add_13ns_13s_13_2_1_U10.din1 ;
wire [12:0] \add_13ns_13s_13_2_1_U10.dout ;
wire \add_13ns_13s_13_2_1_U10.reset ;
wire [12:0] \add_13ns_13s_13_2_1_U10.top_add_13ns_13s_13_2_1_Adder_7_U.a ;
wire [12:0] \add_13ns_13s_13_2_1_U10.top_add_13ns_13s_13_2_1_Adder_7_U.ain_s0 ;
wire [12:0] \add_13ns_13s_13_2_1_U10.top_add_13ns_13s_13_2_1_Adder_7_U.b ;
wire [12:0] \add_13ns_13s_13_2_1_U10.top_add_13ns_13s_13_2_1_Adder_7_U.bin_s0 ;
wire \add_13ns_13s_13_2_1_U10.top_add_13ns_13s_13_2_1_Adder_7_U.ce ;
wire \add_13ns_13s_13_2_1_U10.top_add_13ns_13s_13_2_1_Adder_7_U.clk ;
wire \add_13ns_13s_13_2_1_U10.top_add_13ns_13s_13_2_1_Adder_7_U.facout_s1 ;
wire \add_13ns_13s_13_2_1_U10.top_add_13ns_13s_13_2_1_Adder_7_U.facout_s2 ;
wire [5:0] \add_13ns_13s_13_2_1_U10.top_add_13ns_13s_13_2_1_Adder_7_U.fas_s1 ;
wire [6:0] \add_13ns_13s_13_2_1_U10.top_add_13ns_13s_13_2_1_Adder_7_U.fas_s2 ;
wire \add_13ns_13s_13_2_1_U10.top_add_13ns_13s_13_2_1_Adder_7_U.reset ;
wire [12:0] \add_13ns_13s_13_2_1_U10.top_add_13ns_13s_13_2_1_Adder_7_U.s ;
wire [5:0] \add_13ns_13s_13_2_1_U10.top_add_13ns_13s_13_2_1_Adder_7_U.u1.a ;
wire [5:0] \add_13ns_13s_13_2_1_U10.top_add_13ns_13s_13_2_1_Adder_7_U.u1.b ;
wire \add_13ns_13s_13_2_1_U10.top_add_13ns_13s_13_2_1_Adder_7_U.u1.cin ;
wire \add_13ns_13s_13_2_1_U10.top_add_13ns_13s_13_2_1_Adder_7_U.u1.cout ;
wire [5:0] \add_13ns_13s_13_2_1_U10.top_add_13ns_13s_13_2_1_Adder_7_U.u1.s ;
wire [6:0] \add_13ns_13s_13_2_1_U10.top_add_13ns_13s_13_2_1_Adder_7_U.u2.a ;
wire [6:0] \add_13ns_13s_13_2_1_U10.top_add_13ns_13s_13_2_1_Adder_7_U.u2.b ;
wire \add_13ns_13s_13_2_1_U10.top_add_13ns_13s_13_2_1_Adder_7_U.u2.cin ;
wire \add_13ns_13s_13_2_1_U10.top_add_13ns_13s_13_2_1_Adder_7_U.u2.cout ;
wire [6:0] \add_13ns_13s_13_2_1_U10.top_add_13ns_13s_13_2_1_Adder_7_U.u2.s ;
wire \add_17s_17s_17_2_1_U28.ce ;
wire \add_17s_17s_17_2_1_U28.clk ;
wire [16:0] \add_17s_17s_17_2_1_U28.din0 ;
wire [16:0] \add_17s_17s_17_2_1_U28.din1 ;
wire [16:0] \add_17s_17s_17_2_1_U28.dout ;
wire \add_17s_17s_17_2_1_U28.reset ;
wire [16:0] \add_17s_17s_17_2_1_U28.top_add_17s_17s_17_2_1_Adder_18_U.a ;
wire [16:0] \add_17s_17s_17_2_1_U28.top_add_17s_17s_17_2_1_Adder_18_U.ain_s0 ;
wire [16:0] \add_17s_17s_17_2_1_U28.top_add_17s_17s_17_2_1_Adder_18_U.b ;
wire [16:0] \add_17s_17s_17_2_1_U28.top_add_17s_17s_17_2_1_Adder_18_U.bin_s0 ;
wire \add_17s_17s_17_2_1_U28.top_add_17s_17s_17_2_1_Adder_18_U.ce ;
wire \add_17s_17s_17_2_1_U28.top_add_17s_17s_17_2_1_Adder_18_U.clk ;
wire \add_17s_17s_17_2_1_U28.top_add_17s_17s_17_2_1_Adder_18_U.facout_s1 ;
wire \add_17s_17s_17_2_1_U28.top_add_17s_17s_17_2_1_Adder_18_U.facout_s2 ;
wire [7:0] \add_17s_17s_17_2_1_U28.top_add_17s_17s_17_2_1_Adder_18_U.fas_s1 ;
wire [8:0] \add_17s_17s_17_2_1_U28.top_add_17s_17s_17_2_1_Adder_18_U.fas_s2 ;
wire \add_17s_17s_17_2_1_U28.top_add_17s_17s_17_2_1_Adder_18_U.reset ;
wire [16:0] \add_17s_17s_17_2_1_U28.top_add_17s_17s_17_2_1_Adder_18_U.s ;
wire [7:0] \add_17s_17s_17_2_1_U28.top_add_17s_17s_17_2_1_Adder_18_U.u1.a ;
wire [7:0] \add_17s_17s_17_2_1_U28.top_add_17s_17s_17_2_1_Adder_18_U.u1.b ;
wire \add_17s_17s_17_2_1_U28.top_add_17s_17s_17_2_1_Adder_18_U.u1.cin ;
wire \add_17s_17s_17_2_1_U28.top_add_17s_17s_17_2_1_Adder_18_U.u1.cout ;
wire [7:0] \add_17s_17s_17_2_1_U28.top_add_17s_17s_17_2_1_Adder_18_U.u1.s ;
wire [8:0] \add_17s_17s_17_2_1_U28.top_add_17s_17s_17_2_1_Adder_18_U.u2.a ;
wire [8:0] \add_17s_17s_17_2_1_U28.top_add_17s_17s_17_2_1_Adder_18_U.u2.b ;
wire \add_17s_17s_17_2_1_U28.top_add_17s_17s_17_2_1_Adder_18_U.u2.cin ;
wire \add_17s_17s_17_2_1_U28.top_add_17s_17s_17_2_1_Adder_18_U.u2.cout ;
wire [8:0] \add_17s_17s_17_2_1_U28.top_add_17s_17s_17_2_1_Adder_18_U.u2.s ;
wire \add_24s_24s_24_2_1_U16.ce ;
wire \add_24s_24s_24_2_1_U16.clk ;
wire [23:0] \add_24s_24s_24_2_1_U16.din0 ;
wire [23:0] \add_24s_24s_24_2_1_U16.din1 ;
wire [23:0] \add_24s_24s_24_2_1_U16.dout ;
wire \add_24s_24s_24_2_1_U16.reset ;
wire [23:0] \add_24s_24s_24_2_1_U16.top_add_24s_24s_24_2_1_Adder_12_U.a ;
wire [23:0] \add_24s_24s_24_2_1_U16.top_add_24s_24s_24_2_1_Adder_12_U.ain_s0 ;
wire [23:0] \add_24s_24s_24_2_1_U16.top_add_24s_24s_24_2_1_Adder_12_U.b ;
wire [23:0] \add_24s_24s_24_2_1_U16.top_add_24s_24s_24_2_1_Adder_12_U.bin_s0 ;
wire \add_24s_24s_24_2_1_U16.top_add_24s_24s_24_2_1_Adder_12_U.ce ;
wire \add_24s_24s_24_2_1_U16.top_add_24s_24s_24_2_1_Adder_12_U.clk ;
wire \add_24s_24s_24_2_1_U16.top_add_24s_24s_24_2_1_Adder_12_U.facout_s1 ;
wire \add_24s_24s_24_2_1_U16.top_add_24s_24s_24_2_1_Adder_12_U.facout_s2 ;
wire [11:0] \add_24s_24s_24_2_1_U16.top_add_24s_24s_24_2_1_Adder_12_U.fas_s1 ;
wire [11:0] \add_24s_24s_24_2_1_U16.top_add_24s_24s_24_2_1_Adder_12_U.fas_s2 ;
wire \add_24s_24s_24_2_1_U16.top_add_24s_24s_24_2_1_Adder_12_U.reset ;
wire [23:0] \add_24s_24s_24_2_1_U16.top_add_24s_24s_24_2_1_Adder_12_U.s ;
wire [11:0] \add_24s_24s_24_2_1_U16.top_add_24s_24s_24_2_1_Adder_12_U.u1.a ;
wire [11:0] \add_24s_24s_24_2_1_U16.top_add_24s_24s_24_2_1_Adder_12_U.u1.b ;
wire \add_24s_24s_24_2_1_U16.top_add_24s_24s_24_2_1_Adder_12_U.u1.cin ;
wire \add_24s_24s_24_2_1_U16.top_add_24s_24s_24_2_1_Adder_12_U.u1.cout ;
wire [11:0] \add_24s_24s_24_2_1_U16.top_add_24s_24s_24_2_1_Adder_12_U.u1.s ;
wire [11:0] \add_24s_24s_24_2_1_U16.top_add_24s_24s_24_2_1_Adder_12_U.u2.a ;
wire [11:0] \add_24s_24s_24_2_1_U16.top_add_24s_24s_24_2_1_Adder_12_U.u2.b ;
wire \add_24s_24s_24_2_1_U16.top_add_24s_24s_24_2_1_Adder_12_U.u2.cin ;
wire \add_24s_24s_24_2_1_U16.top_add_24s_24s_24_2_1_Adder_12_U.u2.cout ;
wire [11:0] \add_24s_24s_24_2_1_U16.top_add_24s_24s_24_2_1_Adder_12_U.u2.s ;
wire \add_2ns_2ns_2_2_1_U9.ce ;
wire \add_2ns_2ns_2_2_1_U9.clk ;
wire [1:0] \add_2ns_2ns_2_2_1_U9.din0 ;
wire [1:0] \add_2ns_2ns_2_2_1_U9.din1 ;
wire [1:0] \add_2ns_2ns_2_2_1_U9.dout ;
wire \add_2ns_2ns_2_2_1_U9.reset ;
wire [1:0] \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.a ;
wire [1:0] \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.ain_s0 ;
wire [1:0] \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.b ;
wire [1:0] \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.bin_s0 ;
wire \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.ce ;
wire \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.clk ;
wire \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.facout_s1 ;
wire \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.facout_s2 ;
wire \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.fas_s1 ;
wire \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.fas_s2 ;
wire \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.reset ;
wire [1:0] \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.s ;
wire \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.u1.a ;
wire \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.u1.b ;
wire \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.u1.cin ;
wire \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.u1.cout ;
wire \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.u1.s ;
wire \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.u2.a ;
wire \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.u2.b ;
wire \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.u2.cin ;
wire \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.u2.cout ;
wire \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.u2.s ;
wire \add_32ns_32ns_32_2_1_U20.ce ;
wire \add_32ns_32ns_32_2_1_U20.clk ;
wire [31:0] \add_32ns_32ns_32_2_1_U20.din0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U20.din1 ;
wire [31:0] \add_32ns_32ns_32_2_1_U20.dout ;
wire \add_32ns_32ns_32_2_1_U20.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_15_U.a ;
wire [31:0] \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_15_U.ain_s0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_15_U.b ;
wire [31:0] \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_15_U.bin_s0 ;
wire \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_15_U.ce ;
wire \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_15_U.clk ;
wire \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_15_U.facout_s1 ;
wire \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_15_U.facout_s2 ;
wire [15:0] \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_15_U.fas_s1 ;
wire [15:0] \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_15_U.fas_s2 ;
wire \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_15_U.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_15_U.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.b ;
wire \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.cin ;
wire \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.b ;
wire \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.cin ;
wire \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.s ;
wire \add_32ns_32ns_32_2_1_U22.ce ;
wire \add_32ns_32ns_32_2_1_U22.clk ;
wire [31:0] \add_32ns_32ns_32_2_1_U22.din0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U22.din1 ;
wire [31:0] \add_32ns_32ns_32_2_1_U22.dout ;
wire \add_32ns_32ns_32_2_1_U22.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_15_U.a ;
wire [31:0] \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_15_U.ain_s0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_15_U.b ;
wire [31:0] \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_15_U.bin_s0 ;
wire \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_15_U.ce ;
wire \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_15_U.clk ;
wire \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_15_U.facout_s1 ;
wire \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_15_U.facout_s2 ;
wire [15:0] \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_15_U.fas_s1 ;
wire [15:0] \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_15_U.fas_s2 ;
wire \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_15_U.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_15_U.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.b ;
wire \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.cin ;
wire \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.b ;
wire \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.cin ;
wire \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.s ;
wire \add_32ns_32ns_32_2_1_U23.ce ;
wire \add_32ns_32ns_32_2_1_U23.clk ;
wire [31:0] \add_32ns_32ns_32_2_1_U23.din0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U23.din1 ;
wire [31:0] \add_32ns_32ns_32_2_1_U23.dout ;
wire \add_32ns_32ns_32_2_1_U23.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.a ;
wire [31:0] \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.ain_s0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.b ;
wire [31:0] \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.bin_s0 ;
wire \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.ce ;
wire \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.clk ;
wire \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.facout_s1 ;
wire \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.facout_s2 ;
wire [15:0] \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.fas_s1 ;
wire [15:0] \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.fas_s2 ;
wire \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.b ;
wire \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.cin ;
wire \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.b ;
wire \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.cin ;
wire \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.s ;
wire \add_32ns_32ns_32_2_1_U25.ce ;
wire \add_32ns_32ns_32_2_1_U25.clk ;
wire [31:0] \add_32ns_32ns_32_2_1_U25.din0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U25.din1 ;
wire [31:0] \add_32ns_32ns_32_2_1_U25.dout ;
wire \add_32ns_32ns_32_2_1_U25.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.a ;
wire [31:0] \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.ain_s0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.b ;
wire [31:0] \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.bin_s0 ;
wire \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.ce ;
wire \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.clk ;
wire \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.facout_s1 ;
wire \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.facout_s2 ;
wire [15:0] \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.fas_s1 ;
wire [15:0] \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.fas_s2 ;
wire \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.b ;
wire \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.cin ;
wire \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.b ;
wire \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.cin ;
wire \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.s ;
wire \add_32ns_32ns_32_2_1_U27.ce ;
wire \add_32ns_32ns_32_2_1_U27.clk ;
wire [31:0] \add_32ns_32ns_32_2_1_U27.din0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U27.din1 ;
wire [31:0] \add_32ns_32ns_32_2_1_U27.dout ;
wire \add_32ns_32ns_32_2_1_U27.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U27.top_add_32ns_32ns_32_2_1_Adder_15_U.a ;
wire [31:0] \add_32ns_32ns_32_2_1_U27.top_add_32ns_32ns_32_2_1_Adder_15_U.ain_s0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U27.top_add_32ns_32ns_32_2_1_Adder_15_U.b ;
wire [31:0] \add_32ns_32ns_32_2_1_U27.top_add_32ns_32ns_32_2_1_Adder_15_U.bin_s0 ;
wire \add_32ns_32ns_32_2_1_U27.top_add_32ns_32ns_32_2_1_Adder_15_U.ce ;
wire \add_32ns_32ns_32_2_1_U27.top_add_32ns_32ns_32_2_1_Adder_15_U.clk ;
wire \add_32ns_32ns_32_2_1_U27.top_add_32ns_32ns_32_2_1_Adder_15_U.facout_s1 ;
wire \add_32ns_32ns_32_2_1_U27.top_add_32ns_32ns_32_2_1_Adder_15_U.facout_s2 ;
wire [15:0] \add_32ns_32ns_32_2_1_U27.top_add_32ns_32ns_32_2_1_Adder_15_U.fas_s1 ;
wire [15:0] \add_32ns_32ns_32_2_1_U27.top_add_32ns_32ns_32_2_1_Adder_15_U.fas_s2 ;
wire \add_32ns_32ns_32_2_1_U27.top_add_32ns_32ns_32_2_1_Adder_15_U.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U27.top_add_32ns_32ns_32_2_1_Adder_15_U.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U27.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U27.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.b ;
wire \add_32ns_32ns_32_2_1_U27.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.cin ;
wire \add_32ns_32ns_32_2_1_U27.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U27.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U27.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U27.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.b ;
wire \add_32ns_32ns_32_2_1_U27.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.cin ;
wire \add_32ns_32ns_32_2_1_U27.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U27.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.s ;
wire \add_32s_32ns_32_2_1_U29.ce ;
wire \add_32s_32ns_32_2_1_U29.clk ;
wire [31:0] \add_32s_32ns_32_2_1_U29.din0 ;
wire [31:0] \add_32s_32ns_32_2_1_U29.din1 ;
wire [31:0] \add_32s_32ns_32_2_1_U29.dout ;
wire \add_32s_32ns_32_2_1_U29.reset ;
wire [31:0] \add_32s_32ns_32_2_1_U29.top_add_32s_32ns_32_2_1_Adder_19_U.a ;
wire [31:0] \add_32s_32ns_32_2_1_U29.top_add_32s_32ns_32_2_1_Adder_19_U.ain_s0 ;
wire [31:0] \add_32s_32ns_32_2_1_U29.top_add_32s_32ns_32_2_1_Adder_19_U.b ;
wire [31:0] \add_32s_32ns_32_2_1_U29.top_add_32s_32ns_32_2_1_Adder_19_U.bin_s0 ;
wire \add_32s_32ns_32_2_1_U29.top_add_32s_32ns_32_2_1_Adder_19_U.ce ;
wire \add_32s_32ns_32_2_1_U29.top_add_32s_32ns_32_2_1_Adder_19_U.clk ;
wire \add_32s_32ns_32_2_1_U29.top_add_32s_32ns_32_2_1_Adder_19_U.facout_s1 ;
wire \add_32s_32ns_32_2_1_U29.top_add_32s_32ns_32_2_1_Adder_19_U.facout_s2 ;
wire [15:0] \add_32s_32ns_32_2_1_U29.top_add_32s_32ns_32_2_1_Adder_19_U.fas_s1 ;
wire [15:0] \add_32s_32ns_32_2_1_U29.top_add_32s_32ns_32_2_1_Adder_19_U.fas_s2 ;
wire \add_32s_32ns_32_2_1_U29.top_add_32s_32ns_32_2_1_Adder_19_U.reset ;
wire [31:0] \add_32s_32ns_32_2_1_U29.top_add_32s_32ns_32_2_1_Adder_19_U.s ;
wire [15:0] \add_32s_32ns_32_2_1_U29.top_add_32s_32ns_32_2_1_Adder_19_U.u1.a ;
wire [15:0] \add_32s_32ns_32_2_1_U29.top_add_32s_32ns_32_2_1_Adder_19_U.u1.b ;
wire \add_32s_32ns_32_2_1_U29.top_add_32s_32ns_32_2_1_Adder_19_U.u1.cin ;
wire \add_32s_32ns_32_2_1_U29.top_add_32s_32ns_32_2_1_Adder_19_U.u1.cout ;
wire [15:0] \add_32s_32ns_32_2_1_U29.top_add_32s_32ns_32_2_1_Adder_19_U.u1.s ;
wire [15:0] \add_32s_32ns_32_2_1_U29.top_add_32s_32ns_32_2_1_Adder_19_U.u2.a ;
wire [15:0] \add_32s_32ns_32_2_1_U29.top_add_32s_32ns_32_2_1_Adder_19_U.u2.b ;
wire \add_32s_32ns_32_2_1_U29.top_add_32s_32ns_32_2_1_Adder_19_U.u2.cin ;
wire \add_32s_32ns_32_2_1_U29.top_add_32s_32ns_32_2_1_Adder_19_U.u2.cout ;
wire [15:0] \add_32s_32ns_32_2_1_U29.top_add_32s_32ns_32_2_1_Adder_19_U.u2.s ;
wire \add_34s_34s_34_2_1_U24.ce ;
wire \add_34s_34s_34_2_1_U24.clk ;
wire [33:0] \add_34s_34s_34_2_1_U24.din0 ;
wire [33:0] \add_34s_34s_34_2_1_U24.din1 ;
wire [33:0] \add_34s_34s_34_2_1_U24.dout ;
wire \add_34s_34s_34_2_1_U24.reset ;
wire [33:0] \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_16_U.a ;
wire [33:0] \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_16_U.ain_s0 ;
wire [33:0] \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_16_U.b ;
wire [33:0] \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_16_U.bin_s0 ;
wire \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_16_U.ce ;
wire \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_16_U.clk ;
wire \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_16_U.facout_s1 ;
wire \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_16_U.facout_s2 ;
wire [16:0] \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_16_U.fas_s1 ;
wire [16:0] \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_16_U.fas_s2 ;
wire \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_16_U.reset ;
wire [33:0] \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_16_U.s ;
wire [16:0] \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_16_U.u1.a ;
wire [16:0] \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_16_U.u1.b ;
wire \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_16_U.u1.cin ;
wire \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_16_U.u1.cout ;
wire [16:0] \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_16_U.u1.s ;
wire [16:0] \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_16_U.u2.a ;
wire [16:0] \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_16_U.u2.b ;
wire \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_16_U.u2.cin ;
wire \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_16_U.u2.cout ;
wire [16:0] \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_16_U.u2.s ;
wire \add_35s_35s_35_2_1_U19.ce ;
wire \add_35s_35s_35_2_1_U19.clk ;
wire [34:0] \add_35s_35s_35_2_1_U19.din0 ;
wire [34:0] \add_35s_35s_35_2_1_U19.din1 ;
wire [34:0] \add_35s_35s_35_2_1_U19.dout ;
wire \add_35s_35s_35_2_1_U19.reset ;
wire [34:0] \add_35s_35s_35_2_1_U19.top_add_35s_35s_35_2_1_Adder_14_U.a ;
wire [34:0] \add_35s_35s_35_2_1_U19.top_add_35s_35s_35_2_1_Adder_14_U.ain_s0 ;
wire [34:0] \add_35s_35s_35_2_1_U19.top_add_35s_35s_35_2_1_Adder_14_U.b ;
wire [34:0] \add_35s_35s_35_2_1_U19.top_add_35s_35s_35_2_1_Adder_14_U.bin_s0 ;
wire \add_35s_35s_35_2_1_U19.top_add_35s_35s_35_2_1_Adder_14_U.ce ;
wire \add_35s_35s_35_2_1_U19.top_add_35s_35s_35_2_1_Adder_14_U.clk ;
wire \add_35s_35s_35_2_1_U19.top_add_35s_35s_35_2_1_Adder_14_U.facout_s1 ;
wire \add_35s_35s_35_2_1_U19.top_add_35s_35s_35_2_1_Adder_14_U.facout_s2 ;
wire [16:0] \add_35s_35s_35_2_1_U19.top_add_35s_35s_35_2_1_Adder_14_U.fas_s1 ;
wire [17:0] \add_35s_35s_35_2_1_U19.top_add_35s_35s_35_2_1_Adder_14_U.fas_s2 ;
wire \add_35s_35s_35_2_1_U19.top_add_35s_35s_35_2_1_Adder_14_U.reset ;
wire [34:0] \add_35s_35s_35_2_1_U19.top_add_35s_35s_35_2_1_Adder_14_U.s ;
wire [16:0] \add_35s_35s_35_2_1_U19.top_add_35s_35s_35_2_1_Adder_14_U.u1.a ;
wire [16:0] \add_35s_35s_35_2_1_U19.top_add_35s_35s_35_2_1_Adder_14_U.u1.b ;
wire \add_35s_35s_35_2_1_U19.top_add_35s_35s_35_2_1_Adder_14_U.u1.cin ;
wire \add_35s_35s_35_2_1_U19.top_add_35s_35s_35_2_1_Adder_14_U.u1.cout ;
wire [16:0] \add_35s_35s_35_2_1_U19.top_add_35s_35s_35_2_1_Adder_14_U.u1.s ;
wire [17:0] \add_35s_35s_35_2_1_U19.top_add_35s_35s_35_2_1_Adder_14_U.u2.a ;
wire [17:0] \add_35s_35s_35_2_1_U19.top_add_35s_35s_35_2_1_Adder_14_U.u2.b ;
wire \add_35s_35s_35_2_1_U19.top_add_35s_35s_35_2_1_Adder_14_U.u2.cin ;
wire \add_35s_35s_35_2_1_U19.top_add_35s_35s_35_2_1_Adder_14_U.u2.cout ;
wire [17:0] \add_35s_35s_35_2_1_U19.top_add_35s_35s_35_2_1_Adder_14_U.u2.s ;
wire \add_35s_35s_35_2_1_U21.ce ;
wire \add_35s_35s_35_2_1_U21.clk ;
wire [34:0] \add_35s_35s_35_2_1_U21.din0 ;
wire [34:0] \add_35s_35s_35_2_1_U21.din1 ;
wire [34:0] \add_35s_35s_35_2_1_U21.dout ;
wire \add_35s_35s_35_2_1_U21.reset ;
wire [34:0] \add_35s_35s_35_2_1_U21.top_add_35s_35s_35_2_1_Adder_14_U.a ;
wire [34:0] \add_35s_35s_35_2_1_U21.top_add_35s_35s_35_2_1_Adder_14_U.ain_s0 ;
wire [34:0] \add_35s_35s_35_2_1_U21.top_add_35s_35s_35_2_1_Adder_14_U.b ;
wire [34:0] \add_35s_35s_35_2_1_U21.top_add_35s_35s_35_2_1_Adder_14_U.bin_s0 ;
wire \add_35s_35s_35_2_1_U21.top_add_35s_35s_35_2_1_Adder_14_U.ce ;
wire \add_35s_35s_35_2_1_U21.top_add_35s_35s_35_2_1_Adder_14_U.clk ;
wire \add_35s_35s_35_2_1_U21.top_add_35s_35s_35_2_1_Adder_14_U.facout_s1 ;
wire \add_35s_35s_35_2_1_U21.top_add_35s_35s_35_2_1_Adder_14_U.facout_s2 ;
wire [16:0] \add_35s_35s_35_2_1_U21.top_add_35s_35s_35_2_1_Adder_14_U.fas_s1 ;
wire [17:0] \add_35s_35s_35_2_1_U21.top_add_35s_35s_35_2_1_Adder_14_U.fas_s2 ;
wire \add_35s_35s_35_2_1_U21.top_add_35s_35s_35_2_1_Adder_14_U.reset ;
wire [34:0] \add_35s_35s_35_2_1_U21.top_add_35s_35s_35_2_1_Adder_14_U.s ;
wire [16:0] \add_35s_35s_35_2_1_U21.top_add_35s_35s_35_2_1_Adder_14_U.u1.a ;
wire [16:0] \add_35s_35s_35_2_1_U21.top_add_35s_35s_35_2_1_Adder_14_U.u1.b ;
wire \add_35s_35s_35_2_1_U21.top_add_35s_35s_35_2_1_Adder_14_U.u1.cin ;
wire \add_35s_35s_35_2_1_U21.top_add_35s_35s_35_2_1_Adder_14_U.u1.cout ;
wire [16:0] \add_35s_35s_35_2_1_U21.top_add_35s_35s_35_2_1_Adder_14_U.u1.s ;
wire [17:0] \add_35s_35s_35_2_1_U21.top_add_35s_35s_35_2_1_Adder_14_U.u2.a ;
wire [17:0] \add_35s_35s_35_2_1_U21.top_add_35s_35s_35_2_1_Adder_14_U.u2.b ;
wire \add_35s_35s_35_2_1_U21.top_add_35s_35s_35_2_1_Adder_14_U.u2.cin ;
wire \add_35s_35s_35_2_1_U21.top_add_35s_35s_35_2_1_Adder_14_U.u2.cout ;
wire [17:0] \add_35s_35s_35_2_1_U21.top_add_35s_35s_35_2_1_Adder_14_U.u2.s ;
wire \add_3ns_3ns_3_2_1_U1.ce ;
wire \add_3ns_3ns_3_2_1_U1.clk ;
wire [2:0] \add_3ns_3ns_3_2_1_U1.din0 ;
wire [2:0] \add_3ns_3ns_3_2_1_U1.din1 ;
wire [2:0] \add_3ns_3ns_3_2_1_U1.dout ;
wire \add_3ns_3ns_3_2_1_U1.reset ;
wire [2:0] \add_3ns_3ns_3_2_1_U1.top_add_3ns_3ns_3_2_1_Adder_0_U.a ;
wire [2:0] \add_3ns_3ns_3_2_1_U1.top_add_3ns_3ns_3_2_1_Adder_0_U.ain_s0 ;
wire [2:0] \add_3ns_3ns_3_2_1_U1.top_add_3ns_3ns_3_2_1_Adder_0_U.b ;
wire [2:0] \add_3ns_3ns_3_2_1_U1.top_add_3ns_3ns_3_2_1_Adder_0_U.bin_s0 ;
wire \add_3ns_3ns_3_2_1_U1.top_add_3ns_3ns_3_2_1_Adder_0_U.ce ;
wire \add_3ns_3ns_3_2_1_U1.top_add_3ns_3ns_3_2_1_Adder_0_U.clk ;
wire \add_3ns_3ns_3_2_1_U1.top_add_3ns_3ns_3_2_1_Adder_0_U.facout_s1 ;
wire \add_3ns_3ns_3_2_1_U1.top_add_3ns_3ns_3_2_1_Adder_0_U.facout_s2 ;
wire \add_3ns_3ns_3_2_1_U1.top_add_3ns_3ns_3_2_1_Adder_0_U.fas_s1 ;
wire [1:0] \add_3ns_3ns_3_2_1_U1.top_add_3ns_3ns_3_2_1_Adder_0_U.fas_s2 ;
wire \add_3ns_3ns_3_2_1_U1.top_add_3ns_3ns_3_2_1_Adder_0_U.reset ;
wire [2:0] \add_3ns_3ns_3_2_1_U1.top_add_3ns_3ns_3_2_1_Adder_0_U.s ;
wire \add_3ns_3ns_3_2_1_U1.top_add_3ns_3ns_3_2_1_Adder_0_U.u1.a ;
wire \add_3ns_3ns_3_2_1_U1.top_add_3ns_3ns_3_2_1_Adder_0_U.u1.b ;
wire \add_3ns_3ns_3_2_1_U1.top_add_3ns_3ns_3_2_1_Adder_0_U.u1.cin ;
wire \add_3ns_3ns_3_2_1_U1.top_add_3ns_3ns_3_2_1_Adder_0_U.u1.cout ;
wire \add_3ns_3ns_3_2_1_U1.top_add_3ns_3ns_3_2_1_Adder_0_U.u1.s ;
wire [1:0] \add_3ns_3ns_3_2_1_U1.top_add_3ns_3ns_3_2_1_Adder_0_U.u2.a ;
wire [1:0] \add_3ns_3ns_3_2_1_U1.top_add_3ns_3ns_3_2_1_Adder_0_U.u2.b ;
wire \add_3ns_3ns_3_2_1_U1.top_add_3ns_3ns_3_2_1_Adder_0_U.u2.cin ;
wire \add_3ns_3ns_3_2_1_U1.top_add_3ns_3ns_3_2_1_Adder_0_U.u2.cout ;
wire [1:0] \add_3ns_3ns_3_2_1_U1.top_add_3ns_3ns_3_2_1_Adder_0_U.u2.s ;
wire \add_4ns_4ns_4_2_1_U18.ce ;
wire \add_4ns_4ns_4_2_1_U18.clk ;
wire [3:0] \add_4ns_4ns_4_2_1_U18.din0 ;
wire [3:0] \add_4ns_4ns_4_2_1_U18.din1 ;
wire [3:0] \add_4ns_4ns_4_2_1_U18.dout ;
wire \add_4ns_4ns_4_2_1_U18.reset ;
wire [3:0] \add_4ns_4ns_4_2_1_U18.top_add_4ns_4ns_4_2_1_Adder_5_U.a ;
wire [3:0] \add_4ns_4ns_4_2_1_U18.top_add_4ns_4ns_4_2_1_Adder_5_U.ain_s0 ;
wire [3:0] \add_4ns_4ns_4_2_1_U18.top_add_4ns_4ns_4_2_1_Adder_5_U.b ;
wire [3:0] \add_4ns_4ns_4_2_1_U18.top_add_4ns_4ns_4_2_1_Adder_5_U.bin_s0 ;
wire \add_4ns_4ns_4_2_1_U18.top_add_4ns_4ns_4_2_1_Adder_5_U.ce ;
wire \add_4ns_4ns_4_2_1_U18.top_add_4ns_4ns_4_2_1_Adder_5_U.clk ;
wire \add_4ns_4ns_4_2_1_U18.top_add_4ns_4ns_4_2_1_Adder_5_U.facout_s1 ;
wire \add_4ns_4ns_4_2_1_U18.top_add_4ns_4ns_4_2_1_Adder_5_U.facout_s2 ;
wire [1:0] \add_4ns_4ns_4_2_1_U18.top_add_4ns_4ns_4_2_1_Adder_5_U.fas_s1 ;
wire [1:0] \add_4ns_4ns_4_2_1_U18.top_add_4ns_4ns_4_2_1_Adder_5_U.fas_s2 ;
wire \add_4ns_4ns_4_2_1_U18.top_add_4ns_4ns_4_2_1_Adder_5_U.reset ;
wire [3:0] \add_4ns_4ns_4_2_1_U18.top_add_4ns_4ns_4_2_1_Adder_5_U.s ;
wire [1:0] \add_4ns_4ns_4_2_1_U18.top_add_4ns_4ns_4_2_1_Adder_5_U.u1.a ;
wire [1:0] \add_4ns_4ns_4_2_1_U18.top_add_4ns_4ns_4_2_1_Adder_5_U.u1.b ;
wire \add_4ns_4ns_4_2_1_U18.top_add_4ns_4ns_4_2_1_Adder_5_U.u1.cin ;
wire \add_4ns_4ns_4_2_1_U18.top_add_4ns_4ns_4_2_1_Adder_5_U.u1.cout ;
wire [1:0] \add_4ns_4ns_4_2_1_U18.top_add_4ns_4ns_4_2_1_Adder_5_U.u1.s ;
wire [1:0] \add_4ns_4ns_4_2_1_U18.top_add_4ns_4ns_4_2_1_Adder_5_U.u2.a ;
wire [1:0] \add_4ns_4ns_4_2_1_U18.top_add_4ns_4ns_4_2_1_Adder_5_U.u2.b ;
wire \add_4ns_4ns_4_2_1_U18.top_add_4ns_4ns_4_2_1_Adder_5_U.u2.cin ;
wire \add_4ns_4ns_4_2_1_U18.top_add_4ns_4ns_4_2_1_Adder_5_U.u2.cout ;
wire [1:0] \add_4ns_4ns_4_2_1_U18.top_add_4ns_4ns_4_2_1_Adder_5_U.u2.s ;
wire \add_4ns_4ns_4_2_1_U8.ce ;
wire \add_4ns_4ns_4_2_1_U8.clk ;
wire [3:0] \add_4ns_4ns_4_2_1_U8.din0 ;
wire [3:0] \add_4ns_4ns_4_2_1_U8.din1 ;
wire [3:0] \add_4ns_4ns_4_2_1_U8.dout ;
wire \add_4ns_4ns_4_2_1_U8.reset ;
wire [3:0] \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_5_U.a ;
wire [3:0] \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_5_U.ain_s0 ;
wire [3:0] \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_5_U.b ;
wire [3:0] \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_5_U.bin_s0 ;
wire \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_5_U.ce ;
wire \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_5_U.clk ;
wire \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_5_U.facout_s1 ;
wire \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_5_U.facout_s2 ;
wire [1:0] \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_5_U.fas_s1 ;
wire [1:0] \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_5_U.fas_s2 ;
wire \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_5_U.reset ;
wire [3:0] \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_5_U.s ;
wire [1:0] \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_5_U.u1.a ;
wire [1:0] \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_5_U.u1.b ;
wire \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_5_U.u1.cin ;
wire \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_5_U.u1.cout ;
wire [1:0] \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_5_U.u1.s ;
wire [1:0] \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_5_U.u2.a ;
wire [1:0] \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_5_U.u2.b ;
wire \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_5_U.u2.cin ;
wire \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_5_U.u2.cout ;
wire [1:0] \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_5_U.u2.s ;
wire \add_4s_4ns_4_2_1_U4.ce ;
wire \add_4s_4ns_4_2_1_U4.clk ;
wire [3:0] \add_4s_4ns_4_2_1_U4.din0 ;
wire [3:0] \add_4s_4ns_4_2_1_U4.din1 ;
wire [3:0] \add_4s_4ns_4_2_1_U4.dout ;
wire \add_4s_4ns_4_2_1_U4.reset ;
wire [3:0] \add_4s_4ns_4_2_1_U4.top_add_4s_4ns_4_2_1_Adder_3_U.a ;
wire [3:0] \add_4s_4ns_4_2_1_U4.top_add_4s_4ns_4_2_1_Adder_3_U.ain_s0 ;
wire [3:0] \add_4s_4ns_4_2_1_U4.top_add_4s_4ns_4_2_1_Adder_3_U.b ;
wire [3:0] \add_4s_4ns_4_2_1_U4.top_add_4s_4ns_4_2_1_Adder_3_U.bin_s0 ;
wire \add_4s_4ns_4_2_1_U4.top_add_4s_4ns_4_2_1_Adder_3_U.ce ;
wire \add_4s_4ns_4_2_1_U4.top_add_4s_4ns_4_2_1_Adder_3_U.clk ;
wire \add_4s_4ns_4_2_1_U4.top_add_4s_4ns_4_2_1_Adder_3_U.facout_s1 ;
wire \add_4s_4ns_4_2_1_U4.top_add_4s_4ns_4_2_1_Adder_3_U.facout_s2 ;
wire [1:0] \add_4s_4ns_4_2_1_U4.top_add_4s_4ns_4_2_1_Adder_3_U.fas_s1 ;
wire [1:0] \add_4s_4ns_4_2_1_U4.top_add_4s_4ns_4_2_1_Adder_3_U.fas_s2 ;
wire \add_4s_4ns_4_2_1_U4.top_add_4s_4ns_4_2_1_Adder_3_U.reset ;
wire [3:0] \add_4s_4ns_4_2_1_U4.top_add_4s_4ns_4_2_1_Adder_3_U.s ;
wire [1:0] \add_4s_4ns_4_2_1_U4.top_add_4s_4ns_4_2_1_Adder_3_U.u1.a ;
wire [1:0] \add_4s_4ns_4_2_1_U4.top_add_4s_4ns_4_2_1_Adder_3_U.u1.b ;
wire \add_4s_4ns_4_2_1_U4.top_add_4s_4ns_4_2_1_Adder_3_U.u1.cin ;
wire \add_4s_4ns_4_2_1_U4.top_add_4s_4ns_4_2_1_Adder_3_U.u1.cout ;
wire [1:0] \add_4s_4ns_4_2_1_U4.top_add_4s_4ns_4_2_1_Adder_3_U.u1.s ;
wire [1:0] \add_4s_4ns_4_2_1_U4.top_add_4s_4ns_4_2_1_Adder_3_U.u2.a ;
wire [1:0] \add_4s_4ns_4_2_1_U4.top_add_4s_4ns_4_2_1_Adder_3_U.u2.b ;
wire \add_4s_4ns_4_2_1_U4.top_add_4s_4ns_4_2_1_Adder_3_U.u2.cin ;
wire \add_4s_4ns_4_2_1_U4.top_add_4s_4ns_4_2_1_Adder_3_U.u2.cout ;
wire [1:0] \add_4s_4ns_4_2_1_U4.top_add_4s_4ns_4_2_1_Adder_3_U.u2.s ;
wire \add_5ns_5s_5_2_1_U3.ce ;
wire \add_5ns_5s_5_2_1_U3.clk ;
wire [4:0] \add_5ns_5s_5_2_1_U3.din0 ;
wire [4:0] \add_5ns_5s_5_2_1_U3.din1 ;
wire [4:0] \add_5ns_5s_5_2_1_U3.dout ;
wire \add_5ns_5s_5_2_1_U3.reset ;
wire [4:0] \add_5ns_5s_5_2_1_U3.top_add_5ns_5s_5_2_1_Adder_2_U.a ;
wire [4:0] \add_5ns_5s_5_2_1_U3.top_add_5ns_5s_5_2_1_Adder_2_U.ain_s0 ;
wire [4:0] \add_5ns_5s_5_2_1_U3.top_add_5ns_5s_5_2_1_Adder_2_U.b ;
wire [4:0] \add_5ns_5s_5_2_1_U3.top_add_5ns_5s_5_2_1_Adder_2_U.bin_s0 ;
wire \add_5ns_5s_5_2_1_U3.top_add_5ns_5s_5_2_1_Adder_2_U.ce ;
wire \add_5ns_5s_5_2_1_U3.top_add_5ns_5s_5_2_1_Adder_2_U.clk ;
wire \add_5ns_5s_5_2_1_U3.top_add_5ns_5s_5_2_1_Adder_2_U.facout_s1 ;
wire \add_5ns_5s_5_2_1_U3.top_add_5ns_5s_5_2_1_Adder_2_U.facout_s2 ;
wire [1:0] \add_5ns_5s_5_2_1_U3.top_add_5ns_5s_5_2_1_Adder_2_U.fas_s1 ;
wire [2:0] \add_5ns_5s_5_2_1_U3.top_add_5ns_5s_5_2_1_Adder_2_U.fas_s2 ;
wire \add_5ns_5s_5_2_1_U3.top_add_5ns_5s_5_2_1_Adder_2_U.reset ;
wire [4:0] \add_5ns_5s_5_2_1_U3.top_add_5ns_5s_5_2_1_Adder_2_U.s ;
wire [1:0] \add_5ns_5s_5_2_1_U3.top_add_5ns_5s_5_2_1_Adder_2_U.u1.a ;
wire [1:0] \add_5ns_5s_5_2_1_U3.top_add_5ns_5s_5_2_1_Adder_2_U.u1.b ;
wire \add_5ns_5s_5_2_1_U3.top_add_5ns_5s_5_2_1_Adder_2_U.u1.cin ;
wire \add_5ns_5s_5_2_1_U3.top_add_5ns_5s_5_2_1_Adder_2_U.u1.cout ;
wire [1:0] \add_5ns_5s_5_2_1_U3.top_add_5ns_5s_5_2_1_Adder_2_U.u1.s ;
wire [2:0] \add_5ns_5s_5_2_1_U3.top_add_5ns_5s_5_2_1_Adder_2_U.u2.a ;
wire [2:0] \add_5ns_5s_5_2_1_U3.top_add_5ns_5s_5_2_1_Adder_2_U.u2.b ;
wire \add_5ns_5s_5_2_1_U3.top_add_5ns_5s_5_2_1_Adder_2_U.u2.cin ;
wire \add_5ns_5s_5_2_1_U3.top_add_5ns_5s_5_2_1_Adder_2_U.u2.cout ;
wire [2:0] \add_5ns_5s_5_2_1_U3.top_add_5ns_5s_5_2_1_Adder_2_U.u2.s ;
wire \add_7s_7s_7_2_1_U2.ce ;
wire \add_7s_7s_7_2_1_U2.clk ;
wire [6:0] \add_7s_7s_7_2_1_U2.din0 ;
wire [6:0] \add_7s_7s_7_2_1_U2.din1 ;
wire [6:0] \add_7s_7s_7_2_1_U2.dout ;
wire \add_7s_7s_7_2_1_U2.reset ;
wire [6:0] \add_7s_7s_7_2_1_U2.top_add_7s_7s_7_2_1_Adder_1_U.a ;
wire [6:0] \add_7s_7s_7_2_1_U2.top_add_7s_7s_7_2_1_Adder_1_U.ain_s0 ;
wire [6:0] \add_7s_7s_7_2_1_U2.top_add_7s_7s_7_2_1_Adder_1_U.b ;
wire [6:0] \add_7s_7s_7_2_1_U2.top_add_7s_7s_7_2_1_Adder_1_U.bin_s0 ;
wire \add_7s_7s_7_2_1_U2.top_add_7s_7s_7_2_1_Adder_1_U.ce ;
wire \add_7s_7s_7_2_1_U2.top_add_7s_7s_7_2_1_Adder_1_U.clk ;
wire \add_7s_7s_7_2_1_U2.top_add_7s_7s_7_2_1_Adder_1_U.facout_s1 ;
wire \add_7s_7s_7_2_1_U2.top_add_7s_7s_7_2_1_Adder_1_U.facout_s2 ;
wire [2:0] \add_7s_7s_7_2_1_U2.top_add_7s_7s_7_2_1_Adder_1_U.fas_s1 ;
wire [3:0] \add_7s_7s_7_2_1_U2.top_add_7s_7s_7_2_1_Adder_1_U.fas_s2 ;
wire \add_7s_7s_7_2_1_U2.top_add_7s_7s_7_2_1_Adder_1_U.reset ;
wire [6:0] \add_7s_7s_7_2_1_U2.top_add_7s_7s_7_2_1_Adder_1_U.s ;
wire [2:0] \add_7s_7s_7_2_1_U2.top_add_7s_7s_7_2_1_Adder_1_U.u1.a ;
wire [2:0] \add_7s_7s_7_2_1_U2.top_add_7s_7s_7_2_1_Adder_1_U.u1.b ;
wire \add_7s_7s_7_2_1_U2.top_add_7s_7s_7_2_1_Adder_1_U.u1.cin ;
wire \add_7s_7s_7_2_1_U2.top_add_7s_7s_7_2_1_Adder_1_U.u1.cout ;
wire [2:0] \add_7s_7s_7_2_1_U2.top_add_7s_7s_7_2_1_Adder_1_U.u1.s ;
wire [3:0] \add_7s_7s_7_2_1_U2.top_add_7s_7s_7_2_1_Adder_1_U.u2.a ;
wire [3:0] \add_7s_7s_7_2_1_U2.top_add_7s_7s_7_2_1_Adder_1_U.u2.b ;
wire \add_7s_7s_7_2_1_U2.top_add_7s_7s_7_2_1_Adder_1_U.u2.cin ;
wire \add_7s_7s_7_2_1_U2.top_add_7s_7s_7_2_1_Adder_1_U.u2.cout ;
wire [3:0] \add_7s_7s_7_2_1_U2.top_add_7s_7s_7_2_1_Adder_1_U.u2.s ;
wire \add_9s_9ns_9_2_1_U26.ce ;
wire \add_9s_9ns_9_2_1_U26.clk ;
wire [8:0] \add_9s_9ns_9_2_1_U26.din0 ;
wire [8:0] \add_9s_9ns_9_2_1_U26.din1 ;
wire [8:0] \add_9s_9ns_9_2_1_U26.dout ;
wire \add_9s_9ns_9_2_1_U26.reset ;
wire [8:0] \add_9s_9ns_9_2_1_U26.top_add_9s_9ns_9_2_1_Adder_17_U.a ;
wire [8:0] \add_9s_9ns_9_2_1_U26.top_add_9s_9ns_9_2_1_Adder_17_U.ain_s0 ;
wire [8:0] \add_9s_9ns_9_2_1_U26.top_add_9s_9ns_9_2_1_Adder_17_U.b ;
wire [8:0] \add_9s_9ns_9_2_1_U26.top_add_9s_9ns_9_2_1_Adder_17_U.bin_s0 ;
wire \add_9s_9ns_9_2_1_U26.top_add_9s_9ns_9_2_1_Adder_17_U.ce ;
wire \add_9s_9ns_9_2_1_U26.top_add_9s_9ns_9_2_1_Adder_17_U.clk ;
wire \add_9s_9ns_9_2_1_U26.top_add_9s_9ns_9_2_1_Adder_17_U.facout_s1 ;
wire \add_9s_9ns_9_2_1_U26.top_add_9s_9ns_9_2_1_Adder_17_U.facout_s2 ;
wire [3:0] \add_9s_9ns_9_2_1_U26.top_add_9s_9ns_9_2_1_Adder_17_U.fas_s1 ;
wire [4:0] \add_9s_9ns_9_2_1_U26.top_add_9s_9ns_9_2_1_Adder_17_U.fas_s2 ;
wire \add_9s_9ns_9_2_1_U26.top_add_9s_9ns_9_2_1_Adder_17_U.reset ;
wire [8:0] \add_9s_9ns_9_2_1_U26.top_add_9s_9ns_9_2_1_Adder_17_U.s ;
wire [3:0] \add_9s_9ns_9_2_1_U26.top_add_9s_9ns_9_2_1_Adder_17_U.u1.a ;
wire [3:0] \add_9s_9ns_9_2_1_U26.top_add_9s_9ns_9_2_1_Adder_17_U.u1.b ;
wire \add_9s_9ns_9_2_1_U26.top_add_9s_9ns_9_2_1_Adder_17_U.u1.cin ;
wire \add_9s_9ns_9_2_1_U26.top_add_9s_9ns_9_2_1_Adder_17_U.u1.cout ;
wire [3:0] \add_9s_9ns_9_2_1_U26.top_add_9s_9ns_9_2_1_Adder_17_U.u1.s ;
wire [4:0] \add_9s_9ns_9_2_1_U26.top_add_9s_9ns_9_2_1_Adder_17_U.u2.a ;
wire [4:0] \add_9s_9ns_9_2_1_U26.top_add_9s_9ns_9_2_1_Adder_17_U.u2.b ;
wire \add_9s_9ns_9_2_1_U26.top_add_9s_9ns_9_2_1_Adder_17_U.u2.cin ;
wire \add_9s_9ns_9_2_1_U26.top_add_9s_9ns_9_2_1_Adder_17_U.u2.cout ;
wire [4:0] \add_9s_9ns_9_2_1_U26.top_add_9s_9ns_9_2_1_Adder_17_U.u2.s ;
wire and_ln340_1_fu_572_p2;
wire and_ln340_2_fu_584_p2;
wire and_ln340_3_fu_1152_p2;
wire and_ln340_4_fu_1381_p2;
wire and_ln340_5_fu_1394_p2;
wire and_ln340_fu_332_p2;
wire and_ln412_fu_741_p2;
wire and_ln780_fu_972_p2;
wire and_ln781_fu_1087_p2;
wire and_ln785_10_fu_1247_p2;
wire and_ln785_12_fu_1434_p2;
wire and_ln785_13_fu_1398_p2;
wire and_ln785_1_fu_378_p2;
wire and_ln785_3_fu_614_p2;
wire and_ln785_4_fu_588_p2;
wire and_ln785_6_fu_1206_p2;
wire and_ln785_7_fu_1215_p2;
wire and_ln785_9_fu_1241_p2;
wire and_ln785_fu_372_p2;
wire and_ln786_1_fu_514_p2;
wire and_ln786_2_fu_1292_p2;
wire and_ln786_fu_983_p2;
wire ap_CS_fsm_state1;
wire ap_CS_fsm_state10;
wire ap_CS_fsm_state11;
wire ap_CS_fsm_state12;
wire ap_CS_fsm_state13;
wire ap_CS_fsm_state19;
wire ap_CS_fsm_state2;
wire ap_CS_fsm_state20;
wire ap_CS_fsm_state21;
wire ap_CS_fsm_state22;
wire ap_CS_fsm_state23;
wire ap_CS_fsm_state24;
wire ap_CS_fsm_state25;
wire ap_CS_fsm_state26;
wire ap_CS_fsm_state27;
wire ap_CS_fsm_state28;
wire ap_CS_fsm_state29;
wire ap_CS_fsm_state3;
wire ap_CS_fsm_state30;
wire ap_CS_fsm_state31;
wire ap_CS_fsm_state32;
wire ap_CS_fsm_state33;
wire ap_CS_fsm_state34;
wire ap_CS_fsm_state35;
wire ap_CS_fsm_state36;
wire ap_CS_fsm_state37;
wire ap_CS_fsm_state38;
wire ap_CS_fsm_state39;
wire ap_CS_fsm_state4;
wire ap_CS_fsm_state40;
wire ap_CS_fsm_state41;
wire ap_CS_fsm_state42;
wire ap_CS_fsm_state43;
wire ap_CS_fsm_state44;
wire ap_CS_fsm_state45;
wire ap_CS_fsm_state46;
wire ap_CS_fsm_state47;
wire ap_CS_fsm_state48;
wire ap_CS_fsm_state49;
wire ap_CS_fsm_state5;
wire ap_CS_fsm_state50;
wire ap_CS_fsm_state51;
wire ap_CS_fsm_state52;
wire ap_CS_fsm_state6;
wire ap_CS_fsm_state7;
wire ap_CS_fsm_state8;
wire ap_CS_fsm_state9;
wire [51:0] ap_NS_fsm;
wire ap_clk;
wire ap_done;
wire ap_idle;
wire ap_ready;
wire ap_rst;
wire ap_start;
wire carry_1_fu_895_p2;
wire deleted_ones_fu_977_p3;
wire deleted_zeros_fu_954_p3;
wire [23:0] grp_fu_1181_p0;
wire [23:0] grp_fu_1181_p1;
wire [23:0] grp_fu_1181_p2;
wire [11:0] grp_fu_1314_p0;
wire [11:0] grp_fu_1314_p2;
wire [3:0] grp_fu_1419_p2;
wire [34:0] grp_fu_1510_p0;
wire [34:0] grp_fu_1510_p1;
wire [34:0] grp_fu_1510_p2;
wire [31:0] grp_fu_1531_p2;
wire [34:0] grp_fu_1569_p0;
wire [34:0] grp_fu_1569_p1;
wire [34:0] grp_fu_1569_p2;
wire [31:0] grp_fu_1585_p2;
wire [31:0] grp_fu_1612_p1;
wire [31:0] grp_fu_1612_p2;
wire [33:0] grp_fu_1631_p0;
wire [33:0] grp_fu_1631_p1;
wire [33:0] grp_fu_1631_p2;
wire [31:0] grp_fu_1647_p2;
wire [8:0] grp_fu_1659_p0;
wire [8:0] grp_fu_1659_p1;
wire [8:0] grp_fu_1659_p2;
wire [31:0] grp_fu_1692_p2;
wire [16:0] grp_fu_1700_p0;
wire [16:0] grp_fu_1700_p1;
wire [16:0] grp_fu_1700_p2;
wire [31:0] grp_fu_1709_p0;
wire [31:0] grp_fu_1709_p2;
wire [2:0] grp_fu_279_p0;
wire [2:0] grp_fu_279_p2;
wire [6:0] grp_fu_428_p0;
wire [6:0] grp_fu_428_p1;
wire [6:0] grp_fu_428_p2;
wire [4:0] grp_fu_434_p0;
wire [4:0] grp_fu_434_p1;
wire [4:0] grp_fu_434_p2;
wire [3:0] grp_fu_440_p1;
wire [3:0] grp_fu_440_p2;
wire [31:0] grp_fu_641_p0;
wire [35:0] grp_fu_641_p2;
wire [31:0] grp_fu_650_p0;
wire [35:0] grp_fu_650_p2;
wire [7:0] grp_fu_735_p0;
wire [7:0] grp_fu_735_p1;
wire [7:0] grp_fu_735_p2;
wire [3:0] grp_fu_765_p2;
wire [1:0] grp_fu_773_p1;
wire [1:0] grp_fu_773_p2;
wire [12:0] grp_fu_820_p0;
wire [12:0] grp_fu_820_p1;
wire [12:0] grp_fu_820_p2;
wire [16:0] grp_fu_880_p0;
wire [16:0] grp_fu_880_p1;
wire [16:0] grp_fu_880_p2;
wire [3:0] grp_fu_889_p0;
wire [6:0] grp_fu_889_p00;
wire [6:0] grp_fu_889_p2;
wire [9:0] grp_fu_899_p2;
wire [32:0] grp_fu_940_p0;
wire [32:0] grp_fu_940_p1;
wire [32:0] grp_fu_940_p2;
wire [7:0] grp_fu_949_p1;
wire [7:0] grp_fu_949_p2;
wire icmp_ln768_1_fu_471_p2;
wire icmp_ln768_3_fu_988_p2;
wire icmp_ln768_4_fu_1077_p2;
wire icmp_ln768_fu_273_p2;
wire icmp_ln786_1_fu_476_p2;
wire icmp_ln786_2_fu_993_p2;
wire icmp_ln786_3_fu_1082_p2;
wire icmp_ln786_fu_293_p2;
wire icmp_ln851_1_fu_830_p2;
wire icmp_ln851_2_fu_1191_p2;
wire icmp_ln851_3_fu_1516_p2;
wire icmp_ln851_4_fu_1414_p2;
wire icmp_ln851_fu_760_p2;
wire [5:0] lhs_fu_399_p3;
wire \mul_32ns_4s_36_7_1_U5.ce ;
wire \mul_32ns_4s_36_7_1_U5.clk ;
wire [31:0] \mul_32ns_4s_36_7_1_U5.din0 ;
wire [3:0] \mul_32ns_4s_36_7_1_U5.din1 ;
wire [35:0] \mul_32ns_4s_36_7_1_U5.dout ;
wire \mul_32ns_4s_36_7_1_U5.reset ;
wire [31:0] \mul_32ns_4s_36_7_1_U5.top_mul_32ns_4s_36_7_1_Mul_DSP_0_U.a ;
wire [3:0] \mul_32ns_4s_36_7_1_U5.top_mul_32ns_4s_36_7_1_Mul_DSP_0_U.b ;
wire \mul_32ns_4s_36_7_1_U5.top_mul_32ns_4s_36_7_1_Mul_DSP_0_U.ce ;
wire \mul_32ns_4s_36_7_1_U5.top_mul_32ns_4s_36_7_1_Mul_DSP_0_U.clk ;
wire [35:0] \mul_32ns_4s_36_7_1_U5.top_mul_32ns_4s_36_7_1_Mul_DSP_0_U.p ;
wire [35:0] \mul_32ns_4s_36_7_1_U5.top_mul_32ns_4s_36_7_1_Mul_DSP_0_U.tmp_product ;
wire \mul_32ns_4s_36_7_1_U6.ce ;
wire \mul_32ns_4s_36_7_1_U6.clk ;
wire [31:0] \mul_32ns_4s_36_7_1_U6.din0 ;
wire [3:0] \mul_32ns_4s_36_7_1_U6.din1 ;
wire [35:0] \mul_32ns_4s_36_7_1_U6.dout ;
wire \mul_32ns_4s_36_7_1_U6.reset ;
wire [31:0] \mul_32ns_4s_36_7_1_U6.top_mul_32ns_4s_36_7_1_Mul_DSP_0_U.a ;
wire [3:0] \mul_32ns_4s_36_7_1_U6.top_mul_32ns_4s_36_7_1_Mul_DSP_0_U.b ;
wire \mul_32ns_4s_36_7_1_U6.top_mul_32ns_4s_36_7_1_Mul_DSP_0_U.ce ;
wire \mul_32ns_4s_36_7_1_U6.top_mul_32ns_4s_36_7_1_Mul_DSP_0_U.clk ;
wire [35:0] \mul_32ns_4s_36_7_1_U6.top_mul_32ns_4s_36_7_1_Mul_DSP_0_U.p ;
wire [35:0] \mul_32ns_4s_36_7_1_U6.top_mul_32ns_4s_36_7_1_Mul_DSP_0_U.tmp_product ;
wire \mul_4ns_3s_7_7_1_U12.ce ;
wire \mul_4ns_3s_7_7_1_U12.clk ;
wire [3:0] \mul_4ns_3s_7_7_1_U12.din0 ;
wire [2:0] \mul_4ns_3s_7_7_1_U12.din1 ;
wire [6:0] \mul_4ns_3s_7_7_1_U12.dout ;
wire \mul_4ns_3s_7_7_1_U12.reset ;
wire [3:0] \mul_4ns_3s_7_7_1_U12.top_mul_4ns_3s_7_7_1_Mul_DSP_1_U.a ;
wire [2:0] \mul_4ns_3s_7_7_1_U12.top_mul_4ns_3s_7_7_1_Mul_DSP_1_U.b ;
wire \mul_4ns_3s_7_7_1_U12.top_mul_4ns_3s_7_7_1_Mul_DSP_1_U.ce ;
wire \mul_4ns_3s_7_7_1_U12.top_mul_4ns_3s_7_7_1_Mul_DSP_1_U.clk ;
wire [6:0] \mul_4ns_3s_7_7_1_U12.top_mul_4ns_3s_7_7_1_Mul_DSP_1_U.p ;
wire [6:0] \mul_4ns_3s_7_7_1_U12.top_mul_4ns_3s_7_7_1_Mul_DSP_1_U.tmp_product ;
wire neg_src_fu_1097_p2;
wire [3:0] op_0;
wire [15:0] op_11;
wire [7:0] op_12_V_fu_1452_p3;
wire [15:0] op_13_V_fu_1252_p3;
wire [1:0] op_15_V_fu_1220_p3;
wire [15:0] op_16;
wire [31:0] op_17;
wire [3:0] op_18;
wire [3:0] op_1_V_fu_383_p3;
wire [31:0] op_29;
wire op_29_ap_vld;
wire [3:0] op_3_V_fu_625_p3;
wire [7:0] op_6;
wire [15:0] op_7;
wire [3:0] op_8;
wire or_ln340_1_fu_504_p2;
wire or_ln340_2_fu_1049_p2;
wire or_ln340_3_fu_1141_p2;
wire or_ln340_4_fu_1282_p2;
wire or_ln340_5_fu_1102_p2;
wire or_ln340_fu_321_p2;
wire or_ln785_10_fu_1429_p2;
wire or_ln785_11_fu_1402_p2;
wire or_ln785_1_fu_481_p2;
wire or_ln785_2_fu_1033_p2;
wire or_ln785_3_fu_1061_p2;
wire or_ln785_4_fu_1197_p2;
wire or_ln785_5_fu_367_p2;
wire or_ln785_6_fu_609_p2;
wire or_ln785_7_fu_592_p2;
wire or_ln785_8_fu_1210_p2;
wire or_ln785_9_fu_1236_p2;
wire or_ln785_fu_289_p2;
wire or_ln786_1_fu_499_p2;
wire or_ln786_2_fu_1136_p2;
wire or_ln786_3_fu_1277_p2;
wire or_ln786_fu_316_p2;
wire overflow_1_fu_490_p2;
wire overflow_2_fu_1043_p2;
wire overflow_3_fu_1126_p2;
wire overflow_4_fu_1268_p2;
wire overflow_fu_306_p2;
wire p_Result_13_fu_786_p3;
wire p_Result_14_fu_1054_p3;
wire p_Result_17_fu_1473_p3;
wire p_Result_18_fu_1445_p3;
wire [7:0] p_Result_22_fu_1366_p4;
wire p_Result_23_fu_1536_p3;
wire p_Result_24_fu_1590_p3;
wire p_Result_25_fu_1665_p3;
wire p_Result_26_fu_257_p2;
wire p_Result_29_fu_519_p3;
wire p_Result_31_fu_656_p1;
wire p_Result_38_fu_1327_p3;
wire [3:0] p_Result_7_fu_557_p4;
wire [15:0] p_Val2_10_fu_1114_p3;
wire [7:0] p_Val2_14_fu_1320_p3;
wire [6:0] p_Val2_15_fu_1360_p2;
wire [2:0] p_Val2_3_fu_552_p2;
wire [3:0] p_Val2_s_fu_251_p2;
wire [2:0] ret_V_16_fu_351_p3;
wire [3:0] ret_V_18_fu_798_p3;
wire [3:0] ret_V_20_fu_1489_p3;
wire [31:0] ret_V_24_fu_1602_p3;
wire [31:0] ret_V_26_fu_1681_p3;
wire [2:0] ret_V_fu_263_p4;
wire [10:0] rhs_2_fu_809_p3;
wire [22:0] rhs_3_fu_1170_p3;
wire rhs_4_fu_868_p2;
wire [33:0] rhs_5_fu_1558_p3;
wire [32:0] rhs_7_fu_1620_p3;
wire sel_tmp19_fu_598_p2;
wire sel_tmp51_fu_1408_p2;
wire [3:0] select_ln340_1_fu_577_p3;
wire [1:0] select_ln340_2_fu_1107_p3;
wire [15:0] select_ln340_3_fu_1158_p3;
wire [7:0] select_ln340_4_fu_1386_p3;
wire [3:0] select_ln340_fu_338_p3;
wire [31:0] select_ln353_1_fu_1548_p3;
wire [11:0] select_ln353_fu_1462_p3;
wire [7:0] select_ln785_3_fu_1439_p3;
wire [3:0] select_ln785_fu_619_p3;
wire [3:0] select_ln850_1_fu_793_p3;
wire [3:0] select_ln850_2_fu_1483_p3;
wire [9:0] select_ln850_3_fu_1065_p3;
wire [9:0] select_ln850_4_fu_1070_p3;
wire [11:0] select_ln850_5_fu_1457_p3;
wire [31:0] select_ln850_6_fu_1597_p3;
wire [31:0] select_ln850_7_fu_1675_p3;
wire [31:0] select_ln850_8_fu_1543_p3;
wire [2:0] select_ln850_fu_345_p3;
wire [31:0] sext_ln1116_fu_630_p1;
wire [15:0] sext_ln1192_2_fu_1166_p0;
wire [7:0] sext_ln703_1_fu_805_p0;
wire [7:0] sext_ln727_fu_851_p1;
wire [11:0] sext_ln850_fu_1311_p1;
wire [6:0] shl_ln_fu_857_p3;
wire \sub_17ns_17ns_17_2_1_U11.ce ;
wire \sub_17ns_17ns_17_2_1_U11.clk ;
wire [16:0] \sub_17ns_17ns_17_2_1_U11.din0 ;
wire [16:0] \sub_17ns_17ns_17_2_1_U11.din1 ;
wire [16:0] \sub_17ns_17ns_17_2_1_U11.dout ;
wire \sub_17ns_17ns_17_2_1_U11.reset ;
wire [16:0] \sub_17ns_17ns_17_2_1_U11.top_sub_17ns_17ns_17_2_1_Adder_8_U.a ;
wire [16:0] \sub_17ns_17ns_17_2_1_U11.top_sub_17ns_17ns_17_2_1_Adder_8_U.ain_s0 ;
wire [16:0] \sub_17ns_17ns_17_2_1_U11.top_sub_17ns_17ns_17_2_1_Adder_8_U.b ;
wire [16:0] \sub_17ns_17ns_17_2_1_U11.top_sub_17ns_17ns_17_2_1_Adder_8_U.bin_s0 ;
wire \sub_17ns_17ns_17_2_1_U11.top_sub_17ns_17ns_17_2_1_Adder_8_U.ce ;
wire \sub_17ns_17ns_17_2_1_U11.top_sub_17ns_17ns_17_2_1_Adder_8_U.clk ;
wire \sub_17ns_17ns_17_2_1_U11.top_sub_17ns_17ns_17_2_1_Adder_8_U.facout_s1 ;
wire \sub_17ns_17ns_17_2_1_U11.top_sub_17ns_17ns_17_2_1_Adder_8_U.facout_s2 ;
wire [7:0] \sub_17ns_17ns_17_2_1_U11.top_sub_17ns_17ns_17_2_1_Adder_8_U.fas_s1 ;
wire [8:0] \sub_17ns_17ns_17_2_1_U11.top_sub_17ns_17ns_17_2_1_Adder_8_U.fas_s2 ;
wire \sub_17ns_17ns_17_2_1_U11.top_sub_17ns_17ns_17_2_1_Adder_8_U.reset ;
wire [16:0] \sub_17ns_17ns_17_2_1_U11.top_sub_17ns_17ns_17_2_1_Adder_8_U.s ;
wire [7:0] \sub_17ns_17ns_17_2_1_U11.top_sub_17ns_17ns_17_2_1_Adder_8_U.u1.a ;
wire [7:0] \sub_17ns_17ns_17_2_1_U11.top_sub_17ns_17ns_17_2_1_Adder_8_U.u1.b ;
wire \sub_17ns_17ns_17_2_1_U11.top_sub_17ns_17ns_17_2_1_Adder_8_U.u1.cin ;
wire \sub_17ns_17ns_17_2_1_U11.top_sub_17ns_17ns_17_2_1_Adder_8_U.u1.cout ;
wire [7:0] \sub_17ns_17ns_17_2_1_U11.top_sub_17ns_17ns_17_2_1_Adder_8_U.u1.s ;
wire [8:0] \sub_17ns_17ns_17_2_1_U11.top_sub_17ns_17ns_17_2_1_Adder_8_U.u2.a ;
wire [8:0] \sub_17ns_17ns_17_2_1_U11.top_sub_17ns_17ns_17_2_1_Adder_8_U.u2.b ;
wire \sub_17ns_17ns_17_2_1_U11.top_sub_17ns_17ns_17_2_1_Adder_8_U.u2.cin ;
wire \sub_17ns_17ns_17_2_1_U11.top_sub_17ns_17ns_17_2_1_Adder_8_U.u2.cout ;
wire [8:0] \sub_17ns_17ns_17_2_1_U11.top_sub_17ns_17ns_17_2_1_Adder_8_U.u2.s ;
wire \sub_33ns_33ns_33_2_1_U14.ce ;
wire \sub_33ns_33ns_33_2_1_U14.clk ;
wire [32:0] \sub_33ns_33ns_33_2_1_U14.din0 ;
wire [32:0] \sub_33ns_33ns_33_2_1_U14.din1 ;
wire [32:0] \sub_33ns_33ns_33_2_1_U14.dout ;
wire \sub_33ns_33ns_33_2_1_U14.reset ;
wire [32:0] \sub_33ns_33ns_33_2_1_U14.top_sub_33ns_33ns_33_2_1_Adder_10_U.a ;
wire [32:0] \sub_33ns_33ns_33_2_1_U14.top_sub_33ns_33ns_33_2_1_Adder_10_U.ain_s0 ;
wire [32:0] \sub_33ns_33ns_33_2_1_U14.top_sub_33ns_33ns_33_2_1_Adder_10_U.b ;
wire [32:0] \sub_33ns_33ns_33_2_1_U14.top_sub_33ns_33ns_33_2_1_Adder_10_U.bin_s0 ;
wire \sub_33ns_33ns_33_2_1_U14.top_sub_33ns_33ns_33_2_1_Adder_10_U.ce ;
wire \sub_33ns_33ns_33_2_1_U14.top_sub_33ns_33ns_33_2_1_Adder_10_U.clk ;
wire \sub_33ns_33ns_33_2_1_U14.top_sub_33ns_33ns_33_2_1_Adder_10_U.facout_s1 ;
wire \sub_33ns_33ns_33_2_1_U14.top_sub_33ns_33ns_33_2_1_Adder_10_U.facout_s2 ;
wire [15:0] \sub_33ns_33ns_33_2_1_U14.top_sub_33ns_33ns_33_2_1_Adder_10_U.fas_s1 ;
wire [16:0] \sub_33ns_33ns_33_2_1_U14.top_sub_33ns_33ns_33_2_1_Adder_10_U.fas_s2 ;
wire \sub_33ns_33ns_33_2_1_U14.top_sub_33ns_33ns_33_2_1_Adder_10_U.reset ;
wire [32:0] \sub_33ns_33ns_33_2_1_U14.top_sub_33ns_33ns_33_2_1_Adder_10_U.s ;
wire [15:0] \sub_33ns_33ns_33_2_1_U14.top_sub_33ns_33ns_33_2_1_Adder_10_U.u1.a ;
wire [15:0] \sub_33ns_33ns_33_2_1_U14.top_sub_33ns_33ns_33_2_1_Adder_10_U.u1.b ;
wire \sub_33ns_33ns_33_2_1_U14.top_sub_33ns_33ns_33_2_1_Adder_10_U.u1.cin ;
wire \sub_33ns_33ns_33_2_1_U14.top_sub_33ns_33ns_33_2_1_Adder_10_U.u1.cout ;
wire [15:0] \sub_33ns_33ns_33_2_1_U14.top_sub_33ns_33ns_33_2_1_Adder_10_U.u1.s ;
wire [16:0] \sub_33ns_33ns_33_2_1_U14.top_sub_33ns_33ns_33_2_1_Adder_10_U.u2.a ;
wire [16:0] \sub_33ns_33ns_33_2_1_U14.top_sub_33ns_33ns_33_2_1_Adder_10_U.u2.b ;
wire \sub_33ns_33ns_33_2_1_U14.top_sub_33ns_33ns_33_2_1_Adder_10_U.u2.cin ;
wire \sub_33ns_33ns_33_2_1_U14.top_sub_33ns_33ns_33_2_1_Adder_10_U.u2.cout ;
wire [16:0] \sub_33ns_33ns_33_2_1_U14.top_sub_33ns_33ns_33_2_1_Adder_10_U.u2.s ;
wire \sub_8ns_8ns_8_2_1_U15.ce ;
wire \sub_8ns_8ns_8_2_1_U15.clk ;
wire [7:0] \sub_8ns_8ns_8_2_1_U15.din0 ;
wire [7:0] \sub_8ns_8ns_8_2_1_U15.din1 ;
wire [7:0] \sub_8ns_8ns_8_2_1_U15.dout ;
wire \sub_8ns_8ns_8_2_1_U15.reset ;
wire [7:0] \sub_8ns_8ns_8_2_1_U15.top_sub_8ns_8ns_8_2_1_Adder_11_U.a ;
wire [7:0] \sub_8ns_8ns_8_2_1_U15.top_sub_8ns_8ns_8_2_1_Adder_11_U.ain_s0 ;
wire [7:0] \sub_8ns_8ns_8_2_1_U15.top_sub_8ns_8ns_8_2_1_Adder_11_U.b ;
wire [7:0] \sub_8ns_8ns_8_2_1_U15.top_sub_8ns_8ns_8_2_1_Adder_11_U.bin_s0 ;
wire \sub_8ns_8ns_8_2_1_U15.top_sub_8ns_8ns_8_2_1_Adder_11_U.ce ;
wire \sub_8ns_8ns_8_2_1_U15.top_sub_8ns_8ns_8_2_1_Adder_11_U.clk ;
wire \sub_8ns_8ns_8_2_1_U15.top_sub_8ns_8ns_8_2_1_Adder_11_U.facout_s1 ;
wire \sub_8ns_8ns_8_2_1_U15.top_sub_8ns_8ns_8_2_1_Adder_11_U.facout_s2 ;
wire [3:0] \sub_8ns_8ns_8_2_1_U15.top_sub_8ns_8ns_8_2_1_Adder_11_U.fas_s1 ;
wire [3:0] \sub_8ns_8ns_8_2_1_U15.top_sub_8ns_8ns_8_2_1_Adder_11_U.fas_s2 ;
wire \sub_8ns_8ns_8_2_1_U15.top_sub_8ns_8ns_8_2_1_Adder_11_U.reset ;
wire [7:0] \sub_8ns_8ns_8_2_1_U15.top_sub_8ns_8ns_8_2_1_Adder_11_U.s ;
wire [3:0] \sub_8ns_8ns_8_2_1_U15.top_sub_8ns_8ns_8_2_1_Adder_11_U.u1.a ;
wire [3:0] \sub_8ns_8ns_8_2_1_U15.top_sub_8ns_8ns_8_2_1_Adder_11_U.u1.b ;
wire \sub_8ns_8ns_8_2_1_U15.top_sub_8ns_8ns_8_2_1_Adder_11_U.u1.cin ;
wire \sub_8ns_8ns_8_2_1_U15.top_sub_8ns_8ns_8_2_1_Adder_11_U.u1.cout ;
wire [3:0] \sub_8ns_8ns_8_2_1_U15.top_sub_8ns_8ns_8_2_1_Adder_11_U.u1.s ;
wire [3:0] \sub_8ns_8ns_8_2_1_U15.top_sub_8ns_8ns_8_2_1_Adder_11_U.u2.a ;
wire [3:0] \sub_8ns_8ns_8_2_1_U15.top_sub_8ns_8ns_8_2_1_Adder_11_U.u2.b ;
wire \sub_8ns_8ns_8_2_1_U15.top_sub_8ns_8ns_8_2_1_Adder_11_U.u2.cin ;
wire \sub_8ns_8ns_8_2_1_U15.top_sub_8ns_8ns_8_2_1_Adder_11_U.u2.cout ;
wire [3:0] \sub_8ns_8ns_8_2_1_U15.top_sub_8ns_8ns_8_2_1_Adder_11_U.u2.s ;
wire \sub_8s_8ns_8_2_1_U7.ce ;
wire \sub_8s_8ns_8_2_1_U7.clk ;
wire [7:0] \sub_8s_8ns_8_2_1_U7.din0 ;
wire [7:0] \sub_8s_8ns_8_2_1_U7.din1 ;
wire [7:0] \sub_8s_8ns_8_2_1_U7.dout ;
wire \sub_8s_8ns_8_2_1_U7.reset ;
wire [7:0] \sub_8s_8ns_8_2_1_U7.top_sub_8s_8ns_8_2_1_Adder_4_U.a ;
wire [7:0] \sub_8s_8ns_8_2_1_U7.top_sub_8s_8ns_8_2_1_Adder_4_U.ain_s0 ;
wire [7:0] \sub_8s_8ns_8_2_1_U7.top_sub_8s_8ns_8_2_1_Adder_4_U.b ;
wire [7:0] \sub_8s_8ns_8_2_1_U7.top_sub_8s_8ns_8_2_1_Adder_4_U.bin_s0 ;
wire \sub_8s_8ns_8_2_1_U7.top_sub_8s_8ns_8_2_1_Adder_4_U.ce ;
wire \sub_8s_8ns_8_2_1_U7.top_sub_8s_8ns_8_2_1_Adder_4_U.clk ;
wire \sub_8s_8ns_8_2_1_U7.top_sub_8s_8ns_8_2_1_Adder_4_U.facout_s1 ;
wire \sub_8s_8ns_8_2_1_U7.top_sub_8s_8ns_8_2_1_Adder_4_U.facout_s2 ;
wire [3:0] \sub_8s_8ns_8_2_1_U7.top_sub_8s_8ns_8_2_1_Adder_4_U.fas_s1 ;
wire [3:0] \sub_8s_8ns_8_2_1_U7.top_sub_8s_8ns_8_2_1_Adder_4_U.fas_s2 ;
wire \sub_8s_8ns_8_2_1_U7.top_sub_8s_8ns_8_2_1_Adder_4_U.reset ;
wire [7:0] \sub_8s_8ns_8_2_1_U7.top_sub_8s_8ns_8_2_1_Adder_4_U.s ;
wire [3:0] \sub_8s_8ns_8_2_1_U7.top_sub_8s_8ns_8_2_1_Adder_4_U.u1.a ;
wire [3:0] \sub_8s_8ns_8_2_1_U7.top_sub_8s_8ns_8_2_1_Adder_4_U.u1.b ;
wire \sub_8s_8ns_8_2_1_U7.top_sub_8s_8ns_8_2_1_Adder_4_U.u1.cin ;
wire \sub_8s_8ns_8_2_1_U7.top_sub_8s_8ns_8_2_1_Adder_4_U.u1.cout ;
wire [3:0] \sub_8s_8ns_8_2_1_U7.top_sub_8s_8ns_8_2_1_Adder_4_U.u1.s ;
wire [3:0] \sub_8s_8ns_8_2_1_U7.top_sub_8s_8ns_8_2_1_Adder_4_U.u2.a ;
wire [3:0] \sub_8s_8ns_8_2_1_U7.top_sub_8s_8ns_8_2_1_Adder_4_U.u2.b ;
wire \sub_8s_8ns_8_2_1_U7.top_sub_8s_8ns_8_2_1_Adder_4_U.u2.cin ;
wire \sub_8s_8ns_8_2_1_U7.top_sub_8s_8ns_8_2_1_Adder_4_U.u2.cout ;
wire [3:0] \sub_8s_8ns_8_2_1_U7.top_sub_8s_8ns_8_2_1_Adder_4_U.u2.s ;
wire tmp_13_fu_959_p3;
wire tmp_23_fu_1334_p3;
wire tmp_24_fu_1341_p3;
wire [13:0] tmp_26_fu_1499_p3;
wire tmp_6_fu_526_p3;
wire tmp_7_fu_533_p3;
wire [2:0] trunc_ln1192_fu_285_p1;
wire [7:0] trunc_ln213_fu_731_p1;
wire [13:0] trunc_ln731_1_fu_912_p1;
wire [5:0] trunc_ln731_2_fu_1006_p1;
wire trunc_ln731_fu_298_p1;
wire [7:0] trunc_ln851_1_fu_826_p0;
wire [2:0] trunc_ln851_1_fu_826_p1;
wire trunc_ln851_2_fu_1480_p1;
wire [15:0] trunc_ln851_3_fu_1187_p0;
wire [12:0] trunc_ln851_3_fu_1187_p1;
wire [1:0] trunc_ln851_4_fu_1469_p1;
wire [1:0] trunc_ln851_5_fu_1297_p1;
wire trunc_ln851_6_fu_1672_p1;
wire [2:0] trunc_ln851_fu_724_p1;
wire xor_ln340_1_fu_567_p2;
wire xor_ln340_2_fu_1146_p2;
wire xor_ln340_3_fu_1376_p2;
wire xor_ln340_fu_326_p2;
wire xor_ln365_1_fu_546_p2;
wire xor_ln365_2_fu_1348_p2;
wire xor_ln365_3_fu_1354_p2;
wire xor_ln365_fu_540_p2;
wire xor_ln416_fu_836_p2;
wire xor_ln780_fu_966_p2;
wire xor_ln781_fu_1091_p2;
wire xor_ln785_1_fu_485_p2;
wire xor_ln785_2_fu_1028_p2;
wire xor_ln785_3_fu_1038_p2;
wire xor_ln785_4_fu_1121_p2;
wire xor_ln785_5_fu_1201_p2;
wire xor_ln785_6_fu_362_p2;
wire xor_ln785_7_fu_604_p2;
wire xor_ln785_8_fu_1231_p2;
wire xor_ln785_9_fu_1424_p2;
wire xor_ln785_fu_301_p2;
wire xor_ln786_1_fu_494_p2;
wire xor_ln786_2_fu_1131_p2;
wire xor_ln786_3_fu_1272_p2;
wire xor_ln786_4_fu_357_p2;
wire xor_ln786_5_fu_509_p2;
wire xor_ln786_6_fu_1226_p2;
wire xor_ln786_7_fu_1287_p2;
wire xor_ln786_fu_311_p2;
wire [35:0] zext_ln1116_fu_633_p1;
wire [7:0] zext_ln1499_fu_864_p1;


assign _0124_ = icmp_ln851_2_reg_2305 & ap_CS_fsm[29];
assign _0125_ = icmp_ln851_3_reg_2452 & ap_CS_fsm[34];
assign _0126_ = icmp_ln851_4_reg_2402 & ap_CS_fsm[39];
assign _0127_ = _0132_ & ap_CS_fsm[24];
assign _0128_ = _0133_ & ap_CS_fsm[29];
assign _0129_ = ap_CS_fsm[10] & _0134_;
assign _0130_ = _0135_ & ap_CS_fsm[0];
assign _0131_ = ap_start & ap_CS_fsm[0];
assign and_ln340_1_fu_572_p2 = xor_ln340_1_fu_567_p2 & or_ln786_1_reg_1884;
assign and_ln340_2_fu_584_p2 = or_ln786_1_reg_1884 & or_ln340_1_reg_1890;
assign and_ln340_3_fu_1152_p2 = xor_ln340_2_fu_1146_p2 & or_ln786_2_fu_1136_p2;
assign and_ln340_4_fu_1381_p2 = xor_ln340_3_fu_1376_p2 & or_ln786_3_reg_2343;
assign and_ln340_5_fu_1394_p2 = or_ln786_3_reg_2343 & or_ln340_4_reg_2349;
assign and_ln340_fu_332_p2 = xor_ln340_fu_326_p2 & or_ln786_fu_316_p2;
assign and_ln412_fu_741_p2 = p_Result_31_reg_1949 & p_Result_11_reg_1966;
assign and_ln780_fu_972_p2 = xor_ln780_fu_966_p2 & Range2_all_ones_reg_2025;
assign and_ln781_fu_1087_p2 = carry_1_reg_2141 & Range1_all_ones_reg_2030;
assign and_ln785_10_fu_1247_p2 = p_Result_35_reg_2160 & and_ln785_9_fu_1241_p2;
assign and_ln785_12_fu_1434_p2 = or_ln785_10_fu_1429_p2 & and_ln786_2_reg_2355;
assign and_ln785_13_fu_1398_p2 = xor_ln785_5_reg_2316 & and_ln786_2_reg_2355;
assign and_ln785_1_fu_378_p2 = p_Result_26_reg_1736 & and_ln785_fu_372_p2;
assign and_ln785_3_fu_614_p2 = or_ln785_6_fu_609_p2 & and_ln786_1_reg_1896;
assign and_ln785_4_fu_588_p2 = xor_ln785_1_reg_1878 & and_ln786_1_reg_1896;
assign and_ln785_6_fu_1206_p2 = xor_ln416_reg_2097 & deleted_zeros_reg_2188;
assign and_ln785_7_fu_1215_p2 = or_ln785_8_fu_1210_p2 & and_ln786_reg_2194;
assign and_ln785_9_fu_1241_p2 = xor_ln786_6_fu_1226_p2 & or_ln785_9_fu_1236_p2;
assign and_ln785_fu_372_p2 = xor_ln786_4_fu_357_p2 & or_ln785_5_fu_367_p2;
assign and_ln786_1_fu_514_p2 = xor_ln786_5_fu_509_p2 & p_Result_28_reg_1848;
assign and_ln786_2_fu_1292_p2 = xor_ln786_7_fu_1287_p2 & p_Result_37_reg_2235;
assign and_ln786_fu_983_p2 = p_Result_33_reg_2068 & deleted_ones_fu_977_p3;
assign carry_1_fu_895_p2 = xor_ln416_reg_2097 & p_Result_32_reg_1971;
assign neg_src_fu_1097_p2 = xor_ln781_fu_1091_p2 & p_Result_30_reg_1954;
assign overflow_1_fu_490_p2 = xor_ln785_1_reg_1878 & or_ln785_1_reg_1872;
assign overflow_2_fu_1043_p2 = xor_ln785_3_fu_1038_p2 & or_ln785_2_fu_1033_p2;
assign overflow_3_fu_1126_p2 = xor_ln785_4_fu_1121_p2 & or_ln785_3_reg_2258;
assign overflow_4_fu_1268_p2 = xor_ln785_5_reg_2316 & or_ln785_4_reg_2310;
assign overflow_fu_306_p2 = xor_ln785_fu_301_p2 & or_ln785_reg_1761;
assign sel_tmp19_fu_598_p2 = xor_ln365_1_fu_546_p2 & or_ln785_7_fu_592_p2;
assign sel_tmp51_fu_1408_p2 = xor_ln365_3_fu_1354_p2 & or_ln785_11_fu_1402_p2;
assign xor_ln340_1_fu_567_p2 = ~ or_ln340_1_reg_1890;
assign xor_ln786_2_fu_1131_p2 = ~ p_Result_35_reg_2160;
assign xor_ln785_4_fu_1121_p2 = ~ p_Result_34_reg_2148;
assign xor_ln340_2_fu_1146_p2 = ~ or_ln340_3_fu_1141_p2;
assign xor_ln340_3_fu_1376_p2 = ~ or_ln340_4_reg_2349;
assign xor_ln786_fu_311_p2 = ~ p_Result_26_reg_1736;
assign xor_ln785_fu_301_p2 = ~ p_Result_s_reg_1722;
assign xor_ln340_fu_326_p2 = ~ or_ln340_fu_321_p2;
assign xor_ln780_fu_966_p2 = ~ r_V_5_reg_1944[3];
assign xor_ln785_8_fu_1231_p2 = ~ or_ln785_3_reg_2258;
assign xor_ln786_6_fu_1226_p2 = ~ icmp_ln786_2_reg_2210;
assign xor_ln785_9_fu_1424_p2 = ~ or_ln785_4_reg_2310;
assign xor_ln785_6_fu_362_p2 = ~ or_ln785_reg_1761;
assign xor_ln786_4_fu_357_p2 = ~ icmp_ln786_reg_1767;
assign xor_ln785_7_fu_604_p2 = ~ or_ln785_1_reg_1872;
assign xor_ln786_5_fu_509_p2 = ~ icmp_ln786_1_reg_1866;
assign xor_ln786_7_fu_1287_p2 = ~ icmp_ln786_3_reg_2274;
assign xor_ln781_fu_1091_p2 = ~ and_ln781_fu_1087_p2;
assign xor_ln785_2_fu_1028_p2 = ~ deleted_zeros_reg_2188;
assign xor_ln785_3_fu_1038_p2 = ~ p_Result_30_reg_1954;
assign xor_ln786_1_fu_494_p2 = ~ p_Result_28_reg_1848;
assign xor_ln786_3_fu_1272_p2 = ~ p_Result_37_reg_2235;
assign xor_ln365_1_fu_546_p2 = ~ xor_ln365_fu_540_p2;
assign xor_ln365_3_fu_1354_p2 = ~ xor_ln365_2_fu_1348_p2;
assign xor_ln416_fu_836_p2 = ~ p_Result_33_reg_2068;
assign xor_ln785_1_fu_485_p2 = ~ p_Result_27_reg_1832;
assign xor_ln785_5_fu_1201_p2 = ~ p_Result_36_reg_2223;
assign p_Val2_15_fu_1360_p2 = ~ { trunc_ln731_2_reg_2230[4:0], 2'h0 };
assign p_Val2_3_fu_552_p2 = ~ p_Val2_2_reg_1839[2:0];
assign _0132_ = ~ icmp_ln851_1_reg_2092;
assign _0133_ = ~ sel_tmp51_reg_2397;
assign _0134_ = ~ sel_tmp19_reg_1907;
assign _0135_ = ~ ap_start;
assign _0136_ = p_Result_3_reg_1981 == 33'h1ffffffff;
assign _0137_ = ! p_Result_3_reg_1981;
assign _0138_ = p_Result_1_reg_1976 == 32'd4294967295;
assign _0139_ = ! op_6[2:0];
always @(posedge \add_10ns_10ns_10_2_1_U13.top_add_10ns_10ns_10_2_1_Adder_9_U.clk )
\add_10ns_10ns_10_2_1_U13.top_add_10ns_10ns_10_2_1_Adder_9_U.bin_s1  <= _0141_;
always @(posedge \add_10ns_10ns_10_2_1_U13.top_add_10ns_10ns_10_2_1_Adder_9_U.clk )
\add_10ns_10ns_10_2_1_U13.top_add_10ns_10ns_10_2_1_Adder_9_U.ain_s1  <= _0140_;
always @(posedge \add_10ns_10ns_10_2_1_U13.top_add_10ns_10ns_10_2_1_Adder_9_U.clk )
\add_10ns_10ns_10_2_1_U13.top_add_10ns_10ns_10_2_1_Adder_9_U.sum_s1  <= _0143_;
always @(posedge \add_10ns_10ns_10_2_1_U13.top_add_10ns_10ns_10_2_1_Adder_9_U.clk )
\add_10ns_10ns_10_2_1_U13.top_add_10ns_10ns_10_2_1_Adder_9_U.carry_s1  <= _0142_;
assign _0141_ = \add_10ns_10ns_10_2_1_U13.top_add_10ns_10ns_10_2_1_Adder_9_U.ce  ? \add_10ns_10ns_10_2_1_U13.top_add_10ns_10ns_10_2_1_Adder_9_U.b [9:5] : \add_10ns_10ns_10_2_1_U13.top_add_10ns_10ns_10_2_1_Adder_9_U.bin_s1 ;
assign _0140_ = \add_10ns_10ns_10_2_1_U13.top_add_10ns_10ns_10_2_1_Adder_9_U.ce  ? \add_10ns_10ns_10_2_1_U13.top_add_10ns_10ns_10_2_1_Adder_9_U.a [9:5] : \add_10ns_10ns_10_2_1_U13.top_add_10ns_10ns_10_2_1_Adder_9_U.ain_s1 ;
assign _0142_ = \add_10ns_10ns_10_2_1_U13.top_add_10ns_10ns_10_2_1_Adder_9_U.ce  ? \add_10ns_10ns_10_2_1_U13.top_add_10ns_10ns_10_2_1_Adder_9_U.facout_s1  : \add_10ns_10ns_10_2_1_U13.top_add_10ns_10ns_10_2_1_Adder_9_U.carry_s1 ;
assign _0143_ = \add_10ns_10ns_10_2_1_U13.top_add_10ns_10ns_10_2_1_Adder_9_U.ce  ? \add_10ns_10ns_10_2_1_U13.top_add_10ns_10ns_10_2_1_Adder_9_U.fas_s1  : \add_10ns_10ns_10_2_1_U13.top_add_10ns_10ns_10_2_1_Adder_9_U.sum_s1 ;
assign _0144_ = \add_10ns_10ns_10_2_1_U13.top_add_10ns_10ns_10_2_1_Adder_9_U.u1.a  + \add_10ns_10ns_10_2_1_U13.top_add_10ns_10ns_10_2_1_Adder_9_U.u1.b ;
assign { \add_10ns_10ns_10_2_1_U13.top_add_10ns_10ns_10_2_1_Adder_9_U.u1.cout , \add_10ns_10ns_10_2_1_U13.top_add_10ns_10ns_10_2_1_Adder_9_U.u1.s  } = _0144_ + \add_10ns_10ns_10_2_1_U13.top_add_10ns_10ns_10_2_1_Adder_9_U.u1.cin ;
assign _0145_ = \add_10ns_10ns_10_2_1_U13.top_add_10ns_10ns_10_2_1_Adder_9_U.u2.a  + \add_10ns_10ns_10_2_1_U13.top_add_10ns_10ns_10_2_1_Adder_9_U.u2.b ;
assign { \add_10ns_10ns_10_2_1_U13.top_add_10ns_10ns_10_2_1_Adder_9_U.u2.cout , \add_10ns_10ns_10_2_1_U13.top_add_10ns_10ns_10_2_1_Adder_9_U.u2.s  } = _0145_ + \add_10ns_10ns_10_2_1_U13.top_add_10ns_10ns_10_2_1_Adder_9_U.u2.cin ;
always @(posedge \add_12s_12ns_12_2_1_U17.top_add_12s_12ns_12_2_1_Adder_13_U.clk )
\add_12s_12ns_12_2_1_U17.top_add_12s_12ns_12_2_1_Adder_13_U.bin_s1  <= _0147_;
always @(posedge \add_12s_12ns_12_2_1_U17.top_add_12s_12ns_12_2_1_Adder_13_U.clk )
\add_12s_12ns_12_2_1_U17.top_add_12s_12ns_12_2_1_Adder_13_U.ain_s1  <= _0146_;
always @(posedge \add_12s_12ns_12_2_1_U17.top_add_12s_12ns_12_2_1_Adder_13_U.clk )
\add_12s_12ns_12_2_1_U17.top_add_12s_12ns_12_2_1_Adder_13_U.sum_s1  <= _0149_;
always @(posedge \add_12s_12ns_12_2_1_U17.top_add_12s_12ns_12_2_1_Adder_13_U.clk )
\add_12s_12ns_12_2_1_U17.top_add_12s_12ns_12_2_1_Adder_13_U.carry_s1  <= _0148_;
assign _0147_ = \add_12s_12ns_12_2_1_U17.top_add_12s_12ns_12_2_1_Adder_13_U.ce  ? \add_12s_12ns_12_2_1_U17.top_add_12s_12ns_12_2_1_Adder_13_U.b [11:6] : \add_12s_12ns_12_2_1_U17.top_add_12s_12ns_12_2_1_Adder_13_U.bin_s1 ;
assign _0146_ = \add_12s_12ns_12_2_1_U17.top_add_12s_12ns_12_2_1_Adder_13_U.ce  ? \add_12s_12ns_12_2_1_U17.top_add_12s_12ns_12_2_1_Adder_13_U.a [11:6] : \add_12s_12ns_12_2_1_U17.top_add_12s_12ns_12_2_1_Adder_13_U.ain_s1 ;
assign _0148_ = \add_12s_12ns_12_2_1_U17.top_add_12s_12ns_12_2_1_Adder_13_U.ce  ? \add_12s_12ns_12_2_1_U17.top_add_12s_12ns_12_2_1_Adder_13_U.facout_s1  : \add_12s_12ns_12_2_1_U17.top_add_12s_12ns_12_2_1_Adder_13_U.carry_s1 ;
assign _0149_ = \add_12s_12ns_12_2_1_U17.top_add_12s_12ns_12_2_1_Adder_13_U.ce  ? \add_12s_12ns_12_2_1_U17.top_add_12s_12ns_12_2_1_Adder_13_U.fas_s1  : \add_12s_12ns_12_2_1_U17.top_add_12s_12ns_12_2_1_Adder_13_U.sum_s1 ;
assign _0150_ = \add_12s_12ns_12_2_1_U17.top_add_12s_12ns_12_2_1_Adder_13_U.u1.a  + \add_12s_12ns_12_2_1_U17.top_add_12s_12ns_12_2_1_Adder_13_U.u1.b ;
assign { \add_12s_12ns_12_2_1_U17.top_add_12s_12ns_12_2_1_Adder_13_U.u1.cout , \add_12s_12ns_12_2_1_U17.top_add_12s_12ns_12_2_1_Adder_13_U.u1.s  } = _0150_ + \add_12s_12ns_12_2_1_U17.top_add_12s_12ns_12_2_1_Adder_13_U.u1.cin ;
assign _0151_ = \add_12s_12ns_12_2_1_U17.top_add_12s_12ns_12_2_1_Adder_13_U.u2.a  + \add_12s_12ns_12_2_1_U17.top_add_12s_12ns_12_2_1_Adder_13_U.u2.b ;
assign { \add_12s_12ns_12_2_1_U17.top_add_12s_12ns_12_2_1_Adder_13_U.u2.cout , \add_12s_12ns_12_2_1_U17.top_add_12s_12ns_12_2_1_Adder_13_U.u2.s  } = _0151_ + \add_12s_12ns_12_2_1_U17.top_add_12s_12ns_12_2_1_Adder_13_U.u2.cin ;
always @(posedge \add_13ns_13s_13_2_1_U10.top_add_13ns_13s_13_2_1_Adder_7_U.clk )
\add_13ns_13s_13_2_1_U10.top_add_13ns_13s_13_2_1_Adder_7_U.bin_s1  <= _0153_;
always @(posedge \add_13ns_13s_13_2_1_U10.top_add_13ns_13s_13_2_1_Adder_7_U.clk )
\add_13ns_13s_13_2_1_U10.top_add_13ns_13s_13_2_1_Adder_7_U.ain_s1  <= _0152_;
always @(posedge \add_13ns_13s_13_2_1_U10.top_add_13ns_13s_13_2_1_Adder_7_U.clk )
\add_13ns_13s_13_2_1_U10.top_add_13ns_13s_13_2_1_Adder_7_U.sum_s1  <= _0155_;
always @(posedge \add_13ns_13s_13_2_1_U10.top_add_13ns_13s_13_2_1_Adder_7_U.clk )
\add_13ns_13s_13_2_1_U10.top_add_13ns_13s_13_2_1_Adder_7_U.carry_s1  <= _0154_;
assign _0153_ = \add_13ns_13s_13_2_1_U10.top_add_13ns_13s_13_2_1_Adder_7_U.ce  ? \add_13ns_13s_13_2_1_U10.top_add_13ns_13s_13_2_1_Adder_7_U.b [12:6] : \add_13ns_13s_13_2_1_U10.top_add_13ns_13s_13_2_1_Adder_7_U.bin_s1 ;
assign _0152_ = \add_13ns_13s_13_2_1_U10.top_add_13ns_13s_13_2_1_Adder_7_U.ce  ? \add_13ns_13s_13_2_1_U10.top_add_13ns_13s_13_2_1_Adder_7_U.a [12:6] : \add_13ns_13s_13_2_1_U10.top_add_13ns_13s_13_2_1_Adder_7_U.ain_s1 ;
assign _0154_ = \add_13ns_13s_13_2_1_U10.top_add_13ns_13s_13_2_1_Adder_7_U.ce  ? \add_13ns_13s_13_2_1_U10.top_add_13ns_13s_13_2_1_Adder_7_U.facout_s1  : \add_13ns_13s_13_2_1_U10.top_add_13ns_13s_13_2_1_Adder_7_U.carry_s1 ;
assign _0155_ = \add_13ns_13s_13_2_1_U10.top_add_13ns_13s_13_2_1_Adder_7_U.ce  ? \add_13ns_13s_13_2_1_U10.top_add_13ns_13s_13_2_1_Adder_7_U.fas_s1  : \add_13ns_13s_13_2_1_U10.top_add_13ns_13s_13_2_1_Adder_7_U.sum_s1 ;
assign _0156_ = \add_13ns_13s_13_2_1_U10.top_add_13ns_13s_13_2_1_Adder_7_U.u1.a  + \add_13ns_13s_13_2_1_U10.top_add_13ns_13s_13_2_1_Adder_7_U.u1.b ;
assign { \add_13ns_13s_13_2_1_U10.top_add_13ns_13s_13_2_1_Adder_7_U.u1.cout , \add_13ns_13s_13_2_1_U10.top_add_13ns_13s_13_2_1_Adder_7_U.u1.s  } = _0156_ + \add_13ns_13s_13_2_1_U10.top_add_13ns_13s_13_2_1_Adder_7_U.u1.cin ;
assign _0157_ = \add_13ns_13s_13_2_1_U10.top_add_13ns_13s_13_2_1_Adder_7_U.u2.a  + \add_13ns_13s_13_2_1_U10.top_add_13ns_13s_13_2_1_Adder_7_U.u2.b ;
assign { \add_13ns_13s_13_2_1_U10.top_add_13ns_13s_13_2_1_Adder_7_U.u2.cout , \add_13ns_13s_13_2_1_U10.top_add_13ns_13s_13_2_1_Adder_7_U.u2.s  } = _0157_ + \add_13ns_13s_13_2_1_U10.top_add_13ns_13s_13_2_1_Adder_7_U.u2.cin ;
always @(posedge \add_17s_17s_17_2_1_U28.top_add_17s_17s_17_2_1_Adder_18_U.clk )
\add_17s_17s_17_2_1_U28.top_add_17s_17s_17_2_1_Adder_18_U.bin_s1  <= _0159_;
always @(posedge \add_17s_17s_17_2_1_U28.top_add_17s_17s_17_2_1_Adder_18_U.clk )
\add_17s_17s_17_2_1_U28.top_add_17s_17s_17_2_1_Adder_18_U.ain_s1  <= _0158_;
always @(posedge \add_17s_17s_17_2_1_U28.top_add_17s_17s_17_2_1_Adder_18_U.clk )
\add_17s_17s_17_2_1_U28.top_add_17s_17s_17_2_1_Adder_18_U.sum_s1  <= _0161_;
always @(posedge \add_17s_17s_17_2_1_U28.top_add_17s_17s_17_2_1_Adder_18_U.clk )
\add_17s_17s_17_2_1_U28.top_add_17s_17s_17_2_1_Adder_18_U.carry_s1  <= _0160_;
assign _0159_ = \add_17s_17s_17_2_1_U28.top_add_17s_17s_17_2_1_Adder_18_U.ce  ? \add_17s_17s_17_2_1_U28.top_add_17s_17s_17_2_1_Adder_18_U.b [16:8] : \add_17s_17s_17_2_1_U28.top_add_17s_17s_17_2_1_Adder_18_U.bin_s1 ;
assign _0158_ = \add_17s_17s_17_2_1_U28.top_add_17s_17s_17_2_1_Adder_18_U.ce  ? \add_17s_17s_17_2_1_U28.top_add_17s_17s_17_2_1_Adder_18_U.a [16:8] : \add_17s_17s_17_2_1_U28.top_add_17s_17s_17_2_1_Adder_18_U.ain_s1 ;
assign _0160_ = \add_17s_17s_17_2_1_U28.top_add_17s_17s_17_2_1_Adder_18_U.ce  ? \add_17s_17s_17_2_1_U28.top_add_17s_17s_17_2_1_Adder_18_U.facout_s1  : \add_17s_17s_17_2_1_U28.top_add_17s_17s_17_2_1_Adder_18_U.carry_s1 ;
assign _0161_ = \add_17s_17s_17_2_1_U28.top_add_17s_17s_17_2_1_Adder_18_U.ce  ? \add_17s_17s_17_2_1_U28.top_add_17s_17s_17_2_1_Adder_18_U.fas_s1  : \add_17s_17s_17_2_1_U28.top_add_17s_17s_17_2_1_Adder_18_U.sum_s1 ;
assign _0162_ = \add_17s_17s_17_2_1_U28.top_add_17s_17s_17_2_1_Adder_18_U.u1.a  + \add_17s_17s_17_2_1_U28.top_add_17s_17s_17_2_1_Adder_18_U.u1.b ;
assign { \add_17s_17s_17_2_1_U28.top_add_17s_17s_17_2_1_Adder_18_U.u1.cout , \add_17s_17s_17_2_1_U28.top_add_17s_17s_17_2_1_Adder_18_U.u1.s  } = _0162_ + \add_17s_17s_17_2_1_U28.top_add_17s_17s_17_2_1_Adder_18_U.u1.cin ;
assign _0163_ = \add_17s_17s_17_2_1_U28.top_add_17s_17s_17_2_1_Adder_18_U.u2.a  + \add_17s_17s_17_2_1_U28.top_add_17s_17s_17_2_1_Adder_18_U.u2.b ;
assign { \add_17s_17s_17_2_1_U28.top_add_17s_17s_17_2_1_Adder_18_U.u2.cout , \add_17s_17s_17_2_1_U28.top_add_17s_17s_17_2_1_Adder_18_U.u2.s  } = _0163_ + \add_17s_17s_17_2_1_U28.top_add_17s_17s_17_2_1_Adder_18_U.u2.cin ;
always @(posedge \add_24s_24s_24_2_1_U16.top_add_24s_24s_24_2_1_Adder_12_U.clk )
\add_24s_24s_24_2_1_U16.top_add_24s_24s_24_2_1_Adder_12_U.bin_s1  <= _0165_;
always @(posedge \add_24s_24s_24_2_1_U16.top_add_24s_24s_24_2_1_Adder_12_U.clk )
\add_24s_24s_24_2_1_U16.top_add_24s_24s_24_2_1_Adder_12_U.ain_s1  <= _0164_;
always @(posedge \add_24s_24s_24_2_1_U16.top_add_24s_24s_24_2_1_Adder_12_U.clk )
\add_24s_24s_24_2_1_U16.top_add_24s_24s_24_2_1_Adder_12_U.sum_s1  <= _0167_;
always @(posedge \add_24s_24s_24_2_1_U16.top_add_24s_24s_24_2_1_Adder_12_U.clk )
\add_24s_24s_24_2_1_U16.top_add_24s_24s_24_2_1_Adder_12_U.carry_s1  <= _0166_;
assign _0165_ = \add_24s_24s_24_2_1_U16.top_add_24s_24s_24_2_1_Adder_12_U.ce  ? \add_24s_24s_24_2_1_U16.top_add_24s_24s_24_2_1_Adder_12_U.b [23:12] : \add_24s_24s_24_2_1_U16.top_add_24s_24s_24_2_1_Adder_12_U.bin_s1 ;
assign _0164_ = \add_24s_24s_24_2_1_U16.top_add_24s_24s_24_2_1_Adder_12_U.ce  ? \add_24s_24s_24_2_1_U16.top_add_24s_24s_24_2_1_Adder_12_U.a [23:12] : \add_24s_24s_24_2_1_U16.top_add_24s_24s_24_2_1_Adder_12_U.ain_s1 ;
assign _0166_ = \add_24s_24s_24_2_1_U16.top_add_24s_24s_24_2_1_Adder_12_U.ce  ? \add_24s_24s_24_2_1_U16.top_add_24s_24s_24_2_1_Adder_12_U.facout_s1  : \add_24s_24s_24_2_1_U16.top_add_24s_24s_24_2_1_Adder_12_U.carry_s1 ;
assign _0167_ = \add_24s_24s_24_2_1_U16.top_add_24s_24s_24_2_1_Adder_12_U.ce  ? \add_24s_24s_24_2_1_U16.top_add_24s_24s_24_2_1_Adder_12_U.fas_s1  : \add_24s_24s_24_2_1_U16.top_add_24s_24s_24_2_1_Adder_12_U.sum_s1 ;
assign _0168_ = \add_24s_24s_24_2_1_U16.top_add_24s_24s_24_2_1_Adder_12_U.u1.a  + \add_24s_24s_24_2_1_U16.top_add_24s_24s_24_2_1_Adder_12_U.u1.b ;
assign { \add_24s_24s_24_2_1_U16.top_add_24s_24s_24_2_1_Adder_12_U.u1.cout , \add_24s_24s_24_2_1_U16.top_add_24s_24s_24_2_1_Adder_12_U.u1.s  } = _0168_ + \add_24s_24s_24_2_1_U16.top_add_24s_24s_24_2_1_Adder_12_U.u1.cin ;
assign _0169_ = \add_24s_24s_24_2_1_U16.top_add_24s_24s_24_2_1_Adder_12_U.u2.a  + \add_24s_24s_24_2_1_U16.top_add_24s_24s_24_2_1_Adder_12_U.u2.b ;
assign { \add_24s_24s_24_2_1_U16.top_add_24s_24s_24_2_1_Adder_12_U.u2.cout , \add_24s_24s_24_2_1_U16.top_add_24s_24s_24_2_1_Adder_12_U.u2.s  } = _0169_ + \add_24s_24s_24_2_1_U16.top_add_24s_24s_24_2_1_Adder_12_U.u2.cin ;
always @(posedge \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.clk )
\add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.bin_s1  <= _0171_;
always @(posedge \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.clk )
\add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.ain_s1  <= _0170_;
always @(posedge \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.clk )
\add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.sum_s1  <= _0173_;
always @(posedge \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.clk )
\add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.carry_s1  <= _0172_;
assign _0171_ = \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.ce  ? \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.b [1] : \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.bin_s1 ;
assign _0170_ = \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.ce  ? \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.a [1] : \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.ain_s1 ;
assign _0172_ = \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.ce  ? \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.facout_s1  : \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.carry_s1 ;
assign _0173_ = \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.ce  ? \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.fas_s1  : \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.sum_s1 ;
assign _0174_ = \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.u1.a  + \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.u1.b ;
assign { \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.u1.cout , \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.u1.s  } = _0174_ + \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.u1.cin ;
assign _0175_ = \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.u2.a  + \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.u2.b ;
assign { \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.u2.cout , \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.u2.s  } = _0175_ + \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.u2.cin ;
always @(posedge \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_15_U.clk )
\add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_15_U.bin_s1  <= _0177_;
always @(posedge \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_15_U.clk )
\add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_15_U.ain_s1  <= _0176_;
always @(posedge \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_15_U.clk )
\add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_15_U.sum_s1  <= _0179_;
always @(posedge \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_15_U.clk )
\add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_15_U.carry_s1  <= _0178_;
assign _0177_ = \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_15_U.ce  ? \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_15_U.b [31:16] : \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_15_U.bin_s1 ;
assign _0176_ = \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_15_U.ce  ? \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_15_U.a [31:16] : \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_15_U.ain_s1 ;
assign _0178_ = \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_15_U.ce  ? \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_15_U.facout_s1  : \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_15_U.carry_s1 ;
assign _0179_ = \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_15_U.ce  ? \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_15_U.fas_s1  : \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_15_U.sum_s1 ;
assign _0180_ = \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.a  + \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.b ;
assign { \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.cout , \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.s  } = _0180_ + \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.cin ;
assign _0181_ = \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.a  + \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.b ;
assign { \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.cout , \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.s  } = _0181_ + \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.cin ;
always @(posedge \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_15_U.clk )
\add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_15_U.bin_s1  <= _0183_;
always @(posedge \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_15_U.clk )
\add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_15_U.ain_s1  <= _0182_;
always @(posedge \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_15_U.clk )
\add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_15_U.sum_s1  <= _0185_;
always @(posedge \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_15_U.clk )
\add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_15_U.carry_s1  <= _0184_;
assign _0183_ = \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_15_U.ce  ? \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_15_U.b [31:16] : \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_15_U.bin_s1 ;
assign _0182_ = \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_15_U.ce  ? \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_15_U.a [31:16] : \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_15_U.ain_s1 ;
assign _0184_ = \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_15_U.ce  ? \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_15_U.facout_s1  : \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_15_U.carry_s1 ;
assign _0185_ = \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_15_U.ce  ? \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_15_U.fas_s1  : \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_15_U.sum_s1 ;
assign _0186_ = \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.a  + \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.b ;
assign { \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.cout , \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.s  } = _0186_ + \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.cin ;
assign _0187_ = \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.a  + \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.b ;
assign { \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.cout , \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.s  } = _0187_ + \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.cin ;
always @(posedge \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.clk )
\add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.bin_s1  <= _0189_;
always @(posedge \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.clk )
\add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.ain_s1  <= _0188_;
always @(posedge \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.clk )
\add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.sum_s1  <= _0191_;
always @(posedge \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.clk )
\add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.carry_s1  <= _0190_;
assign _0189_ = \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.ce  ? \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.b [31:16] : \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.bin_s1 ;
assign _0188_ = \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.ce  ? \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.a [31:16] : \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.ain_s1 ;
assign _0190_ = \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.ce  ? \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.facout_s1  : \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.carry_s1 ;
assign _0191_ = \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.ce  ? \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.fas_s1  : \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.sum_s1 ;
assign _0192_ = \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.a  + \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.b ;
assign { \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.cout , \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.s  } = _0192_ + \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.cin ;
assign _0193_ = \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.a  + \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.b ;
assign { \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.cout , \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.s  } = _0193_ + \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.cin ;
always @(posedge \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.clk )
\add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.bin_s1  <= _0195_;
always @(posedge \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.clk )
\add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.ain_s1  <= _0194_;
always @(posedge \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.clk )
\add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.sum_s1  <= _0197_;
always @(posedge \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.clk )
\add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.carry_s1  <= _0196_;
assign _0195_ = \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.ce  ? \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.b [31:16] : \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.bin_s1 ;
assign _0194_ = \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.ce  ? \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.a [31:16] : \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.ain_s1 ;
assign _0196_ = \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.ce  ? \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.facout_s1  : \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.carry_s1 ;
assign _0197_ = \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.ce  ? \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.fas_s1  : \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.sum_s1 ;
assign _0198_ = \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.a  + \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.b ;
assign { \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.cout , \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.s  } = _0198_ + \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.cin ;
assign _0199_ = \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.a  + \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.b ;
assign { \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.cout , \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.s  } = _0199_ + \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.cin ;
always @(posedge \add_32ns_32ns_32_2_1_U27.top_add_32ns_32ns_32_2_1_Adder_15_U.clk )
\add_32ns_32ns_32_2_1_U27.top_add_32ns_32ns_32_2_1_Adder_15_U.bin_s1  <= _0201_;
always @(posedge \add_32ns_32ns_32_2_1_U27.top_add_32ns_32ns_32_2_1_Adder_15_U.clk )
\add_32ns_32ns_32_2_1_U27.top_add_32ns_32ns_32_2_1_Adder_15_U.ain_s1  <= _0200_;
always @(posedge \add_32ns_32ns_32_2_1_U27.top_add_32ns_32ns_32_2_1_Adder_15_U.clk )
\add_32ns_32ns_32_2_1_U27.top_add_32ns_32ns_32_2_1_Adder_15_U.sum_s1  <= _0203_;
always @(posedge \add_32ns_32ns_32_2_1_U27.top_add_32ns_32ns_32_2_1_Adder_15_U.clk )
\add_32ns_32ns_32_2_1_U27.top_add_32ns_32ns_32_2_1_Adder_15_U.carry_s1  <= _0202_;
assign _0201_ = \add_32ns_32ns_32_2_1_U27.top_add_32ns_32ns_32_2_1_Adder_15_U.ce  ? \add_32ns_32ns_32_2_1_U27.top_add_32ns_32ns_32_2_1_Adder_15_U.b [31:16] : \add_32ns_32ns_32_2_1_U27.top_add_32ns_32ns_32_2_1_Adder_15_U.bin_s1 ;
assign _0200_ = \add_32ns_32ns_32_2_1_U27.top_add_32ns_32ns_32_2_1_Adder_15_U.ce  ? \add_32ns_32ns_32_2_1_U27.top_add_32ns_32ns_32_2_1_Adder_15_U.a [31:16] : \add_32ns_32ns_32_2_1_U27.top_add_32ns_32ns_32_2_1_Adder_15_U.ain_s1 ;
assign _0202_ = \add_32ns_32ns_32_2_1_U27.top_add_32ns_32ns_32_2_1_Adder_15_U.ce  ? \add_32ns_32ns_32_2_1_U27.top_add_32ns_32ns_32_2_1_Adder_15_U.facout_s1  : \add_32ns_32ns_32_2_1_U27.top_add_32ns_32ns_32_2_1_Adder_15_U.carry_s1 ;
assign _0203_ = \add_32ns_32ns_32_2_1_U27.top_add_32ns_32ns_32_2_1_Adder_15_U.ce  ? \add_32ns_32ns_32_2_1_U27.top_add_32ns_32ns_32_2_1_Adder_15_U.fas_s1  : \add_32ns_32ns_32_2_1_U27.top_add_32ns_32ns_32_2_1_Adder_15_U.sum_s1 ;
assign _0204_ = \add_32ns_32ns_32_2_1_U27.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.a  + \add_32ns_32ns_32_2_1_U27.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.b ;
assign { \add_32ns_32ns_32_2_1_U27.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.cout , \add_32ns_32ns_32_2_1_U27.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.s  } = _0204_ + \add_32ns_32ns_32_2_1_U27.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.cin ;
assign _0205_ = \add_32ns_32ns_32_2_1_U27.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.a  + \add_32ns_32ns_32_2_1_U27.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.b ;
assign { \add_32ns_32ns_32_2_1_U27.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.cout , \add_32ns_32ns_32_2_1_U27.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.s  } = _0205_ + \add_32ns_32ns_32_2_1_U27.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.cin ;
always @(posedge \add_32s_32ns_32_2_1_U29.top_add_32s_32ns_32_2_1_Adder_19_U.clk )
\add_32s_32ns_32_2_1_U29.top_add_32s_32ns_32_2_1_Adder_19_U.bin_s1  <= _0207_;
always @(posedge \add_32s_32ns_32_2_1_U29.top_add_32s_32ns_32_2_1_Adder_19_U.clk )
\add_32s_32ns_32_2_1_U29.top_add_32s_32ns_32_2_1_Adder_19_U.ain_s1  <= _0206_;
always @(posedge \add_32s_32ns_32_2_1_U29.top_add_32s_32ns_32_2_1_Adder_19_U.clk )
\add_32s_32ns_32_2_1_U29.top_add_32s_32ns_32_2_1_Adder_19_U.sum_s1  <= _0209_;
always @(posedge \add_32s_32ns_32_2_1_U29.top_add_32s_32ns_32_2_1_Adder_19_U.clk )
\add_32s_32ns_32_2_1_U29.top_add_32s_32ns_32_2_1_Adder_19_U.carry_s1  <= _0208_;
assign _0207_ = \add_32s_32ns_32_2_1_U29.top_add_32s_32ns_32_2_1_Adder_19_U.ce  ? \add_32s_32ns_32_2_1_U29.top_add_32s_32ns_32_2_1_Adder_19_U.b [31:16] : \add_32s_32ns_32_2_1_U29.top_add_32s_32ns_32_2_1_Adder_19_U.bin_s1 ;
assign _0206_ = \add_32s_32ns_32_2_1_U29.top_add_32s_32ns_32_2_1_Adder_19_U.ce  ? \add_32s_32ns_32_2_1_U29.top_add_32s_32ns_32_2_1_Adder_19_U.a [31:16] : \add_32s_32ns_32_2_1_U29.top_add_32s_32ns_32_2_1_Adder_19_U.ain_s1 ;
assign _0208_ = \add_32s_32ns_32_2_1_U29.top_add_32s_32ns_32_2_1_Adder_19_U.ce  ? \add_32s_32ns_32_2_1_U29.top_add_32s_32ns_32_2_1_Adder_19_U.facout_s1  : \add_32s_32ns_32_2_1_U29.top_add_32s_32ns_32_2_1_Adder_19_U.carry_s1 ;
assign _0209_ = \add_32s_32ns_32_2_1_U29.top_add_32s_32ns_32_2_1_Adder_19_U.ce  ? \add_32s_32ns_32_2_1_U29.top_add_32s_32ns_32_2_1_Adder_19_U.fas_s1  : \add_32s_32ns_32_2_1_U29.top_add_32s_32ns_32_2_1_Adder_19_U.sum_s1 ;
assign _0210_ = \add_32s_32ns_32_2_1_U29.top_add_32s_32ns_32_2_1_Adder_19_U.u1.a  + \add_32s_32ns_32_2_1_U29.top_add_32s_32ns_32_2_1_Adder_19_U.u1.b ;
assign { \add_32s_32ns_32_2_1_U29.top_add_32s_32ns_32_2_1_Adder_19_U.u1.cout , \add_32s_32ns_32_2_1_U29.top_add_32s_32ns_32_2_1_Adder_19_U.u1.s  } = _0210_ + \add_32s_32ns_32_2_1_U29.top_add_32s_32ns_32_2_1_Adder_19_U.u1.cin ;
assign _0211_ = \add_32s_32ns_32_2_1_U29.top_add_32s_32ns_32_2_1_Adder_19_U.u2.a  + \add_32s_32ns_32_2_1_U29.top_add_32s_32ns_32_2_1_Adder_19_U.u2.b ;
assign { \add_32s_32ns_32_2_1_U29.top_add_32s_32ns_32_2_1_Adder_19_U.u2.cout , \add_32s_32ns_32_2_1_U29.top_add_32s_32ns_32_2_1_Adder_19_U.u2.s  } = _0211_ + \add_32s_32ns_32_2_1_U29.top_add_32s_32ns_32_2_1_Adder_19_U.u2.cin ;
always @(posedge \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_16_U.clk )
\add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_16_U.bin_s1  <= _0213_;
always @(posedge \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_16_U.clk )
\add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_16_U.ain_s1  <= _0212_;
always @(posedge \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_16_U.clk )
\add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_16_U.sum_s1  <= _0215_;
always @(posedge \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_16_U.clk )
\add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_16_U.carry_s1  <= _0214_;
assign _0213_ = \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_16_U.ce  ? \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_16_U.b [33:17] : \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_16_U.bin_s1 ;
assign _0212_ = \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_16_U.ce  ? \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_16_U.a [33:17] : \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_16_U.ain_s1 ;
assign _0214_ = \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_16_U.ce  ? \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_16_U.facout_s1  : \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_16_U.carry_s1 ;
assign _0215_ = \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_16_U.ce  ? \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_16_U.fas_s1  : \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_16_U.sum_s1 ;
assign _0216_ = \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_16_U.u1.a  + \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_16_U.u1.b ;
assign { \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_16_U.u1.cout , \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_16_U.u1.s  } = _0216_ + \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_16_U.u1.cin ;
assign _0217_ = \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_16_U.u2.a  + \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_16_U.u2.b ;
assign { \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_16_U.u2.cout , \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_16_U.u2.s  } = _0217_ + \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_16_U.u2.cin ;
always @(posedge \add_35s_35s_35_2_1_U19.top_add_35s_35s_35_2_1_Adder_14_U.clk )
\add_35s_35s_35_2_1_U19.top_add_35s_35s_35_2_1_Adder_14_U.bin_s1  <= _0219_;
always @(posedge \add_35s_35s_35_2_1_U19.top_add_35s_35s_35_2_1_Adder_14_U.clk )
\add_35s_35s_35_2_1_U19.top_add_35s_35s_35_2_1_Adder_14_U.ain_s1  <= _0218_;
always @(posedge \add_35s_35s_35_2_1_U19.top_add_35s_35s_35_2_1_Adder_14_U.clk )
\add_35s_35s_35_2_1_U19.top_add_35s_35s_35_2_1_Adder_14_U.sum_s1  <= _0221_;
always @(posedge \add_35s_35s_35_2_1_U19.top_add_35s_35s_35_2_1_Adder_14_U.clk )
\add_35s_35s_35_2_1_U19.top_add_35s_35s_35_2_1_Adder_14_U.carry_s1  <= _0220_;
assign _0219_ = \add_35s_35s_35_2_1_U19.top_add_35s_35s_35_2_1_Adder_14_U.ce  ? \add_35s_35s_35_2_1_U19.top_add_35s_35s_35_2_1_Adder_14_U.b [34:17] : \add_35s_35s_35_2_1_U19.top_add_35s_35s_35_2_1_Adder_14_U.bin_s1 ;
assign _0218_ = \add_35s_35s_35_2_1_U19.top_add_35s_35s_35_2_1_Adder_14_U.ce  ? \add_35s_35s_35_2_1_U19.top_add_35s_35s_35_2_1_Adder_14_U.a [34:17] : \add_35s_35s_35_2_1_U19.top_add_35s_35s_35_2_1_Adder_14_U.ain_s1 ;
assign _0220_ = \add_35s_35s_35_2_1_U19.top_add_35s_35s_35_2_1_Adder_14_U.ce  ? \add_35s_35s_35_2_1_U19.top_add_35s_35s_35_2_1_Adder_14_U.facout_s1  : \add_35s_35s_35_2_1_U19.top_add_35s_35s_35_2_1_Adder_14_U.carry_s1 ;
assign _0221_ = \add_35s_35s_35_2_1_U19.top_add_35s_35s_35_2_1_Adder_14_U.ce  ? \add_35s_35s_35_2_1_U19.top_add_35s_35s_35_2_1_Adder_14_U.fas_s1  : \add_35s_35s_35_2_1_U19.top_add_35s_35s_35_2_1_Adder_14_U.sum_s1 ;
assign _0222_ = \add_35s_35s_35_2_1_U19.top_add_35s_35s_35_2_1_Adder_14_U.u1.a  + \add_35s_35s_35_2_1_U19.top_add_35s_35s_35_2_1_Adder_14_U.u1.b ;
assign { \add_35s_35s_35_2_1_U19.top_add_35s_35s_35_2_1_Adder_14_U.u1.cout , \add_35s_35s_35_2_1_U19.top_add_35s_35s_35_2_1_Adder_14_U.u1.s  } = _0222_ + \add_35s_35s_35_2_1_U19.top_add_35s_35s_35_2_1_Adder_14_U.u1.cin ;
assign _0223_ = \add_35s_35s_35_2_1_U19.top_add_35s_35s_35_2_1_Adder_14_U.u2.a  + \add_35s_35s_35_2_1_U19.top_add_35s_35s_35_2_1_Adder_14_U.u2.b ;
assign { \add_35s_35s_35_2_1_U19.top_add_35s_35s_35_2_1_Adder_14_U.u2.cout , \add_35s_35s_35_2_1_U19.top_add_35s_35s_35_2_1_Adder_14_U.u2.s  } = _0223_ + \add_35s_35s_35_2_1_U19.top_add_35s_35s_35_2_1_Adder_14_U.u2.cin ;
always @(posedge \add_35s_35s_35_2_1_U21.top_add_35s_35s_35_2_1_Adder_14_U.clk )
\add_35s_35s_35_2_1_U21.top_add_35s_35s_35_2_1_Adder_14_U.bin_s1  <= _0225_;
always @(posedge \add_35s_35s_35_2_1_U21.top_add_35s_35s_35_2_1_Adder_14_U.clk )
\add_35s_35s_35_2_1_U21.top_add_35s_35s_35_2_1_Adder_14_U.ain_s1  <= _0224_;
always @(posedge \add_35s_35s_35_2_1_U21.top_add_35s_35s_35_2_1_Adder_14_U.clk )
\add_35s_35s_35_2_1_U21.top_add_35s_35s_35_2_1_Adder_14_U.sum_s1  <= _0227_;
always @(posedge \add_35s_35s_35_2_1_U21.top_add_35s_35s_35_2_1_Adder_14_U.clk )
\add_35s_35s_35_2_1_U21.top_add_35s_35s_35_2_1_Adder_14_U.carry_s1  <= _0226_;
assign _0225_ = \add_35s_35s_35_2_1_U21.top_add_35s_35s_35_2_1_Adder_14_U.ce  ? \add_35s_35s_35_2_1_U21.top_add_35s_35s_35_2_1_Adder_14_U.b [34:17] : \add_35s_35s_35_2_1_U21.top_add_35s_35s_35_2_1_Adder_14_U.bin_s1 ;
assign _0224_ = \add_35s_35s_35_2_1_U21.top_add_35s_35s_35_2_1_Adder_14_U.ce  ? \add_35s_35s_35_2_1_U21.top_add_35s_35s_35_2_1_Adder_14_U.a [34:17] : \add_35s_35s_35_2_1_U21.top_add_35s_35s_35_2_1_Adder_14_U.ain_s1 ;
assign _0226_ = \add_35s_35s_35_2_1_U21.top_add_35s_35s_35_2_1_Adder_14_U.ce  ? \add_35s_35s_35_2_1_U21.top_add_35s_35s_35_2_1_Adder_14_U.facout_s1  : \add_35s_35s_35_2_1_U21.top_add_35s_35s_35_2_1_Adder_14_U.carry_s1 ;
assign _0227_ = \add_35s_35s_35_2_1_U21.top_add_35s_35s_35_2_1_Adder_14_U.ce  ? \add_35s_35s_35_2_1_U21.top_add_35s_35s_35_2_1_Adder_14_U.fas_s1  : \add_35s_35s_35_2_1_U21.top_add_35s_35s_35_2_1_Adder_14_U.sum_s1 ;
assign _0228_ = \add_35s_35s_35_2_1_U21.top_add_35s_35s_35_2_1_Adder_14_U.u1.a  + \add_35s_35s_35_2_1_U21.top_add_35s_35s_35_2_1_Adder_14_U.u1.b ;
assign { \add_35s_35s_35_2_1_U21.top_add_35s_35s_35_2_1_Adder_14_U.u1.cout , \add_35s_35s_35_2_1_U21.top_add_35s_35s_35_2_1_Adder_14_U.u1.s  } = _0228_ + \add_35s_35s_35_2_1_U21.top_add_35s_35s_35_2_1_Adder_14_U.u1.cin ;
assign _0229_ = \add_35s_35s_35_2_1_U21.top_add_35s_35s_35_2_1_Adder_14_U.u2.a  + \add_35s_35s_35_2_1_U21.top_add_35s_35s_35_2_1_Adder_14_U.u2.b ;
assign { \add_35s_35s_35_2_1_U21.top_add_35s_35s_35_2_1_Adder_14_U.u2.cout , \add_35s_35s_35_2_1_U21.top_add_35s_35s_35_2_1_Adder_14_U.u2.s  } = _0229_ + \add_35s_35s_35_2_1_U21.top_add_35s_35s_35_2_1_Adder_14_U.u2.cin ;
always @(posedge \add_3ns_3ns_3_2_1_U1.top_add_3ns_3ns_3_2_1_Adder_0_U.clk )
\add_3ns_3ns_3_2_1_U1.top_add_3ns_3ns_3_2_1_Adder_0_U.bin_s1  <= _0231_;
always @(posedge \add_3ns_3ns_3_2_1_U1.top_add_3ns_3ns_3_2_1_Adder_0_U.clk )
\add_3ns_3ns_3_2_1_U1.top_add_3ns_3ns_3_2_1_Adder_0_U.ain_s1  <= _0230_;
always @(posedge \add_3ns_3ns_3_2_1_U1.top_add_3ns_3ns_3_2_1_Adder_0_U.clk )
\add_3ns_3ns_3_2_1_U1.top_add_3ns_3ns_3_2_1_Adder_0_U.sum_s1  <= _0233_;
always @(posedge \add_3ns_3ns_3_2_1_U1.top_add_3ns_3ns_3_2_1_Adder_0_U.clk )
\add_3ns_3ns_3_2_1_U1.top_add_3ns_3ns_3_2_1_Adder_0_U.carry_s1  <= _0232_;
assign _0231_ = \add_3ns_3ns_3_2_1_U1.top_add_3ns_3ns_3_2_1_Adder_0_U.ce  ? \add_3ns_3ns_3_2_1_U1.top_add_3ns_3ns_3_2_1_Adder_0_U.b [2:1] : \add_3ns_3ns_3_2_1_U1.top_add_3ns_3ns_3_2_1_Adder_0_U.bin_s1 ;
assign _0230_ = \add_3ns_3ns_3_2_1_U1.top_add_3ns_3ns_3_2_1_Adder_0_U.ce  ? \add_3ns_3ns_3_2_1_U1.top_add_3ns_3ns_3_2_1_Adder_0_U.a [2:1] : \add_3ns_3ns_3_2_1_U1.top_add_3ns_3ns_3_2_1_Adder_0_U.ain_s1 ;
assign _0232_ = \add_3ns_3ns_3_2_1_U1.top_add_3ns_3ns_3_2_1_Adder_0_U.ce  ? \add_3ns_3ns_3_2_1_U1.top_add_3ns_3ns_3_2_1_Adder_0_U.facout_s1  : \add_3ns_3ns_3_2_1_U1.top_add_3ns_3ns_3_2_1_Adder_0_U.carry_s1 ;
assign _0233_ = \add_3ns_3ns_3_2_1_U1.top_add_3ns_3ns_3_2_1_Adder_0_U.ce  ? \add_3ns_3ns_3_2_1_U1.top_add_3ns_3ns_3_2_1_Adder_0_U.fas_s1  : \add_3ns_3ns_3_2_1_U1.top_add_3ns_3ns_3_2_1_Adder_0_U.sum_s1 ;
assign _0234_ = \add_3ns_3ns_3_2_1_U1.top_add_3ns_3ns_3_2_1_Adder_0_U.u1.a  + \add_3ns_3ns_3_2_1_U1.top_add_3ns_3ns_3_2_1_Adder_0_U.u1.b ;
assign { \add_3ns_3ns_3_2_1_U1.top_add_3ns_3ns_3_2_1_Adder_0_U.u1.cout , \add_3ns_3ns_3_2_1_U1.top_add_3ns_3ns_3_2_1_Adder_0_U.u1.s  } = _0234_ + \add_3ns_3ns_3_2_1_U1.top_add_3ns_3ns_3_2_1_Adder_0_U.u1.cin ;
assign _0235_ = \add_3ns_3ns_3_2_1_U1.top_add_3ns_3ns_3_2_1_Adder_0_U.u2.a  + \add_3ns_3ns_3_2_1_U1.top_add_3ns_3ns_3_2_1_Adder_0_U.u2.b ;
assign { \add_3ns_3ns_3_2_1_U1.top_add_3ns_3ns_3_2_1_Adder_0_U.u2.cout , \add_3ns_3ns_3_2_1_U1.top_add_3ns_3ns_3_2_1_Adder_0_U.u2.s  } = _0235_ + \add_3ns_3ns_3_2_1_U1.top_add_3ns_3ns_3_2_1_Adder_0_U.u2.cin ;
always @(posedge \add_4ns_4ns_4_2_1_U18.top_add_4ns_4ns_4_2_1_Adder_5_U.clk )
\add_4ns_4ns_4_2_1_U18.top_add_4ns_4ns_4_2_1_Adder_5_U.bin_s1  <= _0237_;
always @(posedge \add_4ns_4ns_4_2_1_U18.top_add_4ns_4ns_4_2_1_Adder_5_U.clk )
\add_4ns_4ns_4_2_1_U18.top_add_4ns_4ns_4_2_1_Adder_5_U.ain_s1  <= _0236_;
always @(posedge \add_4ns_4ns_4_2_1_U18.top_add_4ns_4ns_4_2_1_Adder_5_U.clk )
\add_4ns_4ns_4_2_1_U18.top_add_4ns_4ns_4_2_1_Adder_5_U.sum_s1  <= _0239_;
always @(posedge \add_4ns_4ns_4_2_1_U18.top_add_4ns_4ns_4_2_1_Adder_5_U.clk )
\add_4ns_4ns_4_2_1_U18.top_add_4ns_4ns_4_2_1_Adder_5_U.carry_s1  <= _0238_;
assign _0237_ = \add_4ns_4ns_4_2_1_U18.top_add_4ns_4ns_4_2_1_Adder_5_U.ce  ? \add_4ns_4ns_4_2_1_U18.top_add_4ns_4ns_4_2_1_Adder_5_U.b [3:2] : \add_4ns_4ns_4_2_1_U18.top_add_4ns_4ns_4_2_1_Adder_5_U.bin_s1 ;
assign _0236_ = \add_4ns_4ns_4_2_1_U18.top_add_4ns_4ns_4_2_1_Adder_5_U.ce  ? \add_4ns_4ns_4_2_1_U18.top_add_4ns_4ns_4_2_1_Adder_5_U.a [3:2] : \add_4ns_4ns_4_2_1_U18.top_add_4ns_4ns_4_2_1_Adder_5_U.ain_s1 ;
assign _0238_ = \add_4ns_4ns_4_2_1_U18.top_add_4ns_4ns_4_2_1_Adder_5_U.ce  ? \add_4ns_4ns_4_2_1_U18.top_add_4ns_4ns_4_2_1_Adder_5_U.facout_s1  : \add_4ns_4ns_4_2_1_U18.top_add_4ns_4ns_4_2_1_Adder_5_U.carry_s1 ;
assign _0239_ = \add_4ns_4ns_4_2_1_U18.top_add_4ns_4ns_4_2_1_Adder_5_U.ce  ? \add_4ns_4ns_4_2_1_U18.top_add_4ns_4ns_4_2_1_Adder_5_U.fas_s1  : \add_4ns_4ns_4_2_1_U18.top_add_4ns_4ns_4_2_1_Adder_5_U.sum_s1 ;
assign _0240_ = \add_4ns_4ns_4_2_1_U18.top_add_4ns_4ns_4_2_1_Adder_5_U.u1.a  + \add_4ns_4ns_4_2_1_U18.top_add_4ns_4ns_4_2_1_Adder_5_U.u1.b ;
assign { \add_4ns_4ns_4_2_1_U18.top_add_4ns_4ns_4_2_1_Adder_5_U.u1.cout , \add_4ns_4ns_4_2_1_U18.top_add_4ns_4ns_4_2_1_Adder_5_U.u1.s  } = _0240_ + \add_4ns_4ns_4_2_1_U18.top_add_4ns_4ns_4_2_1_Adder_5_U.u1.cin ;
assign _0241_ = \add_4ns_4ns_4_2_1_U18.top_add_4ns_4ns_4_2_1_Adder_5_U.u2.a  + \add_4ns_4ns_4_2_1_U18.top_add_4ns_4ns_4_2_1_Adder_5_U.u2.b ;
assign { \add_4ns_4ns_4_2_1_U18.top_add_4ns_4ns_4_2_1_Adder_5_U.u2.cout , \add_4ns_4ns_4_2_1_U18.top_add_4ns_4ns_4_2_1_Adder_5_U.u2.s  } = _0241_ + \add_4ns_4ns_4_2_1_U18.top_add_4ns_4ns_4_2_1_Adder_5_U.u2.cin ;
always @(posedge \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_5_U.clk )
\add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_5_U.bin_s1  <= _0243_;
always @(posedge \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_5_U.clk )
\add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_5_U.ain_s1  <= _0242_;
always @(posedge \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_5_U.clk )
\add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_5_U.sum_s1  <= _0245_;
always @(posedge \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_5_U.clk )
\add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_5_U.carry_s1  <= _0244_;
assign _0243_ = \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_5_U.ce  ? \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_5_U.b [3:2] : \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_5_U.bin_s1 ;
assign _0242_ = \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_5_U.ce  ? \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_5_U.a [3:2] : \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_5_U.ain_s1 ;
assign _0244_ = \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_5_U.ce  ? \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_5_U.facout_s1  : \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_5_U.carry_s1 ;
assign _0245_ = \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_5_U.ce  ? \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_5_U.fas_s1  : \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_5_U.sum_s1 ;
assign _0246_ = \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_5_U.u1.a  + \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_5_U.u1.b ;
assign { \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_5_U.u1.cout , \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_5_U.u1.s  } = _0246_ + \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_5_U.u1.cin ;
assign _0247_ = \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_5_U.u2.a  + \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_5_U.u2.b ;
assign { \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_5_U.u2.cout , \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_5_U.u2.s  } = _0247_ + \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_5_U.u2.cin ;
always @(posedge \add_4s_4ns_4_2_1_U4.top_add_4s_4ns_4_2_1_Adder_3_U.clk )
\add_4s_4ns_4_2_1_U4.top_add_4s_4ns_4_2_1_Adder_3_U.bin_s1  <= _0249_;
always @(posedge \add_4s_4ns_4_2_1_U4.top_add_4s_4ns_4_2_1_Adder_3_U.clk )
\add_4s_4ns_4_2_1_U4.top_add_4s_4ns_4_2_1_Adder_3_U.ain_s1  <= _0248_;
always @(posedge \add_4s_4ns_4_2_1_U4.top_add_4s_4ns_4_2_1_Adder_3_U.clk )
\add_4s_4ns_4_2_1_U4.top_add_4s_4ns_4_2_1_Adder_3_U.sum_s1  <= _0251_;
always @(posedge \add_4s_4ns_4_2_1_U4.top_add_4s_4ns_4_2_1_Adder_3_U.clk )
\add_4s_4ns_4_2_1_U4.top_add_4s_4ns_4_2_1_Adder_3_U.carry_s1  <= _0250_;
assign _0249_ = \add_4s_4ns_4_2_1_U4.top_add_4s_4ns_4_2_1_Adder_3_U.ce  ? \add_4s_4ns_4_2_1_U4.top_add_4s_4ns_4_2_1_Adder_3_U.b [3:2] : \add_4s_4ns_4_2_1_U4.top_add_4s_4ns_4_2_1_Adder_3_U.bin_s1 ;
assign _0248_ = \add_4s_4ns_4_2_1_U4.top_add_4s_4ns_4_2_1_Adder_3_U.ce  ? \add_4s_4ns_4_2_1_U4.top_add_4s_4ns_4_2_1_Adder_3_U.a [3:2] : \add_4s_4ns_4_2_1_U4.top_add_4s_4ns_4_2_1_Adder_3_U.ain_s1 ;
assign _0250_ = \add_4s_4ns_4_2_1_U4.top_add_4s_4ns_4_2_1_Adder_3_U.ce  ? \add_4s_4ns_4_2_1_U4.top_add_4s_4ns_4_2_1_Adder_3_U.facout_s1  : \add_4s_4ns_4_2_1_U4.top_add_4s_4ns_4_2_1_Adder_3_U.carry_s1 ;
assign _0251_ = \add_4s_4ns_4_2_1_U4.top_add_4s_4ns_4_2_1_Adder_3_U.ce  ? \add_4s_4ns_4_2_1_U4.top_add_4s_4ns_4_2_1_Adder_3_U.fas_s1  : \add_4s_4ns_4_2_1_U4.top_add_4s_4ns_4_2_1_Adder_3_U.sum_s1 ;
assign _0252_ = \add_4s_4ns_4_2_1_U4.top_add_4s_4ns_4_2_1_Adder_3_U.u1.a  + \add_4s_4ns_4_2_1_U4.top_add_4s_4ns_4_2_1_Adder_3_U.u1.b ;
assign { \add_4s_4ns_4_2_1_U4.top_add_4s_4ns_4_2_1_Adder_3_U.u1.cout , \add_4s_4ns_4_2_1_U4.top_add_4s_4ns_4_2_1_Adder_3_U.u1.s  } = _0252_ + \add_4s_4ns_4_2_1_U4.top_add_4s_4ns_4_2_1_Adder_3_U.u1.cin ;
assign _0253_ = \add_4s_4ns_4_2_1_U4.top_add_4s_4ns_4_2_1_Adder_3_U.u2.a  + \add_4s_4ns_4_2_1_U4.top_add_4s_4ns_4_2_1_Adder_3_U.u2.b ;
assign { \add_4s_4ns_4_2_1_U4.top_add_4s_4ns_4_2_1_Adder_3_U.u2.cout , \add_4s_4ns_4_2_1_U4.top_add_4s_4ns_4_2_1_Adder_3_U.u2.s  } = _0253_ + \add_4s_4ns_4_2_1_U4.top_add_4s_4ns_4_2_1_Adder_3_U.u2.cin ;
always @(posedge \add_5ns_5s_5_2_1_U3.top_add_5ns_5s_5_2_1_Adder_2_U.clk )
\add_5ns_5s_5_2_1_U3.top_add_5ns_5s_5_2_1_Adder_2_U.bin_s1  <= _0255_;
always @(posedge \add_5ns_5s_5_2_1_U3.top_add_5ns_5s_5_2_1_Adder_2_U.clk )
\add_5ns_5s_5_2_1_U3.top_add_5ns_5s_5_2_1_Adder_2_U.ain_s1  <= _0254_;
always @(posedge \add_5ns_5s_5_2_1_U3.top_add_5ns_5s_5_2_1_Adder_2_U.clk )
\add_5ns_5s_5_2_1_U3.top_add_5ns_5s_5_2_1_Adder_2_U.sum_s1  <= _0257_;
always @(posedge \add_5ns_5s_5_2_1_U3.top_add_5ns_5s_5_2_1_Adder_2_U.clk )
\add_5ns_5s_5_2_1_U3.top_add_5ns_5s_5_2_1_Adder_2_U.carry_s1  <= _0256_;
assign _0255_ = \add_5ns_5s_5_2_1_U3.top_add_5ns_5s_5_2_1_Adder_2_U.ce  ? \add_5ns_5s_5_2_1_U3.top_add_5ns_5s_5_2_1_Adder_2_U.b [4:2] : \add_5ns_5s_5_2_1_U3.top_add_5ns_5s_5_2_1_Adder_2_U.bin_s1 ;
assign _0254_ = \add_5ns_5s_5_2_1_U3.top_add_5ns_5s_5_2_1_Adder_2_U.ce  ? \add_5ns_5s_5_2_1_U3.top_add_5ns_5s_5_2_1_Adder_2_U.a [4:2] : \add_5ns_5s_5_2_1_U3.top_add_5ns_5s_5_2_1_Adder_2_U.ain_s1 ;
assign _0256_ = \add_5ns_5s_5_2_1_U3.top_add_5ns_5s_5_2_1_Adder_2_U.ce  ? \add_5ns_5s_5_2_1_U3.top_add_5ns_5s_5_2_1_Adder_2_U.facout_s1  : \add_5ns_5s_5_2_1_U3.top_add_5ns_5s_5_2_1_Adder_2_U.carry_s1 ;
assign _0257_ = \add_5ns_5s_5_2_1_U3.top_add_5ns_5s_5_2_1_Adder_2_U.ce  ? \add_5ns_5s_5_2_1_U3.top_add_5ns_5s_5_2_1_Adder_2_U.fas_s1  : \add_5ns_5s_5_2_1_U3.top_add_5ns_5s_5_2_1_Adder_2_U.sum_s1 ;
assign _0258_ = \add_5ns_5s_5_2_1_U3.top_add_5ns_5s_5_2_1_Adder_2_U.u1.a  + \add_5ns_5s_5_2_1_U3.top_add_5ns_5s_5_2_1_Adder_2_U.u1.b ;
assign { \add_5ns_5s_5_2_1_U3.top_add_5ns_5s_5_2_1_Adder_2_U.u1.cout , \add_5ns_5s_5_2_1_U3.top_add_5ns_5s_5_2_1_Adder_2_U.u1.s  } = _0258_ + \add_5ns_5s_5_2_1_U3.top_add_5ns_5s_5_2_1_Adder_2_U.u1.cin ;
assign _0259_ = \add_5ns_5s_5_2_1_U3.top_add_5ns_5s_5_2_1_Adder_2_U.u2.a  + \add_5ns_5s_5_2_1_U3.top_add_5ns_5s_5_2_1_Adder_2_U.u2.b ;
assign { \add_5ns_5s_5_2_1_U3.top_add_5ns_5s_5_2_1_Adder_2_U.u2.cout , \add_5ns_5s_5_2_1_U3.top_add_5ns_5s_5_2_1_Adder_2_U.u2.s  } = _0259_ + \add_5ns_5s_5_2_1_U3.top_add_5ns_5s_5_2_1_Adder_2_U.u2.cin ;
always @(posedge \add_7s_7s_7_2_1_U2.top_add_7s_7s_7_2_1_Adder_1_U.clk )
\add_7s_7s_7_2_1_U2.top_add_7s_7s_7_2_1_Adder_1_U.bin_s1  <= _0261_;
always @(posedge \add_7s_7s_7_2_1_U2.top_add_7s_7s_7_2_1_Adder_1_U.clk )
\add_7s_7s_7_2_1_U2.top_add_7s_7s_7_2_1_Adder_1_U.ain_s1  <= _0260_;
always @(posedge \add_7s_7s_7_2_1_U2.top_add_7s_7s_7_2_1_Adder_1_U.clk )
\add_7s_7s_7_2_1_U2.top_add_7s_7s_7_2_1_Adder_1_U.sum_s1  <= _0263_;
always @(posedge \add_7s_7s_7_2_1_U2.top_add_7s_7s_7_2_1_Adder_1_U.clk )
\add_7s_7s_7_2_1_U2.top_add_7s_7s_7_2_1_Adder_1_U.carry_s1  <= _0262_;
assign _0261_ = \add_7s_7s_7_2_1_U2.top_add_7s_7s_7_2_1_Adder_1_U.ce  ? \add_7s_7s_7_2_1_U2.top_add_7s_7s_7_2_1_Adder_1_U.b [6:3] : \add_7s_7s_7_2_1_U2.top_add_7s_7s_7_2_1_Adder_1_U.bin_s1 ;
assign _0260_ = \add_7s_7s_7_2_1_U2.top_add_7s_7s_7_2_1_Adder_1_U.ce  ? \add_7s_7s_7_2_1_U2.top_add_7s_7s_7_2_1_Adder_1_U.a [6:3] : \add_7s_7s_7_2_1_U2.top_add_7s_7s_7_2_1_Adder_1_U.ain_s1 ;
assign _0262_ = \add_7s_7s_7_2_1_U2.top_add_7s_7s_7_2_1_Adder_1_U.ce  ? \add_7s_7s_7_2_1_U2.top_add_7s_7s_7_2_1_Adder_1_U.facout_s1  : \add_7s_7s_7_2_1_U2.top_add_7s_7s_7_2_1_Adder_1_U.carry_s1 ;
assign _0263_ = \add_7s_7s_7_2_1_U2.top_add_7s_7s_7_2_1_Adder_1_U.ce  ? \add_7s_7s_7_2_1_U2.top_add_7s_7s_7_2_1_Adder_1_U.fas_s1  : \add_7s_7s_7_2_1_U2.top_add_7s_7s_7_2_1_Adder_1_U.sum_s1 ;
assign _0264_ = \add_7s_7s_7_2_1_U2.top_add_7s_7s_7_2_1_Adder_1_U.u1.a  + \add_7s_7s_7_2_1_U2.top_add_7s_7s_7_2_1_Adder_1_U.u1.b ;
assign { \add_7s_7s_7_2_1_U2.top_add_7s_7s_7_2_1_Adder_1_U.u1.cout , \add_7s_7s_7_2_1_U2.top_add_7s_7s_7_2_1_Adder_1_U.u1.s  } = _0264_ + \add_7s_7s_7_2_1_U2.top_add_7s_7s_7_2_1_Adder_1_U.u1.cin ;
assign _0265_ = \add_7s_7s_7_2_1_U2.top_add_7s_7s_7_2_1_Adder_1_U.u2.a  + \add_7s_7s_7_2_1_U2.top_add_7s_7s_7_2_1_Adder_1_U.u2.b ;
assign { \add_7s_7s_7_2_1_U2.top_add_7s_7s_7_2_1_Adder_1_U.u2.cout , \add_7s_7s_7_2_1_U2.top_add_7s_7s_7_2_1_Adder_1_U.u2.s  } = _0265_ + \add_7s_7s_7_2_1_U2.top_add_7s_7s_7_2_1_Adder_1_U.u2.cin ;
always @(posedge \add_9s_9ns_9_2_1_U26.top_add_9s_9ns_9_2_1_Adder_17_U.clk )
\add_9s_9ns_9_2_1_U26.top_add_9s_9ns_9_2_1_Adder_17_U.bin_s1  <= _0267_;
always @(posedge \add_9s_9ns_9_2_1_U26.top_add_9s_9ns_9_2_1_Adder_17_U.clk )
\add_9s_9ns_9_2_1_U26.top_add_9s_9ns_9_2_1_Adder_17_U.ain_s1  <= _0266_;
always @(posedge \add_9s_9ns_9_2_1_U26.top_add_9s_9ns_9_2_1_Adder_17_U.clk )
\add_9s_9ns_9_2_1_U26.top_add_9s_9ns_9_2_1_Adder_17_U.sum_s1  <= _0269_;
always @(posedge \add_9s_9ns_9_2_1_U26.top_add_9s_9ns_9_2_1_Adder_17_U.clk )
\add_9s_9ns_9_2_1_U26.top_add_9s_9ns_9_2_1_Adder_17_U.carry_s1  <= _0268_;
assign _0267_ = \add_9s_9ns_9_2_1_U26.top_add_9s_9ns_9_2_1_Adder_17_U.ce  ? \add_9s_9ns_9_2_1_U26.top_add_9s_9ns_9_2_1_Adder_17_U.b [8:4] : \add_9s_9ns_9_2_1_U26.top_add_9s_9ns_9_2_1_Adder_17_U.bin_s1 ;
assign _0266_ = \add_9s_9ns_9_2_1_U26.top_add_9s_9ns_9_2_1_Adder_17_U.ce  ? \add_9s_9ns_9_2_1_U26.top_add_9s_9ns_9_2_1_Adder_17_U.a [8:4] : \add_9s_9ns_9_2_1_U26.top_add_9s_9ns_9_2_1_Adder_17_U.ain_s1 ;
assign _0268_ = \add_9s_9ns_9_2_1_U26.top_add_9s_9ns_9_2_1_Adder_17_U.ce  ? \add_9s_9ns_9_2_1_U26.top_add_9s_9ns_9_2_1_Adder_17_U.facout_s1  : \add_9s_9ns_9_2_1_U26.top_add_9s_9ns_9_2_1_Adder_17_U.carry_s1 ;
assign _0269_ = \add_9s_9ns_9_2_1_U26.top_add_9s_9ns_9_2_1_Adder_17_U.ce  ? \add_9s_9ns_9_2_1_U26.top_add_9s_9ns_9_2_1_Adder_17_U.fas_s1  : \add_9s_9ns_9_2_1_U26.top_add_9s_9ns_9_2_1_Adder_17_U.sum_s1 ;
assign _0270_ = \add_9s_9ns_9_2_1_U26.top_add_9s_9ns_9_2_1_Adder_17_U.u1.a  + \add_9s_9ns_9_2_1_U26.top_add_9s_9ns_9_2_1_Adder_17_U.u1.b ;
assign { \add_9s_9ns_9_2_1_U26.top_add_9s_9ns_9_2_1_Adder_17_U.u1.cout , \add_9s_9ns_9_2_1_U26.top_add_9s_9ns_9_2_1_Adder_17_U.u1.s  } = _0270_ + \add_9s_9ns_9_2_1_U26.top_add_9s_9ns_9_2_1_Adder_17_U.u1.cin ;
assign _0271_ = \add_9s_9ns_9_2_1_U26.top_add_9s_9ns_9_2_1_Adder_17_U.u2.a  + \add_9s_9ns_9_2_1_U26.top_add_9s_9ns_9_2_1_Adder_17_U.u2.b ;
assign { \add_9s_9ns_9_2_1_U26.top_add_9s_9ns_9_2_1_Adder_17_U.u2.cout , \add_9s_9ns_9_2_1_U26.top_add_9s_9ns_9_2_1_Adder_17_U.u2.s  } = _0271_ + \add_9s_9ns_9_2_1_U26.top_add_9s_9ns_9_2_1_Adder_17_U.u2.cin ;
assign \mul_32ns_4s_36_7_1_U5.top_mul_32ns_4s_36_7_1_Mul_DSP_0_U.tmp_product  = $signed({ 1'h0, \mul_32ns_4s_36_7_1_U5.top_mul_32ns_4s_36_7_1_Mul_DSP_0_U.a_reg0  }) * $signed(\mul_32ns_4s_36_7_1_U5.top_mul_32ns_4s_36_7_1_Mul_DSP_0_U.b_reg0 );
always @(posedge \mul_32ns_4s_36_7_1_U5.top_mul_32ns_4s_36_7_1_Mul_DSP_0_U.clk )
\mul_32ns_4s_36_7_1_U5.top_mul_32ns_4s_36_7_1_Mul_DSP_0_U.a_reg0  <= _0272_;
always @(posedge \mul_32ns_4s_36_7_1_U5.top_mul_32ns_4s_36_7_1_Mul_DSP_0_U.clk )
\mul_32ns_4s_36_7_1_U5.top_mul_32ns_4s_36_7_1_Mul_DSP_0_U.b_reg0  <= _0273_;
always @(posedge \mul_32ns_4s_36_7_1_U5.top_mul_32ns_4s_36_7_1_Mul_DSP_0_U.clk )
\mul_32ns_4s_36_7_1_U5.top_mul_32ns_4s_36_7_1_Mul_DSP_0_U.buff0  <= _0274_;
always @(posedge \mul_32ns_4s_36_7_1_U5.top_mul_32ns_4s_36_7_1_Mul_DSP_0_U.clk )
\mul_32ns_4s_36_7_1_U5.top_mul_32ns_4s_36_7_1_Mul_DSP_0_U.buff1  <= _0275_;
always @(posedge \mul_32ns_4s_36_7_1_U5.top_mul_32ns_4s_36_7_1_Mul_DSP_0_U.clk )
\mul_32ns_4s_36_7_1_U5.top_mul_32ns_4s_36_7_1_Mul_DSP_0_U.buff2  <= _0276_;
always @(posedge \mul_32ns_4s_36_7_1_U5.top_mul_32ns_4s_36_7_1_Mul_DSP_0_U.clk )
\mul_32ns_4s_36_7_1_U5.top_mul_32ns_4s_36_7_1_Mul_DSP_0_U.buff3  <= _0277_;
always @(posedge \mul_32ns_4s_36_7_1_U5.top_mul_32ns_4s_36_7_1_Mul_DSP_0_U.clk )
\mul_32ns_4s_36_7_1_U5.top_mul_32ns_4s_36_7_1_Mul_DSP_0_U.buff4  <= _0278_;
assign _0278_ = \mul_32ns_4s_36_7_1_U5.top_mul_32ns_4s_36_7_1_Mul_DSP_0_U.ce  ? \mul_32ns_4s_36_7_1_U5.top_mul_32ns_4s_36_7_1_Mul_DSP_0_U.buff3  : \mul_32ns_4s_36_7_1_U5.top_mul_32ns_4s_36_7_1_Mul_DSP_0_U.buff4 ;
assign _0277_ = \mul_32ns_4s_36_7_1_U5.top_mul_32ns_4s_36_7_1_Mul_DSP_0_U.ce  ? \mul_32ns_4s_36_7_1_U5.top_mul_32ns_4s_36_7_1_Mul_DSP_0_U.buff2  : \mul_32ns_4s_36_7_1_U5.top_mul_32ns_4s_36_7_1_Mul_DSP_0_U.buff3 ;
assign _0276_ = \mul_32ns_4s_36_7_1_U5.top_mul_32ns_4s_36_7_1_Mul_DSP_0_U.ce  ? \mul_32ns_4s_36_7_1_U5.top_mul_32ns_4s_36_7_1_Mul_DSP_0_U.buff1  : \mul_32ns_4s_36_7_1_U5.top_mul_32ns_4s_36_7_1_Mul_DSP_0_U.buff2 ;
assign _0275_ = \mul_32ns_4s_36_7_1_U5.top_mul_32ns_4s_36_7_1_Mul_DSP_0_U.ce  ? \mul_32ns_4s_36_7_1_U5.top_mul_32ns_4s_36_7_1_Mul_DSP_0_U.buff0  : \mul_32ns_4s_36_7_1_U5.top_mul_32ns_4s_36_7_1_Mul_DSP_0_U.buff1 ;
assign _0274_ = \mul_32ns_4s_36_7_1_U5.top_mul_32ns_4s_36_7_1_Mul_DSP_0_U.ce  ? \mul_32ns_4s_36_7_1_U5.top_mul_32ns_4s_36_7_1_Mul_DSP_0_U.tmp_product  : \mul_32ns_4s_36_7_1_U5.top_mul_32ns_4s_36_7_1_Mul_DSP_0_U.buff0 ;
assign _0273_ = \mul_32ns_4s_36_7_1_U5.top_mul_32ns_4s_36_7_1_Mul_DSP_0_U.ce  ? \mul_32ns_4s_36_7_1_U5.top_mul_32ns_4s_36_7_1_Mul_DSP_0_U.b  : \mul_32ns_4s_36_7_1_U5.top_mul_32ns_4s_36_7_1_Mul_DSP_0_U.b_reg0 ;
assign _0272_ = \mul_32ns_4s_36_7_1_U5.top_mul_32ns_4s_36_7_1_Mul_DSP_0_U.ce  ? \mul_32ns_4s_36_7_1_U5.top_mul_32ns_4s_36_7_1_Mul_DSP_0_U.a  : \mul_32ns_4s_36_7_1_U5.top_mul_32ns_4s_36_7_1_Mul_DSP_0_U.a_reg0 ;
assign \mul_32ns_4s_36_7_1_U6.top_mul_32ns_4s_36_7_1_Mul_DSP_0_U.tmp_product  = $signed({ 1'h0, \mul_32ns_4s_36_7_1_U6.top_mul_32ns_4s_36_7_1_Mul_DSP_0_U.a_reg0  }) * $signed(\mul_32ns_4s_36_7_1_U6.top_mul_32ns_4s_36_7_1_Mul_DSP_0_U.b_reg0 );
always @(posedge \mul_32ns_4s_36_7_1_U6.top_mul_32ns_4s_36_7_1_Mul_DSP_0_U.clk )
\mul_32ns_4s_36_7_1_U6.top_mul_32ns_4s_36_7_1_Mul_DSP_0_U.a_reg0  <= _0279_;
always @(posedge \mul_32ns_4s_36_7_1_U6.top_mul_32ns_4s_36_7_1_Mul_DSP_0_U.clk )
\mul_32ns_4s_36_7_1_U6.top_mul_32ns_4s_36_7_1_Mul_DSP_0_U.b_reg0  <= _0280_;
always @(posedge \mul_32ns_4s_36_7_1_U6.top_mul_32ns_4s_36_7_1_Mul_DSP_0_U.clk )
\mul_32ns_4s_36_7_1_U6.top_mul_32ns_4s_36_7_1_Mul_DSP_0_U.buff0  <= _0281_;
always @(posedge \mul_32ns_4s_36_7_1_U6.top_mul_32ns_4s_36_7_1_Mul_DSP_0_U.clk )
\mul_32ns_4s_36_7_1_U6.top_mul_32ns_4s_36_7_1_Mul_DSP_0_U.buff1  <= _0282_;
always @(posedge \mul_32ns_4s_36_7_1_U6.top_mul_32ns_4s_36_7_1_Mul_DSP_0_U.clk )
\mul_32ns_4s_36_7_1_U6.top_mul_32ns_4s_36_7_1_Mul_DSP_0_U.buff2  <= _0283_;
always @(posedge \mul_32ns_4s_36_7_1_U6.top_mul_32ns_4s_36_7_1_Mul_DSP_0_U.clk )
\mul_32ns_4s_36_7_1_U6.top_mul_32ns_4s_36_7_1_Mul_DSP_0_U.buff3  <= _0284_;
always @(posedge \mul_32ns_4s_36_7_1_U6.top_mul_32ns_4s_36_7_1_Mul_DSP_0_U.clk )
\mul_32ns_4s_36_7_1_U6.top_mul_32ns_4s_36_7_1_Mul_DSP_0_U.buff4  <= _0285_;
assign _0285_ = \mul_32ns_4s_36_7_1_U6.top_mul_32ns_4s_36_7_1_Mul_DSP_0_U.ce  ? \mul_32ns_4s_36_7_1_U6.top_mul_32ns_4s_36_7_1_Mul_DSP_0_U.buff3  : \mul_32ns_4s_36_7_1_U6.top_mul_32ns_4s_36_7_1_Mul_DSP_0_U.buff4 ;
assign _0284_ = \mul_32ns_4s_36_7_1_U6.top_mul_32ns_4s_36_7_1_Mul_DSP_0_U.ce  ? \mul_32ns_4s_36_7_1_U6.top_mul_32ns_4s_36_7_1_Mul_DSP_0_U.buff2  : \mul_32ns_4s_36_7_1_U6.top_mul_32ns_4s_36_7_1_Mul_DSP_0_U.buff3 ;
assign _0283_ = \mul_32ns_4s_36_7_1_U6.top_mul_32ns_4s_36_7_1_Mul_DSP_0_U.ce  ? \mul_32ns_4s_36_7_1_U6.top_mul_32ns_4s_36_7_1_Mul_DSP_0_U.buff1  : \mul_32ns_4s_36_7_1_U6.top_mul_32ns_4s_36_7_1_Mul_DSP_0_U.buff2 ;
assign _0282_ = \mul_32ns_4s_36_7_1_U6.top_mul_32ns_4s_36_7_1_Mul_DSP_0_U.ce  ? \mul_32ns_4s_36_7_1_U6.top_mul_32ns_4s_36_7_1_Mul_DSP_0_U.buff0  : \mul_32ns_4s_36_7_1_U6.top_mul_32ns_4s_36_7_1_Mul_DSP_0_U.buff1 ;
assign _0281_ = \mul_32ns_4s_36_7_1_U6.top_mul_32ns_4s_36_7_1_Mul_DSP_0_U.ce  ? \mul_32ns_4s_36_7_1_U6.top_mul_32ns_4s_36_7_1_Mul_DSP_0_U.tmp_product  : \mul_32ns_4s_36_7_1_U6.top_mul_32ns_4s_36_7_1_Mul_DSP_0_U.buff0 ;
assign _0280_ = \mul_32ns_4s_36_7_1_U6.top_mul_32ns_4s_36_7_1_Mul_DSP_0_U.ce  ? \mul_32ns_4s_36_7_1_U6.top_mul_32ns_4s_36_7_1_Mul_DSP_0_U.b  : \mul_32ns_4s_36_7_1_U6.top_mul_32ns_4s_36_7_1_Mul_DSP_0_U.b_reg0 ;
assign _0279_ = \mul_32ns_4s_36_7_1_U6.top_mul_32ns_4s_36_7_1_Mul_DSP_0_U.ce  ? \mul_32ns_4s_36_7_1_U6.top_mul_32ns_4s_36_7_1_Mul_DSP_0_U.a  : \mul_32ns_4s_36_7_1_U6.top_mul_32ns_4s_36_7_1_Mul_DSP_0_U.a_reg0 ;
assign \mul_4ns_3s_7_7_1_U12.top_mul_4ns_3s_7_7_1_Mul_DSP_1_U.tmp_product  = $signed({ 1'h0, \mul_4ns_3s_7_7_1_U12.top_mul_4ns_3s_7_7_1_Mul_DSP_1_U.a_reg0  }) * $signed(\mul_4ns_3s_7_7_1_U12.top_mul_4ns_3s_7_7_1_Mul_DSP_1_U.b_reg0 );
always @(posedge \mul_4ns_3s_7_7_1_U12.top_mul_4ns_3s_7_7_1_Mul_DSP_1_U.clk )
\mul_4ns_3s_7_7_1_U12.top_mul_4ns_3s_7_7_1_Mul_DSP_1_U.a_reg0  <= _0286_;
always @(posedge \mul_4ns_3s_7_7_1_U12.top_mul_4ns_3s_7_7_1_Mul_DSP_1_U.clk )
\mul_4ns_3s_7_7_1_U12.top_mul_4ns_3s_7_7_1_Mul_DSP_1_U.b_reg0  <= _0287_;
always @(posedge \mul_4ns_3s_7_7_1_U12.top_mul_4ns_3s_7_7_1_Mul_DSP_1_U.clk )
\mul_4ns_3s_7_7_1_U12.top_mul_4ns_3s_7_7_1_Mul_DSP_1_U.buff0  <= _0288_;
always @(posedge \mul_4ns_3s_7_7_1_U12.top_mul_4ns_3s_7_7_1_Mul_DSP_1_U.clk )
\mul_4ns_3s_7_7_1_U12.top_mul_4ns_3s_7_7_1_Mul_DSP_1_U.buff1  <= _0289_;
always @(posedge \mul_4ns_3s_7_7_1_U12.top_mul_4ns_3s_7_7_1_Mul_DSP_1_U.clk )
\mul_4ns_3s_7_7_1_U12.top_mul_4ns_3s_7_7_1_Mul_DSP_1_U.buff2  <= _0290_;
always @(posedge \mul_4ns_3s_7_7_1_U12.top_mul_4ns_3s_7_7_1_Mul_DSP_1_U.clk )
\mul_4ns_3s_7_7_1_U12.top_mul_4ns_3s_7_7_1_Mul_DSP_1_U.buff3  <= _0291_;
always @(posedge \mul_4ns_3s_7_7_1_U12.top_mul_4ns_3s_7_7_1_Mul_DSP_1_U.clk )
\mul_4ns_3s_7_7_1_U12.top_mul_4ns_3s_7_7_1_Mul_DSP_1_U.buff4  <= _0292_;
assign _0292_ = \mul_4ns_3s_7_7_1_U12.top_mul_4ns_3s_7_7_1_Mul_DSP_1_U.ce  ? \mul_4ns_3s_7_7_1_U12.top_mul_4ns_3s_7_7_1_Mul_DSP_1_U.buff3  : \mul_4ns_3s_7_7_1_U12.top_mul_4ns_3s_7_7_1_Mul_DSP_1_U.buff4 ;
assign _0291_ = \mul_4ns_3s_7_7_1_U12.top_mul_4ns_3s_7_7_1_Mul_DSP_1_U.ce  ? \mul_4ns_3s_7_7_1_U12.top_mul_4ns_3s_7_7_1_Mul_DSP_1_U.buff2  : \mul_4ns_3s_7_7_1_U12.top_mul_4ns_3s_7_7_1_Mul_DSP_1_U.buff3 ;
assign _0290_ = \mul_4ns_3s_7_7_1_U12.top_mul_4ns_3s_7_7_1_Mul_DSP_1_U.ce  ? \mul_4ns_3s_7_7_1_U12.top_mul_4ns_3s_7_7_1_Mul_DSP_1_U.buff1  : \mul_4ns_3s_7_7_1_U12.top_mul_4ns_3s_7_7_1_Mul_DSP_1_U.buff2 ;
assign _0289_ = \mul_4ns_3s_7_7_1_U12.top_mul_4ns_3s_7_7_1_Mul_DSP_1_U.ce  ? \mul_4ns_3s_7_7_1_U12.top_mul_4ns_3s_7_7_1_Mul_DSP_1_U.buff0  : \mul_4ns_3s_7_7_1_U12.top_mul_4ns_3s_7_7_1_Mul_DSP_1_U.buff1 ;
assign _0288_ = \mul_4ns_3s_7_7_1_U12.top_mul_4ns_3s_7_7_1_Mul_DSP_1_U.ce  ? \mul_4ns_3s_7_7_1_U12.top_mul_4ns_3s_7_7_1_Mul_DSP_1_U.tmp_product  : \mul_4ns_3s_7_7_1_U12.top_mul_4ns_3s_7_7_1_Mul_DSP_1_U.buff0 ;
assign _0287_ = \mul_4ns_3s_7_7_1_U12.top_mul_4ns_3s_7_7_1_Mul_DSP_1_U.ce  ? \mul_4ns_3s_7_7_1_U12.top_mul_4ns_3s_7_7_1_Mul_DSP_1_U.b  : \mul_4ns_3s_7_7_1_U12.top_mul_4ns_3s_7_7_1_Mul_DSP_1_U.b_reg0 ;
assign _0286_ = \mul_4ns_3s_7_7_1_U12.top_mul_4ns_3s_7_7_1_Mul_DSP_1_U.ce  ? \mul_4ns_3s_7_7_1_U12.top_mul_4ns_3s_7_7_1_Mul_DSP_1_U.a  : \mul_4ns_3s_7_7_1_U12.top_mul_4ns_3s_7_7_1_Mul_DSP_1_U.a_reg0 ;
assign \sub_17ns_17ns_17_2_1_U11.top_sub_17ns_17ns_17_2_1_Adder_8_U.bin_s0  = ~ \sub_17ns_17ns_17_2_1_U11.top_sub_17ns_17ns_17_2_1_Adder_8_U.b ;
always @(posedge \sub_17ns_17ns_17_2_1_U11.top_sub_17ns_17ns_17_2_1_Adder_8_U.clk )
\sub_17ns_17ns_17_2_1_U11.top_sub_17ns_17ns_17_2_1_Adder_8_U.bin_s1  <= _0294_;
always @(posedge \sub_17ns_17ns_17_2_1_U11.top_sub_17ns_17ns_17_2_1_Adder_8_U.clk )
\sub_17ns_17ns_17_2_1_U11.top_sub_17ns_17ns_17_2_1_Adder_8_U.ain_s1  <= _0293_;
always @(posedge \sub_17ns_17ns_17_2_1_U11.top_sub_17ns_17ns_17_2_1_Adder_8_U.clk )
\sub_17ns_17ns_17_2_1_U11.top_sub_17ns_17ns_17_2_1_Adder_8_U.sum_s1  <= _0296_;
always @(posedge \sub_17ns_17ns_17_2_1_U11.top_sub_17ns_17ns_17_2_1_Adder_8_U.clk )
\sub_17ns_17ns_17_2_1_U11.top_sub_17ns_17ns_17_2_1_Adder_8_U.carry_s1  <= _0295_;
assign _0294_ = \sub_17ns_17ns_17_2_1_U11.top_sub_17ns_17ns_17_2_1_Adder_8_U.ce  ? \sub_17ns_17ns_17_2_1_U11.top_sub_17ns_17ns_17_2_1_Adder_8_U.bin_s0 [16:8] : \sub_17ns_17ns_17_2_1_U11.top_sub_17ns_17ns_17_2_1_Adder_8_U.bin_s1 ;
assign _0293_ = \sub_17ns_17ns_17_2_1_U11.top_sub_17ns_17ns_17_2_1_Adder_8_U.ce  ? \sub_17ns_17ns_17_2_1_U11.top_sub_17ns_17ns_17_2_1_Adder_8_U.a [16:8] : \sub_17ns_17ns_17_2_1_U11.top_sub_17ns_17ns_17_2_1_Adder_8_U.ain_s1 ;
assign _0295_ = \sub_17ns_17ns_17_2_1_U11.top_sub_17ns_17ns_17_2_1_Adder_8_U.ce  ? \sub_17ns_17ns_17_2_1_U11.top_sub_17ns_17ns_17_2_1_Adder_8_U.facout_s1  : \sub_17ns_17ns_17_2_1_U11.top_sub_17ns_17ns_17_2_1_Adder_8_U.carry_s1 ;
assign _0296_ = \sub_17ns_17ns_17_2_1_U11.top_sub_17ns_17ns_17_2_1_Adder_8_U.ce  ? \sub_17ns_17ns_17_2_1_U11.top_sub_17ns_17ns_17_2_1_Adder_8_U.fas_s1  : \sub_17ns_17ns_17_2_1_U11.top_sub_17ns_17ns_17_2_1_Adder_8_U.sum_s1 ;
assign _0297_ = \sub_17ns_17ns_17_2_1_U11.top_sub_17ns_17ns_17_2_1_Adder_8_U.u1.a  + \sub_17ns_17ns_17_2_1_U11.top_sub_17ns_17ns_17_2_1_Adder_8_U.u1.b ;
assign { \sub_17ns_17ns_17_2_1_U11.top_sub_17ns_17ns_17_2_1_Adder_8_U.u1.cout , \sub_17ns_17ns_17_2_1_U11.top_sub_17ns_17ns_17_2_1_Adder_8_U.u1.s  } = _0297_ + \sub_17ns_17ns_17_2_1_U11.top_sub_17ns_17ns_17_2_1_Adder_8_U.u1.cin ;
assign _0298_ = \sub_17ns_17ns_17_2_1_U11.top_sub_17ns_17ns_17_2_1_Adder_8_U.u2.a  + \sub_17ns_17ns_17_2_1_U11.top_sub_17ns_17ns_17_2_1_Adder_8_U.u2.b ;
assign { \sub_17ns_17ns_17_2_1_U11.top_sub_17ns_17ns_17_2_1_Adder_8_U.u2.cout , \sub_17ns_17ns_17_2_1_U11.top_sub_17ns_17ns_17_2_1_Adder_8_U.u2.s  } = _0298_ + \sub_17ns_17ns_17_2_1_U11.top_sub_17ns_17ns_17_2_1_Adder_8_U.u2.cin ;
assign \sub_33ns_33ns_33_2_1_U14.top_sub_33ns_33ns_33_2_1_Adder_10_U.bin_s0  = ~ \sub_33ns_33ns_33_2_1_U14.top_sub_33ns_33ns_33_2_1_Adder_10_U.b ;
always @(posedge \sub_33ns_33ns_33_2_1_U14.top_sub_33ns_33ns_33_2_1_Adder_10_U.clk )
\sub_33ns_33ns_33_2_1_U14.top_sub_33ns_33ns_33_2_1_Adder_10_U.bin_s1  <= _0300_;
always @(posedge \sub_33ns_33ns_33_2_1_U14.top_sub_33ns_33ns_33_2_1_Adder_10_U.clk )
\sub_33ns_33ns_33_2_1_U14.top_sub_33ns_33ns_33_2_1_Adder_10_U.ain_s1  <= _0299_;
always @(posedge \sub_33ns_33ns_33_2_1_U14.top_sub_33ns_33ns_33_2_1_Adder_10_U.clk )
\sub_33ns_33ns_33_2_1_U14.top_sub_33ns_33ns_33_2_1_Adder_10_U.sum_s1  <= _0302_;
always @(posedge \sub_33ns_33ns_33_2_1_U14.top_sub_33ns_33ns_33_2_1_Adder_10_U.clk )
\sub_33ns_33ns_33_2_1_U14.top_sub_33ns_33ns_33_2_1_Adder_10_U.carry_s1  <= _0301_;
assign _0300_ = \sub_33ns_33ns_33_2_1_U14.top_sub_33ns_33ns_33_2_1_Adder_10_U.ce  ? \sub_33ns_33ns_33_2_1_U14.top_sub_33ns_33ns_33_2_1_Adder_10_U.bin_s0 [32:16] : \sub_33ns_33ns_33_2_1_U14.top_sub_33ns_33ns_33_2_1_Adder_10_U.bin_s1 ;
assign _0299_ = \sub_33ns_33ns_33_2_1_U14.top_sub_33ns_33ns_33_2_1_Adder_10_U.ce  ? \sub_33ns_33ns_33_2_1_U14.top_sub_33ns_33ns_33_2_1_Adder_10_U.a [32:16] : \sub_33ns_33ns_33_2_1_U14.top_sub_33ns_33ns_33_2_1_Adder_10_U.ain_s1 ;
assign _0301_ = \sub_33ns_33ns_33_2_1_U14.top_sub_33ns_33ns_33_2_1_Adder_10_U.ce  ? \sub_33ns_33ns_33_2_1_U14.top_sub_33ns_33ns_33_2_1_Adder_10_U.facout_s1  : \sub_33ns_33ns_33_2_1_U14.top_sub_33ns_33ns_33_2_1_Adder_10_U.carry_s1 ;
assign _0302_ = \sub_33ns_33ns_33_2_1_U14.top_sub_33ns_33ns_33_2_1_Adder_10_U.ce  ? \sub_33ns_33ns_33_2_1_U14.top_sub_33ns_33ns_33_2_1_Adder_10_U.fas_s1  : \sub_33ns_33ns_33_2_1_U14.top_sub_33ns_33ns_33_2_1_Adder_10_U.sum_s1 ;
assign _0303_ = \sub_33ns_33ns_33_2_1_U14.top_sub_33ns_33ns_33_2_1_Adder_10_U.u1.a  + \sub_33ns_33ns_33_2_1_U14.top_sub_33ns_33ns_33_2_1_Adder_10_U.u1.b ;
assign { \sub_33ns_33ns_33_2_1_U14.top_sub_33ns_33ns_33_2_1_Adder_10_U.u1.cout , \sub_33ns_33ns_33_2_1_U14.top_sub_33ns_33ns_33_2_1_Adder_10_U.u1.s  } = _0303_ + \sub_33ns_33ns_33_2_1_U14.top_sub_33ns_33ns_33_2_1_Adder_10_U.u1.cin ;
assign _0304_ = \sub_33ns_33ns_33_2_1_U14.top_sub_33ns_33ns_33_2_1_Adder_10_U.u2.a  + \sub_33ns_33ns_33_2_1_U14.top_sub_33ns_33ns_33_2_1_Adder_10_U.u2.b ;
assign { \sub_33ns_33ns_33_2_1_U14.top_sub_33ns_33ns_33_2_1_Adder_10_U.u2.cout , \sub_33ns_33ns_33_2_1_U14.top_sub_33ns_33ns_33_2_1_Adder_10_U.u2.s  } = _0304_ + \sub_33ns_33ns_33_2_1_U14.top_sub_33ns_33ns_33_2_1_Adder_10_U.u2.cin ;
assign \sub_8ns_8ns_8_2_1_U15.top_sub_8ns_8ns_8_2_1_Adder_11_U.bin_s0  = ~ \sub_8ns_8ns_8_2_1_U15.top_sub_8ns_8ns_8_2_1_Adder_11_U.b ;
always @(posedge \sub_8ns_8ns_8_2_1_U15.top_sub_8ns_8ns_8_2_1_Adder_11_U.clk )
\sub_8ns_8ns_8_2_1_U15.top_sub_8ns_8ns_8_2_1_Adder_11_U.bin_s1  <= _0306_;
always @(posedge \sub_8ns_8ns_8_2_1_U15.top_sub_8ns_8ns_8_2_1_Adder_11_U.clk )
\sub_8ns_8ns_8_2_1_U15.top_sub_8ns_8ns_8_2_1_Adder_11_U.ain_s1  <= _0305_;
always @(posedge \sub_8ns_8ns_8_2_1_U15.top_sub_8ns_8ns_8_2_1_Adder_11_U.clk )
\sub_8ns_8ns_8_2_1_U15.top_sub_8ns_8ns_8_2_1_Adder_11_U.sum_s1  <= _0308_;
always @(posedge \sub_8ns_8ns_8_2_1_U15.top_sub_8ns_8ns_8_2_1_Adder_11_U.clk )
\sub_8ns_8ns_8_2_1_U15.top_sub_8ns_8ns_8_2_1_Adder_11_U.carry_s1  <= _0307_;
assign _0306_ = \sub_8ns_8ns_8_2_1_U15.top_sub_8ns_8ns_8_2_1_Adder_11_U.ce  ? \sub_8ns_8ns_8_2_1_U15.top_sub_8ns_8ns_8_2_1_Adder_11_U.bin_s0 [7:4] : \sub_8ns_8ns_8_2_1_U15.top_sub_8ns_8ns_8_2_1_Adder_11_U.bin_s1 ;
assign _0305_ = \sub_8ns_8ns_8_2_1_U15.top_sub_8ns_8ns_8_2_1_Adder_11_U.ce  ? \sub_8ns_8ns_8_2_1_U15.top_sub_8ns_8ns_8_2_1_Adder_11_U.a [7:4] : \sub_8ns_8ns_8_2_1_U15.top_sub_8ns_8ns_8_2_1_Adder_11_U.ain_s1 ;
assign _0307_ = \sub_8ns_8ns_8_2_1_U15.top_sub_8ns_8ns_8_2_1_Adder_11_U.ce  ? \sub_8ns_8ns_8_2_1_U15.top_sub_8ns_8ns_8_2_1_Adder_11_U.facout_s1  : \sub_8ns_8ns_8_2_1_U15.top_sub_8ns_8ns_8_2_1_Adder_11_U.carry_s1 ;
assign _0308_ = \sub_8ns_8ns_8_2_1_U15.top_sub_8ns_8ns_8_2_1_Adder_11_U.ce  ? \sub_8ns_8ns_8_2_1_U15.top_sub_8ns_8ns_8_2_1_Adder_11_U.fas_s1  : \sub_8ns_8ns_8_2_1_U15.top_sub_8ns_8ns_8_2_1_Adder_11_U.sum_s1 ;
assign _0309_ = \sub_8ns_8ns_8_2_1_U15.top_sub_8ns_8ns_8_2_1_Adder_11_U.u1.a  + \sub_8ns_8ns_8_2_1_U15.top_sub_8ns_8ns_8_2_1_Adder_11_U.u1.b ;
assign { \sub_8ns_8ns_8_2_1_U15.top_sub_8ns_8ns_8_2_1_Adder_11_U.u1.cout , \sub_8ns_8ns_8_2_1_U15.top_sub_8ns_8ns_8_2_1_Adder_11_U.u1.s  } = _0309_ + \sub_8ns_8ns_8_2_1_U15.top_sub_8ns_8ns_8_2_1_Adder_11_U.u1.cin ;
assign _0310_ = \sub_8ns_8ns_8_2_1_U15.top_sub_8ns_8ns_8_2_1_Adder_11_U.u2.a  + \sub_8ns_8ns_8_2_1_U15.top_sub_8ns_8ns_8_2_1_Adder_11_U.u2.b ;
assign { \sub_8ns_8ns_8_2_1_U15.top_sub_8ns_8ns_8_2_1_Adder_11_U.u2.cout , \sub_8ns_8ns_8_2_1_U15.top_sub_8ns_8ns_8_2_1_Adder_11_U.u2.s  } = _0310_ + \sub_8ns_8ns_8_2_1_U15.top_sub_8ns_8ns_8_2_1_Adder_11_U.u2.cin ;
assign \sub_8s_8ns_8_2_1_U7.top_sub_8s_8ns_8_2_1_Adder_4_U.bin_s0  = ~ \sub_8s_8ns_8_2_1_U7.top_sub_8s_8ns_8_2_1_Adder_4_U.b ;
always @(posedge \sub_8s_8ns_8_2_1_U7.top_sub_8s_8ns_8_2_1_Adder_4_U.clk )
\sub_8s_8ns_8_2_1_U7.top_sub_8s_8ns_8_2_1_Adder_4_U.bin_s1  <= _0312_;
always @(posedge \sub_8s_8ns_8_2_1_U7.top_sub_8s_8ns_8_2_1_Adder_4_U.clk )
\sub_8s_8ns_8_2_1_U7.top_sub_8s_8ns_8_2_1_Adder_4_U.ain_s1  <= _0311_;
always @(posedge \sub_8s_8ns_8_2_1_U7.top_sub_8s_8ns_8_2_1_Adder_4_U.clk )
\sub_8s_8ns_8_2_1_U7.top_sub_8s_8ns_8_2_1_Adder_4_U.sum_s1  <= _0314_;
always @(posedge \sub_8s_8ns_8_2_1_U7.top_sub_8s_8ns_8_2_1_Adder_4_U.clk )
\sub_8s_8ns_8_2_1_U7.top_sub_8s_8ns_8_2_1_Adder_4_U.carry_s1  <= _0313_;
assign _0312_ = \sub_8s_8ns_8_2_1_U7.top_sub_8s_8ns_8_2_1_Adder_4_U.ce  ? \sub_8s_8ns_8_2_1_U7.top_sub_8s_8ns_8_2_1_Adder_4_U.bin_s0 [7:4] : \sub_8s_8ns_8_2_1_U7.top_sub_8s_8ns_8_2_1_Adder_4_U.bin_s1 ;
assign _0311_ = \sub_8s_8ns_8_2_1_U7.top_sub_8s_8ns_8_2_1_Adder_4_U.ce  ? \sub_8s_8ns_8_2_1_U7.top_sub_8s_8ns_8_2_1_Adder_4_U.a [7:4] : \sub_8s_8ns_8_2_1_U7.top_sub_8s_8ns_8_2_1_Adder_4_U.ain_s1 ;
assign _0313_ = \sub_8s_8ns_8_2_1_U7.top_sub_8s_8ns_8_2_1_Adder_4_U.ce  ? \sub_8s_8ns_8_2_1_U7.top_sub_8s_8ns_8_2_1_Adder_4_U.facout_s1  : \sub_8s_8ns_8_2_1_U7.top_sub_8s_8ns_8_2_1_Adder_4_U.carry_s1 ;
assign _0314_ = \sub_8s_8ns_8_2_1_U7.top_sub_8s_8ns_8_2_1_Adder_4_U.ce  ? \sub_8s_8ns_8_2_1_U7.top_sub_8s_8ns_8_2_1_Adder_4_U.fas_s1  : \sub_8s_8ns_8_2_1_U7.top_sub_8s_8ns_8_2_1_Adder_4_U.sum_s1 ;
assign _0315_ = \sub_8s_8ns_8_2_1_U7.top_sub_8s_8ns_8_2_1_Adder_4_U.u1.a  + \sub_8s_8ns_8_2_1_U7.top_sub_8s_8ns_8_2_1_Adder_4_U.u1.b ;
assign { \sub_8s_8ns_8_2_1_U7.top_sub_8s_8ns_8_2_1_Adder_4_U.u1.cout , \sub_8s_8ns_8_2_1_U7.top_sub_8s_8ns_8_2_1_Adder_4_U.u1.s  } = _0315_ + \sub_8s_8ns_8_2_1_U7.top_sub_8s_8ns_8_2_1_Adder_4_U.u1.cin ;
assign _0316_ = \sub_8s_8ns_8_2_1_U7.top_sub_8s_8ns_8_2_1_Adder_4_U.u2.a  + \sub_8s_8ns_8_2_1_U7.top_sub_8s_8ns_8_2_1_Adder_4_U.u2.b ;
assign { \sub_8s_8ns_8_2_1_U7.top_sub_8s_8ns_8_2_1_Adder_4_U.u2.cout , \sub_8s_8ns_8_2_1_U7.top_sub_8s_8ns_8_2_1_Adder_4_U.u2.s  } = _0316_ + \sub_8s_8ns_8_2_1_U7.top_sub_8s_8ns_8_2_1_Adder_4_U.u2.cin ;
assign _0317_ = | p_Result_s_22_reg_1855;
assign _0318_ = | p_Result_4_reg_2167;
assign _0319_ = | tmp_1_reg_2242;
assign _0320_ = | op_0[3:1];
assign _0321_ = p_Result_s_22_reg_1855 != 3'h7;
assign _0322_ = p_Result_4_reg_2167 != 3'h7;
assign _0323_ = tmp_1_reg_2242 != 27'h7ffffff;
assign _0324_ = ret_V_reg_1743 != 3'h7;
assign _0325_ = | op_11[12:0];
assign _0326_ = | trunc_ln851_4_reg_2432;
assign _0327_ = | trunc_ln851_5_reg_2361;
assign _0328_ = | trunc_ln851_reg_1999;
assign _0329_ = { op_3_V_reg_1917[3], op_3_V_reg_1917[3], op_3_V_reg_1917[3], op_3_V_reg_1917[3], op_3_V_reg_1917 } != { ret_V_18_reg_2075, 3'h0 };
assign or_ln340_1_fu_504_p2 = p_Result_27_reg_1832 | overflow_1_fu_490_p2;
assign or_ln340_2_fu_1049_p2 = overflow_2_fu_1043_p2 | and_ln786_reg_2194;
assign or_ln340_3_fu_1141_p2 = p_Result_34_reg_2148 | overflow_3_fu_1126_p2;
assign or_ln340_4_fu_1282_p2 = p_Result_36_reg_2223 | overflow_4_fu_1268_p2;
assign or_ln340_5_fu_1102_p2 = or_ln340_2_reg_2253 | neg_src_fu_1097_p2;
assign or_ln340_fu_321_p2 = p_Result_s_reg_1722 | overflow_fu_306_p2;
assign or_ln785_10_fu_1429_p2 = xor_ln785_9_fu_1424_p2 | p_Result_36_reg_2223;
assign or_ln785_11_fu_1402_p2 = and_ln785_13_fu_1398_p2 | and_ln340_5_fu_1394_p2;
assign or_ln785_1_fu_481_p2 = p_Result_28_reg_1848 | icmp_ln768_1_reg_1861;
assign or_ln785_2_fu_1033_p2 = xor_ln785_2_fu_1028_p2 | p_Result_33_reg_2068;
assign or_ln785_3_fu_1061_p2 = p_Result_35_reg_2160 | icmp_ln768_3_reg_2205;
assign or_ln785_4_fu_1197_p2 = p_Result_37_reg_2235 | icmp_ln768_4_reg_2269;
assign or_ln785_5_fu_367_p2 = xor_ln785_6_fu_362_p2 | p_Result_s_reg_1722;
assign or_ln785_6_fu_609_p2 = xor_ln785_7_fu_604_p2 | p_Result_27_reg_1832;
assign or_ln785_7_fu_592_p2 = and_ln785_4_fu_588_p2 | and_ln340_2_fu_584_p2;
assign or_ln785_8_fu_1210_p2 = p_Result_30_reg_1954 | and_ln785_6_fu_1206_p2;
assign or_ln785_9_fu_1236_p2 = xor_ln785_8_fu_1231_p2 | p_Result_34_reg_2148;
assign or_ln785_fu_289_p2 = p_Result_26_reg_1736 | icmp_ln768_reg_1751;
assign or_ln786_1_fu_499_p2 = xor_ln786_1_fu_494_p2 | icmp_ln786_1_reg_1866;
assign or_ln786_2_fu_1136_p2 = xor_ln786_2_fu_1131_p2 | icmp_ln786_2_reg_2210;
assign or_ln786_3_fu_1277_p2 = xor_ln786_3_fu_1272_p2 | icmp_ln786_3_reg_2274;
assign or_ln786_fu_316_p2 = xor_ln786_fu_311_p2 | icmp_ln786_reg_1767;
always @(posedge ap_clk)
rhs_4_reg_2120 <= _0097_;
always @(posedge ap_clk)
ret_V_22_reg_2457 <= _0086_;
always @(posedge ap_clk)
ret_V_17_cast_reg_2462 <= _0079_;
always @(posedge ap_clk)
select_ln340_reg_1778[3] <= _0104_;
always @(posedge ap_clk)
ret_V_16_reg_1783 <= _0078_;
always @(posedge ap_clk)
r_V_5_reg_1944 <= _0072_;
always @(posedge ap_clk)
p_Result_31_reg_1949 <= _0055_;
always @(posedge ap_clk)
p_Result_30_reg_1954 <= _0054_;
always @(posedge ap_clk)
p_Val2_5_reg_1961 <= _0069_;
always @(posedge ap_clk)
p_Result_11_reg_1966 <= _0049_;
always @(posedge ap_clk)
p_Result_32_reg_1971 <= _0056_;
always @(posedge ap_clk)
p_Result_1_reg_1976 <= _0050_;
always @(posedge ap_clk)
p_Result_3_reg_1981 <= _0062_;
always @(posedge ap_clk)
r_V_6_reg_1987 <= _0073_;
always @(posedge ap_clk)
ret_V_4_cast_reg_1992 <= _0092_;
always @(posedge ap_clk)
trunc_ln851_reg_1999 <= _0119_;
always @(posedge ap_clk)
or_ln785_1_reg_1872 <= _0043_;
always @(posedge ap_clk)
xor_ln785_1_reg_1878 <= _0121_;
always @(posedge ap_clk)
op_3_V_reg_1917 <= _0039_;
always @(posedge ap_clk)
op_24_V_reg_2516 <= _0038_;
always @(posedge ap_clk)
op_1_V_reg_1789[3] <= _0037_;
always @(posedge ap_clk)
r_V_reg_1796 <= _0075_;
always @(posedge ap_clk)
ret_V_8_reg_2417 <= _0095_;
always @(posedge ap_clk)
op_12_V_reg_2422 <= _0033_;
always @(posedge ap_clk)
select_ln353_reg_2427 <= _0106_;
always @(posedge ap_clk)
trunc_ln851_4_reg_2432 <= _0118_;
always @(posedge ap_clk)
r_V_7_reg_2366 <= _0074_;
always @(posedge ap_clk)
ret_V_10_cast_reg_2372 <= _0077_;
always @(posedge ap_clk)
sext_ln850_reg_2379 <= _0111_;
always @(posedge ap_clk)
p_Val2_14_reg_2386[7:2] <= _0067_;
always @(posedge ap_clk)
select_ln340_4_reg_2392 <= _0103_;
always @(posedge ap_clk)
sel_tmp51_reg_2397 <= _0099_;
always @(posedge ap_clk)
icmp_ln851_4_reg_2402 <= _0030_;
always @(posedge ap_clk)
ret_V_20_reg_2437 <= _0084_;
always @(posedge ap_clk)
icmp_ln851_3_reg_2452 <= _0029_;
always @(posedge ap_clk)
select_ln340_2_reg_2280 <= _0101_;
always @(posedge ap_clk)
p_Val2_10_reg_2285[15:2] <= _0066_;
always @(posedge ap_clk)
select_ln340_3_reg_2290[15:2] <= _0102_;
always @(posedge ap_clk)
icmp_ln851_2_reg_2305 <= _0028_;
always @(posedge ap_clk)
or_ln785_4_reg_2310 <= _0045_;
always @(posedge ap_clk)
xor_ln785_5_reg_2316 <= _0122_;
always @(posedge ap_clk)
p_Val2_6_reg_2062 <= _0070_;
always @(posedge ap_clk)
p_Result_33_reg_2068 <= _0057_;
always @(posedge ap_clk)
ret_V_18_reg_2075 <= _0080_;
always @(posedge ap_clk)
icmp_ln851_1_reg_2092 <= _0027_;
always @(posedge ap_clk)
or_ln785_reg_1761 <= _0046_;
always @(posedge ap_clk)
icmp_ln786_reg_1767 <= _0026_;
always @(posedge ap_clk)
ret_V_1_reg_1773 <= _0082_;
always @(posedge ap_clk)
p_Result_s_reg_1722 <= _0065_;
always @(posedge ap_clk)
p_Val2_s_reg_1730[3] <= _0071_;
always @(posedge ap_clk)
p_Result_26_reg_1736 <= _0051_;
always @(posedge ap_clk)
ret_V_reg_1743 <= _0096_;
always @(posedge ap_clk)
icmp_ln768_reg_1751 <= _0022_;
always @(posedge ap_clk)
trunc_ln1192_reg_1756 <= _0114_;
always @(posedge ap_clk)
or_ln340_2_reg_2253 <= _0041_;
always @(posedge ap_clk)
or_ln785_3_reg_2258 <= _0044_;
always @(posedge ap_clk)
select_ln850_4_reg_2264 <= _0109_;
always @(posedge ap_clk)
icmp_ln768_4_reg_2269 <= _0021_;
always @(posedge ap_clk)
icmp_ln786_3_reg_2274 <= _0025_;
always @(posedge ap_clk)
icmp_ln768_1_reg_1861 <= _0019_;
always @(posedge ap_clk)
icmp_ln786_1_reg_1866 <= _0023_;
always @(posedge ap_clk)
carry_1_reg_2141 <= _0017_;
always @(posedge ap_clk)
p_Result_34_reg_2148 <= _0058_;
always @(posedge ap_clk)
trunc_ln731_1_reg_2155 <= _0116_;
always @(posedge ap_clk)
p_Result_35_reg_2160 <= _0059_;
always @(posedge ap_clk)
p_Result_4_reg_2167 <= _0063_;
always @(posedge ap_clk)
deleted_zeros_reg_2188 <= _0018_;
always @(posedge ap_clk)
and_ln786_reg_2194 <= _0015_;
always @(posedge ap_clk)
icmp_ln768_3_reg_2205 <= _0020_;
always @(posedge ap_clk)
icmp_ln786_2_reg_2210 <= _0024_;
always @(posedge ap_clk)
ret_1_reg_2216 <= _0076_;
always @(posedge ap_clk)
p_Result_36_reg_2223 <= _0060_;
always @(posedge ap_clk)
trunc_ln731_2_reg_2230 <= _0117_;
always @(posedge ap_clk)
p_Result_37_reg_2235 <= _0061_;
always @(posedge ap_clk)
tmp_1_reg_2242 <= _0112_;
always @(posedge ap_clk)
op_19_V_reg_2248 <= _0036_;
always @(posedge ap_clk)
op_15_V_reg_2322 <= _0035_;
always @(posedge ap_clk)
op_13_V_reg_2328[15:2] <= _0034_;
always @(posedge ap_clk)
ret_V_21_reg_2333 <= _0085_;
always @(posedge ap_clk)
tmp_reg_2338 <= _0113_;
always @(posedge ap_clk)
or_ln786_3_reg_2343 <= _0048_;
always @(posedge ap_clk)
or_ln340_4_reg_2349 <= _0042_;
always @(posedge ap_clk)
and_ln786_2_reg_2355 <= _0014_;
always @(posedge ap_clk)
or_ln786_1_reg_1884 <= _0047_;
always @(posedge ap_clk)
or_ln340_1_reg_1890 <= _0040_;
always @(posedge ap_clk)
and_ln786_1_reg_1896 <= _0013_;
always @(posedge ap_clk)
add_ln69_reg_2583 <= _0011_;
always @(posedge ap_clk)
add_ln69_2_reg_2588 <= _0010_;
always @(posedge ap_clk)
ret_V_26_reg_2558 <= _0091_;
always @(posedge ap_clk)
add_ln69_1_reg_2563 <= _0009_;
always @(posedge ap_clk)
op_10_V_reg_2047 <= _0032_;
always @(posedge ap_clk)
add_ln691_reg_2057 <= _0008_;
always @(posedge ap_clk)
add_ln691_6_reg_2543 <= _0007_;
always @(posedge ap_clk)
add_ln691_5_reg_2501 <= _0006_;
always @(posedge ap_clk)
add_ln691_4_reg_2469 <= _0005_;
always @(posedge ap_clk)
add_ln691_3_reg_2407 <= _0004_;
always @(posedge ap_clk)
add_ln1192_1_reg_1826 <= _0003_;
always @(posedge ap_clk)
p_Result_27_reg_1832 <= _0052_;
always @(posedge ap_clk)
p_Val2_2_reg_1839 <= _0068_;
always @(posedge ap_clk)
p_Result_28_reg_1848 <= _0053_;
always @(posedge ap_clk)
p_Result_s_22_reg_1855 <= _0064_;
always @(posedge ap_clk)
trunc_ln213_reg_2014 <= _0115_;
always @(posedge ap_clk)
and_ln412_reg_2020 <= _0012_;
always @(posedge ap_clk)
Range2_all_ones_reg_2025 <= _0002_;
always @(posedge ap_clk)
Range1_all_ones_reg_2030 <= _0000_;
always @(posedge ap_clk)
Range1_all_zeros_reg_2037 <= _0001_;
always @(posedge ap_clk)
icmp_ln851_reg_2042 <= _0031_;
always @(posedge ap_clk)
ap_CS_fsm <= _0016_;
always @(posedge ap_clk)
p_Val2_s_reg_1730[2:0] <= 3'h0;
always @(posedge ap_clk)
select_ln340_reg_1778[2:0] <= 3'h0;
always @(posedge ap_clk)
op_1_V_reg_1789[2:0] <= 3'h0;
always @(posedge ap_clk)
p_Val2_10_reg_2285[1:0] <= 2'h0;
always @(posedge ap_clk)
select_ln340_3_reg_2290[1:0] <= 2'h0;
always @(posedge ap_clk)
op_13_V_reg_2328[1:0] <= 2'h0;
always @(posedge ap_clk)
trunc_ln851_5_reg_2361 <= 2'h0;
always @(posedge ap_clk)
p_Val2_14_reg_2386[1:0] <= 2'h0;
always @(posedge ap_clk)
sext_ln1116_reg_1923 <= _0110_;
always @(posedge ap_clk)
select_ln785_reg_1912 <= _0108_;
always @(posedge ap_clk)
select_ln785_3_reg_2412 <= _0107_;
always @(posedge ap_clk)
select_ln353_1_reg_2474 <= _0105_;
always @(posedge ap_clk)
select_ln340_1_reg_1902 <= _0100_;
always @(posedge ap_clk)
sel_tmp19_reg_1907 <= _0098_;
always @(posedge ap_clk)
ret_V_7_reg_2200 <= _0094_;
always @(posedge ap_clk)
ret_V_24_reg_2506 <= _0089_;
always @(posedge ap_clk)
ret_V_25_reg_2531 <= _0090_;
always @(posedge ap_clk)
ret_V_23_cast_reg_2536 <= _0087_;
always @(posedge ap_clk)
ret_V_23_reg_2489 <= _0088_;
always @(posedge ap_clk)
ret_V_20_cast_reg_2494 <= _0083_;
always @(posedge ap_clk)
xor_ln416_reg_2097 <= _0120_;
always @(posedge ap_clk)
ret_V_19_reg_2103 <= _0081_;
always @(posedge ap_clk)
ret_V_6_reg_2108 <= _0093_;
assign _0123_ = _0131_ ? 2'h2 : 2'h1;
assign _0330_ = ap_CS_fsm == 1'h1;
function [51:0] _0987_;
input [51:0] a;
input [2703:0] b;
input [51:0] s;
case (s)
52'b0000000000000000000000000000000000000000000000000001:
_0987_ = b[51:0];
52'b0000000000000000000000000000000000000000000000000010:
_0987_ = b[103:52];
52'b0000000000000000000000000000000000000000000000000100:
_0987_ = b[155:104];
52'b0000000000000000000000000000000000000000000000001000:
_0987_ = b[207:156];
52'b0000000000000000000000000000000000000000000000010000:
_0987_ = b[259:208];
52'b0000000000000000000000000000000000000000000000100000:
_0987_ = b[311:260];
52'b0000000000000000000000000000000000000000000001000000:
_0987_ = b[363:312];
52'b0000000000000000000000000000000000000000000010000000:
_0987_ = b[415:364];
52'b0000000000000000000000000000000000000000000100000000:
_0987_ = b[467:416];
52'b0000000000000000000000000000000000000000001000000000:
_0987_ = b[519:468];
52'b0000000000000000000000000000000000000000010000000000:
_0987_ = b[571:520];
52'b0000000000000000000000000000000000000000100000000000:
_0987_ = b[623:572];
52'b0000000000000000000000000000000000000001000000000000:
_0987_ = b[675:624];
52'b0000000000000000000000000000000000000010000000000000:
_0987_ = b[727:676];
52'b0000000000000000000000000000000000000100000000000000:
_0987_ = b[779:728];
52'b0000000000000000000000000000000000001000000000000000:
_0987_ = b[831:780];
52'b0000000000000000000000000000000000010000000000000000:
_0987_ = b[883:832];
52'b0000000000000000000000000000000000100000000000000000:
_0987_ = b[935:884];
52'b0000000000000000000000000000000001000000000000000000:
_0987_ = b[987:936];
52'b0000000000000000000000000000000010000000000000000000:
_0987_ = b[1039:988];
52'b0000000000000000000000000000000100000000000000000000:
_0987_ = b[1091:1040];
52'b0000000000000000000000000000001000000000000000000000:
_0987_ = b[1143:1092];
52'b0000000000000000000000000000010000000000000000000000:
_0987_ = b[1195:1144];
52'b0000000000000000000000000000100000000000000000000000:
_0987_ = b[1247:1196];
52'b0000000000000000000000000001000000000000000000000000:
_0987_ = b[1299:1248];
52'b0000000000000000000000000010000000000000000000000000:
_0987_ = b[1351:1300];
52'b0000000000000000000000000100000000000000000000000000:
_0987_ = b[1403:1352];
52'b0000000000000000000000001000000000000000000000000000:
_0987_ = b[1455:1404];
52'b0000000000000000000000010000000000000000000000000000:
_0987_ = b[1507:1456];
52'b0000000000000000000000100000000000000000000000000000:
_0987_ = b[1559:1508];
52'b0000000000000000000001000000000000000000000000000000:
_0987_ = b[1611:1560];
52'b0000000000000000000010000000000000000000000000000000:
_0987_ = b[1663:1612];
52'b0000000000000000000100000000000000000000000000000000:
_0987_ = b[1715:1664];
52'b0000000000000000001000000000000000000000000000000000:
_0987_ = b[1767:1716];
52'b0000000000000000010000000000000000000000000000000000:
_0987_ = b[1819:1768];
52'b0000000000000000100000000000000000000000000000000000:
_0987_ = b[1871:1820];
52'b0000000000000001000000000000000000000000000000000000:
_0987_ = b[1923:1872];
52'b0000000000000010000000000000000000000000000000000000:
_0987_ = b[1975:1924];
52'b0000000000000100000000000000000000000000000000000000:
_0987_ = b[2027:1976];
52'b0000000000001000000000000000000000000000000000000000:
_0987_ = b[2079:2028];
52'b0000000000010000000000000000000000000000000000000000:
_0987_ = b[2131:2080];
52'b0000000000100000000000000000000000000000000000000000:
_0987_ = b[2183:2132];
52'b0000000001000000000000000000000000000000000000000000:
_0987_ = b[2235:2184];
52'b0000000010000000000000000000000000000000000000000000:
_0987_ = b[2287:2236];
52'b0000000100000000000000000000000000000000000000000000:
_0987_ = b[2339:2288];
52'b0000001000000000000000000000000000000000000000000000:
_0987_ = b[2391:2340];
52'b0000010000000000000000000000000000000000000000000000:
_0987_ = b[2443:2392];
52'b0000100000000000000000000000000000000000000000000000:
_0987_ = b[2495:2444];
52'b0001000000000000000000000000000000000000000000000000:
_0987_ = b[2547:2496];
52'b0010000000000000000000000000000000000000000000000000:
_0987_ = b[2599:2548];
52'b0100000000000000000000000000000000000000000000000000:
_0987_ = b[2651:2600];
52'b1000000000000000000000000000000000000000000000000000:
_0987_ = b[2703:2652];
52'b0000000000000000000000000000000000000000000000000000:
_0987_ = a;
default:
_0987_ = 52'bx;
endcase
endfunction
assign ap_NS_fsm = _0987_(52'hxxxxxxxxxxxxx, { 50'h0000000000000, _0123_, 2652'h000000000000400000000000080000000000010000000000002000000000000400000000000080000000000010000000000002000000000000400000000000080000000000010000000000002000000000000400000000000080000000000010000000000002000000000000400000000000080000000000010000000000002000000000000400000000000080000000000010000000000002000000000000400000000000080000000000010000000000002000000000000400000000000080000000000010000000000002000000000000400000000000080000000000010000000000002000000000000400000000000080000000000010000000000002000000000000400000000000080000000000010000000000002000000000000400000000000080000000000010000000000002000000000000400000000000080000000000000000000000001 }, { _0330_, _0381_, _0380_, _0379_, _0378_, _0377_, _0376_, _0375_, _0374_, _0373_, _0372_, _0371_, _0370_, _0369_, _0368_, _0367_, _0366_, _0365_, _0364_, _0363_, _0362_, _0361_, _0360_, _0359_, _0358_, _0357_, _0356_, _0355_, _0354_, _0353_, _0352_, _0351_, _0350_, _0349_, _0348_, _0347_, _0346_, _0345_, _0344_, _0343_, _0342_, _0341_, _0340_, _0339_, _0338_, _0337_, _0336_, _0335_, _0334_, _0333_, _0332_, _0331_ });
assign _0331_ = ap_CS_fsm == 52'h8000000000000;
assign _0332_ = ap_CS_fsm == 51'h4000000000000;
assign _0333_ = ap_CS_fsm == 50'h2000000000000;
assign _0334_ = ap_CS_fsm == 49'h1000000000000;
assign _0335_ = ap_CS_fsm == 48'h800000000000;
assign _0336_ = ap_CS_fsm == 47'h400000000000;
assign _0337_ = ap_CS_fsm == 46'h200000000000;
assign _0338_ = ap_CS_fsm == 45'h100000000000;
assign _0339_ = ap_CS_fsm == 44'h80000000000;
assign _0340_ = ap_CS_fsm == 43'h40000000000;
assign _0341_ = ap_CS_fsm == 42'h20000000000;
assign _0342_ = ap_CS_fsm == 41'h10000000000;
assign _0343_ = ap_CS_fsm == 40'h8000000000;
assign _0344_ = ap_CS_fsm == 39'h4000000000;
assign _0345_ = ap_CS_fsm == 38'h2000000000;
assign _0346_ = ap_CS_fsm == 37'h1000000000;
assign _0347_ = ap_CS_fsm == 36'h800000000;
assign _0348_ = ap_CS_fsm == 35'h400000000;
assign _0349_ = ap_CS_fsm == 34'h200000000;
assign _0350_ = ap_CS_fsm == 33'h100000000;
assign _0351_ = ap_CS_fsm == 32'd2147483648;
assign _0352_ = ap_CS_fsm == 31'h40000000;
assign _0353_ = ap_CS_fsm == 30'h20000000;
assign _0354_ = ap_CS_fsm == 29'h10000000;
assign _0355_ = ap_CS_fsm == 28'h8000000;
assign _0356_ = ap_CS_fsm == 27'h4000000;
assign _0357_ = ap_CS_fsm == 26'h2000000;
assign _0358_ = ap_CS_fsm == 25'h1000000;
assign _0359_ = ap_CS_fsm == 24'h800000;
assign _0360_ = ap_CS_fsm == 23'h400000;
assign _0361_ = ap_CS_fsm == 22'h200000;
assign _0362_ = ap_CS_fsm == 21'h100000;
assign _0363_ = ap_CS_fsm == 20'h80000;
assign _0364_ = ap_CS_fsm == 19'h40000;
assign _0365_ = ap_CS_fsm == 18'h20000;
assign _0366_ = ap_CS_fsm == 17'h10000;
assign _0367_ = ap_CS_fsm == 16'h8000;
assign _0368_ = ap_CS_fsm == 15'h4000;
assign _0369_ = ap_CS_fsm == 14'h2000;
assign _0370_ = ap_CS_fsm == 13'h1000;
assign _0371_ = ap_CS_fsm == 12'h800;
assign _0372_ = ap_CS_fsm == 11'h400;
assign _0373_ = ap_CS_fsm == 10'h200;
assign _0374_ = ap_CS_fsm == 9'h100;
assign _0375_ = ap_CS_fsm == 8'h80;
assign _0376_ = ap_CS_fsm == 7'h40;
assign _0377_ = ap_CS_fsm == 6'h20;
assign _0378_ = ap_CS_fsm == 5'h10;
assign _0379_ = ap_CS_fsm == 4'h8;
assign _0380_ = ap_CS_fsm == 3'h4;
assign _0381_ = ap_CS_fsm == 2'h2;
assign op_29_ap_vld = ap_CS_fsm[51] ? 1'h1 : 1'h0;
assign ap_idle = _0130_ ? 1'h1 : 1'h0;
assign _0110_ = ap_CS_fsm[12] ? { ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783 } : sext_ln1116_reg_1923;
assign _0108_ = _0129_ ? select_ln785_fu_619_p3 : select_ln785_reg_1912;
assign _0107_ = _0128_ ? select_ln785_3_fu_1439_p3 : select_ln785_3_reg_2412;
assign _0105_ = ap_CS_fsm[35] ? select_ln353_1_fu_1548_p3 : select_ln353_1_reg_2474;
assign _0098_ = ap_CS_fsm[9] ? sel_tmp19_fu_598_p2 : sel_tmp19_reg_1907;
assign _0100_ = ap_CS_fsm[9] ? select_ln340_1_fu_577_p3 : select_ln340_1_reg_1902;
assign _0094_ = _0127_ ? grp_fu_899_p2 : ret_V_7_reg_2200;
assign _0089_ = ap_CS_fsm[40] ? ret_V_24_fu_1602_p3 : ret_V_24_reg_2506;
assign _0087_ = ap_CS_fsm[44] ? grp_fu_1631_p2[32:1] : ret_V_23_cast_reg_2536;
assign _0090_ = ap_CS_fsm[44] ? grp_fu_1631_p2 : ret_V_25_reg_2531;
assign _0083_ = ap_CS_fsm[37] ? grp_fu_1569_p2[33:2] : ret_V_20_cast_reg_2494;
assign _0088_ = ap_CS_fsm[37] ? grp_fu_1569_p2 : ret_V_23_reg_2489;
assign _0097_ = ap_CS_fsm[22] ? rhs_4_fu_868_p2 : rhs_4_reg_2120;
assign _0093_ = ap_CS_fsm[22] ? grp_fu_820_p2[12:3] : ret_V_6_reg_2108;
assign _0081_ = ap_CS_fsm[22] ? grp_fu_820_p2 : ret_V_19_reg_2103;
assign _0120_ = ap_CS_fsm[22] ? xor_ln416_fu_836_p2 : xor_ln416_reg_2097;
assign _0079_ = ap_CS_fsm[32] ? grp_fu_1510_p2[33:2] : ret_V_17_cast_reg_2462;
assign _0086_ = ap_CS_fsm[32] ? grp_fu_1510_p2 : ret_V_22_reg_2457;
assign _0078_ = ap_CS_fsm[2] ? ret_V_16_fu_351_p3 : ret_V_16_reg_1783;
assign _0104_ = ap_CS_fsm[2] ? select_ln340_fu_338_p3[3] : select_ln340_reg_1778[3];
assign _0119_ = ap_CS_fsm[18] ? grp_fu_650_p2[2:0] : trunc_ln851_reg_1999;
assign _0092_ = ap_CS_fsm[18] ? grp_fu_650_p2[6:3] : ret_V_4_cast_reg_1992;
assign _0073_ = ap_CS_fsm[18] ? grp_fu_650_p2 : r_V_6_reg_1987;
assign _0062_ = ap_CS_fsm[18] ? grp_fu_641_p2[35:3] : p_Result_3_reg_1981;
assign _0050_ = ap_CS_fsm[18] ? grp_fu_641_p2[35:4] : p_Result_1_reg_1976;
assign _0056_ = ap_CS_fsm[18] ? grp_fu_641_p2[2] : p_Result_32_reg_1971;
assign _0049_ = ap_CS_fsm[18] ? grp_fu_641_p2[1] : p_Result_11_reg_1966;
assign _0069_ = ap_CS_fsm[18] ? grp_fu_641_p2[2:1] : p_Val2_5_reg_1961;
assign _0054_ = ap_CS_fsm[18] ? grp_fu_641_p2[35] : p_Result_30_reg_1954;
assign _0055_ = ap_CS_fsm[18] ? grp_fu_641_p2[0] : p_Result_31_reg_1949;
assign _0072_ = ap_CS_fsm[18] ? grp_fu_641_p2 : r_V_5_reg_1944;
assign _0121_ = ap_CS_fsm[7] ? xor_ln785_1_fu_485_p2 : xor_ln785_1_reg_1878;
assign _0043_ = ap_CS_fsm[7] ? or_ln785_1_fu_481_p2 : or_ln785_1_reg_1872;
assign _0039_ = ap_CS_fsm[11] ? op_3_V_fu_625_p3 : op_3_V_reg_1917;
assign _0038_ = ap_CS_fsm[42] ? grp_fu_1612_p2 : op_24_V_reg_2516;
assign _0075_ = ap_CS_fsm[3] ? op_1_V_fu_383_p3[3:1] : r_V_reg_1796;
assign _0037_ = ap_CS_fsm[3] ? op_1_V_fu_383_p3[3] : op_1_V_reg_1789[3];
assign _0118_ = ap_CS_fsm[30] ? op_12_V_fu_1452_p3[1:0] : trunc_ln851_4_reg_2432;
assign _0106_ = ap_CS_fsm[30] ? select_ln353_fu_1462_p3 : select_ln353_reg_2427;
assign _0033_ = ap_CS_fsm[30] ? op_12_V_fu_1452_p3 : op_12_V_reg_2422;
assign _0095_ = ap_CS_fsm[30] ? grp_fu_1419_p2 : ret_V_8_reg_2417;
assign _0030_ = ap_CS_fsm[28] ? icmp_ln851_4_fu_1414_p2 : icmp_ln851_4_reg_2402;
assign _0099_ = ap_CS_fsm[28] ? sel_tmp51_fu_1408_p2 : sel_tmp51_reg_2397;
assign _0103_ = ap_CS_fsm[28] ? select_ln340_4_fu_1386_p3 : select_ln340_4_reg_2392;
assign _0067_ = ap_CS_fsm[28] ? trunc_ln731_2_reg_2230 : p_Val2_14_reg_2386[7:2];
assign _0111_ = ap_CS_fsm[28] ? { tmp_reg_2338[10], tmp_reg_2338 } : sext_ln850_reg_2379;
assign _0077_ = ap_CS_fsm[28] ? grp_fu_889_p2[4:1] : ret_V_10_cast_reg_2372;
assign _0074_ = ap_CS_fsm[28] ? grp_fu_889_p2 : r_V_7_reg_2366;
assign _0029_ = ap_CS_fsm[31] ? icmp_ln851_3_fu_1516_p2 : icmp_ln851_3_reg_2452;
assign _0084_ = ap_CS_fsm[31] ? ret_V_20_fu_1489_p3 : ret_V_20_reg_2437;
assign _0122_ = ap_CS_fsm[26] ? xor_ln785_5_fu_1201_p2 : xor_ln785_5_reg_2316;
assign _0045_ = ap_CS_fsm[26] ? or_ln785_4_fu_1197_p2 : or_ln785_4_reg_2310;
assign _0028_ = ap_CS_fsm[26] ? icmp_ln851_2_fu_1191_p2 : icmp_ln851_2_reg_2305;
assign _0102_ = ap_CS_fsm[26] ? select_ln340_3_fu_1158_p3[15:2] : select_ln340_3_reg_2290[15:2];
assign _0066_ = ap_CS_fsm[26] ? trunc_ln731_1_reg_2155 : p_Val2_10_reg_2285[15:2];
assign _0101_ = ap_CS_fsm[26] ? select_ln340_2_fu_1107_p3 : select_ln340_2_reg_2280;
assign _0027_ = ap_CS_fsm[21] ? icmp_ln851_1_fu_830_p2 : icmp_ln851_1_reg_2092;
assign _0080_ = ap_CS_fsm[21] ? ret_V_18_fu_798_p3 : ret_V_18_reg_2075;
assign _0057_ = ap_CS_fsm[21] ? grp_fu_773_p2[1] : p_Result_33_reg_2068;
assign _0070_ = ap_CS_fsm[21] ? grp_fu_773_p2 : p_Val2_6_reg_2062;
assign _0082_ = ap_CS_fsm[1] ? grp_fu_279_p2 : ret_V_1_reg_1773;
assign _0026_ = ap_CS_fsm[1] ? icmp_ln786_fu_293_p2 : icmp_ln786_reg_1767;
assign _0046_ = ap_CS_fsm[1] ? or_ln785_fu_289_p2 : or_ln785_reg_1761;
assign _0114_ = ap_CS_fsm[0] ? op_0[2:0] : trunc_ln1192_reg_1756;
assign _0022_ = ap_CS_fsm[0] ? icmp_ln768_fu_273_p2 : icmp_ln768_reg_1751;
assign _0096_ = ap_CS_fsm[0] ? op_0[3:1] : ret_V_reg_1743;
assign _0051_ = ap_CS_fsm[0] ? p_Result_26_fu_257_p2 : p_Result_26_reg_1736;
assign _0071_ = ap_CS_fsm[0] ? op_0[0] : p_Val2_s_reg_1730[3];
assign _0065_ = ap_CS_fsm[0] ? op_0[3] : p_Result_s_reg_1722;
assign _0025_ = ap_CS_fsm[25] ? icmp_ln786_3_fu_1082_p2 : icmp_ln786_3_reg_2274;
assign _0021_ = ap_CS_fsm[25] ? icmp_ln768_4_fu_1077_p2 : icmp_ln768_4_reg_2269;
assign _0109_ = ap_CS_fsm[25] ? select_ln850_4_fu_1070_p3 : select_ln850_4_reg_2264;
assign _0044_ = ap_CS_fsm[25] ? or_ln785_3_fu_1061_p2 : or_ln785_3_reg_2258;
assign _0041_ = ap_CS_fsm[25] ? or_ln340_2_fu_1049_p2 : or_ln340_2_reg_2253;
assign _0023_ = ap_CS_fsm[6] ? icmp_ln786_1_fu_476_p2 : icmp_ln786_1_reg_1866;
assign _0019_ = ap_CS_fsm[6] ? icmp_ln768_1_fu_471_p2 : icmp_ln768_1_reg_1861;
assign _0063_ = ap_CS_fsm[23] ? grp_fu_880_p2[16:14] : p_Result_4_reg_2167;
assign _0059_ = ap_CS_fsm[23] ? grp_fu_880_p2[13] : p_Result_35_reg_2160;
assign _0116_ = ap_CS_fsm[23] ? grp_fu_880_p2[13:0] : trunc_ln731_1_reg_2155;
assign _0058_ = ap_CS_fsm[23] ? grp_fu_880_p2[16] : p_Result_34_reg_2148;
assign _0017_ = ap_CS_fsm[23] ? carry_1_fu_895_p2 : carry_1_reg_2141;
assign _0036_ = ap_CS_fsm[24] ? grp_fu_949_p2 : op_19_V_reg_2248;
assign _0112_ = ap_CS_fsm[24] ? grp_fu_940_p2[32:6] : tmp_1_reg_2242;
assign _0061_ = ap_CS_fsm[24] ? grp_fu_940_p2[5] : p_Result_37_reg_2235;
assign _0117_ = ap_CS_fsm[24] ? grp_fu_940_p2[5:0] : trunc_ln731_2_reg_2230;
assign _0060_ = ap_CS_fsm[24] ? grp_fu_940_p2[32] : p_Result_36_reg_2223;
assign _0076_ = ap_CS_fsm[24] ? grp_fu_940_p2 : ret_1_reg_2216;
assign _0024_ = ap_CS_fsm[24] ? icmp_ln786_2_fu_993_p2 : icmp_ln786_2_reg_2210;
assign _0020_ = ap_CS_fsm[24] ? icmp_ln768_3_fu_988_p2 : icmp_ln768_3_reg_2205;
assign _0015_ = ap_CS_fsm[24] ? and_ln786_fu_983_p2 : and_ln786_reg_2194;
assign _0018_ = ap_CS_fsm[24] ? deleted_zeros_fu_954_p3 : deleted_zeros_reg_2188;
assign _0014_ = ap_CS_fsm[27] ? and_ln786_2_fu_1292_p2 : and_ln786_2_reg_2355;
assign _0042_ = ap_CS_fsm[27] ? or_ln340_4_fu_1282_p2 : or_ln340_4_reg_2349;
assign _0048_ = ap_CS_fsm[27] ? or_ln786_3_fu_1277_p2 : or_ln786_3_reg_2343;
assign _0113_ = ap_CS_fsm[27] ? grp_fu_1181_p2[23:13] : tmp_reg_2338;
assign _0085_ = ap_CS_fsm[27] ? grp_fu_1181_p2 : ret_V_21_reg_2333;
assign _0034_ = ap_CS_fsm[27] ? op_13_V_fu_1252_p3[15:2] : op_13_V_reg_2328[15:2];
assign _0035_ = ap_CS_fsm[27] ? op_15_V_fu_1220_p3 : op_15_V_reg_2322;
assign _0013_ = ap_CS_fsm[8] ? and_ln786_1_fu_514_p2 : and_ln786_1_reg_1896;
assign _0040_ = ap_CS_fsm[8] ? or_ln340_1_fu_504_p2 : or_ln340_1_reg_1890;
assign _0047_ = ap_CS_fsm[8] ? or_ln786_1_fu_499_p2 : or_ln786_1_reg_1884;
assign _0010_ = ap_CS_fsm[49] ? grp_fu_1700_p2 : add_ln69_2_reg_2588;
assign _0011_ = ap_CS_fsm[49] ? grp_fu_1692_p2 : add_ln69_reg_2583;
assign _0009_ = ap_CS_fsm[47] ? grp_fu_1659_p2 : add_ln69_1_reg_2563;
assign _0091_ = ap_CS_fsm[47] ? ret_V_26_fu_1681_p3 : ret_V_26_reg_2558;
assign _0008_ = ap_CS_fsm[20] ? grp_fu_765_p2 : add_ln691_reg_2057;
assign _0032_ = ap_CS_fsm[20] ? grp_fu_735_p2 : op_10_V_reg_2047;
assign _0007_ = ap_CS_fsm[46] ? grp_fu_1647_p2 : add_ln691_6_reg_2543;
assign _0006_ = _0126_ ? grp_fu_1585_p2 : add_ln691_5_reg_2501;
assign _0005_ = _0125_ ? grp_fu_1531_p2 : add_ln691_4_reg_2469;
assign _0004_ = _0124_ ? grp_fu_1314_p2 : add_ln691_3_reg_2407;
assign _0064_ = ap_CS_fsm[5] ? grp_fu_428_p2[6:4] : p_Result_s_22_reg_1855;
assign _0053_ = ap_CS_fsm[5] ? grp_fu_440_p2[3] : p_Result_28_reg_1848;
assign _0068_ = ap_CS_fsm[5] ? grp_fu_440_p2 : p_Val2_2_reg_1839;
assign _0052_ = ap_CS_fsm[5] ? grp_fu_428_p2[6] : p_Result_27_reg_1832;
assign _0003_ = ap_CS_fsm[5] ? grp_fu_434_p2 : add_ln1192_1_reg_1826;
assign _0031_ = ap_CS_fsm[19] ? icmp_ln851_fu_760_p2 : icmp_ln851_reg_2042;
assign _0001_ = ap_CS_fsm[19] ? Range1_all_zeros_fu_755_p2 : Range1_all_zeros_reg_2037;
assign _0000_ = ap_CS_fsm[19] ? Range1_all_ones_fu_750_p2 : Range1_all_ones_reg_2030;
assign _0002_ = ap_CS_fsm[19] ? Range2_all_ones_fu_745_p2 : Range2_all_ones_reg_2025;
assign _0012_ = ap_CS_fsm[19] ? and_ln412_fu_741_p2 : and_ln412_reg_2020;
assign _0115_ = ap_CS_fsm[19] ? op_7[7:0] : trunc_ln213_reg_2014;
assign _0016_ = ap_rst ? 52'h0000000000001 : ap_NS_fsm;
assign Range1_all_ones_fu_750_p2 = _0136_ ? 1'h1 : 1'h0;
assign Range1_all_zeros_fu_755_p2 = _0137_ ? 1'h1 : 1'h0;
assign Range2_all_ones_fu_745_p2 = _0138_ ? 1'h1 : 1'h0;
assign deleted_ones_fu_977_p3 = carry_1_reg_2141 ? and_ln780_fu_972_p2 : Range1_all_ones_reg_2030;
assign deleted_zeros_fu_954_p3 = carry_1_reg_2141 ? Range1_all_ones_reg_2030 : Range1_all_zeros_reg_2037;
assign icmp_ln768_1_fu_471_p2 = _0317_ ? 1'h1 : 1'h0;
assign icmp_ln768_3_fu_988_p2 = _0318_ ? 1'h1 : 1'h0;
assign icmp_ln768_4_fu_1077_p2 = _0319_ ? 1'h1 : 1'h0;
assign icmp_ln768_fu_273_p2 = _0320_ ? 1'h1 : 1'h0;
assign icmp_ln786_1_fu_476_p2 = _0321_ ? 1'h1 : 1'h0;
assign icmp_ln786_2_fu_993_p2 = _0322_ ? 1'h1 : 1'h0;
assign icmp_ln786_3_fu_1082_p2 = _0323_ ? 1'h1 : 1'h0;
assign icmp_ln786_fu_293_p2 = _0324_ ? 1'h1 : 1'h0;
assign icmp_ln851_1_fu_830_p2 = _0139_ ? 1'h1 : 1'h0;
assign icmp_ln851_2_fu_1191_p2 = _0325_ ? 1'h1 : 1'h0;
assign icmp_ln851_3_fu_1516_p2 = _0326_ ? 1'h1 : 1'h0;
assign icmp_ln851_4_fu_1414_p2 = _0327_ ? 1'h1 : 1'h0;
assign icmp_ln851_fu_760_p2 = _0328_ ? 1'h1 : 1'h0;
assign op_12_V_fu_1452_p3 = sel_tmp51_reg_2397 ? p_Val2_14_reg_2386 : select_ln785_3_reg_2412;
assign op_13_V_fu_1252_p3 = and_ln785_10_fu_1247_p2 ? p_Val2_10_reg_2285 : select_ln340_3_reg_2290;
assign op_15_V_fu_1220_p3 = and_ln785_7_fu_1215_p2 ? p_Val2_6_reg_2062 : select_ln340_2_reg_2280;
assign op_1_V_fu_383_p3 = and_ln785_1_fu_378_p2 ? p_Val2_s_reg_1730 : select_ln340_reg_1778;
assign op_3_V_fu_625_p3 = sel_tmp19_reg_1907 ? p_Val2_2_reg_1839 : select_ln785_reg_1912;
assign p_Result_26_fu_257_p2 = op_0[0] ? 1'h1 : 1'h0;
assign ret_V_16_fu_351_p3 = p_Result_s_reg_1722 ? select_ln850_fu_345_p3 : ret_V_reg_1743;
assign ret_V_18_fu_798_p3 = r_V_6_reg_1987[35] ? select_ln850_1_fu_793_p3 : ret_V_4_cast_reg_1992;
assign ret_V_20_fu_1489_p3 = r_V_7_reg_2366[6] ? select_ln850_2_fu_1483_p3 : ret_V_10_cast_reg_2372;
assign ret_V_24_fu_1602_p3 = ret_V_23_reg_2489[34] ? select_ln850_6_fu_1597_p3 : ret_V_20_cast_reg_2494;
assign ret_V_26_fu_1681_p3 = ret_V_25_reg_2531[33] ? select_ln850_7_fu_1675_p3 : ret_V_23_cast_reg_2536;
assign rhs_4_fu_868_p2 = _0329_ ? 1'h1 : 1'h0;
assign select_ln340_1_fu_577_p3 = and_ln340_1_fu_572_p2 ? p_Val2_2_reg_1839 : { add_ln1192_1_reg_1826[4], p_Val2_3_fu_552_p2 };
assign select_ln340_2_fu_1107_p3 = or_ln340_5_fu_1102_p2 ? 2'h0 : p_Val2_6_reg_2062;
assign select_ln340_3_fu_1158_p3 = and_ln340_3_fu_1152_p2 ? { trunc_ln731_1_reg_2155, 2'h0 } : 16'h0000;
assign select_ln340_4_fu_1386_p3 = and_ln340_4_fu_1381_p2 ? { trunc_ln731_2_reg_2230, 2'h0 } : { ret_1_reg_2216[6], p_Val2_15_fu_1360_p2 };
assign select_ln340_fu_338_p3 = and_ln340_fu_332_p2 ? p_Val2_s_reg_1730 : 4'h0;
assign select_ln353_1_fu_1548_p3 = ret_V_22_reg_2457[34] ? select_ln850_8_fu_1543_p3 : ret_V_17_cast_reg_2462;
assign select_ln353_fu_1462_p3 = ret_V_21_reg_2333[23] ? select_ln850_5_fu_1457_p3 : sext_ln850_reg_2379;
assign select_ln785_3_fu_1439_p3 = and_ln785_12_fu_1434_p2 ? p_Val2_14_reg_2386 : select_ln340_4_reg_2392;
assign select_ln785_fu_619_p3 = and_ln785_3_fu_614_p2 ? p_Val2_2_reg_1839 : select_ln340_1_reg_1902;
assign select_ln850_1_fu_793_p3 = icmp_ln851_reg_2042 ? add_ln691_reg_2057 : ret_V_4_cast_reg_1992;
assign select_ln850_2_fu_1483_p3 = r_V_7_reg_2366[0] ? ret_V_8_reg_2417 : ret_V_10_cast_reg_2372;
assign select_ln850_3_fu_1065_p3 = icmp_ln851_1_reg_2092 ? ret_V_6_reg_2108 : ret_V_7_reg_2200;
assign select_ln850_4_fu_1070_p3 = ret_V_19_reg_2103[12] ? select_ln850_3_fu_1065_p3 : ret_V_6_reg_2108;
assign select_ln850_5_fu_1457_p3 = icmp_ln851_2_reg_2305 ? add_ln691_3_reg_2407 : sext_ln850_reg_2379;
assign select_ln850_6_fu_1597_p3 = icmp_ln851_4_reg_2402 ? add_ln691_5_reg_2501 : ret_V_20_cast_reg_2494;
assign select_ln850_7_fu_1675_p3 = op_15_V_reg_2322[0] ? add_ln691_6_reg_2543 : ret_V_23_cast_reg_2536;
assign select_ln850_8_fu_1543_p3 = icmp_ln851_3_reg_2452 ? add_ln691_4_reg_2469 : ret_V_17_cast_reg_2462;
assign select_ln850_fu_345_p3 = op_0[0] ? ret_V_1_reg_1773 : ret_V_reg_1743;
assign xor_ln365_2_fu_1348_p2 = ret_1_reg_2216[5] ^ ret_1_reg_2216[6];
assign xor_ln365_fu_540_p2 = p_Val2_2_reg_1839[3] ^ add_ln1192_1_reg_1826[4];
assign ap_CS_fsm_state1 = ap_CS_fsm[0];
assign ap_CS_fsm_state10 = ap_CS_fsm[9];
assign ap_CS_fsm_state11 = ap_CS_fsm[10];
assign ap_CS_fsm_state12 = ap_CS_fsm[11];
assign ap_CS_fsm_state13 = ap_CS_fsm[12];
assign ap_CS_fsm_state19 = ap_CS_fsm[18];
assign ap_CS_fsm_state2 = ap_CS_fsm[1];
assign ap_CS_fsm_state20 = ap_CS_fsm[19];
assign ap_CS_fsm_state21 = ap_CS_fsm[20];
assign ap_CS_fsm_state22 = ap_CS_fsm[21];
assign ap_CS_fsm_state23 = ap_CS_fsm[22];
assign ap_CS_fsm_state24 = ap_CS_fsm[23];
assign ap_CS_fsm_state25 = ap_CS_fsm[24];
assign ap_CS_fsm_state26 = ap_CS_fsm[25];
assign ap_CS_fsm_state27 = ap_CS_fsm[26];
assign ap_CS_fsm_state28 = ap_CS_fsm[27];
assign ap_CS_fsm_state29 = ap_CS_fsm[28];
assign ap_CS_fsm_state3 = ap_CS_fsm[2];
assign ap_CS_fsm_state30 = ap_CS_fsm[29];
assign ap_CS_fsm_state31 = ap_CS_fsm[30];
assign ap_CS_fsm_state32 = ap_CS_fsm[31];
assign ap_CS_fsm_state33 = ap_CS_fsm[32];
assign ap_CS_fsm_state34 = ap_CS_fsm[33];
assign ap_CS_fsm_state35 = ap_CS_fsm[34];
assign ap_CS_fsm_state36 = ap_CS_fsm[35];
assign ap_CS_fsm_state37 = ap_CS_fsm[36];
assign ap_CS_fsm_state38 = ap_CS_fsm[37];
assign ap_CS_fsm_state39 = ap_CS_fsm[38];
assign ap_CS_fsm_state4 = ap_CS_fsm[3];
assign ap_CS_fsm_state40 = ap_CS_fsm[39];
assign ap_CS_fsm_state41 = ap_CS_fsm[40];
assign ap_CS_fsm_state42 = ap_CS_fsm[41];
assign ap_CS_fsm_state43 = ap_CS_fsm[42];
assign ap_CS_fsm_state44 = ap_CS_fsm[43];
assign ap_CS_fsm_state45 = ap_CS_fsm[44];
assign ap_CS_fsm_state46 = ap_CS_fsm[45];
assign ap_CS_fsm_state47 = ap_CS_fsm[46];
assign ap_CS_fsm_state48 = ap_CS_fsm[47];
assign ap_CS_fsm_state49 = ap_CS_fsm[48];
assign ap_CS_fsm_state5 = ap_CS_fsm[4];
assign ap_CS_fsm_state50 = ap_CS_fsm[49];
assign ap_CS_fsm_state51 = ap_CS_fsm[50];
assign ap_CS_fsm_state52 = ap_CS_fsm[51];
assign ap_CS_fsm_state6 = ap_CS_fsm[5];
assign ap_CS_fsm_state7 = ap_CS_fsm[6];
assign ap_CS_fsm_state8 = ap_CS_fsm[7];
assign ap_CS_fsm_state9 = ap_CS_fsm[8];
assign ap_done = op_29_ap_vld;
assign ap_ready = op_29_ap_vld;
assign grp_fu_1181_p0 = { select_ln850_4_reg_2264[9], select_ln850_4_reg_2264, 13'h0000 };
assign grp_fu_1181_p1 = { op_11[15], op_11[15], op_11[15], op_11[15], op_11[15], op_11[15], op_11[15], op_11[15], op_11 };
assign grp_fu_1314_p0 = { tmp_reg_2338[10], tmp_reg_2338 };
assign grp_fu_1510_p0 = { select_ln353_reg_2427[11], select_ln353_reg_2427[11], select_ln353_reg_2427[11], select_ln353_reg_2427[11], select_ln353_reg_2427[11], select_ln353_reg_2427[11], select_ln353_reg_2427[11], select_ln353_reg_2427[11], select_ln353_reg_2427[11], select_ln353_reg_2427[11], select_ln353_reg_2427[11], select_ln353_reg_2427[11], select_ln353_reg_2427[11], select_ln353_reg_2427[11], select_ln353_reg_2427[11], select_ln353_reg_2427[11], select_ln353_reg_2427[11], select_ln353_reg_2427[11], select_ln353_reg_2427[11], select_ln353_reg_2427[11], select_ln353_reg_2427[11], select_ln353_reg_2427, 2'h0 };
assign grp_fu_1510_p1 = { op_12_V_reg_2422[7], op_12_V_reg_2422[7], op_12_V_reg_2422[7], op_12_V_reg_2422[7], op_12_V_reg_2422[7], op_12_V_reg_2422[7], op_12_V_reg_2422[7], op_12_V_reg_2422[7], op_12_V_reg_2422[7], op_12_V_reg_2422[7], op_12_V_reg_2422[7], op_12_V_reg_2422[7], op_12_V_reg_2422[7], op_12_V_reg_2422[7], op_12_V_reg_2422[7], op_12_V_reg_2422[7], op_12_V_reg_2422[7], op_12_V_reg_2422[7], op_12_V_reg_2422[7], op_12_V_reg_2422[7], op_12_V_reg_2422[7], op_12_V_reg_2422[7], op_12_V_reg_2422[7], op_12_V_reg_2422[7], op_12_V_reg_2422[7], op_12_V_reg_2422[7], op_12_V_reg_2422[7], op_12_V_reg_2422 };
assign grp_fu_1569_p0 = { select_ln353_1_reg_2474[31], select_ln353_1_reg_2474, 2'h0 };
assign grp_fu_1569_p1 = { op_13_V_reg_2328[15], op_13_V_reg_2328[15], op_13_V_reg_2328[15], op_13_V_reg_2328[15], op_13_V_reg_2328[15], op_13_V_reg_2328[15], op_13_V_reg_2328[15], op_13_V_reg_2328[15], op_13_V_reg_2328[15], op_13_V_reg_2328[15], op_13_V_reg_2328[15], op_13_V_reg_2328[15], op_13_V_reg_2328[15], op_13_V_reg_2328[15], op_13_V_reg_2328[15], op_13_V_reg_2328[15], op_13_V_reg_2328[15], op_13_V_reg_2328[15], op_13_V_reg_2328[15], op_13_V_reg_2328 };
assign grp_fu_1612_p1 = { 28'h0000000, ret_V_20_reg_2437 };
assign grp_fu_1631_p0 = { op_24_V_reg_2516[31], op_24_V_reg_2516, 1'h0 };
assign grp_fu_1631_p1 = { op_15_V_reg_2322[1], op_15_V_reg_2322[1], op_15_V_reg_2322[1], op_15_V_reg_2322[1], op_15_V_reg_2322[1], op_15_V_reg_2322[1], op_15_V_reg_2322[1], op_15_V_reg_2322[1], op_15_V_reg_2322[1], op_15_V_reg_2322[1], op_15_V_reg_2322[1], op_15_V_reg_2322[1], op_15_V_reg_2322[1], op_15_V_reg_2322[1], op_15_V_reg_2322[1], op_15_V_reg_2322[1], op_15_V_reg_2322[1], op_15_V_reg_2322[1], op_15_V_reg_2322[1], op_15_V_reg_2322[1], op_15_V_reg_2322[1], op_15_V_reg_2322[1], op_15_V_reg_2322[1], op_15_V_reg_2322[1], op_15_V_reg_2322[1], op_15_V_reg_2322[1], op_15_V_reg_2322[1], op_15_V_reg_2322[1], op_15_V_reg_2322[1], op_15_V_reg_2322[1], op_15_V_reg_2322[1], op_15_V_reg_2322[1], op_15_V_reg_2322 };
assign grp_fu_1659_p0 = { op_19_V_reg_2248[7], op_19_V_reg_2248 };
assign grp_fu_1659_p1 = { 5'h00, op_18 };
assign grp_fu_1700_p0 = { add_ln69_1_reg_2563[8], add_ln69_1_reg_2563[8], add_ln69_1_reg_2563[8], add_ln69_1_reg_2563[8], add_ln69_1_reg_2563[8], add_ln69_1_reg_2563[8], add_ln69_1_reg_2563[8], add_ln69_1_reg_2563[8], add_ln69_1_reg_2563 };
assign grp_fu_1700_p1 = { op_16[15], op_16 };
assign grp_fu_1709_p0 = { add_ln69_2_reg_2588[16], add_ln69_2_reg_2588[16], add_ln69_2_reg_2588[16], add_ln69_2_reg_2588[16], add_ln69_2_reg_2588[16], add_ln69_2_reg_2588[16], add_ln69_2_reg_2588[16], add_ln69_2_reg_2588[16], add_ln69_2_reg_2588[16], add_ln69_2_reg_2588[16], add_ln69_2_reg_2588[16], add_ln69_2_reg_2588[16], add_ln69_2_reg_2588[16], add_ln69_2_reg_2588[16], add_ln69_2_reg_2588[16], add_ln69_2_reg_2588 };
assign grp_fu_279_p0 = op_0[3:1];
assign grp_fu_428_p0 = { op_0[3], op_0, 2'h0 };
assign grp_fu_428_p1 = { op_1_V_reg_1789[3], op_1_V_reg_1789[3], op_1_V_reg_1789[3], op_1_V_reg_1789 };
assign grp_fu_434_p0 = { trunc_ln1192_reg_1756, 2'h0 };
assign grp_fu_434_p1 = { op_1_V_reg_1789[3], op_1_V_reg_1789 };
assign grp_fu_440_p1 = { op_0[1:0], 2'h0 };
assign grp_fu_641_p0 = { ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783 };
assign grp_fu_650_p0 = { ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783 };
assign grp_fu_735_p0 = { ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783 };
assign grp_fu_735_p1 = op_7[7:0];
assign grp_fu_773_p1 = { 1'h0, and_ln412_reg_2020 };
assign grp_fu_820_p0 = { 2'h0, op_10_V_reg_2047, 3'h0 };
assign grp_fu_820_p1 = { op_6[7], op_6[7], op_6[7], op_6[7], op_6[7], op_6 };
assign grp_fu_880_p0 = { 13'h0000, ret_V_18_reg_2075 };
assign grp_fu_880_p1 = { 1'h0, op_7 };
assign grp_fu_889_p0 = ret_V_18_reg_2075;
assign grp_fu_889_p00 = { 3'h0, ret_V_18_reg_2075 };
assign grp_fu_940_p0 = { 1'h0, sext_ln1116_reg_1923 };
assign grp_fu_940_p1 = { 32'h00000000, rhs_4_reg_2120 };
assign grp_fu_949_p1 = { 7'h00, rhs_4_reg_2120 };
assign lhs_fu_399_p3 = { op_0, 2'h0 };
assign op_29 = grp_fu_1709_p2;
assign p_Result_13_fu_786_p3 = r_V_6_reg_1987[35];
assign p_Result_14_fu_1054_p3 = ret_V_19_reg_2103[12];
assign p_Result_17_fu_1473_p3 = r_V_7_reg_2366[6];
assign p_Result_18_fu_1445_p3 = ret_V_21_reg_2333[23];
assign p_Result_22_fu_1366_p4 = { ret_1_reg_2216[6], p_Val2_15_fu_1360_p2 };
assign p_Result_23_fu_1536_p3 = ret_V_22_reg_2457[34];
assign p_Result_24_fu_1590_p3 = ret_V_23_reg_2489[34];
assign p_Result_25_fu_1665_p3 = ret_V_25_reg_2531[33];
assign p_Result_29_fu_519_p3 = add_ln1192_1_reg_1826[4];
assign p_Result_31_fu_656_p1 = grp_fu_641_p2[0];
assign p_Result_38_fu_1327_p3 = ret_1_reg_2216[6];
assign p_Result_7_fu_557_p4 = { add_ln1192_1_reg_1826[4], p_Val2_3_fu_552_p2 };
assign p_Val2_10_fu_1114_p3 = { trunc_ln731_1_reg_2155, 2'h0 };
assign p_Val2_14_fu_1320_p3 = { trunc_ln731_2_reg_2230, 2'h0 };
assign p_Val2_s_fu_251_p2 = { op_0[0], 3'h0 };
assign ret_V_fu_263_p4 = op_0[3:1];
assign rhs_2_fu_809_p3 = { op_10_V_reg_2047, 3'h0 };
assign rhs_3_fu_1170_p3 = { select_ln850_4_reg_2264, 13'h0000 };
assign rhs_5_fu_1558_p3 = { select_ln353_1_reg_2474, 2'h0 };
assign rhs_7_fu_1620_p3 = { op_24_V_reg_2516, 1'h0 };
assign sext_ln1116_fu_630_p1 = { ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783 };
assign sext_ln1192_2_fu_1166_p0 = op_11;
assign sext_ln703_1_fu_805_p0 = op_6;
assign sext_ln727_fu_851_p1 = { op_3_V_reg_1917[3], op_3_V_reg_1917[3], op_3_V_reg_1917[3], op_3_V_reg_1917[3], op_3_V_reg_1917 };
assign sext_ln850_fu_1311_p1 = { tmp_reg_2338[10], tmp_reg_2338 };
assign shl_ln_fu_857_p3 = { ret_V_18_reg_2075, 3'h0 };
assign tmp_13_fu_959_p3 = r_V_5_reg_1944[3];
assign tmp_23_fu_1334_p3 = ret_1_reg_2216[6];
assign tmp_24_fu_1341_p3 = ret_1_reg_2216[5];
assign tmp_26_fu_1499_p3 = { select_ln353_reg_2427, 2'h0 };
assign tmp_6_fu_526_p3 = add_ln1192_1_reg_1826[4];
assign tmp_7_fu_533_p3 = p_Val2_2_reg_1839[3];
assign trunc_ln1192_fu_285_p1 = op_0[2:0];
assign trunc_ln213_fu_731_p1 = op_7[7:0];
assign trunc_ln731_1_fu_912_p1 = grp_fu_880_p2[13:0];
assign trunc_ln731_2_fu_1006_p1 = grp_fu_940_p2[5:0];
assign trunc_ln731_fu_298_p1 = op_0[0];
assign trunc_ln851_1_fu_826_p0 = op_6;
assign trunc_ln851_1_fu_826_p1 = op_6[2:0];
assign trunc_ln851_2_fu_1480_p1 = r_V_7_reg_2366[0];
assign trunc_ln851_3_fu_1187_p0 = op_11;
assign trunc_ln851_3_fu_1187_p1 = op_11[12:0];
assign trunc_ln851_4_fu_1469_p1 = op_12_V_fu_1452_p3[1:0];
assign trunc_ln851_5_fu_1297_p1 = op_13_V_fu_1252_p3[1:0];
assign trunc_ln851_6_fu_1672_p1 = op_15_V_reg_2322[0];
assign trunc_ln851_fu_724_p1 = grp_fu_650_p2[2:0];
assign zext_ln1116_fu_633_p1 = { 4'h0, ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783 };
assign zext_ln1499_fu_864_p1 = { 1'h0, ret_V_18_reg_2075, 3'h0 };
assign \sub_8s_8ns_8_2_1_U7.top_sub_8s_8ns_8_2_1_Adder_4_U.ain_s0  = \sub_8s_8ns_8_2_1_U7.top_sub_8s_8ns_8_2_1_Adder_4_U.a ;
assign \sub_8s_8ns_8_2_1_U7.top_sub_8s_8ns_8_2_1_Adder_4_U.s  = { \sub_8s_8ns_8_2_1_U7.top_sub_8s_8ns_8_2_1_Adder_4_U.fas_s2 , \sub_8s_8ns_8_2_1_U7.top_sub_8s_8ns_8_2_1_Adder_4_U.sum_s1  };
assign \sub_8s_8ns_8_2_1_U7.top_sub_8s_8ns_8_2_1_Adder_4_U.u2.a  = \sub_8s_8ns_8_2_1_U7.top_sub_8s_8ns_8_2_1_Adder_4_U.ain_s1 ;
assign \sub_8s_8ns_8_2_1_U7.top_sub_8s_8ns_8_2_1_Adder_4_U.u2.b  = \sub_8s_8ns_8_2_1_U7.top_sub_8s_8ns_8_2_1_Adder_4_U.bin_s1 ;
assign \sub_8s_8ns_8_2_1_U7.top_sub_8s_8ns_8_2_1_Adder_4_U.u2.cin  = \sub_8s_8ns_8_2_1_U7.top_sub_8s_8ns_8_2_1_Adder_4_U.carry_s1 ;
assign \sub_8s_8ns_8_2_1_U7.top_sub_8s_8ns_8_2_1_Adder_4_U.facout_s2  = \sub_8s_8ns_8_2_1_U7.top_sub_8s_8ns_8_2_1_Adder_4_U.u2.cout ;
assign \sub_8s_8ns_8_2_1_U7.top_sub_8s_8ns_8_2_1_Adder_4_U.fas_s2  = \sub_8s_8ns_8_2_1_U7.top_sub_8s_8ns_8_2_1_Adder_4_U.u2.s ;
assign \sub_8s_8ns_8_2_1_U7.top_sub_8s_8ns_8_2_1_Adder_4_U.u1.a  = \sub_8s_8ns_8_2_1_U7.top_sub_8s_8ns_8_2_1_Adder_4_U.a [3:0];
assign \sub_8s_8ns_8_2_1_U7.top_sub_8s_8ns_8_2_1_Adder_4_U.u1.b  = \sub_8s_8ns_8_2_1_U7.top_sub_8s_8ns_8_2_1_Adder_4_U.bin_s0 [3:0];
assign \sub_8s_8ns_8_2_1_U7.top_sub_8s_8ns_8_2_1_Adder_4_U.u1.cin  = 1'h1;
assign \sub_8s_8ns_8_2_1_U7.top_sub_8s_8ns_8_2_1_Adder_4_U.facout_s1  = \sub_8s_8ns_8_2_1_U7.top_sub_8s_8ns_8_2_1_Adder_4_U.u1.cout ;
assign \sub_8s_8ns_8_2_1_U7.top_sub_8s_8ns_8_2_1_Adder_4_U.fas_s1  = \sub_8s_8ns_8_2_1_U7.top_sub_8s_8ns_8_2_1_Adder_4_U.u1.s ;
assign \sub_8s_8ns_8_2_1_U7.top_sub_8s_8ns_8_2_1_Adder_4_U.a  = \sub_8s_8ns_8_2_1_U7.din0 ;
assign \sub_8s_8ns_8_2_1_U7.top_sub_8s_8ns_8_2_1_Adder_4_U.b  = \sub_8s_8ns_8_2_1_U7.din1 ;
assign \sub_8s_8ns_8_2_1_U7.top_sub_8s_8ns_8_2_1_Adder_4_U.ce  = \sub_8s_8ns_8_2_1_U7.ce ;
assign \sub_8s_8ns_8_2_1_U7.top_sub_8s_8ns_8_2_1_Adder_4_U.clk  = \sub_8s_8ns_8_2_1_U7.clk ;
assign \sub_8s_8ns_8_2_1_U7.top_sub_8s_8ns_8_2_1_Adder_4_U.reset  = \sub_8s_8ns_8_2_1_U7.reset ;
assign \sub_8s_8ns_8_2_1_U7.dout  = \sub_8s_8ns_8_2_1_U7.top_sub_8s_8ns_8_2_1_Adder_4_U.s ;
assign \sub_8s_8ns_8_2_1_U7.ce  = 1'h1;
assign \sub_8s_8ns_8_2_1_U7.clk  = ap_clk;
assign \sub_8s_8ns_8_2_1_U7.din0  = { ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783 };
assign \sub_8s_8ns_8_2_1_U7.din1  = op_7[7:0];
assign grp_fu_735_p2 = \sub_8s_8ns_8_2_1_U7.dout ;
assign \sub_8s_8ns_8_2_1_U7.reset  = ap_rst;
assign \sub_8ns_8ns_8_2_1_U15.top_sub_8ns_8ns_8_2_1_Adder_11_U.ain_s0  = \sub_8ns_8ns_8_2_1_U15.top_sub_8ns_8ns_8_2_1_Adder_11_U.a ;
assign \sub_8ns_8ns_8_2_1_U15.top_sub_8ns_8ns_8_2_1_Adder_11_U.s  = { \sub_8ns_8ns_8_2_1_U15.top_sub_8ns_8ns_8_2_1_Adder_11_U.fas_s2 , \sub_8ns_8ns_8_2_1_U15.top_sub_8ns_8ns_8_2_1_Adder_11_U.sum_s1  };
assign \sub_8ns_8ns_8_2_1_U15.top_sub_8ns_8ns_8_2_1_Adder_11_U.u2.a  = \sub_8ns_8ns_8_2_1_U15.top_sub_8ns_8ns_8_2_1_Adder_11_U.ain_s1 ;
assign \sub_8ns_8ns_8_2_1_U15.top_sub_8ns_8ns_8_2_1_Adder_11_U.u2.b  = \sub_8ns_8ns_8_2_1_U15.top_sub_8ns_8ns_8_2_1_Adder_11_U.bin_s1 ;
assign \sub_8ns_8ns_8_2_1_U15.top_sub_8ns_8ns_8_2_1_Adder_11_U.u2.cin  = \sub_8ns_8ns_8_2_1_U15.top_sub_8ns_8ns_8_2_1_Adder_11_U.carry_s1 ;
assign \sub_8ns_8ns_8_2_1_U15.top_sub_8ns_8ns_8_2_1_Adder_11_U.facout_s2  = \sub_8ns_8ns_8_2_1_U15.top_sub_8ns_8ns_8_2_1_Adder_11_U.u2.cout ;
assign \sub_8ns_8ns_8_2_1_U15.top_sub_8ns_8ns_8_2_1_Adder_11_U.fas_s2  = \sub_8ns_8ns_8_2_1_U15.top_sub_8ns_8ns_8_2_1_Adder_11_U.u2.s ;
assign \sub_8ns_8ns_8_2_1_U15.top_sub_8ns_8ns_8_2_1_Adder_11_U.u1.a  = \sub_8ns_8ns_8_2_1_U15.top_sub_8ns_8ns_8_2_1_Adder_11_U.a [3:0];
assign \sub_8ns_8ns_8_2_1_U15.top_sub_8ns_8ns_8_2_1_Adder_11_U.u1.b  = \sub_8ns_8ns_8_2_1_U15.top_sub_8ns_8ns_8_2_1_Adder_11_U.bin_s0 [3:0];
assign \sub_8ns_8ns_8_2_1_U15.top_sub_8ns_8ns_8_2_1_Adder_11_U.u1.cin  = 1'h1;
assign \sub_8ns_8ns_8_2_1_U15.top_sub_8ns_8ns_8_2_1_Adder_11_U.facout_s1  = \sub_8ns_8ns_8_2_1_U15.top_sub_8ns_8ns_8_2_1_Adder_11_U.u1.cout ;
assign \sub_8ns_8ns_8_2_1_U15.top_sub_8ns_8ns_8_2_1_Adder_11_U.fas_s1  = \sub_8ns_8ns_8_2_1_U15.top_sub_8ns_8ns_8_2_1_Adder_11_U.u1.s ;
assign \sub_8ns_8ns_8_2_1_U15.top_sub_8ns_8ns_8_2_1_Adder_11_U.a  = \sub_8ns_8ns_8_2_1_U15.din0 ;
assign \sub_8ns_8ns_8_2_1_U15.top_sub_8ns_8ns_8_2_1_Adder_11_U.b  = \sub_8ns_8ns_8_2_1_U15.din1 ;
assign \sub_8ns_8ns_8_2_1_U15.top_sub_8ns_8ns_8_2_1_Adder_11_U.ce  = \sub_8ns_8ns_8_2_1_U15.ce ;
assign \sub_8ns_8ns_8_2_1_U15.top_sub_8ns_8ns_8_2_1_Adder_11_U.clk  = \sub_8ns_8ns_8_2_1_U15.clk ;
assign \sub_8ns_8ns_8_2_1_U15.top_sub_8ns_8ns_8_2_1_Adder_11_U.reset  = \sub_8ns_8ns_8_2_1_U15.reset ;
assign \sub_8ns_8ns_8_2_1_U15.dout  = \sub_8ns_8ns_8_2_1_U15.top_sub_8ns_8ns_8_2_1_Adder_11_U.s ;
assign \sub_8ns_8ns_8_2_1_U15.ce  = 1'h1;
assign \sub_8ns_8ns_8_2_1_U15.clk  = ap_clk;
assign \sub_8ns_8ns_8_2_1_U15.din0  = trunc_ln213_reg_2014;
assign \sub_8ns_8ns_8_2_1_U15.din1  = { 7'h00, rhs_4_reg_2120 };
assign grp_fu_949_p2 = \sub_8ns_8ns_8_2_1_U15.dout ;
assign \sub_8ns_8ns_8_2_1_U15.reset  = ap_rst;
assign \sub_33ns_33ns_33_2_1_U14.top_sub_33ns_33ns_33_2_1_Adder_10_U.ain_s0  = \sub_33ns_33ns_33_2_1_U14.top_sub_33ns_33ns_33_2_1_Adder_10_U.a ;
assign \sub_33ns_33ns_33_2_1_U14.top_sub_33ns_33ns_33_2_1_Adder_10_U.s  = { \sub_33ns_33ns_33_2_1_U14.top_sub_33ns_33ns_33_2_1_Adder_10_U.fas_s2 , \sub_33ns_33ns_33_2_1_U14.top_sub_33ns_33ns_33_2_1_Adder_10_U.sum_s1  };
assign \sub_33ns_33ns_33_2_1_U14.top_sub_33ns_33ns_33_2_1_Adder_10_U.u2.a  = \sub_33ns_33ns_33_2_1_U14.top_sub_33ns_33ns_33_2_1_Adder_10_U.ain_s1 ;
assign \sub_33ns_33ns_33_2_1_U14.top_sub_33ns_33ns_33_2_1_Adder_10_U.u2.b  = \sub_33ns_33ns_33_2_1_U14.top_sub_33ns_33ns_33_2_1_Adder_10_U.bin_s1 ;
assign \sub_33ns_33ns_33_2_1_U14.top_sub_33ns_33ns_33_2_1_Adder_10_U.u2.cin  = \sub_33ns_33ns_33_2_1_U14.top_sub_33ns_33ns_33_2_1_Adder_10_U.carry_s1 ;
assign \sub_33ns_33ns_33_2_1_U14.top_sub_33ns_33ns_33_2_1_Adder_10_U.facout_s2  = \sub_33ns_33ns_33_2_1_U14.top_sub_33ns_33ns_33_2_1_Adder_10_U.u2.cout ;
assign \sub_33ns_33ns_33_2_1_U14.top_sub_33ns_33ns_33_2_1_Adder_10_U.fas_s2  = \sub_33ns_33ns_33_2_1_U14.top_sub_33ns_33ns_33_2_1_Adder_10_U.u2.s ;
assign \sub_33ns_33ns_33_2_1_U14.top_sub_33ns_33ns_33_2_1_Adder_10_U.u1.a  = \sub_33ns_33ns_33_2_1_U14.top_sub_33ns_33ns_33_2_1_Adder_10_U.a [15:0];
assign \sub_33ns_33ns_33_2_1_U14.top_sub_33ns_33ns_33_2_1_Adder_10_U.u1.b  = \sub_33ns_33ns_33_2_1_U14.top_sub_33ns_33ns_33_2_1_Adder_10_U.bin_s0 [15:0];
assign \sub_33ns_33ns_33_2_1_U14.top_sub_33ns_33ns_33_2_1_Adder_10_U.u1.cin  = 1'h1;
assign \sub_33ns_33ns_33_2_1_U14.top_sub_33ns_33ns_33_2_1_Adder_10_U.facout_s1  = \sub_33ns_33ns_33_2_1_U14.top_sub_33ns_33ns_33_2_1_Adder_10_U.u1.cout ;
assign \sub_33ns_33ns_33_2_1_U14.top_sub_33ns_33ns_33_2_1_Adder_10_U.fas_s1  = \sub_33ns_33ns_33_2_1_U14.top_sub_33ns_33ns_33_2_1_Adder_10_U.u1.s ;
assign \sub_33ns_33ns_33_2_1_U14.top_sub_33ns_33ns_33_2_1_Adder_10_U.a  = \sub_33ns_33ns_33_2_1_U14.din0 ;
assign \sub_33ns_33ns_33_2_1_U14.top_sub_33ns_33ns_33_2_1_Adder_10_U.b  = \sub_33ns_33ns_33_2_1_U14.din1 ;
assign \sub_33ns_33ns_33_2_1_U14.top_sub_33ns_33ns_33_2_1_Adder_10_U.ce  = \sub_33ns_33ns_33_2_1_U14.ce ;
assign \sub_33ns_33ns_33_2_1_U14.top_sub_33ns_33ns_33_2_1_Adder_10_U.clk  = \sub_33ns_33ns_33_2_1_U14.clk ;
assign \sub_33ns_33ns_33_2_1_U14.top_sub_33ns_33ns_33_2_1_Adder_10_U.reset  = \sub_33ns_33ns_33_2_1_U14.reset ;
assign \sub_33ns_33ns_33_2_1_U14.dout  = \sub_33ns_33ns_33_2_1_U14.top_sub_33ns_33ns_33_2_1_Adder_10_U.s ;
assign \sub_33ns_33ns_33_2_1_U14.ce  = 1'h1;
assign \sub_33ns_33ns_33_2_1_U14.clk  = ap_clk;
assign \sub_33ns_33ns_33_2_1_U14.din0  = { 1'h0, sext_ln1116_reg_1923 };
assign \sub_33ns_33ns_33_2_1_U14.din1  = { 32'h00000000, rhs_4_reg_2120 };
assign grp_fu_940_p2 = \sub_33ns_33ns_33_2_1_U14.dout ;
assign \sub_33ns_33ns_33_2_1_U14.reset  = ap_rst;
assign \sub_17ns_17ns_17_2_1_U11.top_sub_17ns_17ns_17_2_1_Adder_8_U.ain_s0  = \sub_17ns_17ns_17_2_1_U11.top_sub_17ns_17ns_17_2_1_Adder_8_U.a ;
assign \sub_17ns_17ns_17_2_1_U11.top_sub_17ns_17ns_17_2_1_Adder_8_U.s  = { \sub_17ns_17ns_17_2_1_U11.top_sub_17ns_17ns_17_2_1_Adder_8_U.fas_s2 , \sub_17ns_17ns_17_2_1_U11.top_sub_17ns_17ns_17_2_1_Adder_8_U.sum_s1  };
assign \sub_17ns_17ns_17_2_1_U11.top_sub_17ns_17ns_17_2_1_Adder_8_U.u2.a  = \sub_17ns_17ns_17_2_1_U11.top_sub_17ns_17ns_17_2_1_Adder_8_U.ain_s1 ;
assign \sub_17ns_17ns_17_2_1_U11.top_sub_17ns_17ns_17_2_1_Adder_8_U.u2.b  = \sub_17ns_17ns_17_2_1_U11.top_sub_17ns_17ns_17_2_1_Adder_8_U.bin_s1 ;
assign \sub_17ns_17ns_17_2_1_U11.top_sub_17ns_17ns_17_2_1_Adder_8_U.u2.cin  = \sub_17ns_17ns_17_2_1_U11.top_sub_17ns_17ns_17_2_1_Adder_8_U.carry_s1 ;
assign \sub_17ns_17ns_17_2_1_U11.top_sub_17ns_17ns_17_2_1_Adder_8_U.facout_s2  = \sub_17ns_17ns_17_2_1_U11.top_sub_17ns_17ns_17_2_1_Adder_8_U.u2.cout ;
assign \sub_17ns_17ns_17_2_1_U11.top_sub_17ns_17ns_17_2_1_Adder_8_U.fas_s2  = \sub_17ns_17ns_17_2_1_U11.top_sub_17ns_17ns_17_2_1_Adder_8_U.u2.s ;
assign \sub_17ns_17ns_17_2_1_U11.top_sub_17ns_17ns_17_2_1_Adder_8_U.u1.a  = \sub_17ns_17ns_17_2_1_U11.top_sub_17ns_17ns_17_2_1_Adder_8_U.a [7:0];
assign \sub_17ns_17ns_17_2_1_U11.top_sub_17ns_17ns_17_2_1_Adder_8_U.u1.b  = \sub_17ns_17ns_17_2_1_U11.top_sub_17ns_17ns_17_2_1_Adder_8_U.bin_s0 [7:0];
assign \sub_17ns_17ns_17_2_1_U11.top_sub_17ns_17ns_17_2_1_Adder_8_U.u1.cin  = 1'h1;
assign \sub_17ns_17ns_17_2_1_U11.top_sub_17ns_17ns_17_2_1_Adder_8_U.facout_s1  = \sub_17ns_17ns_17_2_1_U11.top_sub_17ns_17ns_17_2_1_Adder_8_U.u1.cout ;
assign \sub_17ns_17ns_17_2_1_U11.top_sub_17ns_17ns_17_2_1_Adder_8_U.fas_s1  = \sub_17ns_17ns_17_2_1_U11.top_sub_17ns_17ns_17_2_1_Adder_8_U.u1.s ;
assign \sub_17ns_17ns_17_2_1_U11.top_sub_17ns_17ns_17_2_1_Adder_8_U.a  = \sub_17ns_17ns_17_2_1_U11.din0 ;
assign \sub_17ns_17ns_17_2_1_U11.top_sub_17ns_17ns_17_2_1_Adder_8_U.b  = \sub_17ns_17ns_17_2_1_U11.din1 ;
assign \sub_17ns_17ns_17_2_1_U11.top_sub_17ns_17ns_17_2_1_Adder_8_U.ce  = \sub_17ns_17ns_17_2_1_U11.ce ;
assign \sub_17ns_17ns_17_2_1_U11.top_sub_17ns_17ns_17_2_1_Adder_8_U.clk  = \sub_17ns_17ns_17_2_1_U11.clk ;
assign \sub_17ns_17ns_17_2_1_U11.top_sub_17ns_17ns_17_2_1_Adder_8_U.reset  = \sub_17ns_17ns_17_2_1_U11.reset ;
assign \sub_17ns_17ns_17_2_1_U11.dout  = \sub_17ns_17ns_17_2_1_U11.top_sub_17ns_17ns_17_2_1_Adder_8_U.s ;
assign \sub_17ns_17ns_17_2_1_U11.ce  = 1'h1;
assign \sub_17ns_17ns_17_2_1_U11.clk  = ap_clk;
assign \sub_17ns_17ns_17_2_1_U11.din0  = { 13'h0000, ret_V_18_reg_2075 };
assign \sub_17ns_17ns_17_2_1_U11.din1  = { 1'h0, op_7 };
assign grp_fu_880_p2 = \sub_17ns_17ns_17_2_1_U11.dout ;
assign \sub_17ns_17ns_17_2_1_U11.reset  = ap_rst;
assign \mul_4ns_3s_7_7_1_U12.top_mul_4ns_3s_7_7_1_Mul_DSP_1_U.p  = \mul_4ns_3s_7_7_1_U12.top_mul_4ns_3s_7_7_1_Mul_DSP_1_U.buff4 ;
assign \mul_4ns_3s_7_7_1_U12.top_mul_4ns_3s_7_7_1_Mul_DSP_1_U.a  = \mul_4ns_3s_7_7_1_U12.din0 ;
assign \mul_4ns_3s_7_7_1_U12.top_mul_4ns_3s_7_7_1_Mul_DSP_1_U.b  = \mul_4ns_3s_7_7_1_U12.din1 ;
assign \mul_4ns_3s_7_7_1_U12.top_mul_4ns_3s_7_7_1_Mul_DSP_1_U.ce  = \mul_4ns_3s_7_7_1_U12.ce ;
assign \mul_4ns_3s_7_7_1_U12.top_mul_4ns_3s_7_7_1_Mul_DSP_1_U.clk  = \mul_4ns_3s_7_7_1_U12.clk ;
assign \mul_4ns_3s_7_7_1_U12.dout  = \mul_4ns_3s_7_7_1_U12.top_mul_4ns_3s_7_7_1_Mul_DSP_1_U.p ;
assign \mul_4ns_3s_7_7_1_U12.ce  = 1'h1;
assign \mul_4ns_3s_7_7_1_U12.clk  = ap_clk;
assign \mul_4ns_3s_7_7_1_U12.din0  = ret_V_18_reg_2075;
assign \mul_4ns_3s_7_7_1_U12.din1  = r_V_reg_1796;
assign grp_fu_889_p2 = \mul_4ns_3s_7_7_1_U12.dout ;
assign \mul_4ns_3s_7_7_1_U12.reset  = ap_rst;
assign \mul_32ns_4s_36_7_1_U6.top_mul_32ns_4s_36_7_1_Mul_DSP_0_U.p  = \mul_32ns_4s_36_7_1_U6.top_mul_32ns_4s_36_7_1_Mul_DSP_0_U.buff4 ;
assign \mul_32ns_4s_36_7_1_U6.top_mul_32ns_4s_36_7_1_Mul_DSP_0_U.a  = \mul_32ns_4s_36_7_1_U6.din0 ;
assign \mul_32ns_4s_36_7_1_U6.top_mul_32ns_4s_36_7_1_Mul_DSP_0_U.b  = \mul_32ns_4s_36_7_1_U6.din1 ;
assign \mul_32ns_4s_36_7_1_U6.top_mul_32ns_4s_36_7_1_Mul_DSP_0_U.ce  = \mul_32ns_4s_36_7_1_U6.ce ;
assign \mul_32ns_4s_36_7_1_U6.top_mul_32ns_4s_36_7_1_Mul_DSP_0_U.clk  = \mul_32ns_4s_36_7_1_U6.clk ;
assign \mul_32ns_4s_36_7_1_U6.dout  = \mul_32ns_4s_36_7_1_U6.top_mul_32ns_4s_36_7_1_Mul_DSP_0_U.p ;
assign \mul_32ns_4s_36_7_1_U6.ce  = 1'h1;
assign \mul_32ns_4s_36_7_1_U6.clk  = ap_clk;
assign \mul_32ns_4s_36_7_1_U6.din0  = { ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783 };
assign \mul_32ns_4s_36_7_1_U6.din1  = op_3_V_reg_1917;
assign grp_fu_650_p2 = \mul_32ns_4s_36_7_1_U6.dout ;
assign \mul_32ns_4s_36_7_1_U6.reset  = ap_rst;
assign \mul_32ns_4s_36_7_1_U5.top_mul_32ns_4s_36_7_1_Mul_DSP_0_U.p  = \mul_32ns_4s_36_7_1_U5.top_mul_32ns_4s_36_7_1_Mul_DSP_0_U.buff4 ;
assign \mul_32ns_4s_36_7_1_U5.top_mul_32ns_4s_36_7_1_Mul_DSP_0_U.a  = \mul_32ns_4s_36_7_1_U5.din0 ;
assign \mul_32ns_4s_36_7_1_U5.top_mul_32ns_4s_36_7_1_Mul_DSP_0_U.b  = \mul_32ns_4s_36_7_1_U5.din1 ;
assign \mul_32ns_4s_36_7_1_U5.top_mul_32ns_4s_36_7_1_Mul_DSP_0_U.ce  = \mul_32ns_4s_36_7_1_U5.ce ;
assign \mul_32ns_4s_36_7_1_U5.top_mul_32ns_4s_36_7_1_Mul_DSP_0_U.clk  = \mul_32ns_4s_36_7_1_U5.clk ;
assign \mul_32ns_4s_36_7_1_U5.dout  = \mul_32ns_4s_36_7_1_U5.top_mul_32ns_4s_36_7_1_Mul_DSP_0_U.p ;
assign \mul_32ns_4s_36_7_1_U5.ce  = 1'h1;
assign \mul_32ns_4s_36_7_1_U5.clk  = ap_clk;
assign \mul_32ns_4s_36_7_1_U5.din0  = { ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783[2], ret_V_16_reg_1783 };
assign \mul_32ns_4s_36_7_1_U5.din1  = op_8;
assign grp_fu_641_p2 = \mul_32ns_4s_36_7_1_U5.dout ;
assign \mul_32ns_4s_36_7_1_U5.reset  = ap_rst;
assign \add_9s_9ns_9_2_1_U26.top_add_9s_9ns_9_2_1_Adder_17_U.ain_s0  = \add_9s_9ns_9_2_1_U26.top_add_9s_9ns_9_2_1_Adder_17_U.a ;
assign \add_9s_9ns_9_2_1_U26.top_add_9s_9ns_9_2_1_Adder_17_U.bin_s0  = \add_9s_9ns_9_2_1_U26.top_add_9s_9ns_9_2_1_Adder_17_U.b ;
assign \add_9s_9ns_9_2_1_U26.top_add_9s_9ns_9_2_1_Adder_17_U.s  = { \add_9s_9ns_9_2_1_U26.top_add_9s_9ns_9_2_1_Adder_17_U.fas_s2 , \add_9s_9ns_9_2_1_U26.top_add_9s_9ns_9_2_1_Adder_17_U.sum_s1  };
assign \add_9s_9ns_9_2_1_U26.top_add_9s_9ns_9_2_1_Adder_17_U.u2.a  = \add_9s_9ns_9_2_1_U26.top_add_9s_9ns_9_2_1_Adder_17_U.ain_s1 ;
assign \add_9s_9ns_9_2_1_U26.top_add_9s_9ns_9_2_1_Adder_17_U.u2.b  = \add_9s_9ns_9_2_1_U26.top_add_9s_9ns_9_2_1_Adder_17_U.bin_s1 ;
assign \add_9s_9ns_9_2_1_U26.top_add_9s_9ns_9_2_1_Adder_17_U.u2.cin  = \add_9s_9ns_9_2_1_U26.top_add_9s_9ns_9_2_1_Adder_17_U.carry_s1 ;
assign \add_9s_9ns_9_2_1_U26.top_add_9s_9ns_9_2_1_Adder_17_U.facout_s2  = \add_9s_9ns_9_2_1_U26.top_add_9s_9ns_9_2_1_Adder_17_U.u2.cout ;
assign \add_9s_9ns_9_2_1_U26.top_add_9s_9ns_9_2_1_Adder_17_U.fas_s2  = \add_9s_9ns_9_2_1_U26.top_add_9s_9ns_9_2_1_Adder_17_U.u2.s ;
assign \add_9s_9ns_9_2_1_U26.top_add_9s_9ns_9_2_1_Adder_17_U.u1.a  = \add_9s_9ns_9_2_1_U26.top_add_9s_9ns_9_2_1_Adder_17_U.a [3:0];
assign \add_9s_9ns_9_2_1_U26.top_add_9s_9ns_9_2_1_Adder_17_U.u1.b  = \add_9s_9ns_9_2_1_U26.top_add_9s_9ns_9_2_1_Adder_17_U.b [3:0];
assign \add_9s_9ns_9_2_1_U26.top_add_9s_9ns_9_2_1_Adder_17_U.u1.cin  = 1'h0;
assign \add_9s_9ns_9_2_1_U26.top_add_9s_9ns_9_2_1_Adder_17_U.facout_s1  = \add_9s_9ns_9_2_1_U26.top_add_9s_9ns_9_2_1_Adder_17_U.u1.cout ;
assign \add_9s_9ns_9_2_1_U26.top_add_9s_9ns_9_2_1_Adder_17_U.fas_s1  = \add_9s_9ns_9_2_1_U26.top_add_9s_9ns_9_2_1_Adder_17_U.u1.s ;
assign \add_9s_9ns_9_2_1_U26.top_add_9s_9ns_9_2_1_Adder_17_U.a  = \add_9s_9ns_9_2_1_U26.din0 ;
assign \add_9s_9ns_9_2_1_U26.top_add_9s_9ns_9_2_1_Adder_17_U.b  = \add_9s_9ns_9_2_1_U26.din1 ;
assign \add_9s_9ns_9_2_1_U26.top_add_9s_9ns_9_2_1_Adder_17_U.ce  = \add_9s_9ns_9_2_1_U26.ce ;
assign \add_9s_9ns_9_2_1_U26.top_add_9s_9ns_9_2_1_Adder_17_U.clk  = \add_9s_9ns_9_2_1_U26.clk ;
assign \add_9s_9ns_9_2_1_U26.top_add_9s_9ns_9_2_1_Adder_17_U.reset  = \add_9s_9ns_9_2_1_U26.reset ;
assign \add_9s_9ns_9_2_1_U26.dout  = \add_9s_9ns_9_2_1_U26.top_add_9s_9ns_9_2_1_Adder_17_U.s ;
assign \add_9s_9ns_9_2_1_U26.ce  = 1'h1;
assign \add_9s_9ns_9_2_1_U26.clk  = ap_clk;
assign \add_9s_9ns_9_2_1_U26.din0  = { op_19_V_reg_2248[7], op_19_V_reg_2248 };
assign \add_9s_9ns_9_2_1_U26.din1  = { 5'h00, op_18 };
assign grp_fu_1659_p2 = \add_9s_9ns_9_2_1_U26.dout ;
assign \add_9s_9ns_9_2_1_U26.reset  = ap_rst;
assign \add_7s_7s_7_2_1_U2.top_add_7s_7s_7_2_1_Adder_1_U.ain_s0  = \add_7s_7s_7_2_1_U2.top_add_7s_7s_7_2_1_Adder_1_U.a ;
assign \add_7s_7s_7_2_1_U2.top_add_7s_7s_7_2_1_Adder_1_U.bin_s0  = \add_7s_7s_7_2_1_U2.top_add_7s_7s_7_2_1_Adder_1_U.b ;
assign \add_7s_7s_7_2_1_U2.top_add_7s_7s_7_2_1_Adder_1_U.s  = { \add_7s_7s_7_2_1_U2.top_add_7s_7s_7_2_1_Adder_1_U.fas_s2 , \add_7s_7s_7_2_1_U2.top_add_7s_7s_7_2_1_Adder_1_U.sum_s1  };
assign \add_7s_7s_7_2_1_U2.top_add_7s_7s_7_2_1_Adder_1_U.u2.a  = \add_7s_7s_7_2_1_U2.top_add_7s_7s_7_2_1_Adder_1_U.ain_s1 ;
assign \add_7s_7s_7_2_1_U2.top_add_7s_7s_7_2_1_Adder_1_U.u2.b  = \add_7s_7s_7_2_1_U2.top_add_7s_7s_7_2_1_Adder_1_U.bin_s1 ;
assign \add_7s_7s_7_2_1_U2.top_add_7s_7s_7_2_1_Adder_1_U.u2.cin  = \add_7s_7s_7_2_1_U2.top_add_7s_7s_7_2_1_Adder_1_U.carry_s1 ;
assign \add_7s_7s_7_2_1_U2.top_add_7s_7s_7_2_1_Adder_1_U.facout_s2  = \add_7s_7s_7_2_1_U2.top_add_7s_7s_7_2_1_Adder_1_U.u2.cout ;
assign \add_7s_7s_7_2_1_U2.top_add_7s_7s_7_2_1_Adder_1_U.fas_s2  = \add_7s_7s_7_2_1_U2.top_add_7s_7s_7_2_1_Adder_1_U.u2.s ;
assign \add_7s_7s_7_2_1_U2.top_add_7s_7s_7_2_1_Adder_1_U.u1.a  = \add_7s_7s_7_2_1_U2.top_add_7s_7s_7_2_1_Adder_1_U.a [2:0];
assign \add_7s_7s_7_2_1_U2.top_add_7s_7s_7_2_1_Adder_1_U.u1.b  = \add_7s_7s_7_2_1_U2.top_add_7s_7s_7_2_1_Adder_1_U.b [2:0];
assign \add_7s_7s_7_2_1_U2.top_add_7s_7s_7_2_1_Adder_1_U.u1.cin  = 1'h0;
assign \add_7s_7s_7_2_1_U2.top_add_7s_7s_7_2_1_Adder_1_U.facout_s1  = \add_7s_7s_7_2_1_U2.top_add_7s_7s_7_2_1_Adder_1_U.u1.cout ;
assign \add_7s_7s_7_2_1_U2.top_add_7s_7s_7_2_1_Adder_1_U.fas_s1  = \add_7s_7s_7_2_1_U2.top_add_7s_7s_7_2_1_Adder_1_U.u1.s ;
assign \add_7s_7s_7_2_1_U2.top_add_7s_7s_7_2_1_Adder_1_U.a  = \add_7s_7s_7_2_1_U2.din0 ;
assign \add_7s_7s_7_2_1_U2.top_add_7s_7s_7_2_1_Adder_1_U.b  = \add_7s_7s_7_2_1_U2.din1 ;
assign \add_7s_7s_7_2_1_U2.top_add_7s_7s_7_2_1_Adder_1_U.ce  = \add_7s_7s_7_2_1_U2.ce ;
assign \add_7s_7s_7_2_1_U2.top_add_7s_7s_7_2_1_Adder_1_U.clk  = \add_7s_7s_7_2_1_U2.clk ;
assign \add_7s_7s_7_2_1_U2.top_add_7s_7s_7_2_1_Adder_1_U.reset  = \add_7s_7s_7_2_1_U2.reset ;
assign \add_7s_7s_7_2_1_U2.dout  = \add_7s_7s_7_2_1_U2.top_add_7s_7s_7_2_1_Adder_1_U.s ;
assign \add_7s_7s_7_2_1_U2.ce  = 1'h1;
assign \add_7s_7s_7_2_1_U2.clk  = ap_clk;
assign \add_7s_7s_7_2_1_U2.din0  = { op_0[3], op_0, 2'h0 };
assign \add_7s_7s_7_2_1_U2.din1  = { op_1_V_reg_1789[3], op_1_V_reg_1789[3], op_1_V_reg_1789[3], op_1_V_reg_1789 };
assign grp_fu_428_p2 = \add_7s_7s_7_2_1_U2.dout ;
assign \add_7s_7s_7_2_1_U2.reset  = ap_rst;
assign \add_5ns_5s_5_2_1_U3.top_add_5ns_5s_5_2_1_Adder_2_U.ain_s0  = \add_5ns_5s_5_2_1_U3.top_add_5ns_5s_5_2_1_Adder_2_U.a ;
assign \add_5ns_5s_5_2_1_U3.top_add_5ns_5s_5_2_1_Adder_2_U.bin_s0  = \add_5ns_5s_5_2_1_U3.top_add_5ns_5s_5_2_1_Adder_2_U.b ;
assign \add_5ns_5s_5_2_1_U3.top_add_5ns_5s_5_2_1_Adder_2_U.s  = { \add_5ns_5s_5_2_1_U3.top_add_5ns_5s_5_2_1_Adder_2_U.fas_s2 , \add_5ns_5s_5_2_1_U3.top_add_5ns_5s_5_2_1_Adder_2_U.sum_s1  };
assign \add_5ns_5s_5_2_1_U3.top_add_5ns_5s_5_2_1_Adder_2_U.u2.a  = \add_5ns_5s_5_2_1_U3.top_add_5ns_5s_5_2_1_Adder_2_U.ain_s1 ;
assign \add_5ns_5s_5_2_1_U3.top_add_5ns_5s_5_2_1_Adder_2_U.u2.b  = \add_5ns_5s_5_2_1_U3.top_add_5ns_5s_5_2_1_Adder_2_U.bin_s1 ;
assign \add_5ns_5s_5_2_1_U3.top_add_5ns_5s_5_2_1_Adder_2_U.u2.cin  = \add_5ns_5s_5_2_1_U3.top_add_5ns_5s_5_2_1_Adder_2_U.carry_s1 ;
assign \add_5ns_5s_5_2_1_U3.top_add_5ns_5s_5_2_1_Adder_2_U.facout_s2  = \add_5ns_5s_5_2_1_U3.top_add_5ns_5s_5_2_1_Adder_2_U.u2.cout ;
assign \add_5ns_5s_5_2_1_U3.top_add_5ns_5s_5_2_1_Adder_2_U.fas_s2  = \add_5ns_5s_5_2_1_U3.top_add_5ns_5s_5_2_1_Adder_2_U.u2.s ;
assign \add_5ns_5s_5_2_1_U3.top_add_5ns_5s_5_2_1_Adder_2_U.u1.a  = \add_5ns_5s_5_2_1_U3.top_add_5ns_5s_5_2_1_Adder_2_U.a [1:0];
assign \add_5ns_5s_5_2_1_U3.top_add_5ns_5s_5_2_1_Adder_2_U.u1.b  = \add_5ns_5s_5_2_1_U3.top_add_5ns_5s_5_2_1_Adder_2_U.b [1:0];
assign \add_5ns_5s_5_2_1_U3.top_add_5ns_5s_5_2_1_Adder_2_U.u1.cin  = 1'h0;
assign \add_5ns_5s_5_2_1_U3.top_add_5ns_5s_5_2_1_Adder_2_U.facout_s1  = \add_5ns_5s_5_2_1_U3.top_add_5ns_5s_5_2_1_Adder_2_U.u1.cout ;
assign \add_5ns_5s_5_2_1_U3.top_add_5ns_5s_5_2_1_Adder_2_U.fas_s1  = \add_5ns_5s_5_2_1_U3.top_add_5ns_5s_5_2_1_Adder_2_U.u1.s ;
assign \add_5ns_5s_5_2_1_U3.top_add_5ns_5s_5_2_1_Adder_2_U.a  = \add_5ns_5s_5_2_1_U3.din0 ;
assign \add_5ns_5s_5_2_1_U3.top_add_5ns_5s_5_2_1_Adder_2_U.b  = \add_5ns_5s_5_2_1_U3.din1 ;
assign \add_5ns_5s_5_2_1_U3.top_add_5ns_5s_5_2_1_Adder_2_U.ce  = \add_5ns_5s_5_2_1_U3.ce ;
assign \add_5ns_5s_5_2_1_U3.top_add_5ns_5s_5_2_1_Adder_2_U.clk  = \add_5ns_5s_5_2_1_U3.clk ;
assign \add_5ns_5s_5_2_1_U3.top_add_5ns_5s_5_2_1_Adder_2_U.reset  = \add_5ns_5s_5_2_1_U3.reset ;
assign \add_5ns_5s_5_2_1_U3.dout  = \add_5ns_5s_5_2_1_U3.top_add_5ns_5s_5_2_1_Adder_2_U.s ;
assign \add_5ns_5s_5_2_1_U3.ce  = 1'h1;
assign \add_5ns_5s_5_2_1_U3.clk  = ap_clk;
assign \add_5ns_5s_5_2_1_U3.din0  = { trunc_ln1192_reg_1756, 2'h0 };
assign \add_5ns_5s_5_2_1_U3.din1  = { op_1_V_reg_1789[3], op_1_V_reg_1789 };
assign grp_fu_434_p2 = \add_5ns_5s_5_2_1_U3.dout ;
assign \add_5ns_5s_5_2_1_U3.reset  = ap_rst;
assign \add_4s_4ns_4_2_1_U4.top_add_4s_4ns_4_2_1_Adder_3_U.ain_s0  = \add_4s_4ns_4_2_1_U4.top_add_4s_4ns_4_2_1_Adder_3_U.a ;
assign \add_4s_4ns_4_2_1_U4.top_add_4s_4ns_4_2_1_Adder_3_U.bin_s0  = \add_4s_4ns_4_2_1_U4.top_add_4s_4ns_4_2_1_Adder_3_U.b ;
assign \add_4s_4ns_4_2_1_U4.top_add_4s_4ns_4_2_1_Adder_3_U.s  = { \add_4s_4ns_4_2_1_U4.top_add_4s_4ns_4_2_1_Adder_3_U.fas_s2 , \add_4s_4ns_4_2_1_U4.top_add_4s_4ns_4_2_1_Adder_3_U.sum_s1  };
assign \add_4s_4ns_4_2_1_U4.top_add_4s_4ns_4_2_1_Adder_3_U.u2.a  = \add_4s_4ns_4_2_1_U4.top_add_4s_4ns_4_2_1_Adder_3_U.ain_s1 ;
assign \add_4s_4ns_4_2_1_U4.top_add_4s_4ns_4_2_1_Adder_3_U.u2.b  = \add_4s_4ns_4_2_1_U4.top_add_4s_4ns_4_2_1_Adder_3_U.bin_s1 ;
assign \add_4s_4ns_4_2_1_U4.top_add_4s_4ns_4_2_1_Adder_3_U.u2.cin  = \add_4s_4ns_4_2_1_U4.top_add_4s_4ns_4_2_1_Adder_3_U.carry_s1 ;
assign \add_4s_4ns_4_2_1_U4.top_add_4s_4ns_4_2_1_Adder_3_U.facout_s2  = \add_4s_4ns_4_2_1_U4.top_add_4s_4ns_4_2_1_Adder_3_U.u2.cout ;
assign \add_4s_4ns_4_2_1_U4.top_add_4s_4ns_4_2_1_Adder_3_U.fas_s2  = \add_4s_4ns_4_2_1_U4.top_add_4s_4ns_4_2_1_Adder_3_U.u2.s ;
assign \add_4s_4ns_4_2_1_U4.top_add_4s_4ns_4_2_1_Adder_3_U.u1.a  = \add_4s_4ns_4_2_1_U4.top_add_4s_4ns_4_2_1_Adder_3_U.a [1:0];
assign \add_4s_4ns_4_2_1_U4.top_add_4s_4ns_4_2_1_Adder_3_U.u1.b  = \add_4s_4ns_4_2_1_U4.top_add_4s_4ns_4_2_1_Adder_3_U.b [1:0];
assign \add_4s_4ns_4_2_1_U4.top_add_4s_4ns_4_2_1_Adder_3_U.u1.cin  = 1'h0;
assign \add_4s_4ns_4_2_1_U4.top_add_4s_4ns_4_2_1_Adder_3_U.facout_s1  = \add_4s_4ns_4_2_1_U4.top_add_4s_4ns_4_2_1_Adder_3_U.u1.cout ;
assign \add_4s_4ns_4_2_1_U4.top_add_4s_4ns_4_2_1_Adder_3_U.fas_s1  = \add_4s_4ns_4_2_1_U4.top_add_4s_4ns_4_2_1_Adder_3_U.u1.s ;
assign \add_4s_4ns_4_2_1_U4.top_add_4s_4ns_4_2_1_Adder_3_U.a  = \add_4s_4ns_4_2_1_U4.din0 ;
assign \add_4s_4ns_4_2_1_U4.top_add_4s_4ns_4_2_1_Adder_3_U.b  = \add_4s_4ns_4_2_1_U4.din1 ;
assign \add_4s_4ns_4_2_1_U4.top_add_4s_4ns_4_2_1_Adder_3_U.ce  = \add_4s_4ns_4_2_1_U4.ce ;
assign \add_4s_4ns_4_2_1_U4.top_add_4s_4ns_4_2_1_Adder_3_U.clk  = \add_4s_4ns_4_2_1_U4.clk ;
assign \add_4s_4ns_4_2_1_U4.top_add_4s_4ns_4_2_1_Adder_3_U.reset  = \add_4s_4ns_4_2_1_U4.reset ;
assign \add_4s_4ns_4_2_1_U4.dout  = \add_4s_4ns_4_2_1_U4.top_add_4s_4ns_4_2_1_Adder_3_U.s ;
assign \add_4s_4ns_4_2_1_U4.ce  = 1'h1;
assign \add_4s_4ns_4_2_1_U4.clk  = ap_clk;
assign \add_4s_4ns_4_2_1_U4.din0  = op_1_V_reg_1789;
assign \add_4s_4ns_4_2_1_U4.din1  = { op_0[1:0], 2'h0 };
assign grp_fu_440_p2 = \add_4s_4ns_4_2_1_U4.dout ;
assign \add_4s_4ns_4_2_1_U4.reset  = ap_rst;
assign \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_5_U.ain_s0  = \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_5_U.a ;
assign \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_5_U.bin_s0  = \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_5_U.b ;
assign \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_5_U.s  = { \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_5_U.fas_s2 , \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_5_U.sum_s1  };
assign \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_5_U.u2.a  = \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_5_U.ain_s1 ;
assign \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_5_U.u2.b  = \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_5_U.bin_s1 ;
assign \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_5_U.u2.cin  = \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_5_U.carry_s1 ;
assign \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_5_U.facout_s2  = \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_5_U.u2.cout ;
assign \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_5_U.fas_s2  = \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_5_U.u2.s ;
assign \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_5_U.u1.a  = \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_5_U.a [1:0];
assign \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_5_U.u1.b  = \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_5_U.b [1:0];
assign \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_5_U.u1.cin  = 1'h0;
assign \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_5_U.facout_s1  = \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_5_U.u1.cout ;
assign \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_5_U.fas_s1  = \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_5_U.u1.s ;
assign \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_5_U.a  = \add_4ns_4ns_4_2_1_U8.din0 ;
assign \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_5_U.b  = \add_4ns_4ns_4_2_1_U8.din1 ;
assign \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_5_U.ce  = \add_4ns_4ns_4_2_1_U8.ce ;
assign \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_5_U.clk  = \add_4ns_4ns_4_2_1_U8.clk ;
assign \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_5_U.reset  = \add_4ns_4ns_4_2_1_U8.reset ;
assign \add_4ns_4ns_4_2_1_U8.dout  = \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_5_U.s ;
assign \add_4ns_4ns_4_2_1_U8.ce  = 1'h1;
assign \add_4ns_4ns_4_2_1_U8.clk  = ap_clk;
assign \add_4ns_4ns_4_2_1_U8.din0  = ret_V_4_cast_reg_1992;
assign \add_4ns_4ns_4_2_1_U8.din1  = 4'h1;
assign grp_fu_765_p2 = \add_4ns_4ns_4_2_1_U8.dout ;
assign \add_4ns_4ns_4_2_1_U8.reset  = ap_rst;
assign \add_4ns_4ns_4_2_1_U18.top_add_4ns_4ns_4_2_1_Adder_5_U.ain_s0  = \add_4ns_4ns_4_2_1_U18.top_add_4ns_4ns_4_2_1_Adder_5_U.a ;
assign \add_4ns_4ns_4_2_1_U18.top_add_4ns_4ns_4_2_1_Adder_5_U.bin_s0  = \add_4ns_4ns_4_2_1_U18.top_add_4ns_4ns_4_2_1_Adder_5_U.b ;
assign \add_4ns_4ns_4_2_1_U18.top_add_4ns_4ns_4_2_1_Adder_5_U.s  = { \add_4ns_4ns_4_2_1_U18.top_add_4ns_4ns_4_2_1_Adder_5_U.fas_s2 , \add_4ns_4ns_4_2_1_U18.top_add_4ns_4ns_4_2_1_Adder_5_U.sum_s1  };
assign \add_4ns_4ns_4_2_1_U18.top_add_4ns_4ns_4_2_1_Adder_5_U.u2.a  = \add_4ns_4ns_4_2_1_U18.top_add_4ns_4ns_4_2_1_Adder_5_U.ain_s1 ;
assign \add_4ns_4ns_4_2_1_U18.top_add_4ns_4ns_4_2_1_Adder_5_U.u2.b  = \add_4ns_4ns_4_2_1_U18.top_add_4ns_4ns_4_2_1_Adder_5_U.bin_s1 ;
assign \add_4ns_4ns_4_2_1_U18.top_add_4ns_4ns_4_2_1_Adder_5_U.u2.cin  = \add_4ns_4ns_4_2_1_U18.top_add_4ns_4ns_4_2_1_Adder_5_U.carry_s1 ;
assign \add_4ns_4ns_4_2_1_U18.top_add_4ns_4ns_4_2_1_Adder_5_U.facout_s2  = \add_4ns_4ns_4_2_1_U18.top_add_4ns_4ns_4_2_1_Adder_5_U.u2.cout ;
assign \add_4ns_4ns_4_2_1_U18.top_add_4ns_4ns_4_2_1_Adder_5_U.fas_s2  = \add_4ns_4ns_4_2_1_U18.top_add_4ns_4ns_4_2_1_Adder_5_U.u2.s ;
assign \add_4ns_4ns_4_2_1_U18.top_add_4ns_4ns_4_2_1_Adder_5_U.u1.a  = \add_4ns_4ns_4_2_1_U18.top_add_4ns_4ns_4_2_1_Adder_5_U.a [1:0];
assign \add_4ns_4ns_4_2_1_U18.top_add_4ns_4ns_4_2_1_Adder_5_U.u1.b  = \add_4ns_4ns_4_2_1_U18.top_add_4ns_4ns_4_2_1_Adder_5_U.b [1:0];
assign \add_4ns_4ns_4_2_1_U18.top_add_4ns_4ns_4_2_1_Adder_5_U.u1.cin  = 1'h0;
assign \add_4ns_4ns_4_2_1_U18.top_add_4ns_4ns_4_2_1_Adder_5_U.facout_s1  = \add_4ns_4ns_4_2_1_U18.top_add_4ns_4ns_4_2_1_Adder_5_U.u1.cout ;
assign \add_4ns_4ns_4_2_1_U18.top_add_4ns_4ns_4_2_1_Adder_5_U.fas_s1  = \add_4ns_4ns_4_2_1_U18.top_add_4ns_4ns_4_2_1_Adder_5_U.u1.s ;
assign \add_4ns_4ns_4_2_1_U18.top_add_4ns_4ns_4_2_1_Adder_5_U.a  = \add_4ns_4ns_4_2_1_U18.din0 ;
assign \add_4ns_4ns_4_2_1_U18.top_add_4ns_4ns_4_2_1_Adder_5_U.b  = \add_4ns_4ns_4_2_1_U18.din1 ;
assign \add_4ns_4ns_4_2_1_U18.top_add_4ns_4ns_4_2_1_Adder_5_U.ce  = \add_4ns_4ns_4_2_1_U18.ce ;
assign \add_4ns_4ns_4_2_1_U18.top_add_4ns_4ns_4_2_1_Adder_5_U.clk  = \add_4ns_4ns_4_2_1_U18.clk ;
assign \add_4ns_4ns_4_2_1_U18.top_add_4ns_4ns_4_2_1_Adder_5_U.reset  = \add_4ns_4ns_4_2_1_U18.reset ;
assign \add_4ns_4ns_4_2_1_U18.dout  = \add_4ns_4ns_4_2_1_U18.top_add_4ns_4ns_4_2_1_Adder_5_U.s ;
assign \add_4ns_4ns_4_2_1_U18.ce  = 1'h1;
assign \add_4ns_4ns_4_2_1_U18.clk  = ap_clk;
assign \add_4ns_4ns_4_2_1_U18.din0  = ret_V_10_cast_reg_2372;
assign \add_4ns_4ns_4_2_1_U18.din1  = 4'h1;
assign grp_fu_1419_p2 = \add_4ns_4ns_4_2_1_U18.dout ;
assign \add_4ns_4ns_4_2_1_U18.reset  = ap_rst;
assign \add_3ns_3ns_3_2_1_U1.top_add_3ns_3ns_3_2_1_Adder_0_U.ain_s0  = \add_3ns_3ns_3_2_1_U1.top_add_3ns_3ns_3_2_1_Adder_0_U.a ;
assign \add_3ns_3ns_3_2_1_U1.top_add_3ns_3ns_3_2_1_Adder_0_U.bin_s0  = \add_3ns_3ns_3_2_1_U1.top_add_3ns_3ns_3_2_1_Adder_0_U.b ;
assign \add_3ns_3ns_3_2_1_U1.top_add_3ns_3ns_3_2_1_Adder_0_U.s  = { \add_3ns_3ns_3_2_1_U1.top_add_3ns_3ns_3_2_1_Adder_0_U.fas_s2 , \add_3ns_3ns_3_2_1_U1.top_add_3ns_3ns_3_2_1_Adder_0_U.sum_s1  };
assign \add_3ns_3ns_3_2_1_U1.top_add_3ns_3ns_3_2_1_Adder_0_U.u2.a  = \add_3ns_3ns_3_2_1_U1.top_add_3ns_3ns_3_2_1_Adder_0_U.ain_s1 ;
assign \add_3ns_3ns_3_2_1_U1.top_add_3ns_3ns_3_2_1_Adder_0_U.u2.b  = \add_3ns_3ns_3_2_1_U1.top_add_3ns_3ns_3_2_1_Adder_0_U.bin_s1 ;
assign \add_3ns_3ns_3_2_1_U1.top_add_3ns_3ns_3_2_1_Adder_0_U.u2.cin  = \add_3ns_3ns_3_2_1_U1.top_add_3ns_3ns_3_2_1_Adder_0_U.carry_s1 ;
assign \add_3ns_3ns_3_2_1_U1.top_add_3ns_3ns_3_2_1_Adder_0_U.facout_s2  = \add_3ns_3ns_3_2_1_U1.top_add_3ns_3ns_3_2_1_Adder_0_U.u2.cout ;
assign \add_3ns_3ns_3_2_1_U1.top_add_3ns_3ns_3_2_1_Adder_0_U.fas_s2  = \add_3ns_3ns_3_2_1_U1.top_add_3ns_3ns_3_2_1_Adder_0_U.u2.s ;
assign \add_3ns_3ns_3_2_1_U1.top_add_3ns_3ns_3_2_1_Adder_0_U.u1.a  = \add_3ns_3ns_3_2_1_U1.top_add_3ns_3ns_3_2_1_Adder_0_U.a [0];
assign \add_3ns_3ns_3_2_1_U1.top_add_3ns_3ns_3_2_1_Adder_0_U.u1.b  = \add_3ns_3ns_3_2_1_U1.top_add_3ns_3ns_3_2_1_Adder_0_U.b [0];
assign \add_3ns_3ns_3_2_1_U1.top_add_3ns_3ns_3_2_1_Adder_0_U.u1.cin  = 1'h0;
assign \add_3ns_3ns_3_2_1_U1.top_add_3ns_3ns_3_2_1_Adder_0_U.facout_s1  = \add_3ns_3ns_3_2_1_U1.top_add_3ns_3ns_3_2_1_Adder_0_U.u1.cout ;
assign \add_3ns_3ns_3_2_1_U1.top_add_3ns_3ns_3_2_1_Adder_0_U.fas_s1  = \add_3ns_3ns_3_2_1_U1.top_add_3ns_3ns_3_2_1_Adder_0_U.u1.s ;
assign \add_3ns_3ns_3_2_1_U1.top_add_3ns_3ns_3_2_1_Adder_0_U.a  = \add_3ns_3ns_3_2_1_U1.din0 ;
assign \add_3ns_3ns_3_2_1_U1.top_add_3ns_3ns_3_2_1_Adder_0_U.b  = \add_3ns_3ns_3_2_1_U1.din1 ;
assign \add_3ns_3ns_3_2_1_U1.top_add_3ns_3ns_3_2_1_Adder_0_U.ce  = \add_3ns_3ns_3_2_1_U1.ce ;
assign \add_3ns_3ns_3_2_1_U1.top_add_3ns_3ns_3_2_1_Adder_0_U.clk  = \add_3ns_3ns_3_2_1_U1.clk ;
assign \add_3ns_3ns_3_2_1_U1.top_add_3ns_3ns_3_2_1_Adder_0_U.reset  = \add_3ns_3ns_3_2_1_U1.reset ;
assign \add_3ns_3ns_3_2_1_U1.dout  = \add_3ns_3ns_3_2_1_U1.top_add_3ns_3ns_3_2_1_Adder_0_U.s ;
assign \add_3ns_3ns_3_2_1_U1.ce  = 1'h1;
assign \add_3ns_3ns_3_2_1_U1.clk  = ap_clk;
assign \add_3ns_3ns_3_2_1_U1.din0  = op_0[3:1];
assign \add_3ns_3ns_3_2_1_U1.din1  = 3'h1;
assign grp_fu_279_p2 = \add_3ns_3ns_3_2_1_U1.dout ;
assign \add_3ns_3ns_3_2_1_U1.reset  = ap_rst;
assign \add_35s_35s_35_2_1_U21.top_add_35s_35s_35_2_1_Adder_14_U.ain_s0  = \add_35s_35s_35_2_1_U21.top_add_35s_35s_35_2_1_Adder_14_U.a ;
assign \add_35s_35s_35_2_1_U21.top_add_35s_35s_35_2_1_Adder_14_U.bin_s0  = \add_35s_35s_35_2_1_U21.top_add_35s_35s_35_2_1_Adder_14_U.b ;
assign \add_35s_35s_35_2_1_U21.top_add_35s_35s_35_2_1_Adder_14_U.s  = { \add_35s_35s_35_2_1_U21.top_add_35s_35s_35_2_1_Adder_14_U.fas_s2 , \add_35s_35s_35_2_1_U21.top_add_35s_35s_35_2_1_Adder_14_U.sum_s1  };
assign \add_35s_35s_35_2_1_U21.top_add_35s_35s_35_2_1_Adder_14_U.u2.a  = \add_35s_35s_35_2_1_U21.top_add_35s_35s_35_2_1_Adder_14_U.ain_s1 ;
assign \add_35s_35s_35_2_1_U21.top_add_35s_35s_35_2_1_Adder_14_U.u2.b  = \add_35s_35s_35_2_1_U21.top_add_35s_35s_35_2_1_Adder_14_U.bin_s1 ;
assign \add_35s_35s_35_2_1_U21.top_add_35s_35s_35_2_1_Adder_14_U.u2.cin  = \add_35s_35s_35_2_1_U21.top_add_35s_35s_35_2_1_Adder_14_U.carry_s1 ;
assign \add_35s_35s_35_2_1_U21.top_add_35s_35s_35_2_1_Adder_14_U.facout_s2  = \add_35s_35s_35_2_1_U21.top_add_35s_35s_35_2_1_Adder_14_U.u2.cout ;
assign \add_35s_35s_35_2_1_U21.top_add_35s_35s_35_2_1_Adder_14_U.fas_s2  = \add_35s_35s_35_2_1_U21.top_add_35s_35s_35_2_1_Adder_14_U.u2.s ;
assign \add_35s_35s_35_2_1_U21.top_add_35s_35s_35_2_1_Adder_14_U.u1.a  = \add_35s_35s_35_2_1_U21.top_add_35s_35s_35_2_1_Adder_14_U.a [16:0];
assign \add_35s_35s_35_2_1_U21.top_add_35s_35s_35_2_1_Adder_14_U.u1.b  = \add_35s_35s_35_2_1_U21.top_add_35s_35s_35_2_1_Adder_14_U.b [16:0];
assign \add_35s_35s_35_2_1_U21.top_add_35s_35s_35_2_1_Adder_14_U.u1.cin  = 1'h0;
assign \add_35s_35s_35_2_1_U21.top_add_35s_35s_35_2_1_Adder_14_U.facout_s1  = \add_35s_35s_35_2_1_U21.top_add_35s_35s_35_2_1_Adder_14_U.u1.cout ;
assign \add_35s_35s_35_2_1_U21.top_add_35s_35s_35_2_1_Adder_14_U.fas_s1  = \add_35s_35s_35_2_1_U21.top_add_35s_35s_35_2_1_Adder_14_U.u1.s ;
assign \add_35s_35s_35_2_1_U21.top_add_35s_35s_35_2_1_Adder_14_U.a  = \add_35s_35s_35_2_1_U21.din0 ;
assign \add_35s_35s_35_2_1_U21.top_add_35s_35s_35_2_1_Adder_14_U.b  = \add_35s_35s_35_2_1_U21.din1 ;
assign \add_35s_35s_35_2_1_U21.top_add_35s_35s_35_2_1_Adder_14_U.ce  = \add_35s_35s_35_2_1_U21.ce ;
assign \add_35s_35s_35_2_1_U21.top_add_35s_35s_35_2_1_Adder_14_U.clk  = \add_35s_35s_35_2_1_U21.clk ;
assign \add_35s_35s_35_2_1_U21.top_add_35s_35s_35_2_1_Adder_14_U.reset  = \add_35s_35s_35_2_1_U21.reset ;
assign \add_35s_35s_35_2_1_U21.dout  = \add_35s_35s_35_2_1_U21.top_add_35s_35s_35_2_1_Adder_14_U.s ;
assign \add_35s_35s_35_2_1_U21.ce  = 1'h1;
assign \add_35s_35s_35_2_1_U21.clk  = ap_clk;
assign \add_35s_35s_35_2_1_U21.din0  = { select_ln353_1_reg_2474[31], select_ln353_1_reg_2474, 2'h0 };
assign \add_35s_35s_35_2_1_U21.din1  = { op_13_V_reg_2328[15], op_13_V_reg_2328[15], op_13_V_reg_2328[15], op_13_V_reg_2328[15], op_13_V_reg_2328[15], op_13_V_reg_2328[15], op_13_V_reg_2328[15], op_13_V_reg_2328[15], op_13_V_reg_2328[15], op_13_V_reg_2328[15], op_13_V_reg_2328[15], op_13_V_reg_2328[15], op_13_V_reg_2328[15], op_13_V_reg_2328[15], op_13_V_reg_2328[15], op_13_V_reg_2328[15], op_13_V_reg_2328[15], op_13_V_reg_2328[15], op_13_V_reg_2328[15], op_13_V_reg_2328 };
assign grp_fu_1569_p2 = \add_35s_35s_35_2_1_U21.dout ;
assign \add_35s_35s_35_2_1_U21.reset  = ap_rst;
assign \add_35s_35s_35_2_1_U19.top_add_35s_35s_35_2_1_Adder_14_U.ain_s0  = \add_35s_35s_35_2_1_U19.top_add_35s_35s_35_2_1_Adder_14_U.a ;
assign \add_35s_35s_35_2_1_U19.top_add_35s_35s_35_2_1_Adder_14_U.bin_s0  = \add_35s_35s_35_2_1_U19.top_add_35s_35s_35_2_1_Adder_14_U.b ;
assign \add_35s_35s_35_2_1_U19.top_add_35s_35s_35_2_1_Adder_14_U.s  = { \add_35s_35s_35_2_1_U19.top_add_35s_35s_35_2_1_Adder_14_U.fas_s2 , \add_35s_35s_35_2_1_U19.top_add_35s_35s_35_2_1_Adder_14_U.sum_s1  };
assign \add_35s_35s_35_2_1_U19.top_add_35s_35s_35_2_1_Adder_14_U.u2.a  = \add_35s_35s_35_2_1_U19.top_add_35s_35s_35_2_1_Adder_14_U.ain_s1 ;
assign \add_35s_35s_35_2_1_U19.top_add_35s_35s_35_2_1_Adder_14_U.u2.b  = \add_35s_35s_35_2_1_U19.top_add_35s_35s_35_2_1_Adder_14_U.bin_s1 ;
assign \add_35s_35s_35_2_1_U19.top_add_35s_35s_35_2_1_Adder_14_U.u2.cin  = \add_35s_35s_35_2_1_U19.top_add_35s_35s_35_2_1_Adder_14_U.carry_s1 ;
assign \add_35s_35s_35_2_1_U19.top_add_35s_35s_35_2_1_Adder_14_U.facout_s2  = \add_35s_35s_35_2_1_U19.top_add_35s_35s_35_2_1_Adder_14_U.u2.cout ;
assign \add_35s_35s_35_2_1_U19.top_add_35s_35s_35_2_1_Adder_14_U.fas_s2  = \add_35s_35s_35_2_1_U19.top_add_35s_35s_35_2_1_Adder_14_U.u2.s ;
assign \add_35s_35s_35_2_1_U19.top_add_35s_35s_35_2_1_Adder_14_U.u1.a  = \add_35s_35s_35_2_1_U19.top_add_35s_35s_35_2_1_Adder_14_U.a [16:0];
assign \add_35s_35s_35_2_1_U19.top_add_35s_35s_35_2_1_Adder_14_U.u1.b  = \add_35s_35s_35_2_1_U19.top_add_35s_35s_35_2_1_Adder_14_U.b [16:0];
assign \add_35s_35s_35_2_1_U19.top_add_35s_35s_35_2_1_Adder_14_U.u1.cin  = 1'h0;
assign \add_35s_35s_35_2_1_U19.top_add_35s_35s_35_2_1_Adder_14_U.facout_s1  = \add_35s_35s_35_2_1_U19.top_add_35s_35s_35_2_1_Adder_14_U.u1.cout ;
assign \add_35s_35s_35_2_1_U19.top_add_35s_35s_35_2_1_Adder_14_U.fas_s1  = \add_35s_35s_35_2_1_U19.top_add_35s_35s_35_2_1_Adder_14_U.u1.s ;
assign \add_35s_35s_35_2_1_U19.top_add_35s_35s_35_2_1_Adder_14_U.a  = \add_35s_35s_35_2_1_U19.din0 ;
assign \add_35s_35s_35_2_1_U19.top_add_35s_35s_35_2_1_Adder_14_U.b  = \add_35s_35s_35_2_1_U19.din1 ;
assign \add_35s_35s_35_2_1_U19.top_add_35s_35s_35_2_1_Adder_14_U.ce  = \add_35s_35s_35_2_1_U19.ce ;
assign \add_35s_35s_35_2_1_U19.top_add_35s_35s_35_2_1_Adder_14_U.clk  = \add_35s_35s_35_2_1_U19.clk ;
assign \add_35s_35s_35_2_1_U19.top_add_35s_35s_35_2_1_Adder_14_U.reset  = \add_35s_35s_35_2_1_U19.reset ;
assign \add_35s_35s_35_2_1_U19.dout  = \add_35s_35s_35_2_1_U19.top_add_35s_35s_35_2_1_Adder_14_U.s ;
assign \add_35s_35s_35_2_1_U19.ce  = 1'h1;
assign \add_35s_35s_35_2_1_U19.clk  = ap_clk;
assign \add_35s_35s_35_2_1_U19.din0  = { select_ln353_reg_2427[11], select_ln353_reg_2427[11], select_ln353_reg_2427[11], select_ln353_reg_2427[11], select_ln353_reg_2427[11], select_ln353_reg_2427[11], select_ln353_reg_2427[11], select_ln353_reg_2427[11], select_ln353_reg_2427[11], select_ln353_reg_2427[11], select_ln353_reg_2427[11], select_ln353_reg_2427[11], select_ln353_reg_2427[11], select_ln353_reg_2427[11], select_ln353_reg_2427[11], select_ln353_reg_2427[11], select_ln353_reg_2427[11], select_ln353_reg_2427[11], select_ln353_reg_2427[11], select_ln353_reg_2427[11], select_ln353_reg_2427[11], select_ln353_reg_2427, 2'h0 };
assign \add_35s_35s_35_2_1_U19.din1  = { op_12_V_reg_2422[7], op_12_V_reg_2422[7], op_12_V_reg_2422[7], op_12_V_reg_2422[7], op_12_V_reg_2422[7], op_12_V_reg_2422[7], op_12_V_reg_2422[7], op_12_V_reg_2422[7], op_12_V_reg_2422[7], op_12_V_reg_2422[7], op_12_V_reg_2422[7], op_12_V_reg_2422[7], op_12_V_reg_2422[7], op_12_V_reg_2422[7], op_12_V_reg_2422[7], op_12_V_reg_2422[7], op_12_V_reg_2422[7], op_12_V_reg_2422[7], op_12_V_reg_2422[7], op_12_V_reg_2422[7], op_12_V_reg_2422[7], op_12_V_reg_2422[7], op_12_V_reg_2422[7], op_12_V_reg_2422[7], op_12_V_reg_2422[7], op_12_V_reg_2422[7], op_12_V_reg_2422[7], op_12_V_reg_2422 };
assign grp_fu_1510_p2 = \add_35s_35s_35_2_1_U19.dout ;
assign \add_35s_35s_35_2_1_U19.reset  = ap_rst;
assign \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_16_U.ain_s0  = \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_16_U.a ;
assign \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_16_U.bin_s0  = \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_16_U.b ;
assign \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_16_U.s  = { \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_16_U.fas_s2 , \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_16_U.sum_s1  };
assign \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_16_U.u2.a  = \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_16_U.ain_s1 ;
assign \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_16_U.u2.b  = \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_16_U.bin_s1 ;
assign \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_16_U.u2.cin  = \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_16_U.carry_s1 ;
assign \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_16_U.facout_s2  = \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_16_U.u2.cout ;
assign \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_16_U.fas_s2  = \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_16_U.u2.s ;
assign \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_16_U.u1.a  = \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_16_U.a [16:0];
assign \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_16_U.u1.b  = \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_16_U.b [16:0];
assign \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_16_U.u1.cin  = 1'h0;
assign \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_16_U.facout_s1  = \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_16_U.u1.cout ;
assign \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_16_U.fas_s1  = \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_16_U.u1.s ;
assign \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_16_U.a  = \add_34s_34s_34_2_1_U24.din0 ;
assign \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_16_U.b  = \add_34s_34s_34_2_1_U24.din1 ;
assign \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_16_U.ce  = \add_34s_34s_34_2_1_U24.ce ;
assign \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_16_U.clk  = \add_34s_34s_34_2_1_U24.clk ;
assign \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_16_U.reset  = \add_34s_34s_34_2_1_U24.reset ;
assign \add_34s_34s_34_2_1_U24.dout  = \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_16_U.s ;
assign \add_34s_34s_34_2_1_U24.ce  = 1'h1;
assign \add_34s_34s_34_2_1_U24.clk  = ap_clk;
assign \add_34s_34s_34_2_1_U24.din0  = { op_24_V_reg_2516[31], op_24_V_reg_2516, 1'h0 };
assign \add_34s_34s_34_2_1_U24.din1  = { op_15_V_reg_2322[1], op_15_V_reg_2322[1], op_15_V_reg_2322[1], op_15_V_reg_2322[1], op_15_V_reg_2322[1], op_15_V_reg_2322[1], op_15_V_reg_2322[1], op_15_V_reg_2322[1], op_15_V_reg_2322[1], op_15_V_reg_2322[1], op_15_V_reg_2322[1], op_15_V_reg_2322[1], op_15_V_reg_2322[1], op_15_V_reg_2322[1], op_15_V_reg_2322[1], op_15_V_reg_2322[1], op_15_V_reg_2322[1], op_15_V_reg_2322[1], op_15_V_reg_2322[1], op_15_V_reg_2322[1], op_15_V_reg_2322[1], op_15_V_reg_2322[1], op_15_V_reg_2322[1], op_15_V_reg_2322[1], op_15_V_reg_2322[1], op_15_V_reg_2322[1], op_15_V_reg_2322[1], op_15_V_reg_2322[1], op_15_V_reg_2322[1], op_15_V_reg_2322[1], op_15_V_reg_2322[1], op_15_V_reg_2322[1], op_15_V_reg_2322 };
assign grp_fu_1631_p2 = \add_34s_34s_34_2_1_U24.dout ;
assign \add_34s_34s_34_2_1_U24.reset  = ap_rst;
assign \add_32s_32ns_32_2_1_U29.top_add_32s_32ns_32_2_1_Adder_19_U.ain_s0  = \add_32s_32ns_32_2_1_U29.top_add_32s_32ns_32_2_1_Adder_19_U.a ;
assign \add_32s_32ns_32_2_1_U29.top_add_32s_32ns_32_2_1_Adder_19_U.bin_s0  = \add_32s_32ns_32_2_1_U29.top_add_32s_32ns_32_2_1_Adder_19_U.b ;
assign \add_32s_32ns_32_2_1_U29.top_add_32s_32ns_32_2_1_Adder_19_U.s  = { \add_32s_32ns_32_2_1_U29.top_add_32s_32ns_32_2_1_Adder_19_U.fas_s2 , \add_32s_32ns_32_2_1_U29.top_add_32s_32ns_32_2_1_Adder_19_U.sum_s1  };
assign \add_32s_32ns_32_2_1_U29.top_add_32s_32ns_32_2_1_Adder_19_U.u2.a  = \add_32s_32ns_32_2_1_U29.top_add_32s_32ns_32_2_1_Adder_19_U.ain_s1 ;
assign \add_32s_32ns_32_2_1_U29.top_add_32s_32ns_32_2_1_Adder_19_U.u2.b  = \add_32s_32ns_32_2_1_U29.top_add_32s_32ns_32_2_1_Adder_19_U.bin_s1 ;
assign \add_32s_32ns_32_2_1_U29.top_add_32s_32ns_32_2_1_Adder_19_U.u2.cin  = \add_32s_32ns_32_2_1_U29.top_add_32s_32ns_32_2_1_Adder_19_U.carry_s1 ;
assign \add_32s_32ns_32_2_1_U29.top_add_32s_32ns_32_2_1_Adder_19_U.facout_s2  = \add_32s_32ns_32_2_1_U29.top_add_32s_32ns_32_2_1_Adder_19_U.u2.cout ;
assign \add_32s_32ns_32_2_1_U29.top_add_32s_32ns_32_2_1_Adder_19_U.fas_s2  = \add_32s_32ns_32_2_1_U29.top_add_32s_32ns_32_2_1_Adder_19_U.u2.s ;
assign \add_32s_32ns_32_2_1_U29.top_add_32s_32ns_32_2_1_Adder_19_U.u1.a  = \add_32s_32ns_32_2_1_U29.top_add_32s_32ns_32_2_1_Adder_19_U.a [15:0];
assign \add_32s_32ns_32_2_1_U29.top_add_32s_32ns_32_2_1_Adder_19_U.u1.b  = \add_32s_32ns_32_2_1_U29.top_add_32s_32ns_32_2_1_Adder_19_U.b [15:0];
assign \add_32s_32ns_32_2_1_U29.top_add_32s_32ns_32_2_1_Adder_19_U.u1.cin  = 1'h0;
assign \add_32s_32ns_32_2_1_U29.top_add_32s_32ns_32_2_1_Adder_19_U.facout_s1  = \add_32s_32ns_32_2_1_U29.top_add_32s_32ns_32_2_1_Adder_19_U.u1.cout ;
assign \add_32s_32ns_32_2_1_U29.top_add_32s_32ns_32_2_1_Adder_19_U.fas_s1  = \add_32s_32ns_32_2_1_U29.top_add_32s_32ns_32_2_1_Adder_19_U.u1.s ;
assign \add_32s_32ns_32_2_1_U29.top_add_32s_32ns_32_2_1_Adder_19_U.a  = \add_32s_32ns_32_2_1_U29.din0 ;
assign \add_32s_32ns_32_2_1_U29.top_add_32s_32ns_32_2_1_Adder_19_U.b  = \add_32s_32ns_32_2_1_U29.din1 ;
assign \add_32s_32ns_32_2_1_U29.top_add_32s_32ns_32_2_1_Adder_19_U.ce  = \add_32s_32ns_32_2_1_U29.ce ;
assign \add_32s_32ns_32_2_1_U29.top_add_32s_32ns_32_2_1_Adder_19_U.clk  = \add_32s_32ns_32_2_1_U29.clk ;
assign \add_32s_32ns_32_2_1_U29.top_add_32s_32ns_32_2_1_Adder_19_U.reset  = \add_32s_32ns_32_2_1_U29.reset ;
assign \add_32s_32ns_32_2_1_U29.dout  = \add_32s_32ns_32_2_1_U29.top_add_32s_32ns_32_2_1_Adder_19_U.s ;
assign \add_32s_32ns_32_2_1_U29.ce  = 1'h1;
assign \add_32s_32ns_32_2_1_U29.clk  = ap_clk;
assign \add_32s_32ns_32_2_1_U29.din0  = { add_ln69_2_reg_2588[16], add_ln69_2_reg_2588[16], add_ln69_2_reg_2588[16], add_ln69_2_reg_2588[16], add_ln69_2_reg_2588[16], add_ln69_2_reg_2588[16], add_ln69_2_reg_2588[16], add_ln69_2_reg_2588[16], add_ln69_2_reg_2588[16], add_ln69_2_reg_2588[16], add_ln69_2_reg_2588[16], add_ln69_2_reg_2588[16], add_ln69_2_reg_2588[16], add_ln69_2_reg_2588[16], add_ln69_2_reg_2588[16], add_ln69_2_reg_2588 };
assign \add_32s_32ns_32_2_1_U29.din1  = add_ln69_reg_2583;
assign grp_fu_1709_p2 = \add_32s_32ns_32_2_1_U29.dout ;
assign \add_32s_32ns_32_2_1_U29.reset  = ap_rst;
assign \add_32ns_32ns_32_2_1_U27.top_add_32ns_32ns_32_2_1_Adder_15_U.ain_s0  = \add_32ns_32ns_32_2_1_U27.top_add_32ns_32ns_32_2_1_Adder_15_U.a ;
assign \add_32ns_32ns_32_2_1_U27.top_add_32ns_32ns_32_2_1_Adder_15_U.bin_s0  = \add_32ns_32ns_32_2_1_U27.top_add_32ns_32ns_32_2_1_Adder_15_U.b ;
assign \add_32ns_32ns_32_2_1_U27.top_add_32ns_32ns_32_2_1_Adder_15_U.s  = { \add_32ns_32ns_32_2_1_U27.top_add_32ns_32ns_32_2_1_Adder_15_U.fas_s2 , \add_32ns_32ns_32_2_1_U27.top_add_32ns_32ns_32_2_1_Adder_15_U.sum_s1  };
assign \add_32ns_32ns_32_2_1_U27.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.a  = \add_32ns_32ns_32_2_1_U27.top_add_32ns_32ns_32_2_1_Adder_15_U.ain_s1 ;
assign \add_32ns_32ns_32_2_1_U27.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.b  = \add_32ns_32ns_32_2_1_U27.top_add_32ns_32ns_32_2_1_Adder_15_U.bin_s1 ;
assign \add_32ns_32ns_32_2_1_U27.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.cin  = \add_32ns_32ns_32_2_1_U27.top_add_32ns_32ns_32_2_1_Adder_15_U.carry_s1 ;
assign \add_32ns_32ns_32_2_1_U27.top_add_32ns_32ns_32_2_1_Adder_15_U.facout_s2  = \add_32ns_32ns_32_2_1_U27.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.cout ;
assign \add_32ns_32ns_32_2_1_U27.top_add_32ns_32ns_32_2_1_Adder_15_U.fas_s2  = \add_32ns_32ns_32_2_1_U27.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.s ;
assign \add_32ns_32ns_32_2_1_U27.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.a  = \add_32ns_32ns_32_2_1_U27.top_add_32ns_32ns_32_2_1_Adder_15_U.a [15:0];
assign \add_32ns_32ns_32_2_1_U27.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.b  = \add_32ns_32ns_32_2_1_U27.top_add_32ns_32ns_32_2_1_Adder_15_U.b [15:0];
assign \add_32ns_32ns_32_2_1_U27.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.cin  = 1'h0;
assign \add_32ns_32ns_32_2_1_U27.top_add_32ns_32ns_32_2_1_Adder_15_U.facout_s1  = \add_32ns_32ns_32_2_1_U27.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.cout ;
assign \add_32ns_32ns_32_2_1_U27.top_add_32ns_32ns_32_2_1_Adder_15_U.fas_s1  = \add_32ns_32ns_32_2_1_U27.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.s ;
assign \add_32ns_32ns_32_2_1_U27.top_add_32ns_32ns_32_2_1_Adder_15_U.a  = \add_32ns_32ns_32_2_1_U27.din0 ;
assign \add_32ns_32ns_32_2_1_U27.top_add_32ns_32ns_32_2_1_Adder_15_U.b  = \add_32ns_32ns_32_2_1_U27.din1 ;
assign \add_32ns_32ns_32_2_1_U27.top_add_32ns_32ns_32_2_1_Adder_15_U.ce  = \add_32ns_32ns_32_2_1_U27.ce ;
assign \add_32ns_32ns_32_2_1_U27.top_add_32ns_32ns_32_2_1_Adder_15_U.clk  = \add_32ns_32ns_32_2_1_U27.clk ;
assign \add_32ns_32ns_32_2_1_U27.top_add_32ns_32ns_32_2_1_Adder_15_U.reset  = \add_32ns_32ns_32_2_1_U27.reset ;
assign \add_32ns_32ns_32_2_1_U27.dout  = \add_32ns_32ns_32_2_1_U27.top_add_32ns_32ns_32_2_1_Adder_15_U.s ;
assign \add_32ns_32ns_32_2_1_U27.ce  = 1'h1;
assign \add_32ns_32ns_32_2_1_U27.clk  = ap_clk;
assign \add_32ns_32ns_32_2_1_U27.din0  = ret_V_26_reg_2558;
assign \add_32ns_32ns_32_2_1_U27.din1  = op_17;
assign grp_fu_1692_p2 = \add_32ns_32ns_32_2_1_U27.dout ;
assign \add_32ns_32ns_32_2_1_U27.reset  = ap_rst;
assign \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.ain_s0  = \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.a ;
assign \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.bin_s0  = \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.b ;
assign \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.s  = { \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.fas_s2 , \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.sum_s1  };
assign \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.a  = \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.ain_s1 ;
assign \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.b  = \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.bin_s1 ;
assign \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.cin  = \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.carry_s1 ;
assign \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.facout_s2  = \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.cout ;
assign \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.fas_s2  = \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.s ;
assign \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.a  = \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.a [15:0];
assign \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.b  = \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.b [15:0];
assign \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.cin  = 1'h0;
assign \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.facout_s1  = \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.cout ;
assign \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.fas_s1  = \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.s ;
assign \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.a  = \add_32ns_32ns_32_2_1_U25.din0 ;
assign \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.b  = \add_32ns_32ns_32_2_1_U25.din1 ;
assign \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.ce  = \add_32ns_32ns_32_2_1_U25.ce ;
assign \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.clk  = \add_32ns_32ns_32_2_1_U25.clk ;
assign \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.reset  = \add_32ns_32ns_32_2_1_U25.reset ;
assign \add_32ns_32ns_32_2_1_U25.dout  = \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.s ;
assign \add_32ns_32ns_32_2_1_U25.ce  = 1'h1;
assign \add_32ns_32ns_32_2_1_U25.clk  = ap_clk;
assign \add_32ns_32ns_32_2_1_U25.din0  = ret_V_23_cast_reg_2536;
assign \add_32ns_32ns_32_2_1_U25.din1  = 32'd1;
assign grp_fu_1647_p2 = \add_32ns_32ns_32_2_1_U25.dout ;
assign \add_32ns_32ns_32_2_1_U25.reset  = ap_rst;
assign \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.ain_s0  = \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.a ;
assign \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.bin_s0  = \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.b ;
assign \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.s  = { \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.fas_s2 , \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.sum_s1  };
assign \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.a  = \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.ain_s1 ;
assign \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.b  = \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.bin_s1 ;
assign \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.cin  = \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.carry_s1 ;
assign \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.facout_s2  = \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.cout ;
assign \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.fas_s2  = \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.s ;
assign \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.a  = \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.a [15:0];
assign \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.b  = \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.b [15:0];
assign \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.cin  = 1'h0;
assign \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.facout_s1  = \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.cout ;
assign \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.fas_s1  = \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.s ;
assign \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.a  = \add_32ns_32ns_32_2_1_U23.din0 ;
assign \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.b  = \add_32ns_32ns_32_2_1_U23.din1 ;
assign \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.ce  = \add_32ns_32ns_32_2_1_U23.ce ;
assign \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.clk  = \add_32ns_32ns_32_2_1_U23.clk ;
assign \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.reset  = \add_32ns_32ns_32_2_1_U23.reset ;
assign \add_32ns_32ns_32_2_1_U23.dout  = \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.s ;
assign \add_32ns_32ns_32_2_1_U23.ce  = 1'h1;
assign \add_32ns_32ns_32_2_1_U23.clk  = ap_clk;
assign \add_32ns_32ns_32_2_1_U23.din0  = ret_V_24_reg_2506;
assign \add_32ns_32ns_32_2_1_U23.din1  = { 28'h0000000, ret_V_20_reg_2437 };
assign grp_fu_1612_p2 = \add_32ns_32ns_32_2_1_U23.dout ;
assign \add_32ns_32ns_32_2_1_U23.reset  = ap_rst;
assign \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_15_U.ain_s0  = \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_15_U.a ;
assign \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_15_U.bin_s0  = \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_15_U.b ;
assign \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_15_U.s  = { \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_15_U.fas_s2 , \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_15_U.sum_s1  };
assign \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.a  = \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_15_U.ain_s1 ;
assign \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.b  = \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_15_U.bin_s1 ;
assign \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.cin  = \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_15_U.carry_s1 ;
assign \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_15_U.facout_s2  = \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.cout ;
assign \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_15_U.fas_s2  = \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.s ;
assign \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.a  = \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_15_U.a [15:0];
assign \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.b  = \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_15_U.b [15:0];
assign \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.cin  = 1'h0;
assign \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_15_U.facout_s1  = \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.cout ;
assign \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_15_U.fas_s1  = \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.s ;
assign \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_15_U.a  = \add_32ns_32ns_32_2_1_U22.din0 ;
assign \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_15_U.b  = \add_32ns_32ns_32_2_1_U22.din1 ;
assign \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_15_U.ce  = \add_32ns_32ns_32_2_1_U22.ce ;
assign \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_15_U.clk  = \add_32ns_32ns_32_2_1_U22.clk ;
assign \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_15_U.reset  = \add_32ns_32ns_32_2_1_U22.reset ;
assign \add_32ns_32ns_32_2_1_U22.dout  = \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_15_U.s ;
assign \add_32ns_32ns_32_2_1_U22.ce  = 1'h1;
assign \add_32ns_32ns_32_2_1_U22.clk  = ap_clk;
assign \add_32ns_32ns_32_2_1_U22.din0  = ret_V_20_cast_reg_2494;
assign \add_32ns_32ns_32_2_1_U22.din1  = 32'd1;
assign grp_fu_1585_p2 = \add_32ns_32ns_32_2_1_U22.dout ;
assign \add_32ns_32ns_32_2_1_U22.reset  = ap_rst;
assign \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_15_U.ain_s0  = \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_15_U.a ;
assign \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_15_U.bin_s0  = \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_15_U.b ;
assign \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_15_U.s  = { \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_15_U.fas_s2 , \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_15_U.sum_s1  };
assign \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.a  = \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_15_U.ain_s1 ;
assign \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.b  = \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_15_U.bin_s1 ;
assign \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.cin  = \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_15_U.carry_s1 ;
assign \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_15_U.facout_s2  = \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.cout ;
assign \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_15_U.fas_s2  = \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.s ;
assign \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.a  = \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_15_U.a [15:0];
assign \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.b  = \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_15_U.b [15:0];
assign \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.cin  = 1'h0;
assign \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_15_U.facout_s1  = \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.cout ;
assign \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_15_U.fas_s1  = \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.s ;
assign \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_15_U.a  = \add_32ns_32ns_32_2_1_U20.din0 ;
assign \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_15_U.b  = \add_32ns_32ns_32_2_1_U20.din1 ;
assign \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_15_U.ce  = \add_32ns_32ns_32_2_1_U20.ce ;
assign \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_15_U.clk  = \add_32ns_32ns_32_2_1_U20.clk ;
assign \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_15_U.reset  = \add_32ns_32ns_32_2_1_U20.reset ;
assign \add_32ns_32ns_32_2_1_U20.dout  = \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_15_U.s ;
assign \add_32ns_32ns_32_2_1_U20.ce  = 1'h1;
assign \add_32ns_32ns_32_2_1_U20.clk  = ap_clk;
assign \add_32ns_32ns_32_2_1_U20.din0  = ret_V_17_cast_reg_2462;
assign \add_32ns_32ns_32_2_1_U20.din1  = 32'd1;
assign grp_fu_1531_p2 = \add_32ns_32ns_32_2_1_U20.dout ;
assign \add_32ns_32ns_32_2_1_U20.reset  = ap_rst;
assign \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.ain_s0  = \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.a ;
assign \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.bin_s0  = \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.b ;
assign \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.s  = { \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.fas_s2 , \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.sum_s1  };
assign \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.u2.a  = \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.ain_s1 ;
assign \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.u2.b  = \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.bin_s1 ;
assign \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.u2.cin  = \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.carry_s1 ;
assign \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.facout_s2  = \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.u2.cout ;
assign \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.fas_s2  = \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.u2.s ;
assign \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.u1.a  = \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.a [0];
assign \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.u1.b  = \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.b [0];
assign \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.u1.cin  = 1'h0;
assign \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.facout_s1  = \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.u1.cout ;
assign \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.fas_s1  = \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.u1.s ;
assign \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.a  = \add_2ns_2ns_2_2_1_U9.din0 ;
assign \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.b  = \add_2ns_2ns_2_2_1_U9.din1 ;
assign \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.ce  = \add_2ns_2ns_2_2_1_U9.ce ;
assign \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.clk  = \add_2ns_2ns_2_2_1_U9.clk ;
assign \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.reset  = \add_2ns_2ns_2_2_1_U9.reset ;
assign \add_2ns_2ns_2_2_1_U9.dout  = \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_6_U.s ;
assign \add_2ns_2ns_2_2_1_U9.ce  = 1'h1;
assign \add_2ns_2ns_2_2_1_U9.clk  = ap_clk;
assign \add_2ns_2ns_2_2_1_U9.din0  = p_Val2_5_reg_1961;
assign \add_2ns_2ns_2_2_1_U9.din1  = { 1'h0, and_ln412_reg_2020 };
assign grp_fu_773_p2 = \add_2ns_2ns_2_2_1_U9.dout ;
assign \add_2ns_2ns_2_2_1_U9.reset  = ap_rst;
assign \add_24s_24s_24_2_1_U16.top_add_24s_24s_24_2_1_Adder_12_U.ain_s0  = \add_24s_24s_24_2_1_U16.top_add_24s_24s_24_2_1_Adder_12_U.a ;
assign \add_24s_24s_24_2_1_U16.top_add_24s_24s_24_2_1_Adder_12_U.bin_s0  = \add_24s_24s_24_2_1_U16.top_add_24s_24s_24_2_1_Adder_12_U.b ;
assign \add_24s_24s_24_2_1_U16.top_add_24s_24s_24_2_1_Adder_12_U.s  = { \add_24s_24s_24_2_1_U16.top_add_24s_24s_24_2_1_Adder_12_U.fas_s2 , \add_24s_24s_24_2_1_U16.top_add_24s_24s_24_2_1_Adder_12_U.sum_s1  };
assign \add_24s_24s_24_2_1_U16.top_add_24s_24s_24_2_1_Adder_12_U.u2.a  = \add_24s_24s_24_2_1_U16.top_add_24s_24s_24_2_1_Adder_12_U.ain_s1 ;
assign \add_24s_24s_24_2_1_U16.top_add_24s_24s_24_2_1_Adder_12_U.u2.b  = \add_24s_24s_24_2_1_U16.top_add_24s_24s_24_2_1_Adder_12_U.bin_s1 ;
assign \add_24s_24s_24_2_1_U16.top_add_24s_24s_24_2_1_Adder_12_U.u2.cin  = \add_24s_24s_24_2_1_U16.top_add_24s_24s_24_2_1_Adder_12_U.carry_s1 ;
assign \add_24s_24s_24_2_1_U16.top_add_24s_24s_24_2_1_Adder_12_U.facout_s2  = \add_24s_24s_24_2_1_U16.top_add_24s_24s_24_2_1_Adder_12_U.u2.cout ;
assign \add_24s_24s_24_2_1_U16.top_add_24s_24s_24_2_1_Adder_12_U.fas_s2  = \add_24s_24s_24_2_1_U16.top_add_24s_24s_24_2_1_Adder_12_U.u2.s ;
assign \add_24s_24s_24_2_1_U16.top_add_24s_24s_24_2_1_Adder_12_U.u1.a  = \add_24s_24s_24_2_1_U16.top_add_24s_24s_24_2_1_Adder_12_U.a [11:0];
assign \add_24s_24s_24_2_1_U16.top_add_24s_24s_24_2_1_Adder_12_U.u1.b  = \add_24s_24s_24_2_1_U16.top_add_24s_24s_24_2_1_Adder_12_U.b [11:0];
assign \add_24s_24s_24_2_1_U16.top_add_24s_24s_24_2_1_Adder_12_U.u1.cin  = 1'h0;
assign \add_24s_24s_24_2_1_U16.top_add_24s_24s_24_2_1_Adder_12_U.facout_s1  = \add_24s_24s_24_2_1_U16.top_add_24s_24s_24_2_1_Adder_12_U.u1.cout ;
assign \add_24s_24s_24_2_1_U16.top_add_24s_24s_24_2_1_Adder_12_U.fas_s1  = \add_24s_24s_24_2_1_U16.top_add_24s_24s_24_2_1_Adder_12_U.u1.s ;
assign \add_24s_24s_24_2_1_U16.top_add_24s_24s_24_2_1_Adder_12_U.a  = \add_24s_24s_24_2_1_U16.din0 ;
assign \add_24s_24s_24_2_1_U16.top_add_24s_24s_24_2_1_Adder_12_U.b  = \add_24s_24s_24_2_1_U16.din1 ;
assign \add_24s_24s_24_2_1_U16.top_add_24s_24s_24_2_1_Adder_12_U.ce  = \add_24s_24s_24_2_1_U16.ce ;
assign \add_24s_24s_24_2_1_U16.top_add_24s_24s_24_2_1_Adder_12_U.clk  = \add_24s_24s_24_2_1_U16.clk ;
assign \add_24s_24s_24_2_1_U16.top_add_24s_24s_24_2_1_Adder_12_U.reset  = \add_24s_24s_24_2_1_U16.reset ;
assign \add_24s_24s_24_2_1_U16.dout  = \add_24s_24s_24_2_1_U16.top_add_24s_24s_24_2_1_Adder_12_U.s ;
assign \add_24s_24s_24_2_1_U16.ce  = 1'h1;
assign \add_24s_24s_24_2_1_U16.clk  = ap_clk;
assign \add_24s_24s_24_2_1_U16.din0  = { select_ln850_4_reg_2264[9], select_ln850_4_reg_2264, 13'h0000 };
assign \add_24s_24s_24_2_1_U16.din1  = { op_11[15], op_11[15], op_11[15], op_11[15], op_11[15], op_11[15], op_11[15], op_11[15], op_11 };
assign grp_fu_1181_p2 = \add_24s_24s_24_2_1_U16.dout ;
assign \add_24s_24s_24_2_1_U16.reset  = ap_rst;
assign \add_17s_17s_17_2_1_U28.top_add_17s_17s_17_2_1_Adder_18_U.ain_s0  = \add_17s_17s_17_2_1_U28.top_add_17s_17s_17_2_1_Adder_18_U.a ;
assign \add_17s_17s_17_2_1_U28.top_add_17s_17s_17_2_1_Adder_18_U.bin_s0  = \add_17s_17s_17_2_1_U28.top_add_17s_17s_17_2_1_Adder_18_U.b ;
assign \add_17s_17s_17_2_1_U28.top_add_17s_17s_17_2_1_Adder_18_U.s  = { \add_17s_17s_17_2_1_U28.top_add_17s_17s_17_2_1_Adder_18_U.fas_s2 , \add_17s_17s_17_2_1_U28.top_add_17s_17s_17_2_1_Adder_18_U.sum_s1  };
assign \add_17s_17s_17_2_1_U28.top_add_17s_17s_17_2_1_Adder_18_U.u2.a  = \add_17s_17s_17_2_1_U28.top_add_17s_17s_17_2_1_Adder_18_U.ain_s1 ;
assign \add_17s_17s_17_2_1_U28.top_add_17s_17s_17_2_1_Adder_18_U.u2.b  = \add_17s_17s_17_2_1_U28.top_add_17s_17s_17_2_1_Adder_18_U.bin_s1 ;
assign \add_17s_17s_17_2_1_U28.top_add_17s_17s_17_2_1_Adder_18_U.u2.cin  = \add_17s_17s_17_2_1_U28.top_add_17s_17s_17_2_1_Adder_18_U.carry_s1 ;
assign \add_17s_17s_17_2_1_U28.top_add_17s_17s_17_2_1_Adder_18_U.facout_s2  = \add_17s_17s_17_2_1_U28.top_add_17s_17s_17_2_1_Adder_18_U.u2.cout ;
assign \add_17s_17s_17_2_1_U28.top_add_17s_17s_17_2_1_Adder_18_U.fas_s2  = \add_17s_17s_17_2_1_U28.top_add_17s_17s_17_2_1_Adder_18_U.u2.s ;
assign \add_17s_17s_17_2_1_U28.top_add_17s_17s_17_2_1_Adder_18_U.u1.a  = \add_17s_17s_17_2_1_U28.top_add_17s_17s_17_2_1_Adder_18_U.a [7:0];
assign \add_17s_17s_17_2_1_U28.top_add_17s_17s_17_2_1_Adder_18_U.u1.b  = \add_17s_17s_17_2_1_U28.top_add_17s_17s_17_2_1_Adder_18_U.b [7:0];
assign \add_17s_17s_17_2_1_U28.top_add_17s_17s_17_2_1_Adder_18_U.u1.cin  = 1'h0;
assign \add_17s_17s_17_2_1_U28.top_add_17s_17s_17_2_1_Adder_18_U.facout_s1  = \add_17s_17s_17_2_1_U28.top_add_17s_17s_17_2_1_Adder_18_U.u1.cout ;
assign \add_17s_17s_17_2_1_U28.top_add_17s_17s_17_2_1_Adder_18_U.fas_s1  = \add_17s_17s_17_2_1_U28.top_add_17s_17s_17_2_1_Adder_18_U.u1.s ;
assign \add_17s_17s_17_2_1_U28.top_add_17s_17s_17_2_1_Adder_18_U.a  = \add_17s_17s_17_2_1_U28.din0 ;
assign \add_17s_17s_17_2_1_U28.top_add_17s_17s_17_2_1_Adder_18_U.b  = \add_17s_17s_17_2_1_U28.din1 ;
assign \add_17s_17s_17_2_1_U28.top_add_17s_17s_17_2_1_Adder_18_U.ce  = \add_17s_17s_17_2_1_U28.ce ;
assign \add_17s_17s_17_2_1_U28.top_add_17s_17s_17_2_1_Adder_18_U.clk  = \add_17s_17s_17_2_1_U28.clk ;
assign \add_17s_17s_17_2_1_U28.top_add_17s_17s_17_2_1_Adder_18_U.reset  = \add_17s_17s_17_2_1_U28.reset ;
assign \add_17s_17s_17_2_1_U28.dout  = \add_17s_17s_17_2_1_U28.top_add_17s_17s_17_2_1_Adder_18_U.s ;
assign \add_17s_17s_17_2_1_U28.ce  = 1'h1;
assign \add_17s_17s_17_2_1_U28.clk  = ap_clk;
assign \add_17s_17s_17_2_1_U28.din0  = { add_ln69_1_reg_2563[8], add_ln69_1_reg_2563[8], add_ln69_1_reg_2563[8], add_ln69_1_reg_2563[8], add_ln69_1_reg_2563[8], add_ln69_1_reg_2563[8], add_ln69_1_reg_2563[8], add_ln69_1_reg_2563[8], add_ln69_1_reg_2563 };
assign \add_17s_17s_17_2_1_U28.din1  = { op_16[15], op_16 };
assign grp_fu_1700_p2 = \add_17s_17s_17_2_1_U28.dout ;
assign \add_17s_17s_17_2_1_U28.reset  = ap_rst;
assign \add_13ns_13s_13_2_1_U10.top_add_13ns_13s_13_2_1_Adder_7_U.ain_s0  = \add_13ns_13s_13_2_1_U10.top_add_13ns_13s_13_2_1_Adder_7_U.a ;
assign \add_13ns_13s_13_2_1_U10.top_add_13ns_13s_13_2_1_Adder_7_U.bin_s0  = \add_13ns_13s_13_2_1_U10.top_add_13ns_13s_13_2_1_Adder_7_U.b ;
assign \add_13ns_13s_13_2_1_U10.top_add_13ns_13s_13_2_1_Adder_7_U.s  = { \add_13ns_13s_13_2_1_U10.top_add_13ns_13s_13_2_1_Adder_7_U.fas_s2 , \add_13ns_13s_13_2_1_U10.top_add_13ns_13s_13_2_1_Adder_7_U.sum_s1  };
assign \add_13ns_13s_13_2_1_U10.top_add_13ns_13s_13_2_1_Adder_7_U.u2.a  = \add_13ns_13s_13_2_1_U10.top_add_13ns_13s_13_2_1_Adder_7_U.ain_s1 ;
assign \add_13ns_13s_13_2_1_U10.top_add_13ns_13s_13_2_1_Adder_7_U.u2.b  = \add_13ns_13s_13_2_1_U10.top_add_13ns_13s_13_2_1_Adder_7_U.bin_s1 ;
assign \add_13ns_13s_13_2_1_U10.top_add_13ns_13s_13_2_1_Adder_7_U.u2.cin  = \add_13ns_13s_13_2_1_U10.top_add_13ns_13s_13_2_1_Adder_7_U.carry_s1 ;
assign \add_13ns_13s_13_2_1_U10.top_add_13ns_13s_13_2_1_Adder_7_U.facout_s2  = \add_13ns_13s_13_2_1_U10.top_add_13ns_13s_13_2_1_Adder_7_U.u2.cout ;
assign \add_13ns_13s_13_2_1_U10.top_add_13ns_13s_13_2_1_Adder_7_U.fas_s2  = \add_13ns_13s_13_2_1_U10.top_add_13ns_13s_13_2_1_Adder_7_U.u2.s ;
assign \add_13ns_13s_13_2_1_U10.top_add_13ns_13s_13_2_1_Adder_7_U.u1.a  = \add_13ns_13s_13_2_1_U10.top_add_13ns_13s_13_2_1_Adder_7_U.a [5:0];
assign \add_13ns_13s_13_2_1_U10.top_add_13ns_13s_13_2_1_Adder_7_U.u1.b  = \add_13ns_13s_13_2_1_U10.top_add_13ns_13s_13_2_1_Adder_7_U.b [5:0];
assign \add_13ns_13s_13_2_1_U10.top_add_13ns_13s_13_2_1_Adder_7_U.u1.cin  = 1'h0;
assign \add_13ns_13s_13_2_1_U10.top_add_13ns_13s_13_2_1_Adder_7_U.facout_s1  = \add_13ns_13s_13_2_1_U10.top_add_13ns_13s_13_2_1_Adder_7_U.u1.cout ;
assign \add_13ns_13s_13_2_1_U10.top_add_13ns_13s_13_2_1_Adder_7_U.fas_s1  = \add_13ns_13s_13_2_1_U10.top_add_13ns_13s_13_2_1_Adder_7_U.u1.s ;
assign \add_13ns_13s_13_2_1_U10.top_add_13ns_13s_13_2_1_Adder_7_U.a  = \add_13ns_13s_13_2_1_U10.din0 ;
assign \add_13ns_13s_13_2_1_U10.top_add_13ns_13s_13_2_1_Adder_7_U.b  = \add_13ns_13s_13_2_1_U10.din1 ;
assign \add_13ns_13s_13_2_1_U10.top_add_13ns_13s_13_2_1_Adder_7_U.ce  = \add_13ns_13s_13_2_1_U10.ce ;
assign \add_13ns_13s_13_2_1_U10.top_add_13ns_13s_13_2_1_Adder_7_U.clk  = \add_13ns_13s_13_2_1_U10.clk ;
assign \add_13ns_13s_13_2_1_U10.top_add_13ns_13s_13_2_1_Adder_7_U.reset  = \add_13ns_13s_13_2_1_U10.reset ;
assign \add_13ns_13s_13_2_1_U10.dout  = \add_13ns_13s_13_2_1_U10.top_add_13ns_13s_13_2_1_Adder_7_U.s ;
assign \add_13ns_13s_13_2_1_U10.ce  = 1'h1;
assign \add_13ns_13s_13_2_1_U10.clk  = ap_clk;
assign \add_13ns_13s_13_2_1_U10.din0  = { 2'h0, op_10_V_reg_2047, 3'h0 };
assign \add_13ns_13s_13_2_1_U10.din1  = { op_6[7], op_6[7], op_6[7], op_6[7], op_6[7], op_6 };
assign grp_fu_820_p2 = \add_13ns_13s_13_2_1_U10.dout ;
assign \add_13ns_13s_13_2_1_U10.reset  = ap_rst;
assign \add_12s_12ns_12_2_1_U17.top_add_12s_12ns_12_2_1_Adder_13_U.ain_s0  = \add_12s_12ns_12_2_1_U17.top_add_12s_12ns_12_2_1_Adder_13_U.a ;
assign \add_12s_12ns_12_2_1_U17.top_add_12s_12ns_12_2_1_Adder_13_U.bin_s0  = \add_12s_12ns_12_2_1_U17.top_add_12s_12ns_12_2_1_Adder_13_U.b ;
assign \add_12s_12ns_12_2_1_U17.top_add_12s_12ns_12_2_1_Adder_13_U.s  = { \add_12s_12ns_12_2_1_U17.top_add_12s_12ns_12_2_1_Adder_13_U.fas_s2 , \add_12s_12ns_12_2_1_U17.top_add_12s_12ns_12_2_1_Adder_13_U.sum_s1  };
assign \add_12s_12ns_12_2_1_U17.top_add_12s_12ns_12_2_1_Adder_13_U.u2.a  = \add_12s_12ns_12_2_1_U17.top_add_12s_12ns_12_2_1_Adder_13_U.ain_s1 ;
assign \add_12s_12ns_12_2_1_U17.top_add_12s_12ns_12_2_1_Adder_13_U.u2.b  = \add_12s_12ns_12_2_1_U17.top_add_12s_12ns_12_2_1_Adder_13_U.bin_s1 ;
assign \add_12s_12ns_12_2_1_U17.top_add_12s_12ns_12_2_1_Adder_13_U.u2.cin  = \add_12s_12ns_12_2_1_U17.top_add_12s_12ns_12_2_1_Adder_13_U.carry_s1 ;
assign \add_12s_12ns_12_2_1_U17.top_add_12s_12ns_12_2_1_Adder_13_U.facout_s2  = \add_12s_12ns_12_2_1_U17.top_add_12s_12ns_12_2_1_Adder_13_U.u2.cout ;
assign \add_12s_12ns_12_2_1_U17.top_add_12s_12ns_12_2_1_Adder_13_U.fas_s2  = \add_12s_12ns_12_2_1_U17.top_add_12s_12ns_12_2_1_Adder_13_U.u2.s ;
assign \add_12s_12ns_12_2_1_U17.top_add_12s_12ns_12_2_1_Adder_13_U.u1.a  = \add_12s_12ns_12_2_1_U17.top_add_12s_12ns_12_2_1_Adder_13_U.a [5:0];
assign \add_12s_12ns_12_2_1_U17.top_add_12s_12ns_12_2_1_Adder_13_U.u1.b  = \add_12s_12ns_12_2_1_U17.top_add_12s_12ns_12_2_1_Adder_13_U.b [5:0];
assign \add_12s_12ns_12_2_1_U17.top_add_12s_12ns_12_2_1_Adder_13_U.u1.cin  = 1'h0;
assign \add_12s_12ns_12_2_1_U17.top_add_12s_12ns_12_2_1_Adder_13_U.facout_s1  = \add_12s_12ns_12_2_1_U17.top_add_12s_12ns_12_2_1_Adder_13_U.u1.cout ;
assign \add_12s_12ns_12_2_1_U17.top_add_12s_12ns_12_2_1_Adder_13_U.fas_s1  = \add_12s_12ns_12_2_1_U17.top_add_12s_12ns_12_2_1_Adder_13_U.u1.s ;
assign \add_12s_12ns_12_2_1_U17.top_add_12s_12ns_12_2_1_Adder_13_U.a  = \add_12s_12ns_12_2_1_U17.din0 ;
assign \add_12s_12ns_12_2_1_U17.top_add_12s_12ns_12_2_1_Adder_13_U.b  = \add_12s_12ns_12_2_1_U17.din1 ;
assign \add_12s_12ns_12_2_1_U17.top_add_12s_12ns_12_2_1_Adder_13_U.ce  = \add_12s_12ns_12_2_1_U17.ce ;
assign \add_12s_12ns_12_2_1_U17.top_add_12s_12ns_12_2_1_Adder_13_U.clk  = \add_12s_12ns_12_2_1_U17.clk ;
assign \add_12s_12ns_12_2_1_U17.top_add_12s_12ns_12_2_1_Adder_13_U.reset  = \add_12s_12ns_12_2_1_U17.reset ;
assign \add_12s_12ns_12_2_1_U17.dout  = \add_12s_12ns_12_2_1_U17.top_add_12s_12ns_12_2_1_Adder_13_U.s ;
assign \add_12s_12ns_12_2_1_U17.ce  = 1'h1;
assign \add_12s_12ns_12_2_1_U17.clk  = ap_clk;
assign \add_12s_12ns_12_2_1_U17.din0  = { tmp_reg_2338[10], tmp_reg_2338 };
assign \add_12s_12ns_12_2_1_U17.din1  = 12'h001;
assign grp_fu_1314_p2 = \add_12s_12ns_12_2_1_U17.dout ;
assign \add_12s_12ns_12_2_1_U17.reset  = ap_rst;
assign \add_10ns_10ns_10_2_1_U13.top_add_10ns_10ns_10_2_1_Adder_9_U.ain_s0  = \add_10ns_10ns_10_2_1_U13.top_add_10ns_10ns_10_2_1_Adder_9_U.a ;
assign \add_10ns_10ns_10_2_1_U13.top_add_10ns_10ns_10_2_1_Adder_9_U.bin_s0  = \add_10ns_10ns_10_2_1_U13.top_add_10ns_10ns_10_2_1_Adder_9_U.b ;
assign \add_10ns_10ns_10_2_1_U13.top_add_10ns_10ns_10_2_1_Adder_9_U.s  = { \add_10ns_10ns_10_2_1_U13.top_add_10ns_10ns_10_2_1_Adder_9_U.fas_s2 , \add_10ns_10ns_10_2_1_U13.top_add_10ns_10ns_10_2_1_Adder_9_U.sum_s1  };
assign \add_10ns_10ns_10_2_1_U13.top_add_10ns_10ns_10_2_1_Adder_9_U.u2.a  = \add_10ns_10ns_10_2_1_U13.top_add_10ns_10ns_10_2_1_Adder_9_U.ain_s1 ;
assign \add_10ns_10ns_10_2_1_U13.top_add_10ns_10ns_10_2_1_Adder_9_U.u2.b  = \add_10ns_10ns_10_2_1_U13.top_add_10ns_10ns_10_2_1_Adder_9_U.bin_s1 ;
assign \add_10ns_10ns_10_2_1_U13.top_add_10ns_10ns_10_2_1_Adder_9_U.u2.cin  = \add_10ns_10ns_10_2_1_U13.top_add_10ns_10ns_10_2_1_Adder_9_U.carry_s1 ;
assign \add_10ns_10ns_10_2_1_U13.top_add_10ns_10ns_10_2_1_Adder_9_U.facout_s2  = \add_10ns_10ns_10_2_1_U13.top_add_10ns_10ns_10_2_1_Adder_9_U.u2.cout ;
assign \add_10ns_10ns_10_2_1_U13.top_add_10ns_10ns_10_2_1_Adder_9_U.fas_s2  = \add_10ns_10ns_10_2_1_U13.top_add_10ns_10ns_10_2_1_Adder_9_U.u2.s ;
assign \add_10ns_10ns_10_2_1_U13.top_add_10ns_10ns_10_2_1_Adder_9_U.u1.a  = \add_10ns_10ns_10_2_1_U13.top_add_10ns_10ns_10_2_1_Adder_9_U.a [4:0];
assign \add_10ns_10ns_10_2_1_U13.top_add_10ns_10ns_10_2_1_Adder_9_U.u1.b  = \add_10ns_10ns_10_2_1_U13.top_add_10ns_10ns_10_2_1_Adder_9_U.b [4:0];
assign \add_10ns_10ns_10_2_1_U13.top_add_10ns_10ns_10_2_1_Adder_9_U.u1.cin  = 1'h0;
assign \add_10ns_10ns_10_2_1_U13.top_add_10ns_10ns_10_2_1_Adder_9_U.facout_s1  = \add_10ns_10ns_10_2_1_U13.top_add_10ns_10ns_10_2_1_Adder_9_U.u1.cout ;
assign \add_10ns_10ns_10_2_1_U13.top_add_10ns_10ns_10_2_1_Adder_9_U.fas_s1  = \add_10ns_10ns_10_2_1_U13.top_add_10ns_10ns_10_2_1_Adder_9_U.u1.s ;
assign \add_10ns_10ns_10_2_1_U13.top_add_10ns_10ns_10_2_1_Adder_9_U.a  = \add_10ns_10ns_10_2_1_U13.din0 ;
assign \add_10ns_10ns_10_2_1_U13.top_add_10ns_10ns_10_2_1_Adder_9_U.b  = \add_10ns_10ns_10_2_1_U13.din1 ;
assign \add_10ns_10ns_10_2_1_U13.top_add_10ns_10ns_10_2_1_Adder_9_U.ce  = \add_10ns_10ns_10_2_1_U13.ce ;
assign \add_10ns_10ns_10_2_1_U13.top_add_10ns_10ns_10_2_1_Adder_9_U.clk  = \add_10ns_10ns_10_2_1_U13.clk ;
assign \add_10ns_10ns_10_2_1_U13.top_add_10ns_10ns_10_2_1_Adder_9_U.reset  = \add_10ns_10ns_10_2_1_U13.reset ;
assign \add_10ns_10ns_10_2_1_U13.dout  = \add_10ns_10ns_10_2_1_U13.top_add_10ns_10ns_10_2_1_Adder_9_U.s ;
assign \add_10ns_10ns_10_2_1_U13.ce  = 1'h1;
assign \add_10ns_10ns_10_2_1_U13.clk  = ap_clk;
assign \add_10ns_10ns_10_2_1_U13.din0  = ret_V_6_reg_2108;
assign \add_10ns_10ns_10_2_1_U13.din1  = 10'h001;
assign grp_fu_899_p2 = \add_10ns_10ns_10_2_1_U13.dout ;
assign \add_10ns_10ns_10_2_1_U13.reset  = ap_rst;
endmodule


// Machine B:
// Processed by function `add_clk_enable_signal` in `verilog_tricks.py`.
// Processed by function `remove_reset_signal` in `verilog_tricks.py`.
module top_B (
  ap_clk,
  ap_start,
  ap_done,
  ap_idle,
  ap_ready,
  op_0,
  op_6,
  op_7,
  op_8,
  op_11,
  op_16,
  op_17,
  op_18,
  op_29,
  op_29_ap_vld,
clk_enable
);
input clk_enable;


input ap_clk;
wire ap_rst;
assign ap_rst = op_29_ap_vld;
input ap_start;
input [3:0] op_0;
input [15:0] op_11;
input [15:0] op_16;
input [31:0] op_17;
input [3:0] op_18;
input [7:0] op_6;
input [15:0] op_7;
input [3:0] op_8;
output ap_done;
output ap_idle;
output ap_ready;
output [31:0] op_29;
output op_29_ap_vld;


reg [11:0] add_ln691_3_reg_2086;
reg [8:0] add_ln69_1_reg_2123;
reg and_ln786_reg_1986;
reg [10:0] ap_CS_fsm = 11'h001;
reg deleted_zeros_reg_1981;
reg icmp_ln768_1_reg_1880;
reg icmp_ln768_4_reg_2049;
reg icmp_ln786_1_reg_1885;
reg icmp_ln786_3_reg_2054;
reg icmp_ln851_2_reg_2081;
reg icmp_ln851_3_reg_2096;
reg icmp_ln851_4_reg_2065;
reg [35:0] \mul_32ns_4s_36_2_1_U1.top_mul_32ns_4s_36_2_1_Multiplier_0_U.p ;
reg [35:0] \mul_32ns_4s_36_2_1_U2.top_mul_32ns_4s_36_2_1_Multiplier_0_U.p ;
reg [7:0] op_10_V_reg_2008;
reg [7:0] op_12_V_reg_2091;
reg [15:0] op_13_V_reg_2013;
reg [7:0] op_19_V_reg_2060;
reg [3:0] op_1_V_reg_1856;
reg [31:0] op_24_V_reg_2113;
reg [3:0] op_3_V_reg_1896;
reg [31:0] p_Result_1_reg_1943;
reg p_Result_27_reg_1873;
reg p_Result_30_reg_1931;
reg p_Result_32_reg_1938;
reg p_Result_36_reg_2030;
reg p_Result_37_reg_2042;
reg [32:0] p_Result_3_reg_1948;
reg [1:0] p_Val2_6_reg_1971;
reg [35:0] r_V_5_reg_1923;
reg [35:0] r_V_6_reg_1954;
reg [2:0] r_V_reg_1891;
reg [32:0] ret_1_reg_2023;
reg [2:0] ret_V_16_reg_1862;
reg [3:0] ret_V_18_reg_1996;
reg [31:0] ret_V_20_cast_reg_2106;
reg [3:0] ret_V_20_reg_2018;
reg [23:0] ret_V_21_reg_2070;
reg [31:0] ret_V_26_reg_2118;
reg [3:0] ret_V_4_cast_reg_1959;
reg rhs_4_reg_2002;
reg [1:0] select_ln340_2_reg_1991;
reg [31:0] sext_ln1116_reg_1902;
reg [11:0] sext_ln850_reg_2075;
reg [2:0] trunc_ln1192_reg_1868;
reg [5:0] trunc_ln731_2_reg_2037;
reg [2:0] trunc_ln851_reg_1966;
reg xor_ln416_reg_1976;
reg [32:0] _215_;
wire [11:0] _000_;
wire [8:0] _001_;
wire _002_;
wire [10:0] _003_;
wire _004_;
wire _005_;
wire _006_;
wire _007_;
wire _008_;
wire _009_;
wire _010_;
wire _011_;
wire [7:0] _012_;
wire [7:0] _013_;
wire [13:0] _014_;
wire [7:0] _015_;
wire _016_;
wire [31:0] _017_;
wire [3:0] _018_;
wire [31:0] _019_;
wire _020_;
wire _021_;
wire _022_;
wire _023_;
wire _024_;
wire [32:0] _025_;
wire [1:0] _026_;
wire [35:0] _027_;
wire [35:0] _028_;
wire [2:0] _029_;
wire [32:0] _030_;
wire [2:0] _031_;
wire [3:0] _032_;
wire [31:0] _033_;
wire [3:0] _034_;
wire [23:0] _035_;
wire [32:0] _036_;
wire [31:0] _037_;
wire [3:0] _038_;
wire _039_;
wire [1:0] _040_;
wire [31:0] _041_;
wire [11:0] _042_;
wire [2:0] _043_;
wire [5:0] _044_;
wire [2:0] _045_;
wire _046_;
wire [1:0] _047_;
wire _048_;
wire _049_;
wire _050_;
wire _051_;
wire _052_;
wire _053_;
wire _054_;
wire [35:0] _055_;
wire [35:0] _056_;
wire _057_;
wire _058_;
wire _059_;
wire _060_;
wire _061_;
wire _062_;
wire _063_;
wire _064_;
wire _065_;
wire _066_;
wire _067_;
wire _068_;
wire _069_;
wire _070_;
wire _071_;
wire _072_;
wire _073_;
wire _074_;
wire _075_;
wire _076_;
wire _077_;
wire _078_;
wire _079_;
wire _080_;
wire Range1_all_ones_fu_812_p2;
wire Range1_all_zeros_fu_817_p2;
wire Range2_all_ones_fu_807_p2;
wire [4:0] add_ln1192_1_fu_486_p2;
wire [11:0] add_ln691_3_fu_1391_p2;
wire [31:0] add_ln691_4_fu_1638_p2;
wire [31:0] add_ln691_5_fu_1697_p2;
wire [31:0] add_ln691_6_fu_1787_p2;
wire [3:0] add_ln691_fu_935_p2;
wire [8:0] add_ln69_1_fu_1816_p2;
wire [16:0] add_ln69_2_fu_1834_p2;
wire [31:0] add_ln69_fu_1826_p2;
wire and_ln340_1_fu_595_p2;
wire and_ln340_2_fu_645_p2;
wire and_ln340_3_fu_1096_p2;
wire and_ln340_4_fu_1489_p2;
wire and_ln340_5_fu_1538_p2;
wire and_ln340_fu_331_p2;
wire and_ln412_fu_772_p2;
wire and_ln780_fu_843_p2;
wire and_ln781_fu_857_p2;
wire and_ln785_10_fu_1134_p2;
wire and_ln785_12_fu_1524_p2;
wire and_ln785_13_fu_1544_p2;
wire and_ln785_1_fu_369_p2;
wire and_ln785_3_fu_631_p2;
wire and_ln785_4_fu_651_p2;
wire and_ln785_6_fu_1724_p2;
wire and_ln785_7_fu_1733_p2;
wire and_ln785_9_fu_1128_p2;
wire and_ln785_fu_363_p2;
wire and_ln786_1_fu_614_p2;
wire and_ln786_2_fu_1508_p2;
wire and_ln786_fu_897_p2;
wire ap_CS_fsm_state1;
wire ap_CS_fsm_state10;
wire ap_CS_fsm_state11;
wire ap_CS_fsm_state2;
wire ap_CS_fsm_state3;
wire ap_CS_fsm_state4;
wire ap_CS_fsm_state5;
wire ap_CS_fsm_state6;
wire ap_CS_fsm_state7;
wire ap_CS_fsm_state8;
wire ap_CS_fsm_state9;
wire [10:0] ap_NS_fsm;
wire ap_clk;
wire ap_done;
wire ap_idle;
wire ap_ready;
wire ap_rst;
wire ap_start;
wire carry_1_fu_802_p2;
wire deleted_ones_fu_849_p3;
wire deleted_zeros_fu_822_p3;
wire [31:0] grp_fu_688_p0;
wire [35:0] grp_fu_688_p2;
wire [31:0] grp_fu_697_p0;
wire [35:0] grp_fu_697_p2;
wire icmp_ln768_1_fu_449_p2;
wire icmp_ln768_3_fu_1042_p2;
wire icmp_ln768_4_fu_1243_p2;
wire icmp_ln768_fu_277_p2;
wire icmp_ln786_1_fu_455_p2;
wire icmp_ln786_2_fu_1072_p2;
wire icmp_ln786_3_fu_1249_p2;
wire icmp_ln786_fu_307_p2;
wire icmp_ln851_1_fu_1317_p2;
wire icmp_ln851_2_fu_1385_p2;
wire icmp_ln851_3_fu_1574_p2;
wire icmp_ln851_4_fu_1268_p2;
wire icmp_ln851_fu_930_p2;
wire [5:0] lhs_fu_405_p3;
wire \mul_32ns_4s_36_2_1_U1.ce ;
wire \mul_32ns_4s_36_2_1_U1.clk ;
wire [31:0] \mul_32ns_4s_36_2_1_U1.din0 ;
wire [3:0] \mul_32ns_4s_36_2_1_U1.din1 ;
wire [35:0] \mul_32ns_4s_36_2_1_U1.dout ;
wire \mul_32ns_4s_36_2_1_U1.reset ;
wire [31:0] \mul_32ns_4s_36_2_1_U1.top_mul_32ns_4s_36_2_1_Multiplier_0_U.a ;
wire [3:0] \mul_32ns_4s_36_2_1_U1.top_mul_32ns_4s_36_2_1_Multiplier_0_U.b ;
wire \mul_32ns_4s_36_2_1_U1.top_mul_32ns_4s_36_2_1_Multiplier_0_U.ce ;
wire \mul_32ns_4s_36_2_1_U1.top_mul_32ns_4s_36_2_1_Multiplier_0_U.clk ;
wire [35:0] \mul_32ns_4s_36_2_1_U1.top_mul_32ns_4s_36_2_1_Multiplier_0_U.tmp_product ;
wire \mul_32ns_4s_36_2_1_U2.ce ;
wire \mul_32ns_4s_36_2_1_U2.clk ;
wire [31:0] \mul_32ns_4s_36_2_1_U2.din0 ;
wire [3:0] \mul_32ns_4s_36_2_1_U2.din1 ;
wire [35:0] \mul_32ns_4s_36_2_1_U2.dout ;
wire \mul_32ns_4s_36_2_1_U2.reset ;
wire [31:0] \mul_32ns_4s_36_2_1_U2.top_mul_32ns_4s_36_2_1_Multiplier_0_U.a ;
wire [3:0] \mul_32ns_4s_36_2_1_U2.top_mul_32ns_4s_36_2_1_Multiplier_0_U.b ;
wire \mul_32ns_4s_36_2_1_U2.top_mul_32ns_4s_36_2_1_Multiplier_0_U.ce ;
wire \mul_32ns_4s_36_2_1_U2.top_mul_32ns_4s_36_2_1_Multiplier_0_U.clk ;
wire [35:0] \mul_32ns_4s_36_2_1_U2.top_mul_32ns_4s_36_2_1_Multiplier_0_U.tmp_product ;
wire [3:0] \mul_4ns_3s_7_1_1_U3.din0 ;
wire [2:0] \mul_4ns_3s_7_1_1_U3.din1 ;
wire [6:0] \mul_4ns_3s_7_1_1_U3.dout ;
wire [3:0] \mul_4ns_3s_7_1_1_U3.top_mul_4ns_3s_7_1_1_Multiplier_1_U.a ;
wire [2:0] \mul_4ns_3s_7_1_1_U3.top_mul_4ns_3s_7_1_1_Multiplier_1_U.b ;
wire [6:0] \mul_4ns_3s_7_1_1_U3.top_mul_4ns_3s_7_1_1_Multiplier_1_U.p ;
wire neg_src_fu_869_p2;
wire [3:0] op_0;
wire [7:0] op_10_V_fu_982_p2;
wire [15:0] op_11;
wire [7:0] op_12_V_fu_1562_p3;
wire [15:0] op_13_V_fu_1140_p3;
wire [1:0] op_15_V_fu_1738_p3;
wire [15:0] op_16;
wire [31:0] op_17;
wire [3:0] op_18;
wire [7:0] op_19_V_fu_1258_p2;
wire [3:0] op_1_V_fu_375_p3;
wire [31:0] op_24_V_fu_1718_p2;
wire [31:0] op_29;
wire op_29_ap_vld;
wire [3:0] op_3_V_fu_669_p3;
wire [7:0] op_6;
wire [15:0] op_7;
wire [3:0] op_8;
wire or_ln340_1_fu_540_p2;
wire or_ln340_2_fu_903_p2;
wire or_ln340_3_fu_1084_p2;
wire or_ln340_4_fu_1436_p2;
wire or_ln340_5_fu_909_p2;
wire or_ln340_fu_319_p2;
wire or_ln785_10_fu_1519_p2;
wire or_ln785_11_fu_1550_p2;
wire or_ln785_1_fu_513_p2;
wire or_ln785_2_fu_880_p2;
wire or_ln785_3_fu_1048_p2;
wire or_ln785_4_fu_1411_p2;
wire or_ln785_5_fu_357_p2;
wire or_ln785_6_fu_626_p2;
wire or_ln785_7_fu_657_p2;
wire or_ln785_8_fu_1728_p2;
wire or_ln785_9_fu_1122_p2;
wire or_ln785_fu_283_p2;
wire or_ln786_1_fu_535_p2;
wire or_ln786_2_fu_1078_p2;
wire or_ln786_3_fu_1431_p2;
wire or_ln786_fu_313_p2;
wire overflow_1_fu_523_p2;
wire overflow_2_fu_891_p2;
wire overflow_3_fu_1060_p2;
wire overflow_4_fu_1420_p2;
wire overflow_fu_295_p2;
wire p_Result_11_fu_765_p3;
wire p_Result_13_fu_923_p3;
wire p_Result_14_fu_1305_p3;
wire p_Result_17_fu_1167_p3;
wire p_Result_18_fu_1580_p3;
wire [7:0] p_Result_22_fu_1473_p4;
wire p_Result_23_fu_1630_p3;
wire p_Result_24_fu_1690_p3;
wire p_Result_25_fu_1775_p3;
wire p_Result_26_fu_261_p2;
wire p_Result_28_fu_497_p3;
wire p_Result_29_fu_505_p3;
wire p_Result_31_fu_753_p1;
wire p_Result_33_fu_788_p3;
wire p_Result_34_fu_1004_p3;
wire p_Result_35_fu_1024_p3;
wire p_Result_38_fu_1404_p3;
wire [2:0] p_Result_4_fu_1032_p4;
wire [3:0] p_Result_7_fu_579_p4;
wire [2:0] p_Result_s_22_fu_439_p4;
wire p_Result_s_fu_243_p3;
wire [15:0] p_Val2_10_fu_1016_p3;
wire [7:0] p_Val2_14_fu_1397_p3;
wire [6:0] p_Val2_15_fu_1467_p2;
wire [3:0] p_Val2_2_fu_492_p2;
wire [2:0] p_Val2_3_fu_573_p2;
wire [1:0] p_Val2_5_fu_756_p4;
wire [1:0] p_Val2_6_fu_782_p2;
wire [3:0] p_Val2_s_fu_255_p2;
wire [3:0] r_V_7_fu_1151_p0;
wire [6:0] r_V_7_fu_1151_p00;
wire [6:0] r_V_7_fu_1151_p2;
wire [32:0] ret_1_fu_1207_p2;
wire [3:0] ret_V_10_cast_fu_1157_p4;
wire [2:0] ret_V_16_fu_397_p3;
wire [31:0] ret_V_17_cast_fu_1620_p4;
wire [6:0] ret_V_17_fu_425_p2;
wire [3:0] ret_V_18_fu_947_p3;
wire [12:0] ret_V_19_fu_1289_p2;
wire [2:0] ret_V_1_fu_383_p2;
wire [3:0] ret_V_20_fu_1193_p3;
wire [23:0] ret_V_21_fu_1361_p2;
wire [34:0] ret_V_22_fu_1614_p2;
wire [31:0] ret_V_23_cast_fu_1765_p4;
wire [34:0] ret_V_23_fu_1674_p2;
wire [34:0] ret_V_23_reg_2101;
wire [31:0] ret_V_24_fu_1708_p3;
wire [33:0] ret_V_25_fu_1759_p2;
wire [31:0] ret_V_26_fu_1801_p3;
wire [9:0] ret_V_6_fu_1295_p4;
wire [9:0] ret_V_7_fu_1323_p2;
wire [3:0] ret_V_8_fu_1179_p2;
wire [2:0] ret_V_fu_267_p4;
wire [16:0] ret_fu_998_p2;
wire [10:0] rhs_2_fu_1278_p3;
wire [22:0] rhs_3_fu_1349_p3;
wire rhs_4_fu_969_p2;
wire [33:0] rhs_5_fu_1662_p3;
wire [32:0] rhs_7_fu_1748_p3;
wire sel_tmp19_fu_663_p2;
wire sel_tmp51_fu_1556_p2;
wire [3:0] select_ln340_1_fu_601_p3;
wire [1:0] select_ln340_2_fu_915_p3;
wire [15:0] select_ln340_3_fu_1102_p3;
wire [7:0] select_ln340_4_fu_1495_p3;
wire [3:0] select_ln340_fu_337_p3;
wire [31:0] select_ln353_1_fu_1654_p3;
wire [11:0] select_ln353_fu_1595_p3;
wire [7:0] select_ln785_3_fu_1530_p3;
wire [3:0] select_ln785_fu_637_p3;
wire [3:0] select_ln850_1_fu_940_p3;
wire [3:0] select_ln850_2_fu_1185_p3;
wire [9:0] select_ln850_3_fu_1333_p3;
wire [9:0] select_ln850_4_fu_1341_p3;
wire [11:0] select_ln850_5_fu_1590_p3;
wire [31:0] select_ln850_6_fu_1702_p3;
wire [31:0] select_ln850_7_fu_1793_p3;
wire [31:0] select_ln850_8_fu_1647_p3;
wire [2:0] select_ln850_fu_389_p3;
wire [31:0] sext_ln1116_fu_677_p1;
wire [4:0] sext_ln1192_1_fu_476_p1;
wire [15:0] sext_ln1192_2_fu_1329_p0;
wire [23:0] sext_ln1192_2_fu_1329_p1;
wire [23:0] sext_ln1192_3_fu_1357_p1;
wire [34:0] sext_ln1192_4_fu_1610_p1;
wire [34:0] sext_ln1192_5_fu_1670_p1;
wire [33:0] sext_ln1192_6_fu_1755_p1;
wire [6:0] sext_ln1192_fu_413_p1;
wire [7:0] sext_ln213_fu_975_p1;
wire [8:0] sext_ln69_1_fu_1813_p1;
wire [16:0] sext_ln69_2_fu_1831_p1;
wire [31:0] sext_ln69_3_fu_1840_p1;
wire [16:0] sext_ln69_fu_1822_p1;
wire [7:0] sext_ln703_1_fu_1274_p0;
wire [12:0] sext_ln703_1_fu_1274_p1;
wire [34:0] sext_ln703_2_fu_1587_p1;
wire [34:0] sext_ln703_3_fu_1644_p1;
wire [33:0] sext_ln703_4_fu_1744_p1;
wire [6:0] sext_ln703_fu_417_p1;
wire [7:0] sext_ln727_fu_954_p1;
wire [11:0] sext_ln850_fu_1377_p1;
wire [3:0] shl_ln1192_fu_471_p2;
wire [6:0] shl_ln_fu_957_p3;
wire tmp_13_fu_830_p3;
wire [26:0] tmp_1_fu_1233_p4;
wire tmp_23_fu_1441_p3;
wire tmp_24_fu_1448_p3;
wire [13:0] tmp_26_fu_1602_p3;
wire tmp_6_fu_545_p3;
wire tmp_7_fu_553_p3;
wire [10:0] tmp_fu_1367_p4;
wire [4:0] trunc_ln1192_1_fu_479_p3;
wire [2:0] trunc_ln1192_fu_421_p1;
wire [7:0] trunc_ln213_fu_978_p1;
wire [13:0] trunc_ln731_1_fu_1012_p1;
wire [5:0] trunc_ln731_2_fu_1221_p1;
wire trunc_ln731_fu_251_p1;
wire [7:0] trunc_ln851_1_fu_1313_p0;
wire [2:0] trunc_ln851_1_fu_1313_p1;
wire trunc_ln851_2_fu_1175_p1;
wire [15:0] trunc_ln851_3_fu_1381_p0;
wire [12:0] trunc_ln851_3_fu_1381_p1;
wire [1:0] trunc_ln851_4_fu_1570_p1;
wire [1:0] trunc_ln851_5_fu_1264_p1;
wire trunc_ln851_6_fu_1783_p1;
wire [2:0] trunc_ln851_fu_749_p1;
wire xor_ln340_1_fu_589_p2;
wire xor_ln340_2_fu_1090_p2;
wire xor_ln340_3_fu_1483_p2;
wire xor_ln340_fu_325_p2;
wire xor_ln365_1_fu_567_p2;
wire xor_ln365_2_fu_1455_p2;
wire xor_ln365_3_fu_1461_p2;
wire xor_ln365_fu_561_p2;
wire xor_ln416_fu_796_p2;
wire xor_ln780_fu_837_p2;
wire xor_ln781_fu_863_p2;
wire xor_ln785_1_fu_518_p2;
wire xor_ln785_2_fu_874_p2;
wire xor_ln785_3_fu_886_p2;
wire xor_ln785_4_fu_1054_p2;
wire xor_ln785_5_fu_1415_p2;
wire xor_ln785_6_fu_351_p2;
wire xor_ln785_7_fu_620_p2;
wire xor_ln785_8_fu_1116_p2;
wire xor_ln785_9_fu_1513_p2;
wire xor_ln785_fu_289_p2;
wire xor_ln786_1_fu_529_p2;
wire xor_ln786_2_fu_1066_p2;
wire xor_ln786_3_fu_1426_p2;
wire xor_ln786_4_fu_345_p2;
wire xor_ln786_5_fu_609_p2;
wire xor_ln786_6_fu_1110_p2;
wire xor_ln786_7_fu_1503_p2;
wire xor_ln786_fu_301_p2;
wire [35:0] zext_ln1116_fu_680_p1;
wire [12:0] zext_ln1192_fu_1285_p1;
wire [32:0] zext_ln1347_1_fu_1204_p1;
wire [32:0] zext_ln1347_fu_1201_p1;
wire [7:0] zext_ln1499_fu_965_p1;
wire [16:0] zext_ln215_1_fu_994_p1;
wire [16:0] zext_ln215_fu_991_p1;
wire [1:0] zext_ln415_fu_778_p1;
wire [31:0] zext_ln69_1_fu_1715_p1;
wire [8:0] zext_ln69_2_fu_1809_p1;
wire [7:0] zext_ln69_fu_1255_p1;


assign ret_V_7_fu_1323_p2 = ret_V_19_fu_1289_p2[12:3] + 1'h1;
assign ret_V_8_fu_1179_p2 = r_V_7_fu_1151_p2[4:1] + 1'h1;
assign add_ln1192_1_fu_486_p2 = $signed({ trunc_ln1192_reg_1868, 2'h0 }) + $signed(op_1_V_reg_1856);
assign add_ln691_3_fu_1391_p2 = $signed(ret_V_21_fu_1361_p2[23:13]) + $signed(2'h1);
assign add_ln691_4_fu_1638_p2 = { ret_V_22_fu_1614_p2[34], ret_V_22_fu_1614_p2[34], ret_V_22_fu_1614_p2[34], ret_V_22_fu_1614_p2[34], ret_V_22_fu_1614_p2[34], ret_V_22_fu_1614_p2[34], ret_V_22_fu_1614_p2[34], ret_V_22_fu_1614_p2[34], ret_V_22_fu_1614_p2[34], ret_V_22_fu_1614_p2[34], ret_V_22_fu_1614_p2[34], ret_V_22_fu_1614_p2[34], ret_V_22_fu_1614_p2[34], ret_V_22_fu_1614_p2[34], ret_V_22_fu_1614_p2[34], ret_V_22_fu_1614_p2[34], ret_V_22_fu_1614_p2[34], ret_V_22_fu_1614_p2[34], ret_V_22_fu_1614_p2[34], ret_V_22_fu_1614_p2[34], ret_V_22_fu_1614_p2[13:2] } + 1'h1;
assign add_ln691_5_fu_1697_p2 = ret_V_20_cast_reg_2106 + 1'h1;
assign add_ln691_6_fu_1787_p2 = ret_V_25_fu_1759_p2[32:1] + 1'h1;
assign add_ln691_fu_935_p2 = ret_V_4_cast_reg_1959 + 1'h1;
assign add_ln69_1_fu_1816_p2 = $signed(op_19_V_reg_2060) + $signed({ 1'h0, op_18 });
assign add_ln69_2_fu_1834_p2 = $signed(add_ln69_1_reg_2123) + $signed(op_16);
assign add_ln69_fu_1826_p2 = ret_V_26_reg_2118 + op_17;
assign op_24_V_fu_1718_p2 = ret_V_24_fu_1708_p3 + ret_V_20_reg_2018;
assign op_29 = $signed(add_ln69_2_fu_1834_p2) + $signed(add_ln69_fu_1826_p2);
assign p_Val2_2_fu_492_p2 = $signed(op_1_V_reg_1856) + $signed({ op_0[1:0], 2'h0 });
assign p_Val2_6_fu_782_p2 = r_V_5_reg_1923[2:1] + and_ln412_fu_772_p2;
assign ret_V_17_fu_425_p2 = $signed({ op_0, 2'h0 }) + $signed(op_1_V_fu_375_p3);
assign ret_V_19_fu_1289_p2 = $signed({ 1'h0, op_10_V_reg_2008, 3'h0 }) + $signed(op_6);
assign ret_V_1_fu_383_p2 = op_0[3:1] + 1'h1;
assign ret_V_21_fu_1361_p2 = $signed({ select_ln850_4_fu_1341_p3, 13'h0000 }) + $signed(op_11);
assign { ret_V_22_fu_1614_p2[34], ret_V_22_fu_1614_p2[13:0] } = $signed({ select_ln353_fu_1595_p3, 2'h0 }) + $signed(op_12_V_reg_2091);
assign ret_V_23_fu_1674_p2 = $signed({ select_ln353_1_fu_1654_p3, 2'h0 }) + $signed(op_13_V_reg_2013);
assign ret_V_25_fu_1759_p2 = $signed({ op_24_V_reg_2113, 1'h0 }) + $signed(op_15_V_fu_1738_p3);
assign sel_tmp19_fu_663_p2 = xor_ln365_1_fu_567_p2 & or_ln785_7_fu_657_p2;
assign sel_tmp51_fu_1556_p2 = xor_ln365_3_fu_1461_p2 & or_ln785_11_fu_1550_p2;
assign _048_ = ap_CS_fsm[0] & _050_;
assign _049_ = ap_CS_fsm[0] & ap_start;
assign and_ln340_1_fu_595_p2 = xor_ln340_1_fu_589_p2 & or_ln786_1_fu_535_p2;
assign and_ln340_2_fu_645_p2 = or_ln786_1_fu_535_p2 & or_ln340_1_fu_540_p2;
assign and_ln340_3_fu_1096_p2 = xor_ln340_2_fu_1090_p2 & or_ln786_2_fu_1078_p2;
assign and_ln340_4_fu_1489_p2 = xor_ln340_3_fu_1483_p2 & or_ln786_3_fu_1431_p2;
assign and_ln340_5_fu_1538_p2 = or_ln786_3_fu_1431_p2 & or_ln340_4_fu_1436_p2;
assign and_ln340_fu_331_p2 = xor_ln340_fu_325_p2 & or_ln786_fu_313_p2;
assign and_ln412_fu_772_p2 = r_V_5_reg_1923[0] & r_V_5_reg_1923[1];
assign and_ln780_fu_843_p2 = xor_ln780_fu_837_p2 & Range2_all_ones_fu_807_p2;
assign and_ln781_fu_857_p2 = carry_1_fu_802_p2 & Range1_all_ones_fu_812_p2;
assign and_ln785_10_fu_1134_p2 = ret_fu_998_p2[13] & and_ln785_9_fu_1128_p2;
assign and_ln785_12_fu_1524_p2 = or_ln785_10_fu_1519_p2 & and_ln786_2_fu_1508_p2;
assign and_ln785_13_fu_1544_p2 = xor_ln785_5_fu_1415_p2 & and_ln786_2_fu_1508_p2;
assign and_ln785_1_fu_369_p2 = p_Result_26_fu_261_p2 & and_ln785_fu_363_p2;
assign and_ln785_3_fu_631_p2 = or_ln785_6_fu_626_p2 & and_ln786_1_fu_614_p2;
assign and_ln785_4_fu_651_p2 = xor_ln785_1_fu_518_p2 & and_ln786_1_fu_614_p2;
assign and_ln785_6_fu_1724_p2 = xor_ln416_reg_1976 & deleted_zeros_reg_1981;
assign and_ln785_7_fu_1733_p2 = or_ln785_8_fu_1728_p2 & and_ln786_reg_1986;
assign and_ln785_9_fu_1128_p2 = xor_ln786_6_fu_1110_p2 & or_ln785_9_fu_1122_p2;
assign and_ln785_fu_363_p2 = xor_ln786_4_fu_345_p2 & or_ln785_5_fu_357_p2;
assign and_ln786_1_fu_614_p2 = xor_ln786_5_fu_609_p2 & p_Val2_2_fu_492_p2[3];
assign and_ln786_2_fu_1508_p2 = xor_ln786_7_fu_1503_p2 & p_Result_37_reg_2042;
assign and_ln786_fu_897_p2 = p_Val2_6_fu_782_p2[1] & deleted_ones_fu_849_p3;
assign carry_1_fu_802_p2 = xor_ln416_fu_796_p2 & p_Result_32_reg_1938;
assign neg_src_fu_869_p2 = xor_ln781_fu_863_p2 & p_Result_30_reg_1931;
assign overflow_1_fu_523_p2 = xor_ln785_1_fu_518_p2 & or_ln785_1_fu_513_p2;
assign overflow_2_fu_891_p2 = xor_ln785_3_fu_886_p2 & or_ln785_2_fu_880_p2;
assign overflow_3_fu_1060_p2 = xor_ln785_4_fu_1054_p2 & or_ln785_3_fu_1048_p2;
assign overflow_4_fu_1420_p2 = xor_ln785_5_fu_1415_p2 & or_ln785_4_fu_1411_p2;
assign overflow_fu_295_p2 = xor_ln785_fu_289_p2 & or_ln785_fu_283_p2;
assign xor_ln786_1_fu_529_p2 = ~ p_Val2_2_fu_492_p2[3];
assign xor_ln785_1_fu_518_p2 = ~ p_Result_27_reg_1873;
assign xor_ln340_1_fu_589_p2 = ~ or_ln340_1_fu_540_p2;
assign xor_ln786_2_fu_1066_p2 = ~ ret_fu_998_p2[13];
assign xor_ln785_4_fu_1054_p2 = ~ ret_fu_998_p2[16];
assign xor_ln340_2_fu_1090_p2 = ~ or_ln340_3_fu_1084_p2;
assign xor_ln786_3_fu_1426_p2 = ~ p_Result_37_reg_2042;
assign xor_ln785_5_fu_1415_p2 = ~ p_Result_36_reg_2030;
assign xor_ln340_3_fu_1483_p2 = ~ or_ln340_4_fu_1436_p2;
assign xor_ln786_fu_301_p2 = ~ p_Result_26_fu_261_p2;
assign xor_ln785_fu_289_p2 = ~ op_0[3];
assign xor_ln340_fu_325_p2 = ~ or_ln340_fu_319_p2;
assign xor_ln780_fu_837_p2 = ~ r_V_5_reg_1923[3];
assign xor_ln416_fu_796_p2 = ~ p_Val2_6_fu_782_p2[1];
assign xor_ln785_8_fu_1116_p2 = ~ or_ln785_3_fu_1048_p2;
assign xor_ln786_6_fu_1110_p2 = ~ icmp_ln786_2_fu_1072_p2;
assign xor_ln786_7_fu_1503_p2 = ~ icmp_ln786_3_reg_2054;
assign xor_ln785_9_fu_1513_p2 = ~ or_ln785_4_fu_1411_p2;
assign xor_ln785_6_fu_351_p2 = ~ or_ln785_fu_283_p2;
assign xor_ln786_4_fu_345_p2 = ~ icmp_ln786_fu_307_p2;
assign xor_ln786_5_fu_609_p2 = ~ icmp_ln786_1_reg_1885;
assign xor_ln785_7_fu_620_p2 = ~ or_ln785_1_fu_513_p2;
assign xor_ln365_3_fu_1461_p2 = ~ xor_ln365_2_fu_1455_p2;
assign xor_ln781_fu_863_p2 = ~ and_ln781_fu_857_p2;
assign xor_ln365_1_fu_567_p2 = ~ xor_ln365_fu_561_p2;
assign xor_ln785_2_fu_874_p2 = ~ deleted_zeros_fu_822_p3;
assign xor_ln785_3_fu_886_p2 = ~ p_Result_30_reg_1931;
assign p_Val2_15_fu_1467_p2 = ~ { trunc_ln731_2_reg_2037[4:0], 2'h0 };
assign p_Val2_3_fu_573_p2 = ~ p_Val2_2_fu_492_p2[2:0];
assign _050_ = ~ ap_start;
assign _051_ = p_Result_3_reg_1948 == 33'h1ffffffff;
assign _052_ = ! p_Result_3_reg_1948;
assign _053_ = p_Result_1_reg_1943 == 32'd4294967295;
assign _054_ = ! op_6[2:0];
assign \mul_32ns_4s_36_2_1_U1.top_mul_32ns_4s_36_2_1_Multiplier_0_U.tmp_product  = $signed({ 1'h0, \mul_32ns_4s_36_2_1_U1.top_mul_32ns_4s_36_2_1_Multiplier_0_U.a  }) * $signed(\mul_32ns_4s_36_2_1_U1.top_mul_32ns_4s_36_2_1_Multiplier_0_U.b );
always @(posedge \mul_32ns_4s_36_2_1_U1.top_mul_32ns_4s_36_2_1_Multiplier_0_U.clk )
\mul_32ns_4s_36_2_1_U1.top_mul_32ns_4s_36_2_1_Multiplier_0_U.p  <= _055_;
assign _055_ = \mul_32ns_4s_36_2_1_U1.top_mul_32ns_4s_36_2_1_Multiplier_0_U.ce  ? \mul_32ns_4s_36_2_1_U1.top_mul_32ns_4s_36_2_1_Multiplier_0_U.tmp_product  : \mul_32ns_4s_36_2_1_U1.top_mul_32ns_4s_36_2_1_Multiplier_0_U.p ;
assign \mul_32ns_4s_36_2_1_U2.top_mul_32ns_4s_36_2_1_Multiplier_0_U.tmp_product  = $signed({ 1'h0, \mul_32ns_4s_36_2_1_U2.top_mul_32ns_4s_36_2_1_Multiplier_0_U.a  }) * $signed(\mul_32ns_4s_36_2_1_U2.top_mul_32ns_4s_36_2_1_Multiplier_0_U.b );
always @(posedge \mul_32ns_4s_36_2_1_U2.top_mul_32ns_4s_36_2_1_Multiplier_0_U.clk )
\mul_32ns_4s_36_2_1_U2.top_mul_32ns_4s_36_2_1_Multiplier_0_U.p  <= _056_;
assign _056_ = \mul_32ns_4s_36_2_1_U2.top_mul_32ns_4s_36_2_1_Multiplier_0_U.ce  ? \mul_32ns_4s_36_2_1_U2.top_mul_32ns_4s_36_2_1_Multiplier_0_U.tmp_product  : \mul_32ns_4s_36_2_1_U2.top_mul_32ns_4s_36_2_1_Multiplier_0_U.p ;
assign \mul_4ns_3s_7_1_1_U3.top_mul_4ns_3s_7_1_1_Multiplier_1_U.p  = $signed({ 1'h0, \mul_4ns_3s_7_1_1_U3.top_mul_4ns_3s_7_1_1_Multiplier_1_U.a  }) * $signed(\mul_4ns_3s_7_1_1_U3.top_mul_4ns_3s_7_1_1_Multiplier_1_U.b );
assign _057_ = { op_3_V_reg_1896[3], op_3_V_reg_1896[3], op_3_V_reg_1896[3], op_3_V_reg_1896[3], op_3_V_reg_1896 } != { ret_V_18_fu_947_p3, 3'h0 };
assign _058_ = | ret_V_17_fu_425_p2[6:4];
assign _059_ = | ret_fu_998_p2[16:14];
assign _060_ = | ret_1_fu_1207_p2[32:6];
assign _061_ = | op_0[3:1];
assign _062_ = ret_V_17_fu_425_p2[6:4] != 3'h7;
assign _063_ = ret_fu_998_p2[16:14] != 3'h7;
assign _064_ = ret_1_fu_1207_p2[32:6] != 27'h7ffffff;
assign _065_ = op_0[3:1] != 3'h7;
assign _066_ = | op_11[12:0];
assign _067_ = | op_12_V_fu_1562_p3[1:0];
assign _068_ = | op_13_V_fu_1140_p3[1:0];
assign _069_ = | trunc_ln851_reg_1966;
assign or_ln340_1_fu_540_p2 = p_Result_27_reg_1873 | overflow_1_fu_523_p2;
assign or_ln340_2_fu_903_p2 = overflow_2_fu_891_p2 | and_ln786_fu_897_p2;
assign or_ln340_3_fu_1084_p2 = ret_fu_998_p2[16] | overflow_3_fu_1060_p2;
assign or_ln340_4_fu_1436_p2 = p_Result_36_reg_2030 | overflow_4_fu_1420_p2;
assign or_ln340_5_fu_909_p2 = or_ln340_2_fu_903_p2 | neg_src_fu_869_p2;
assign or_ln340_fu_319_p2 = op_0[3] | overflow_fu_295_p2;
assign or_ln785_10_fu_1519_p2 = xor_ln785_9_fu_1513_p2 | p_Result_36_reg_2030;
assign or_ln785_11_fu_1550_p2 = and_ln785_13_fu_1544_p2 | and_ln340_5_fu_1538_p2;
assign or_ln785_1_fu_513_p2 = p_Val2_2_fu_492_p2[3] | icmp_ln768_1_reg_1880;
assign or_ln785_2_fu_880_p2 = xor_ln785_2_fu_874_p2 | p_Val2_6_fu_782_p2[1];
assign or_ln785_3_fu_1048_p2 = ret_fu_998_p2[13] | icmp_ln768_3_fu_1042_p2;
assign or_ln785_4_fu_1411_p2 = p_Result_37_reg_2042 | icmp_ln768_4_reg_2049;
assign or_ln785_5_fu_357_p2 = xor_ln785_6_fu_351_p2 | op_0[3];
assign or_ln785_6_fu_626_p2 = xor_ln785_7_fu_620_p2 | p_Result_27_reg_1873;
assign or_ln785_7_fu_657_p2 = and_ln785_4_fu_651_p2 | and_ln340_2_fu_645_p2;
assign or_ln785_8_fu_1728_p2 = p_Result_30_reg_1931 | and_ln785_6_fu_1724_p2;
assign or_ln785_9_fu_1122_p2 = xor_ln785_8_fu_1116_p2 | ret_fu_998_p2[16];
assign or_ln785_fu_283_p2 = p_Result_26_fu_261_p2 | icmp_ln768_fu_277_p2;
assign or_ln786_1_fu_535_p2 = xor_ln786_1_fu_529_p2 | icmp_ln786_1_reg_1885;
assign or_ln786_2_fu_1078_p2 = xor_ln786_2_fu_1066_p2 | icmp_ln786_2_fu_1072_p2;
assign or_ln786_3_fu_1431_p2 = xor_ln786_3_fu_1426_p2 | icmp_ln786_3_reg_2054;
assign or_ln786_fu_313_p2 = xor_ln786_fu_301_p2 | icmp_ln786_fu_307_p2;
always @(posedge ap_clk)
op_1_V_reg_1856[2:0] <= 3'h0;
always @(posedge ap_clk)
op_13_V_reg_2013[1:0] <= 2'h0;
always @(posedge ap_clk)
sext_ln1116_reg_1902 <= _041_;
always @(posedge ap_clk)
_215_ <= _036_;
assign ret_V_23_reg_2101[34:2] = _215_;
always @(posedge ap_clk)
ret_V_20_cast_reg_2106 <= _033_;
always @(posedge ap_clk)
r_V_5_reg_1923 <= _027_;
always @(posedge ap_clk)
p_Result_30_reg_1931 <= _021_;
always @(posedge ap_clk)
p_Result_32_reg_1938 <= _022_;
always @(posedge ap_clk)
p_Result_1_reg_1943 <= _019_;
always @(posedge ap_clk)
p_Result_3_reg_1948 <= _025_;
always @(posedge ap_clk)
r_V_6_reg_1954 <= _028_;
always @(posedge ap_clk)
ret_V_4_cast_reg_1959 <= _038_;
always @(posedge ap_clk)
trunc_ln851_reg_1966 <= _045_;
always @(posedge ap_clk)
op_3_V_reg_1896 <= _018_;
always @(posedge ap_clk)
op_24_V_reg_2113 <= _017_;
always @(posedge ap_clk)
op_10_V_reg_2008 <= _012_;
always @(posedge ap_clk)
op_13_V_reg_2013[15:2] <= _014_;
always @(posedge ap_clk)
ret_V_20_reg_2018 <= _034_;
always @(posedge ap_clk)
ret_1_reg_2023 <= _030_;
always @(posedge ap_clk)
p_Result_36_reg_2030 <= _023_;
always @(posedge ap_clk)
trunc_ln731_2_reg_2037 <= _044_;
always @(posedge ap_clk)
p_Result_37_reg_2042 <= _024_;
always @(posedge ap_clk)
icmp_ln768_4_reg_2049 <= _006_;
always @(posedge ap_clk)
icmp_ln786_3_reg_2054 <= _008_;
always @(posedge ap_clk)
op_19_V_reg_2060 <= _015_;
always @(posedge ap_clk)
icmp_ln851_4_reg_2065 <= _011_;
always @(posedge ap_clk)
op_1_V_reg_1856[3] <= _016_;
always @(posedge ap_clk)
ret_V_16_reg_1862 <= _031_;
always @(posedge ap_clk)
trunc_ln1192_reg_1868 <= _043_;
always @(posedge ap_clk)
p_Result_27_reg_1873 <= _020_;
always @(posedge ap_clk)
icmp_ln768_1_reg_1880 <= _005_;
always @(posedge ap_clk)
icmp_ln786_1_reg_1885 <= _007_;
always @(posedge ap_clk)
r_V_reg_1891 <= _029_;
always @(posedge ap_clk)
p_Val2_6_reg_1971 <= _026_;
always @(posedge ap_clk)
xor_ln416_reg_1976 <= _046_;
always @(posedge ap_clk)
deleted_zeros_reg_1981 <= _004_;
always @(posedge ap_clk)
and_ln786_reg_1986 <= _002_;
always @(posedge ap_clk)
select_ln340_2_reg_1991 <= _040_;
always @(posedge ap_clk)
ret_V_18_reg_1996 <= _032_;
always @(posedge ap_clk)
rhs_4_reg_2002 <= _039_;
always @(posedge ap_clk)
ret_V_26_reg_2118 <= _037_;
always @(posedge ap_clk)
add_ln69_1_reg_2123 <= _001_;
always @(posedge ap_clk)
ret_V_21_reg_2070 <= _035_;
always @(posedge ap_clk)
sext_ln850_reg_2075 <= _042_;
always @(posedge ap_clk)
icmp_ln851_2_reg_2081 <= _009_;
always @(posedge ap_clk)
add_ln691_3_reg_2086 <= _000_;
always @(posedge ap_clk)
op_12_V_reg_2091 <= _013_;
always @(posedge ap_clk)
icmp_ln851_3_reg_2096 <= _010_;
always @(posedge ap_clk)
ap_CS_fsm <= _003_;
assign _047_ = _049_ ? 2'h2 : 2'h1;
assign _070_ = ap_CS_fsm == 1'h1;
function [10:0] _263_;
input [10:0] a;
input [120:0] b;
input [10:0] s;
case (s)
11'b00000000001:
_263_ = b[10:0];
11'b00000000010:
_263_ = b[21:11];
11'b00000000100:
_263_ = b[32:22];
11'b00000001000:
_263_ = b[43:33];
11'b00000010000:
_263_ = b[54:44];
11'b00000100000:
_263_ = b[65:55];
11'b00001000000:
_263_ = b[76:66];
11'b00010000000:
_263_ = b[87:77];
11'b00100000000:
_263_ = b[98:88];
11'b01000000000:
_263_ = b[109:99];
11'b10000000000:
_263_ = b[120:110];
11'b00000000000:
_263_ = a;
default:
_263_ = 11'bx;
endcase
endfunction
assign ap_NS_fsm = _263_(11'hxxx, { 9'h000, _047_, 110'h0020080200802008020080200001 }, { _070_, _080_, _079_, _078_, _077_, _076_, _075_, _074_, _073_, _072_, _071_ });
assign _071_ = ap_CS_fsm == 11'h400;
assign _072_ = ap_CS_fsm == 10'h200;
assign _073_ = ap_CS_fsm == 9'h100;
assign _074_ = ap_CS_fsm == 8'h80;
assign _075_ = ap_CS_fsm == 7'h40;
assign _076_ = ap_CS_fsm == 6'h20;
assign _077_ = ap_CS_fsm == 5'h10;
assign _078_ = ap_CS_fsm == 4'h8;
assign _079_ = ap_CS_fsm == 3'h4;
assign _080_ = ap_CS_fsm == 2'h2;
assign op_29_ap_vld = ap_CS_fsm[10] ? 1'h1 : 1'h0;
assign ap_idle = _048_ ? 1'h1 : 1'h0;
assign _041_ = ap_CS_fsm[2] ? { ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862 } : sext_ln1116_reg_1902;
assign _033_ = ap_CS_fsm[7] ? ret_V_23_fu_1674_p2[33:2] : ret_V_20_cast_reg_2106;
assign _036_ = ap_CS_fsm[7] ? ret_V_23_fu_1674_p2[34:2] : ret_V_23_reg_2101[34:2];
assign _045_ = ap_CS_fsm[3] ? grp_fu_697_p2[2:0] : trunc_ln851_reg_1966;
assign _038_ = ap_CS_fsm[3] ? grp_fu_697_p2[6:3] : ret_V_4_cast_reg_1959;
assign _028_ = ap_CS_fsm[3] ? grp_fu_697_p2 : r_V_6_reg_1954;
assign _025_ = ap_CS_fsm[3] ? grp_fu_688_p2[35:3] : p_Result_3_reg_1948;
assign _019_ = ap_CS_fsm[3] ? grp_fu_688_p2[35:4] : p_Result_1_reg_1943;
assign _022_ = ap_CS_fsm[3] ? grp_fu_688_p2[2] : p_Result_32_reg_1938;
assign _021_ = ap_CS_fsm[3] ? grp_fu_688_p2[35] : p_Result_30_reg_1931;
assign _027_ = ap_CS_fsm[3] ? grp_fu_688_p2 : r_V_5_reg_1923;
assign _018_ = ap_CS_fsm[1] ? op_3_V_fu_669_p3 : op_3_V_reg_1896;
assign _017_ = ap_CS_fsm[8] ? op_24_V_fu_1718_p2 : op_24_V_reg_2113;
assign _011_ = ap_CS_fsm[5] ? icmp_ln851_4_fu_1268_p2 : icmp_ln851_4_reg_2065;
assign _015_ = ap_CS_fsm[5] ? op_19_V_fu_1258_p2 : op_19_V_reg_2060;
assign _008_ = ap_CS_fsm[5] ? icmp_ln786_3_fu_1249_p2 : icmp_ln786_3_reg_2054;
assign _006_ = ap_CS_fsm[5] ? icmp_ln768_4_fu_1243_p2 : icmp_ln768_4_reg_2049;
assign _024_ = ap_CS_fsm[5] ? ret_1_fu_1207_p2[5] : p_Result_37_reg_2042;
assign _044_ = ap_CS_fsm[5] ? ret_1_fu_1207_p2[5:0] : trunc_ln731_2_reg_2037;
assign _023_ = ap_CS_fsm[5] ? ret_1_fu_1207_p2[32] : p_Result_36_reg_2030;
assign _030_ = ap_CS_fsm[5] ? ret_1_fu_1207_p2 : ret_1_reg_2023;
assign _034_ = ap_CS_fsm[5] ? ret_V_20_fu_1193_p3 : ret_V_20_reg_2018;
assign _014_ = ap_CS_fsm[5] ? op_13_V_fu_1140_p3[15:2] : op_13_V_reg_2013[15:2];
assign _012_ = ap_CS_fsm[5] ? op_10_V_fu_982_p2 : op_10_V_reg_2008;
assign _029_ = ap_CS_fsm[0] ? op_1_V_fu_375_p3[3:1] : r_V_reg_1891;
assign _007_ = ap_CS_fsm[0] ? icmp_ln786_1_fu_455_p2 : icmp_ln786_1_reg_1885;
assign _005_ = ap_CS_fsm[0] ? icmp_ln768_1_fu_449_p2 : icmp_ln768_1_reg_1880;
assign _020_ = ap_CS_fsm[0] ? ret_V_17_fu_425_p2[6] : p_Result_27_reg_1873;
assign _043_ = ap_CS_fsm[0] ? op_0[2:0] : trunc_ln1192_reg_1868;
assign _031_ = ap_CS_fsm[0] ? ret_V_16_fu_397_p3 : ret_V_16_reg_1862;
assign _016_ = ap_CS_fsm[0] ? op_1_V_fu_375_p3[3] : op_1_V_reg_1856[3];
assign _039_ = ap_CS_fsm[4] ? rhs_4_fu_969_p2 : rhs_4_reg_2002;
assign _032_ = ap_CS_fsm[4] ? ret_V_18_fu_947_p3 : ret_V_18_reg_1996;
assign _040_ = ap_CS_fsm[4] ? select_ln340_2_fu_915_p3 : select_ln340_2_reg_1991;
assign _002_ = ap_CS_fsm[4] ? and_ln786_fu_897_p2 : and_ln786_reg_1986;
assign _004_ = ap_CS_fsm[4] ? deleted_zeros_fu_822_p3 : deleted_zeros_reg_1981;
assign _046_ = ap_CS_fsm[4] ? xor_ln416_fu_796_p2 : xor_ln416_reg_1976;
assign _026_ = ap_CS_fsm[4] ? p_Val2_6_fu_782_p2 : p_Val2_6_reg_1971;
assign _001_ = ap_CS_fsm[9] ? add_ln69_1_fu_1816_p2 : add_ln69_1_reg_2123;
assign _037_ = ap_CS_fsm[9] ? ret_V_26_fu_1801_p3 : ret_V_26_reg_2118;
assign _010_ = ap_CS_fsm[6] ? icmp_ln851_3_fu_1574_p2 : icmp_ln851_3_reg_2096;
assign _013_ = ap_CS_fsm[6] ? op_12_V_fu_1562_p3 : op_12_V_reg_2091;
assign _000_ = ap_CS_fsm[6] ? add_ln691_3_fu_1391_p2 : add_ln691_3_reg_2086;
assign _009_ = ap_CS_fsm[6] ? icmp_ln851_2_fu_1385_p2 : icmp_ln851_2_reg_2081;
assign _042_ = ap_CS_fsm[6] ? { ret_V_21_fu_1361_p2[23], ret_V_21_fu_1361_p2[23:13] } : sext_ln850_reg_2075;
assign _035_ = ap_CS_fsm[6] ? ret_V_21_fu_1361_p2 : ret_V_21_reg_2070;
assign _003_ = ap_rst ? 11'h001 : ap_NS_fsm;
assign ret_fu_998_p2 = ret_V_18_reg_1996 - op_7;
assign op_10_V_fu_982_p2 = $signed(ret_V_16_reg_1862) - $signed(op_7[7:0]);
assign op_19_V_fu_1258_p2 = op_7[7:0] - rhs_4_reg_2002;
assign ret_1_fu_1207_p2 = sext_ln1116_reg_1902 - rhs_4_reg_2002;
assign rhs_4_fu_969_p2 = _057_ ? 1'h1 : 1'h0;
assign select_ln340_1_fu_601_p3 = and_ln340_1_fu_595_p2 ? p_Val2_2_fu_492_p2 : { add_ln1192_1_fu_486_p2[4], p_Val2_3_fu_573_p2 };
assign select_ln340_2_fu_915_p3 = or_ln340_5_fu_909_p2 ? 2'h0 : p_Val2_6_fu_782_p2;
assign select_ln340_3_fu_1102_p3 = and_ln340_3_fu_1096_p2 ? { ret_fu_998_p2[13:0], 2'h0 } : 16'h0000;
assign select_ln340_4_fu_1495_p3 = and_ln340_4_fu_1489_p2 ? { trunc_ln731_2_reg_2037, 2'h0 } : { ret_1_reg_2023[6], p_Val2_15_fu_1467_p2 };
assign select_ln340_fu_337_p3 = and_ln340_fu_331_p2 ? { op_0[0], 3'h0 } : 4'h0;
assign select_ln353_1_fu_1654_p3 = ret_V_22_fu_1614_p2[34] ? select_ln850_8_fu_1647_p3 : { ret_V_22_fu_1614_p2[34], ret_V_22_fu_1614_p2[34], ret_V_22_fu_1614_p2[34], ret_V_22_fu_1614_p2[34], ret_V_22_fu_1614_p2[34], ret_V_22_fu_1614_p2[34], ret_V_22_fu_1614_p2[34], ret_V_22_fu_1614_p2[34], ret_V_22_fu_1614_p2[34], ret_V_22_fu_1614_p2[34], ret_V_22_fu_1614_p2[34], ret_V_22_fu_1614_p2[34], ret_V_22_fu_1614_p2[34], ret_V_22_fu_1614_p2[34], ret_V_22_fu_1614_p2[34], ret_V_22_fu_1614_p2[34], ret_V_22_fu_1614_p2[34], ret_V_22_fu_1614_p2[34], ret_V_22_fu_1614_p2[34], ret_V_22_fu_1614_p2[34], ret_V_22_fu_1614_p2[13:2] };
assign select_ln353_fu_1595_p3 = ret_V_21_reg_2070[23] ? select_ln850_5_fu_1590_p3 : sext_ln850_reg_2075;
assign select_ln785_3_fu_1530_p3 = and_ln785_12_fu_1524_p2 ? { trunc_ln731_2_reg_2037, 2'h0 } : select_ln340_4_fu_1495_p3;
assign select_ln785_fu_637_p3 = and_ln785_3_fu_631_p2 ? p_Val2_2_fu_492_p2 : select_ln340_1_fu_601_p3;
assign select_ln850_1_fu_940_p3 = icmp_ln851_fu_930_p2 ? add_ln691_fu_935_p2 : ret_V_4_cast_reg_1959;
assign select_ln850_2_fu_1185_p3 = r_V_7_fu_1151_p2[0] ? ret_V_8_fu_1179_p2 : r_V_7_fu_1151_p2[4:1];
assign select_ln850_3_fu_1333_p3 = icmp_ln851_1_fu_1317_p2 ? { 1'h1, ret_V_19_fu_1289_p2[11:3] } : ret_V_7_fu_1323_p2;
assign select_ln850_4_fu_1341_p3 = ret_V_19_fu_1289_p2[12] ? select_ln850_3_fu_1333_p3 : { 1'h0, ret_V_19_fu_1289_p2[11:3] };
assign select_ln850_5_fu_1590_p3 = icmp_ln851_2_reg_2081 ? add_ln691_3_reg_2086 : sext_ln850_reg_2075;
assign select_ln850_6_fu_1702_p3 = icmp_ln851_4_reg_2065 ? add_ln691_5_fu_1697_p2 : ret_V_20_cast_reg_2106;
assign select_ln850_7_fu_1793_p3 = op_15_V_fu_1738_p3[0] ? add_ln691_6_fu_1787_p2 : ret_V_25_fu_1759_p2[32:1];
assign select_ln850_8_fu_1647_p3 = icmp_ln851_3_reg_2096 ? add_ln691_4_fu_1638_p2 : { ret_V_22_fu_1614_p2[34], ret_V_22_fu_1614_p2[34], ret_V_22_fu_1614_p2[34], ret_V_22_fu_1614_p2[34], ret_V_22_fu_1614_p2[34], ret_V_22_fu_1614_p2[34], ret_V_22_fu_1614_p2[34], ret_V_22_fu_1614_p2[34], ret_V_22_fu_1614_p2[34], ret_V_22_fu_1614_p2[34], ret_V_22_fu_1614_p2[34], ret_V_22_fu_1614_p2[34], ret_V_22_fu_1614_p2[34], ret_V_22_fu_1614_p2[34], ret_V_22_fu_1614_p2[34], ret_V_22_fu_1614_p2[34], ret_V_22_fu_1614_p2[34], ret_V_22_fu_1614_p2[34], ret_V_22_fu_1614_p2[34], ret_V_22_fu_1614_p2[34], ret_V_22_fu_1614_p2[13:2] };
assign select_ln850_fu_389_p3 = op_0[0] ? ret_V_1_fu_383_p2 : { 1'h1, op_0[2:1] };
assign Range1_all_ones_fu_812_p2 = _051_ ? 1'h1 : 1'h0;
assign Range1_all_zeros_fu_817_p2 = _052_ ? 1'h1 : 1'h0;
assign Range2_all_ones_fu_807_p2 = _053_ ? 1'h1 : 1'h0;
assign deleted_ones_fu_849_p3 = carry_1_fu_802_p2 ? and_ln780_fu_843_p2 : Range1_all_ones_fu_812_p2;
assign deleted_zeros_fu_822_p3 = carry_1_fu_802_p2 ? Range1_all_ones_fu_812_p2 : Range1_all_zeros_fu_817_p2;
assign icmp_ln768_1_fu_449_p2 = _058_ ? 1'h1 : 1'h0;
assign icmp_ln768_3_fu_1042_p2 = _059_ ? 1'h1 : 1'h0;
assign icmp_ln768_4_fu_1243_p2 = _060_ ? 1'h1 : 1'h0;
assign icmp_ln768_fu_277_p2 = _061_ ? 1'h1 : 1'h0;
assign icmp_ln786_1_fu_455_p2 = _062_ ? 1'h1 : 1'h0;
assign icmp_ln786_2_fu_1072_p2 = _063_ ? 1'h1 : 1'h0;
assign icmp_ln786_3_fu_1249_p2 = _064_ ? 1'h1 : 1'h0;
assign icmp_ln786_fu_307_p2 = _065_ ? 1'h1 : 1'h0;
assign icmp_ln851_1_fu_1317_p2 = _054_ ? 1'h1 : 1'h0;
assign icmp_ln851_2_fu_1385_p2 = _066_ ? 1'h1 : 1'h0;
assign icmp_ln851_3_fu_1574_p2 = _067_ ? 1'h1 : 1'h0;
assign icmp_ln851_4_fu_1268_p2 = _068_ ? 1'h1 : 1'h0;
assign icmp_ln851_fu_930_p2 = _069_ ? 1'h1 : 1'h0;
assign op_12_V_fu_1562_p3 = sel_tmp51_fu_1556_p2 ? { trunc_ln731_2_reg_2037, 2'h0 } : select_ln785_3_fu_1530_p3;
assign op_13_V_fu_1140_p3 = and_ln785_10_fu_1134_p2 ? { ret_fu_998_p2[13:0], 2'h0 } : select_ln340_3_fu_1102_p3;
assign op_15_V_fu_1738_p3 = and_ln785_7_fu_1733_p2 ? p_Val2_6_reg_1971 : select_ln340_2_reg_1991;
assign op_1_V_fu_375_p3 = and_ln785_1_fu_369_p2 ? { op_0[0], 3'h0 } : select_ln340_fu_337_p3;
assign op_3_V_fu_669_p3 = sel_tmp19_fu_663_p2 ? p_Val2_2_fu_492_p2 : select_ln785_fu_637_p3;
assign p_Result_26_fu_261_p2 = op_0[0] ? 1'h1 : 1'h0;
assign ret_V_16_fu_397_p3 = op_0[3] ? select_ln850_fu_389_p3 : { 1'h0, op_0[2:1] };
assign ret_V_18_fu_947_p3 = r_V_6_reg_1954[35] ? select_ln850_1_fu_940_p3 : ret_V_4_cast_reg_1959;
assign ret_V_20_fu_1193_p3 = r_V_7_fu_1151_p2[6] ? select_ln850_2_fu_1185_p3 : r_V_7_fu_1151_p2[4:1];
assign ret_V_24_fu_1708_p3 = ret_V_23_reg_2101[34] ? select_ln850_6_fu_1702_p3 : ret_V_20_cast_reg_2106;
assign ret_V_26_fu_1801_p3 = ret_V_25_fu_1759_p2[33] ? select_ln850_7_fu_1793_p3 : ret_V_25_fu_1759_p2[32:1];
assign xor_ln365_2_fu_1455_p2 = ret_1_reg_2023[5] ^ ret_1_reg_2023[6];
assign xor_ln365_fu_561_p2 = p_Val2_2_fu_492_p2[3] ^ add_ln1192_1_fu_486_p2[4];
assign ap_CS_fsm_state1 = ap_CS_fsm[0];
assign ap_CS_fsm_state10 = ap_CS_fsm[9];
assign ap_CS_fsm_state11 = ap_CS_fsm[10];
assign ap_CS_fsm_state2 = ap_CS_fsm[1];
assign ap_CS_fsm_state3 = ap_CS_fsm[2];
assign ap_CS_fsm_state4 = ap_CS_fsm[3];
assign ap_CS_fsm_state5 = ap_CS_fsm[4];
assign ap_CS_fsm_state6 = ap_CS_fsm[5];
assign ap_CS_fsm_state7 = ap_CS_fsm[6];
assign ap_CS_fsm_state8 = ap_CS_fsm[7];
assign ap_CS_fsm_state9 = ap_CS_fsm[8];
assign ap_done = op_29_ap_vld;
assign ap_ready = op_29_ap_vld;
assign grp_fu_688_p0 = { ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862 };
assign grp_fu_697_p0 = { ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862 };
assign lhs_fu_405_p3 = { op_0, 2'h0 };
assign p_Result_11_fu_765_p3 = r_V_5_reg_1923[1];
assign p_Result_13_fu_923_p3 = r_V_6_reg_1954[35];
assign p_Result_14_fu_1305_p3 = ret_V_19_fu_1289_p2[12];
assign p_Result_17_fu_1167_p3 = r_V_7_fu_1151_p2[6];
assign p_Result_18_fu_1580_p3 = ret_V_21_reg_2070[23];
assign p_Result_22_fu_1473_p4 = { ret_1_reg_2023[6], p_Val2_15_fu_1467_p2 };
assign p_Result_23_fu_1630_p3 = ret_V_22_fu_1614_p2[34];
assign p_Result_24_fu_1690_p3 = ret_V_23_reg_2101[34];
assign p_Result_25_fu_1775_p3 = ret_V_25_fu_1759_p2[33];
assign p_Result_28_fu_497_p3 = p_Val2_2_fu_492_p2[3];
assign p_Result_29_fu_505_p3 = add_ln1192_1_fu_486_p2[4];
assign p_Result_31_fu_753_p1 = r_V_5_reg_1923[0];
assign p_Result_33_fu_788_p3 = p_Val2_6_fu_782_p2[1];
assign p_Result_34_fu_1004_p3 = ret_fu_998_p2[16];
assign p_Result_35_fu_1024_p3 = ret_fu_998_p2[13];
assign p_Result_38_fu_1404_p3 = ret_1_reg_2023[6];
assign p_Result_4_fu_1032_p4 = ret_fu_998_p2[16:14];
assign p_Result_7_fu_579_p4 = { add_ln1192_1_fu_486_p2[4], p_Val2_3_fu_573_p2 };
assign p_Result_s_22_fu_439_p4 = ret_V_17_fu_425_p2[6:4];
assign p_Result_s_fu_243_p3 = op_0[3];
assign p_Val2_10_fu_1016_p3 = { ret_fu_998_p2[13:0], 2'h0 };
assign p_Val2_14_fu_1397_p3 = { trunc_ln731_2_reg_2037, 2'h0 };
assign p_Val2_5_fu_756_p4 = r_V_5_reg_1923[2:1];
assign p_Val2_s_fu_255_p2 = { op_0[0], 3'h0 };
assign r_V_7_fu_1151_p0 = ret_V_18_reg_1996;
assign r_V_7_fu_1151_p00 = { 3'h0, ret_V_18_reg_1996 };
assign ret_V_10_cast_fu_1157_p4 = r_V_7_fu_1151_p2[4:1];
assign ret_V_17_cast_fu_1620_p4 = { ret_V_22_fu_1614_p2[34], ret_V_22_fu_1614_p2[34], ret_V_22_fu_1614_p2[34], ret_V_22_fu_1614_p2[34], ret_V_22_fu_1614_p2[34], ret_V_22_fu_1614_p2[34], ret_V_22_fu_1614_p2[34], ret_V_22_fu_1614_p2[34], ret_V_22_fu_1614_p2[34], ret_V_22_fu_1614_p2[34], ret_V_22_fu_1614_p2[34], ret_V_22_fu_1614_p2[34], ret_V_22_fu_1614_p2[34], ret_V_22_fu_1614_p2[34], ret_V_22_fu_1614_p2[34], ret_V_22_fu_1614_p2[34], ret_V_22_fu_1614_p2[34], ret_V_22_fu_1614_p2[34], ret_V_22_fu_1614_p2[34], ret_V_22_fu_1614_p2[34], ret_V_22_fu_1614_p2[13:2] };
assign ret_V_22_fu_1614_p2[33:14] = { ret_V_22_fu_1614_p2[34], ret_V_22_fu_1614_p2[34], ret_V_22_fu_1614_p2[34], ret_V_22_fu_1614_p2[34], ret_V_22_fu_1614_p2[34], ret_V_22_fu_1614_p2[34], ret_V_22_fu_1614_p2[34], ret_V_22_fu_1614_p2[34], ret_V_22_fu_1614_p2[34], ret_V_22_fu_1614_p2[34], ret_V_22_fu_1614_p2[34], ret_V_22_fu_1614_p2[34], ret_V_22_fu_1614_p2[34], ret_V_22_fu_1614_p2[34], ret_V_22_fu_1614_p2[34], ret_V_22_fu_1614_p2[34], ret_V_22_fu_1614_p2[34], ret_V_22_fu_1614_p2[34], ret_V_22_fu_1614_p2[34], ret_V_22_fu_1614_p2[34] };
assign ret_V_23_cast_fu_1765_p4 = ret_V_25_fu_1759_p2[32:1];
assign ret_V_6_fu_1295_p4 = ret_V_19_fu_1289_p2[12:3];
assign ret_V_fu_267_p4 = op_0[3:1];
assign rhs_2_fu_1278_p3 = { op_10_V_reg_2008, 3'h0 };
assign rhs_3_fu_1349_p3 = { select_ln850_4_fu_1341_p3, 13'h0000 };
assign rhs_5_fu_1662_p3 = { select_ln353_1_fu_1654_p3, 2'h0 };
assign rhs_7_fu_1748_p3 = { op_24_V_reg_2113, 1'h0 };
assign sext_ln1116_fu_677_p1 = { ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862 };
assign sext_ln1192_1_fu_476_p1 = { op_1_V_reg_1856[3], op_1_V_reg_1856 };
assign sext_ln1192_2_fu_1329_p0 = op_11;
assign sext_ln1192_2_fu_1329_p1 = { op_11[15], op_11[15], op_11[15], op_11[15], op_11[15], op_11[15], op_11[15], op_11[15], op_11 };
assign sext_ln1192_3_fu_1357_p1 = { select_ln850_4_fu_1341_p3[9], select_ln850_4_fu_1341_p3, 13'h0000 };
assign sext_ln1192_4_fu_1610_p1 = { select_ln353_fu_1595_p3[11], select_ln353_fu_1595_p3[11], select_ln353_fu_1595_p3[11], select_ln353_fu_1595_p3[11], select_ln353_fu_1595_p3[11], select_ln353_fu_1595_p3[11], select_ln353_fu_1595_p3[11], select_ln353_fu_1595_p3[11], select_ln353_fu_1595_p3[11], select_ln353_fu_1595_p3[11], select_ln353_fu_1595_p3[11], select_ln353_fu_1595_p3[11], select_ln353_fu_1595_p3[11], select_ln353_fu_1595_p3[11], select_ln353_fu_1595_p3[11], select_ln353_fu_1595_p3[11], select_ln353_fu_1595_p3[11], select_ln353_fu_1595_p3[11], select_ln353_fu_1595_p3[11], select_ln353_fu_1595_p3[11], select_ln353_fu_1595_p3[11], select_ln353_fu_1595_p3, 2'h0 };
assign sext_ln1192_5_fu_1670_p1 = { select_ln353_1_fu_1654_p3[31], select_ln353_1_fu_1654_p3, 2'h0 };
assign sext_ln1192_6_fu_1755_p1 = { op_24_V_reg_2113[31], op_24_V_reg_2113, 1'h0 };
assign sext_ln1192_fu_413_p1 = { op_0[3], op_0, 2'h0 };
assign sext_ln213_fu_975_p1 = { ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862 };
assign sext_ln69_1_fu_1813_p1 = { op_19_V_reg_2060[7], op_19_V_reg_2060 };
assign sext_ln69_2_fu_1831_p1 = { add_ln69_1_reg_2123[8], add_ln69_1_reg_2123[8], add_ln69_1_reg_2123[8], add_ln69_1_reg_2123[8], add_ln69_1_reg_2123[8], add_ln69_1_reg_2123[8], add_ln69_1_reg_2123[8], add_ln69_1_reg_2123[8], add_ln69_1_reg_2123 };
assign sext_ln69_3_fu_1840_p1 = { add_ln69_2_fu_1834_p2[16], add_ln69_2_fu_1834_p2[16], add_ln69_2_fu_1834_p2[16], add_ln69_2_fu_1834_p2[16], add_ln69_2_fu_1834_p2[16], add_ln69_2_fu_1834_p2[16], add_ln69_2_fu_1834_p2[16], add_ln69_2_fu_1834_p2[16], add_ln69_2_fu_1834_p2[16], add_ln69_2_fu_1834_p2[16], add_ln69_2_fu_1834_p2[16], add_ln69_2_fu_1834_p2[16], add_ln69_2_fu_1834_p2[16], add_ln69_2_fu_1834_p2[16], add_ln69_2_fu_1834_p2[16], add_ln69_2_fu_1834_p2 };
assign sext_ln69_fu_1822_p1 = { op_16[15], op_16 };
assign sext_ln703_1_fu_1274_p0 = op_6;
assign sext_ln703_1_fu_1274_p1 = { op_6[7], op_6[7], op_6[7], op_6[7], op_6[7], op_6 };
assign sext_ln703_2_fu_1587_p1 = { op_12_V_reg_2091[7], op_12_V_reg_2091[7], op_12_V_reg_2091[7], op_12_V_reg_2091[7], op_12_V_reg_2091[7], op_12_V_reg_2091[7], op_12_V_reg_2091[7], op_12_V_reg_2091[7], op_12_V_reg_2091[7], op_12_V_reg_2091[7], op_12_V_reg_2091[7], op_12_V_reg_2091[7], op_12_V_reg_2091[7], op_12_V_reg_2091[7], op_12_V_reg_2091[7], op_12_V_reg_2091[7], op_12_V_reg_2091[7], op_12_V_reg_2091[7], op_12_V_reg_2091[7], op_12_V_reg_2091[7], op_12_V_reg_2091[7], op_12_V_reg_2091[7], op_12_V_reg_2091[7], op_12_V_reg_2091[7], op_12_V_reg_2091[7], op_12_V_reg_2091[7], op_12_V_reg_2091[7], op_12_V_reg_2091 };
assign sext_ln703_3_fu_1644_p1 = { op_13_V_reg_2013[15], op_13_V_reg_2013[15], op_13_V_reg_2013[15], op_13_V_reg_2013[15], op_13_V_reg_2013[15], op_13_V_reg_2013[15], op_13_V_reg_2013[15], op_13_V_reg_2013[15], op_13_V_reg_2013[15], op_13_V_reg_2013[15], op_13_V_reg_2013[15], op_13_V_reg_2013[15], op_13_V_reg_2013[15], op_13_V_reg_2013[15], op_13_V_reg_2013[15], op_13_V_reg_2013[15], op_13_V_reg_2013[15], op_13_V_reg_2013[15], op_13_V_reg_2013[15], op_13_V_reg_2013 };
assign sext_ln703_4_fu_1744_p1 = { op_15_V_fu_1738_p3[1], op_15_V_fu_1738_p3[1], op_15_V_fu_1738_p3[1], op_15_V_fu_1738_p3[1], op_15_V_fu_1738_p3[1], op_15_V_fu_1738_p3[1], op_15_V_fu_1738_p3[1], op_15_V_fu_1738_p3[1], op_15_V_fu_1738_p3[1], op_15_V_fu_1738_p3[1], op_15_V_fu_1738_p3[1], op_15_V_fu_1738_p3[1], op_15_V_fu_1738_p3[1], op_15_V_fu_1738_p3[1], op_15_V_fu_1738_p3[1], op_15_V_fu_1738_p3[1], op_15_V_fu_1738_p3[1], op_15_V_fu_1738_p3[1], op_15_V_fu_1738_p3[1], op_15_V_fu_1738_p3[1], op_15_V_fu_1738_p3[1], op_15_V_fu_1738_p3[1], op_15_V_fu_1738_p3[1], op_15_V_fu_1738_p3[1], op_15_V_fu_1738_p3[1], op_15_V_fu_1738_p3[1], op_15_V_fu_1738_p3[1], op_15_V_fu_1738_p3[1], op_15_V_fu_1738_p3[1], op_15_V_fu_1738_p3[1], op_15_V_fu_1738_p3[1], op_15_V_fu_1738_p3[1], op_15_V_fu_1738_p3 };
assign sext_ln703_fu_417_p1 = { op_1_V_fu_375_p3[3], op_1_V_fu_375_p3[3], op_1_V_fu_375_p3[3], op_1_V_fu_375_p3 };
assign sext_ln727_fu_954_p1 = { op_3_V_reg_1896[3], op_3_V_reg_1896[3], op_3_V_reg_1896[3], op_3_V_reg_1896[3], op_3_V_reg_1896 };
assign sext_ln850_fu_1377_p1 = { ret_V_21_fu_1361_p2[23], ret_V_21_fu_1361_p2[23:13] };
assign shl_ln1192_fu_471_p2 = { op_0[1:0], 2'h0 };
assign shl_ln_fu_957_p3 = { ret_V_18_fu_947_p3, 3'h0 };
assign tmp_13_fu_830_p3 = r_V_5_reg_1923[3];
assign tmp_1_fu_1233_p4 = ret_1_fu_1207_p2[32:6];
assign tmp_23_fu_1441_p3 = ret_1_reg_2023[6];
assign tmp_24_fu_1448_p3 = ret_1_reg_2023[5];
assign tmp_26_fu_1602_p3 = { select_ln353_fu_1595_p3, 2'h0 };
assign tmp_6_fu_545_p3 = add_ln1192_1_fu_486_p2[4];
assign tmp_7_fu_553_p3 = p_Val2_2_fu_492_p2[3];
assign tmp_fu_1367_p4 = ret_V_21_fu_1361_p2[23:13];
assign trunc_ln1192_1_fu_479_p3 = { trunc_ln1192_reg_1868, 2'h0 };
assign trunc_ln1192_fu_421_p1 = op_0[2:0];
assign trunc_ln213_fu_978_p1 = op_7[7:0];
assign trunc_ln731_1_fu_1012_p1 = ret_fu_998_p2[13:0];
assign trunc_ln731_2_fu_1221_p1 = ret_1_fu_1207_p2[5:0];
assign trunc_ln731_fu_251_p1 = op_0[0];
assign trunc_ln851_1_fu_1313_p0 = op_6;
assign trunc_ln851_1_fu_1313_p1 = op_6[2:0];
assign trunc_ln851_2_fu_1175_p1 = r_V_7_fu_1151_p2[0];
assign trunc_ln851_3_fu_1381_p0 = op_11;
assign trunc_ln851_3_fu_1381_p1 = op_11[12:0];
assign trunc_ln851_4_fu_1570_p1 = op_12_V_fu_1562_p3[1:0];
assign trunc_ln851_5_fu_1264_p1 = op_13_V_fu_1140_p3[1:0];
assign trunc_ln851_6_fu_1783_p1 = op_15_V_fu_1738_p3[0];
assign trunc_ln851_fu_749_p1 = grp_fu_697_p2[2:0];
assign zext_ln1116_fu_680_p1 = { 4'h0, ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862 };
assign zext_ln1192_fu_1285_p1 = { 2'h0, op_10_V_reg_2008, 3'h0 };
assign zext_ln1347_1_fu_1204_p1 = { 32'h00000000, rhs_4_reg_2002 };
assign zext_ln1347_fu_1201_p1 = { 1'h0, sext_ln1116_reg_1902 };
assign zext_ln1499_fu_965_p1 = { 1'h0, ret_V_18_fu_947_p3, 3'h0 };
assign zext_ln215_1_fu_994_p1 = { 1'h0, op_7 };
assign zext_ln215_fu_991_p1 = { 13'h0000, ret_V_18_reg_1996 };
assign zext_ln415_fu_778_p1 = { 1'h0, and_ln412_fu_772_p2 };
assign zext_ln69_1_fu_1715_p1 = { 28'h0000000, ret_V_20_reg_2018 };
assign zext_ln69_2_fu_1809_p1 = { 5'h00, op_18 };
assign zext_ln69_fu_1255_p1 = { 7'h00, rhs_4_reg_2002 };
assign \mul_4ns_3s_7_1_1_U3.top_mul_4ns_3s_7_1_1_Multiplier_1_U.a  = \mul_4ns_3s_7_1_1_U3.din0 ;
assign \mul_4ns_3s_7_1_1_U3.top_mul_4ns_3s_7_1_1_Multiplier_1_U.b  = \mul_4ns_3s_7_1_1_U3.din1 ;
assign \mul_4ns_3s_7_1_1_U3.dout  = \mul_4ns_3s_7_1_1_U3.top_mul_4ns_3s_7_1_1_Multiplier_1_U.p ;
assign \mul_4ns_3s_7_1_1_U3.din0  = ret_V_18_reg_1996;
assign \mul_4ns_3s_7_1_1_U3.din1  = r_V_reg_1891;
assign r_V_7_fu_1151_p2 = \mul_4ns_3s_7_1_1_U3.dout ;
assign \mul_32ns_4s_36_2_1_U2.top_mul_32ns_4s_36_2_1_Multiplier_0_U.a  = \mul_32ns_4s_36_2_1_U2.din0 ;
assign \mul_32ns_4s_36_2_1_U2.top_mul_32ns_4s_36_2_1_Multiplier_0_U.b  = \mul_32ns_4s_36_2_1_U2.din1 ;
assign \mul_32ns_4s_36_2_1_U2.top_mul_32ns_4s_36_2_1_Multiplier_0_U.ce  = \mul_32ns_4s_36_2_1_U2.ce ;
assign \mul_32ns_4s_36_2_1_U2.top_mul_32ns_4s_36_2_1_Multiplier_0_U.clk  = \mul_32ns_4s_36_2_1_U2.clk ;
assign \mul_32ns_4s_36_2_1_U2.dout  = \mul_32ns_4s_36_2_1_U2.top_mul_32ns_4s_36_2_1_Multiplier_0_U.p ;
assign \mul_32ns_4s_36_2_1_U2.ce  = 1'h1;
assign \mul_32ns_4s_36_2_1_U2.clk  = ap_clk;
assign \mul_32ns_4s_36_2_1_U2.din0  = { ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862 };
assign \mul_32ns_4s_36_2_1_U2.din1  = op_3_V_reg_1896;
assign grp_fu_697_p2 = \mul_32ns_4s_36_2_1_U2.dout ;
assign \mul_32ns_4s_36_2_1_U2.reset  = ap_rst;
assign \mul_32ns_4s_36_2_1_U1.top_mul_32ns_4s_36_2_1_Multiplier_0_U.a  = \mul_32ns_4s_36_2_1_U1.din0 ;
assign \mul_32ns_4s_36_2_1_U1.top_mul_32ns_4s_36_2_1_Multiplier_0_U.b  = \mul_32ns_4s_36_2_1_U1.din1 ;
assign \mul_32ns_4s_36_2_1_U1.top_mul_32ns_4s_36_2_1_Multiplier_0_U.ce  = \mul_32ns_4s_36_2_1_U1.ce ;
assign \mul_32ns_4s_36_2_1_U1.top_mul_32ns_4s_36_2_1_Multiplier_0_U.clk  = \mul_32ns_4s_36_2_1_U1.clk ;
assign \mul_32ns_4s_36_2_1_U1.dout  = \mul_32ns_4s_36_2_1_U1.top_mul_32ns_4s_36_2_1_Multiplier_0_U.p ;
assign \mul_32ns_4s_36_2_1_U1.ce  = 1'h1;
assign \mul_32ns_4s_36_2_1_U1.clk  = ap_clk;
assign \mul_32ns_4s_36_2_1_U1.din0  = { ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862[2], ret_V_16_reg_1862 };
assign \mul_32ns_4s_36_2_1_U1.din1  = op_8;
assign grp_fu_688_p2 = \mul_32ns_4s_36_2_1_U1.dout ;
assign \mul_32ns_4s_36_2_1_U1.reset  = ap_rst;
endmodule


// Product machine:
module top_A_times_top_B (ap_start, op_0, op_11, op_16, op_17, op_18, op_6, op_7, op_8, ap_clk, unsafe_signal);
input ap_start;
input [3:0] op_0;
input [15:0] op_11;
input [15:0] op_16;
input [31:0] op_17;
input [3:0] op_18;
input [7:0] op_6;
input [15:0] op_7;
input [3:0] op_8;
input ap_clk;
output unsafe_signal;
reg _setup;
initial _setup = 1'b0;
always @ (posedge ap_clk) _setup <= 1'b1;
reg ap_start_internal;
always @ (posedge ap_clk) if (!_setup) ap_start_internal <= ap_start;
reg [3:0] op_0_internal;
always @ (posedge ap_clk) if (!_setup) op_0_internal <= op_0;
reg [15:0] op_11_internal;
always @ (posedge ap_clk) if (!_setup) op_11_internal <= op_11;
reg [15:0] op_16_internal;
always @ (posedge ap_clk) if (!_setup) op_16_internal <= op_16;
reg [31:0] op_17_internal;
always @ (posedge ap_clk) if (!_setup) op_17_internal <= op_17;
reg [3:0] op_18_internal;
always @ (posedge ap_clk) if (!_setup) op_18_internal <= op_18;
reg [7:0] op_6_internal;
always @ (posedge ap_clk) if (!_setup) op_6_internal <= op_6;
reg [15:0] op_7_internal;
always @ (posedge ap_clk) if (!_setup) op_7_internal <= op_7;
reg [3:0] op_8_internal;
always @ (posedge ap_clk) if (!_setup) op_8_internal <= op_8;
wire ap_done_A;
wire ap_done_B;
wire ap_done_eq;
assign ap_done_eq = ap_done_A == ap_done_B;
wire ap_idle_A;
wire ap_idle_B;
wire ap_idle_eq;
assign ap_idle_eq = ap_idle_A == ap_idle_B;
wire ap_ready_A;
wire ap_ready_B;
wire ap_ready_eq;
assign ap_ready_eq = ap_ready_A == ap_ready_B;
wire [31:0] op_29_A;
wire [31:0] op_29_B;
wire op_29_eq;
assign op_29_eq = op_29_A == op_29_B;
wire op_29_ap_vld_A;
wire op_29_ap_vld_B;
wire clk_enable_A;
wire clk_enable_B;
assign clk_enable_A = _setup & (~op_29_ap_vld_A | op_29_ap_vld_B);
assign clk_enable_B = _setup;
wire divergent;
assign divergent = ~(ap_done_eq & ap_idle_eq & ap_ready_eq & op_29_eq);
assign unsafe_signal = op_29_ap_vld_A & op_29_ap_vld_B & divergent;
top_A instance_A (
    .ap_clk(ap_clk),
    .clk_enable(clk_enable_A),
    .ap_start(ap_start_internal),
    .op_0(op_0_internal),
    .op_11(op_11_internal),
    .op_16(op_16_internal),
    .op_17(op_17_internal),
    .op_18(op_18_internal),
    .op_6(op_6_internal),
    .op_7(op_7_internal),
    .op_8(op_8_internal),
    .ap_done(ap_done_A),
    .ap_idle(ap_idle_A),
    .ap_ready(ap_ready_A),
    .op_29(op_29_A),
    .op_29_ap_vld(op_29_ap_vld_A)
);
top_B instance_B (
    .ap_clk(ap_clk),
    .clk_enable(clk_enable_B),
    .ap_start(ap_start_internal),
    .op_0(op_0_internal),
    .op_11(op_11_internal),
    .op_16(op_16_internal),
    .op_17(op_17_internal),
    .op_18(op_18_internal),
    .op_6(op_6_internal),
    .op_7(op_7_internal),
    .op_8(op_8_internal),
    .ap_done(ap_done_B),
    .ap_idle(ap_idle_B),
    .ap_ready(ap_ready_B),
    .op_29(op_29_B),
    .op_29_ap_vld(op_29_ap_vld_B)
);
endmodule
