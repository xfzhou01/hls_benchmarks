// Processed by function `construct_kairos` in `verilog_tricks.py`.
// Machine A:
// Processed by function `add_clk_enable_signal` in `verilog_tricks.py`.
// Processed by function `remove_reset_signal` in `verilog_tricks.py`.
module top_A (
  ap_clk,
  ap_start,
  ap_done,
  ap_idle,
  ap_ready,
  op_0,
  op_2,
  op_3,
  op_5,
  op_10,
  op_11,
  op_12,
  op_13,
  op_16,
  op_17,
  op_19,
  op_30,
  op_30_ap_vld,
clk_enable
);
input clk_enable;


input ap_clk;
wire ap_rst;
assign ap_rst = op_30_ap_vld;
input ap_start;
input [31:0] op_0;
input [1:0] op_10;
input [31:0] op_11;
input [31:0] op_12;
input op_13;
input [7:0] op_16;
input [31:0] op_17;
input [31:0] op_19;
input [3:0] op_2;
input [1:0] op_3;
input op_5;
output ap_done;
output ap_idle;
output ap_ready;
output [31:0] op_30;
output op_30_ap_vld;


reg [14:0] \add_29ns_29ns_29_2_1_U5.top_add_29ns_29ns_29_2_1_Adder_2_U.ain_s1 ;
reg [14:0] \add_29ns_29ns_29_2_1_U5.top_add_29ns_29ns_29_2_1_Adder_2_U.bin_s1 ;
reg \add_29ns_29ns_29_2_1_U5.top_add_29ns_29ns_29_2_1_Adder_2_U.carry_s1 ;
reg [13:0] \add_29ns_29ns_29_2_1_U5.top_add_29ns_29ns_29_2_1_Adder_2_U.sum_s1 ;
reg [14:0] \add_29ns_29ns_29_2_1_U6.top_add_29ns_29ns_29_2_1_Adder_2_U.ain_s1 ;
reg [14:0] \add_29ns_29ns_29_2_1_U6.top_add_29ns_29ns_29_2_1_Adder_2_U.bin_s1 ;
reg \add_29ns_29ns_29_2_1_U6.top_add_29ns_29ns_29_2_1_Adder_2_U.carry_s1 ;
reg [13:0] \add_29ns_29ns_29_2_1_U6.top_add_29ns_29ns_29_2_1_Adder_2_U.sum_s1 ;
reg [14:0] \add_29ns_29ns_29_2_1_U7.top_add_29ns_29ns_29_2_1_Adder_2_U.ain_s1 ;
reg [14:0] \add_29ns_29ns_29_2_1_U7.top_add_29ns_29ns_29_2_1_Adder_2_U.bin_s1 ;
reg \add_29ns_29ns_29_2_1_U7.top_add_29ns_29ns_29_2_1_Adder_2_U.carry_s1 ;
reg [13:0] \add_29ns_29ns_29_2_1_U7.top_add_29ns_29ns_29_2_1_Adder_2_U.sum_s1 ;
reg [14:0] \add_29ns_29s_29_2_1_U8.top_add_29ns_29s_29_2_1_Adder_3_U.ain_s1 ;
reg [14:0] \add_29ns_29s_29_2_1_U8.top_add_29ns_29s_29_2_1_Adder_3_U.bin_s1 ;
reg \add_29ns_29s_29_2_1_U8.top_add_29ns_29s_29_2_1_Adder_3_U.carry_s1 ;
reg [13:0] \add_29ns_29s_29_2_1_U8.top_add_29ns_29s_29_2_1_Adder_3_U.sum_s1 ;
reg [14:0] \add_29s_29ns_29_2_1_U4.top_add_29s_29ns_29_2_1_Adder_1_U.ain_s1 ;
reg [14:0] \add_29s_29ns_29_2_1_U4.top_add_29s_29ns_29_2_1_Adder_1_U.bin_s1 ;
reg \add_29s_29ns_29_2_1_U4.top_add_29s_29ns_29_2_1_Adder_1_U.carry_s1 ;
reg [13:0] \add_29s_29ns_29_2_1_U4.top_add_29s_29ns_29_2_1_Adder_1_U.sum_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_5_U.ain_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_5_U.bin_s1 ;
reg \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_5_U.carry_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_5_U.sum_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.ain_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.bin_s1 ;
reg \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.carry_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.sum_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_5_U.ain_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_5_U.bin_s1 ;
reg \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_5_U.carry_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_5_U.sum_s1 ;
reg [16:0] \add_33s_33s_33_2_1_U3.top_add_33s_33s_33_2_1_Adder_0_U.ain_s1 ;
reg [16:0] \add_33s_33s_33_2_1_U3.top_add_33s_33s_33_2_1_Adder_0_U.bin_s1 ;
reg \add_33s_33s_33_2_1_U3.top_add_33s_33s_33_2_1_Adder_0_U.carry_s1 ;
reg [15:0] \add_33s_33s_33_2_1_U3.top_add_33s_33s_33_2_1_Adder_0_U.sum_s1 ;
reg [17:0] \add_35s_35s_35_2_1_U11.top_add_35s_35s_35_2_1_Adder_6_U.ain_s1 ;
reg [17:0] \add_35s_35s_35_2_1_U11.top_add_35s_35s_35_2_1_Adder_6_U.bin_s1 ;
reg \add_35s_35s_35_2_1_U11.top_add_35s_35s_35_2_1_Adder_6_U.carry_s1 ;
reg [16:0] \add_35s_35s_35_2_1_U11.top_add_35s_35s_35_2_1_Adder_6_U.sum_s1 ;
reg [21:0] \add_43s_43s_43_2_1_U9.top_add_43s_43s_43_2_1_Adder_4_U.ain_s1 ;
reg [21:0] \add_43s_43s_43_2_1_U9.top_add_43s_43s_43_2_1_Adder_4_U.bin_s1 ;
reg \add_43s_43s_43_2_1_U9.top_add_43s_43s_43_2_1_Adder_4_U.carry_s1 ;
reg [20:0] \add_43s_43s_43_2_1_U9.top_add_43s_43s_43_2_1_Adder_4_U.sum_s1 ;
reg [31:0] add_ln691_1_reg_861;
reg [31:0] add_ln691_2_reg_908;
reg [28:0] add_ln691_reg_737;
reg [2:0] add_ln69_reg_680;
reg [29:0] ap_CS_fsm = 30'h00000001;
reg icmp_ln851_1_reg_812;
reg icmp_ln851_2_reg_891;
reg icmp_ln851_reg_715;
reg lhs_V_reg_772;
reg [3:0] \mul_4ns_4ns_8_4_1_U1.top_mul_4ns_4ns_8_4_1_Mul_DSP_0_U.a_reg0 ;
reg [3:0] \mul_4ns_4ns_8_4_1_U1.top_mul_4ns_4ns_8_4_1_Mul_DSP_0_U.b_reg0 ;
reg [7:0] \mul_4ns_4ns_8_4_1_U1.top_mul_4ns_4ns_8_4_1_Mul_DSP_0_U.buff0 ;
reg [7:0] \mul_4ns_4ns_8_4_1_U1.top_mul_4ns_4ns_8_4_1_Mul_DSP_0_U.buff1 ;
reg [3:0] op_18_V_reg_866;
reg [8:0] op_22_V_reg_700;
reg [28:0] op_25_V_reg_777;
reg [28:0] op_27_V_reg_797;
reg [1:0] op_6_V_reg_670;
reg or_ln785_reg_855;
reg p_Result_4_reg_829;
reg p_Result_5_reg_841;
reg [32:0] ret_V_1_reg_720;
reg [28:0] ret_V_2_reg_742;
reg [28:0] ret_V_3_reg_757;
reg [28:0] ret_V_4_reg_787;
reg [31:0] ret_V_5_cast_reg_822;
reg [42:0] ret_V_5_reg_817;
reg [34:0] ret_V_6_reg_896;
reg [31:0] ret_V_7_reg_913;
reg [31:0] ret_V_8_cast_reg_901;
reg [7:0] ret_reg_685;
reg [28:0] select_ln1192_reg_747;
reg [31:0] select_ln353_reg_871;
reg [15:0] select_ln546_reg_690;
reg [28:0] select_ln69_1_reg_762;
reg [2:0] select_ln69_reg_675;
reg [28:0] sext_ln850_reg_730;
reg [3:0] \shl_16ns_4ns_16_7_1_U2.din1_cast_array[0] ;
reg [3:0] \shl_16ns_4ns_16_7_1_U2.din1_cast_array[1] ;
reg [3:0] \shl_16ns_4ns_16_7_1_U2.din1_cast_array[2] ;
reg [3:0] \shl_16ns_4ns_16_7_1_U2.din1_cast_array[3] ;
reg [3:0] \shl_16ns_4ns_16_7_1_U2.din1_cast_array[4] ;
reg [3:0] \shl_16ns_4ns_16_7_1_U2.din1_cast_array[5] ;
reg [15:0] \shl_16ns_4ns_16_7_1_U2.dout_array[0] ;
reg [15:0] \shl_16ns_4ns_16_7_1_U2.dout_array[1] ;
reg [15:0] \shl_16ns_4ns_16_7_1_U2.dout_array[2] ;
reg [15:0] \shl_16ns_4ns_16_7_1_U2.dout_array[3] ;
reg [15:0] \shl_16ns_4ns_16_7_1_U2.dout_array[4] ;
reg [15:0] \shl_16ns_4ns_16_7_1_U2.dout_array[5] ;
reg [15:0] shl_ln781_reg_752;
reg tmp_5_reg_848;
reg [27:0] tmp_reg_725;
reg [1:0] trunc_ln731_reg_836;
reg [1:0] trunc_ln851_2_reg_876;
wire [31:0] _000_;
wire [31:0] _001_;
wire [28:0] _002_;
wire [2:0] _003_;
wire [29:0] _004_;
wire _005_;
wire _006_;
wire _007_;
wire _008_;
wire [1:0] _009_;
wire [8:0] _010_;
wire [28:0] _011_;
wire [28:0] _012_;
wire [1:0] _013_;
wire _014_;
wire _015_;
wire _016_;
wire [32:0] _017_;
wire [28:0] _018_;
wire [28:0] _019_;
wire [28:0] _020_;
wire [31:0] _021_;
wire [42:0] _022_;
wire [34:0] _023_;
wire [31:0] _024_;
wire [31:0] _025_;
wire [7:0] _026_;
wire [28:0] _027_;
wire [31:0] _028_;
wire [15:0] _029_;
wire [28:0] _030_;
wire [2:0] _031_;
wire [28:0] _032_;
wire [15:0] _033_;
wire _034_;
wire [27:0] _035_;
wire [1:0] _036_;
wire [1:0] _037_;
wire _038_;
wire _039_;
wire _040_;
wire _041_;
wire _042_;
wire _043_;
wire [14:0] _044_;
wire [14:0] _045_;
wire _046_;
wire [13:0] _047_;
wire [14:0] _048_;
wire [15:0] _049_;
wire [14:0] _050_;
wire [14:0] _051_;
wire _052_;
wire [13:0] _053_;
wire [14:0] _054_;
wire [15:0] _055_;
wire [14:0] _056_;
wire [14:0] _057_;
wire _058_;
wire [13:0] _059_;
wire [14:0] _060_;
wire [15:0] _061_;
wire [14:0] _062_;
wire [14:0] _063_;
wire _064_;
wire [13:0] _065_;
wire [14:0] _066_;
wire [15:0] _067_;
wire [14:0] _068_;
wire [14:0] _069_;
wire _070_;
wire [13:0] _071_;
wire [14:0] _072_;
wire [15:0] _073_;
wire [15:0] _074_;
wire [15:0] _075_;
wire _076_;
wire [15:0] _077_;
wire [16:0] _078_;
wire [16:0] _079_;
wire [15:0] _080_;
wire [15:0] _081_;
wire _082_;
wire [15:0] _083_;
wire [16:0] _084_;
wire [16:0] _085_;
wire [15:0] _086_;
wire [15:0] _087_;
wire _088_;
wire [15:0] _089_;
wire [16:0] _090_;
wire [16:0] _091_;
wire [16:0] _092_;
wire [16:0] _093_;
wire _094_;
wire [15:0] _095_;
wire [16:0] _096_;
wire [17:0] _097_;
wire [17:0] _098_;
wire [17:0] _099_;
wire _100_;
wire [16:0] _101_;
wire [17:0] _102_;
wire [18:0] _103_;
wire [21:0] _104_;
wire [21:0] _105_;
wire _106_;
wire [20:0] _107_;
wire [21:0] _108_;
wire [22:0] _109_;
wire [3:0] _110_;
wire [3:0] _111_;
wire [7:0] _112_;
wire [7:0] _113_;
wire [3:0] _114_;
wire [3:0] _115_;
wire [3:0] _116_;
wire [3:0] _117_;
wire [3:0] _118_;
wire [3:0] _119_;
wire [15:0] _120_;
wire [15:0] _121_;
wire [15:0] _122_;
wire [15:0] _123_;
wire [15:0] _124_;
wire [15:0] _125_;
wire [3:0] _126_;
wire [15:0] _127_;
wire [3:0] _128_;
wire [15:0] _129_;
wire [3:0] _130_;
wire [15:0] _131_;
wire [3:0] _132_;
wire [15:0] _133_;
wire [3:0] _134_;
wire [15:0] _135_;
wire [3:0] _136_;
wire [15:0] _137_;
wire [15:0] _138_;
wire [15:0] _139_;
wire [15:0] _140_;
wire _141_;
wire _142_;
wire _143_;
wire _144_;
wire _145_;
wire _146_;
wire _147_;
wire _148_;
wire _149_;
wire _150_;
wire _151_;
wire _152_;
wire _153_;
wire _154_;
wire _155_;
wire _156_;
wire _157_;
wire _158_;
wire _159_;
wire _160_;
wire _161_;
wire _162_;
wire _163_;
wire _164_;
wire _165_;
wire _166_;
wire _167_;
wire _168_;
wire _169_;
wire _170_;
wire _171_;
wire _172_;
wire _173_;
wire _174_;
wire \add_29ns_29ns_29_2_1_U5.ce ;
wire \add_29ns_29ns_29_2_1_U5.clk ;
wire [28:0] \add_29ns_29ns_29_2_1_U5.din0 ;
wire [28:0] \add_29ns_29ns_29_2_1_U5.din1 ;
wire [28:0] \add_29ns_29ns_29_2_1_U5.dout ;
wire \add_29ns_29ns_29_2_1_U5.reset ;
wire [28:0] \add_29ns_29ns_29_2_1_U5.top_add_29ns_29ns_29_2_1_Adder_2_U.a ;
wire [28:0] \add_29ns_29ns_29_2_1_U5.top_add_29ns_29ns_29_2_1_Adder_2_U.ain_s0 ;
wire [28:0] \add_29ns_29ns_29_2_1_U5.top_add_29ns_29ns_29_2_1_Adder_2_U.b ;
wire [28:0] \add_29ns_29ns_29_2_1_U5.top_add_29ns_29ns_29_2_1_Adder_2_U.bin_s0 ;
wire \add_29ns_29ns_29_2_1_U5.top_add_29ns_29ns_29_2_1_Adder_2_U.ce ;
wire \add_29ns_29ns_29_2_1_U5.top_add_29ns_29ns_29_2_1_Adder_2_U.clk ;
wire \add_29ns_29ns_29_2_1_U5.top_add_29ns_29ns_29_2_1_Adder_2_U.facout_s1 ;
wire \add_29ns_29ns_29_2_1_U5.top_add_29ns_29ns_29_2_1_Adder_2_U.facout_s2 ;
wire [13:0] \add_29ns_29ns_29_2_1_U5.top_add_29ns_29ns_29_2_1_Adder_2_U.fas_s1 ;
wire [14:0] \add_29ns_29ns_29_2_1_U5.top_add_29ns_29ns_29_2_1_Adder_2_U.fas_s2 ;
wire \add_29ns_29ns_29_2_1_U5.top_add_29ns_29ns_29_2_1_Adder_2_U.reset ;
wire [28:0] \add_29ns_29ns_29_2_1_U5.top_add_29ns_29ns_29_2_1_Adder_2_U.s ;
wire [13:0] \add_29ns_29ns_29_2_1_U5.top_add_29ns_29ns_29_2_1_Adder_2_U.u1.a ;
wire [13:0] \add_29ns_29ns_29_2_1_U5.top_add_29ns_29ns_29_2_1_Adder_2_U.u1.b ;
wire \add_29ns_29ns_29_2_1_U5.top_add_29ns_29ns_29_2_1_Adder_2_U.u1.cin ;
wire \add_29ns_29ns_29_2_1_U5.top_add_29ns_29ns_29_2_1_Adder_2_U.u1.cout ;
wire [13:0] \add_29ns_29ns_29_2_1_U5.top_add_29ns_29ns_29_2_1_Adder_2_U.u1.s ;
wire [14:0] \add_29ns_29ns_29_2_1_U5.top_add_29ns_29ns_29_2_1_Adder_2_U.u2.a ;
wire [14:0] \add_29ns_29ns_29_2_1_U5.top_add_29ns_29ns_29_2_1_Adder_2_U.u2.b ;
wire \add_29ns_29ns_29_2_1_U5.top_add_29ns_29ns_29_2_1_Adder_2_U.u2.cin ;
wire \add_29ns_29ns_29_2_1_U5.top_add_29ns_29ns_29_2_1_Adder_2_U.u2.cout ;
wire [14:0] \add_29ns_29ns_29_2_1_U5.top_add_29ns_29ns_29_2_1_Adder_2_U.u2.s ;
wire \add_29ns_29ns_29_2_1_U6.ce ;
wire \add_29ns_29ns_29_2_1_U6.clk ;
wire [28:0] \add_29ns_29ns_29_2_1_U6.din0 ;
wire [28:0] \add_29ns_29ns_29_2_1_U6.din1 ;
wire [28:0] \add_29ns_29ns_29_2_1_U6.dout ;
wire \add_29ns_29ns_29_2_1_U6.reset ;
wire [28:0] \add_29ns_29ns_29_2_1_U6.top_add_29ns_29ns_29_2_1_Adder_2_U.a ;
wire [28:0] \add_29ns_29ns_29_2_1_U6.top_add_29ns_29ns_29_2_1_Adder_2_U.ain_s0 ;
wire [28:0] \add_29ns_29ns_29_2_1_U6.top_add_29ns_29ns_29_2_1_Adder_2_U.b ;
wire [28:0] \add_29ns_29ns_29_2_1_U6.top_add_29ns_29ns_29_2_1_Adder_2_U.bin_s0 ;
wire \add_29ns_29ns_29_2_1_U6.top_add_29ns_29ns_29_2_1_Adder_2_U.ce ;
wire \add_29ns_29ns_29_2_1_U6.top_add_29ns_29ns_29_2_1_Adder_2_U.clk ;
wire \add_29ns_29ns_29_2_1_U6.top_add_29ns_29ns_29_2_1_Adder_2_U.facout_s1 ;
wire \add_29ns_29ns_29_2_1_U6.top_add_29ns_29ns_29_2_1_Adder_2_U.facout_s2 ;
wire [13:0] \add_29ns_29ns_29_2_1_U6.top_add_29ns_29ns_29_2_1_Adder_2_U.fas_s1 ;
wire [14:0] \add_29ns_29ns_29_2_1_U6.top_add_29ns_29ns_29_2_1_Adder_2_U.fas_s2 ;
wire \add_29ns_29ns_29_2_1_U6.top_add_29ns_29ns_29_2_1_Adder_2_U.reset ;
wire [28:0] \add_29ns_29ns_29_2_1_U6.top_add_29ns_29ns_29_2_1_Adder_2_U.s ;
wire [13:0] \add_29ns_29ns_29_2_1_U6.top_add_29ns_29ns_29_2_1_Adder_2_U.u1.a ;
wire [13:0] \add_29ns_29ns_29_2_1_U6.top_add_29ns_29ns_29_2_1_Adder_2_U.u1.b ;
wire \add_29ns_29ns_29_2_1_U6.top_add_29ns_29ns_29_2_1_Adder_2_U.u1.cin ;
wire \add_29ns_29ns_29_2_1_U6.top_add_29ns_29ns_29_2_1_Adder_2_U.u1.cout ;
wire [13:0] \add_29ns_29ns_29_2_1_U6.top_add_29ns_29ns_29_2_1_Adder_2_U.u1.s ;
wire [14:0] \add_29ns_29ns_29_2_1_U6.top_add_29ns_29ns_29_2_1_Adder_2_U.u2.a ;
wire [14:0] \add_29ns_29ns_29_2_1_U6.top_add_29ns_29ns_29_2_1_Adder_2_U.u2.b ;
wire \add_29ns_29ns_29_2_1_U6.top_add_29ns_29ns_29_2_1_Adder_2_U.u2.cin ;
wire \add_29ns_29ns_29_2_1_U6.top_add_29ns_29ns_29_2_1_Adder_2_U.u2.cout ;
wire [14:0] \add_29ns_29ns_29_2_1_U6.top_add_29ns_29ns_29_2_1_Adder_2_U.u2.s ;
wire \add_29ns_29ns_29_2_1_U7.ce ;
wire \add_29ns_29ns_29_2_1_U7.clk ;
wire [28:0] \add_29ns_29ns_29_2_1_U7.din0 ;
wire [28:0] \add_29ns_29ns_29_2_1_U7.din1 ;
wire [28:0] \add_29ns_29ns_29_2_1_U7.dout ;
wire \add_29ns_29ns_29_2_1_U7.reset ;
wire [28:0] \add_29ns_29ns_29_2_1_U7.top_add_29ns_29ns_29_2_1_Adder_2_U.a ;
wire [28:0] \add_29ns_29ns_29_2_1_U7.top_add_29ns_29ns_29_2_1_Adder_2_U.ain_s0 ;
wire [28:0] \add_29ns_29ns_29_2_1_U7.top_add_29ns_29ns_29_2_1_Adder_2_U.b ;
wire [28:0] \add_29ns_29ns_29_2_1_U7.top_add_29ns_29ns_29_2_1_Adder_2_U.bin_s0 ;
wire \add_29ns_29ns_29_2_1_U7.top_add_29ns_29ns_29_2_1_Adder_2_U.ce ;
wire \add_29ns_29ns_29_2_1_U7.top_add_29ns_29ns_29_2_1_Adder_2_U.clk ;
wire \add_29ns_29ns_29_2_1_U7.top_add_29ns_29ns_29_2_1_Adder_2_U.facout_s1 ;
wire \add_29ns_29ns_29_2_1_U7.top_add_29ns_29ns_29_2_1_Adder_2_U.facout_s2 ;
wire [13:0] \add_29ns_29ns_29_2_1_U7.top_add_29ns_29ns_29_2_1_Adder_2_U.fas_s1 ;
wire [14:0] \add_29ns_29ns_29_2_1_U7.top_add_29ns_29ns_29_2_1_Adder_2_U.fas_s2 ;
wire \add_29ns_29ns_29_2_1_U7.top_add_29ns_29ns_29_2_1_Adder_2_U.reset ;
wire [28:0] \add_29ns_29ns_29_2_1_U7.top_add_29ns_29ns_29_2_1_Adder_2_U.s ;
wire [13:0] \add_29ns_29ns_29_2_1_U7.top_add_29ns_29ns_29_2_1_Adder_2_U.u1.a ;
wire [13:0] \add_29ns_29ns_29_2_1_U7.top_add_29ns_29ns_29_2_1_Adder_2_U.u1.b ;
wire \add_29ns_29ns_29_2_1_U7.top_add_29ns_29ns_29_2_1_Adder_2_U.u1.cin ;
wire \add_29ns_29ns_29_2_1_U7.top_add_29ns_29ns_29_2_1_Adder_2_U.u1.cout ;
wire [13:0] \add_29ns_29ns_29_2_1_U7.top_add_29ns_29ns_29_2_1_Adder_2_U.u1.s ;
wire [14:0] \add_29ns_29ns_29_2_1_U7.top_add_29ns_29ns_29_2_1_Adder_2_U.u2.a ;
wire [14:0] \add_29ns_29ns_29_2_1_U7.top_add_29ns_29ns_29_2_1_Adder_2_U.u2.b ;
wire \add_29ns_29ns_29_2_1_U7.top_add_29ns_29ns_29_2_1_Adder_2_U.u2.cin ;
wire \add_29ns_29ns_29_2_1_U7.top_add_29ns_29ns_29_2_1_Adder_2_U.u2.cout ;
wire [14:0] \add_29ns_29ns_29_2_1_U7.top_add_29ns_29ns_29_2_1_Adder_2_U.u2.s ;
wire \add_29ns_29s_29_2_1_U8.ce ;
wire \add_29ns_29s_29_2_1_U8.clk ;
wire [28:0] \add_29ns_29s_29_2_1_U8.din0 ;
wire [28:0] \add_29ns_29s_29_2_1_U8.din1 ;
wire [28:0] \add_29ns_29s_29_2_1_U8.dout ;
wire \add_29ns_29s_29_2_1_U8.reset ;
wire [28:0] \add_29ns_29s_29_2_1_U8.top_add_29ns_29s_29_2_1_Adder_3_U.a ;
wire [28:0] \add_29ns_29s_29_2_1_U8.top_add_29ns_29s_29_2_1_Adder_3_U.ain_s0 ;
wire [28:0] \add_29ns_29s_29_2_1_U8.top_add_29ns_29s_29_2_1_Adder_3_U.b ;
wire [28:0] \add_29ns_29s_29_2_1_U8.top_add_29ns_29s_29_2_1_Adder_3_U.bin_s0 ;
wire \add_29ns_29s_29_2_1_U8.top_add_29ns_29s_29_2_1_Adder_3_U.ce ;
wire \add_29ns_29s_29_2_1_U8.top_add_29ns_29s_29_2_1_Adder_3_U.clk ;
wire \add_29ns_29s_29_2_1_U8.top_add_29ns_29s_29_2_1_Adder_3_U.facout_s1 ;
wire \add_29ns_29s_29_2_1_U8.top_add_29ns_29s_29_2_1_Adder_3_U.facout_s2 ;
wire [13:0] \add_29ns_29s_29_2_1_U8.top_add_29ns_29s_29_2_1_Adder_3_U.fas_s1 ;
wire [14:0] \add_29ns_29s_29_2_1_U8.top_add_29ns_29s_29_2_1_Adder_3_U.fas_s2 ;
wire \add_29ns_29s_29_2_1_U8.top_add_29ns_29s_29_2_1_Adder_3_U.reset ;
wire [28:0] \add_29ns_29s_29_2_1_U8.top_add_29ns_29s_29_2_1_Adder_3_U.s ;
wire [13:0] \add_29ns_29s_29_2_1_U8.top_add_29ns_29s_29_2_1_Adder_3_U.u1.a ;
wire [13:0] \add_29ns_29s_29_2_1_U8.top_add_29ns_29s_29_2_1_Adder_3_U.u1.b ;
wire \add_29ns_29s_29_2_1_U8.top_add_29ns_29s_29_2_1_Adder_3_U.u1.cin ;
wire \add_29ns_29s_29_2_1_U8.top_add_29ns_29s_29_2_1_Adder_3_U.u1.cout ;
wire [13:0] \add_29ns_29s_29_2_1_U8.top_add_29ns_29s_29_2_1_Adder_3_U.u1.s ;
wire [14:0] \add_29ns_29s_29_2_1_U8.top_add_29ns_29s_29_2_1_Adder_3_U.u2.a ;
wire [14:0] \add_29ns_29s_29_2_1_U8.top_add_29ns_29s_29_2_1_Adder_3_U.u2.b ;
wire \add_29ns_29s_29_2_1_U8.top_add_29ns_29s_29_2_1_Adder_3_U.u2.cin ;
wire \add_29ns_29s_29_2_1_U8.top_add_29ns_29s_29_2_1_Adder_3_U.u2.cout ;
wire [14:0] \add_29ns_29s_29_2_1_U8.top_add_29ns_29s_29_2_1_Adder_3_U.u2.s ;
wire \add_29s_29ns_29_2_1_U4.ce ;
wire \add_29s_29ns_29_2_1_U4.clk ;
wire [28:0] \add_29s_29ns_29_2_1_U4.din0 ;
wire [28:0] \add_29s_29ns_29_2_1_U4.din1 ;
wire [28:0] \add_29s_29ns_29_2_1_U4.dout ;
wire \add_29s_29ns_29_2_1_U4.reset ;
wire [28:0] \add_29s_29ns_29_2_1_U4.top_add_29s_29ns_29_2_1_Adder_1_U.a ;
wire [28:0] \add_29s_29ns_29_2_1_U4.top_add_29s_29ns_29_2_1_Adder_1_U.ain_s0 ;
wire [28:0] \add_29s_29ns_29_2_1_U4.top_add_29s_29ns_29_2_1_Adder_1_U.b ;
wire [28:0] \add_29s_29ns_29_2_1_U4.top_add_29s_29ns_29_2_1_Adder_1_U.bin_s0 ;
wire \add_29s_29ns_29_2_1_U4.top_add_29s_29ns_29_2_1_Adder_1_U.ce ;
wire \add_29s_29ns_29_2_1_U4.top_add_29s_29ns_29_2_1_Adder_1_U.clk ;
wire \add_29s_29ns_29_2_1_U4.top_add_29s_29ns_29_2_1_Adder_1_U.facout_s1 ;
wire \add_29s_29ns_29_2_1_U4.top_add_29s_29ns_29_2_1_Adder_1_U.facout_s2 ;
wire [13:0] \add_29s_29ns_29_2_1_U4.top_add_29s_29ns_29_2_1_Adder_1_U.fas_s1 ;
wire [14:0] \add_29s_29ns_29_2_1_U4.top_add_29s_29ns_29_2_1_Adder_1_U.fas_s2 ;
wire \add_29s_29ns_29_2_1_U4.top_add_29s_29ns_29_2_1_Adder_1_U.reset ;
wire [28:0] \add_29s_29ns_29_2_1_U4.top_add_29s_29ns_29_2_1_Adder_1_U.s ;
wire [13:0] \add_29s_29ns_29_2_1_U4.top_add_29s_29ns_29_2_1_Adder_1_U.u1.a ;
wire [13:0] \add_29s_29ns_29_2_1_U4.top_add_29s_29ns_29_2_1_Adder_1_U.u1.b ;
wire \add_29s_29ns_29_2_1_U4.top_add_29s_29ns_29_2_1_Adder_1_U.u1.cin ;
wire \add_29s_29ns_29_2_1_U4.top_add_29s_29ns_29_2_1_Adder_1_U.u1.cout ;
wire [13:0] \add_29s_29ns_29_2_1_U4.top_add_29s_29ns_29_2_1_Adder_1_U.u1.s ;
wire [14:0] \add_29s_29ns_29_2_1_U4.top_add_29s_29ns_29_2_1_Adder_1_U.u2.a ;
wire [14:0] \add_29s_29ns_29_2_1_U4.top_add_29s_29ns_29_2_1_Adder_1_U.u2.b ;
wire \add_29s_29ns_29_2_1_U4.top_add_29s_29ns_29_2_1_Adder_1_U.u2.cin ;
wire \add_29s_29ns_29_2_1_U4.top_add_29s_29ns_29_2_1_Adder_1_U.u2.cout ;
wire [14:0] \add_29s_29ns_29_2_1_U4.top_add_29s_29ns_29_2_1_Adder_1_U.u2.s ;
wire \add_32ns_32ns_32_2_1_U10.ce ;
wire \add_32ns_32ns_32_2_1_U10.clk ;
wire [31:0] \add_32ns_32ns_32_2_1_U10.din0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U10.din1 ;
wire [31:0] \add_32ns_32ns_32_2_1_U10.dout ;
wire \add_32ns_32ns_32_2_1_U10.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_5_U.a ;
wire [31:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_5_U.ain_s0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_5_U.b ;
wire [31:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_5_U.bin_s0 ;
wire \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_5_U.ce ;
wire \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_5_U.clk ;
wire \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_5_U.facout_s1 ;
wire \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_5_U.facout_s2 ;
wire [15:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_5_U.fas_s1 ;
wire [15:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_5_U.fas_s2 ;
wire \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_5_U.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_5_U.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.b ;
wire \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.cin ;
wire \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.b ;
wire \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.cin ;
wire \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.s ;
wire \add_32ns_32ns_32_2_1_U12.ce ;
wire \add_32ns_32ns_32_2_1_U12.clk ;
wire [31:0] \add_32ns_32ns_32_2_1_U12.din0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U12.din1 ;
wire [31:0] \add_32ns_32ns_32_2_1_U12.dout ;
wire \add_32ns_32ns_32_2_1_U12.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.a ;
wire [31:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.ain_s0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.b ;
wire [31:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.bin_s0 ;
wire \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.ce ;
wire \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.clk ;
wire \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.facout_s1 ;
wire \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.facout_s2 ;
wire [15:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.fas_s1 ;
wire [15:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.fas_s2 ;
wire \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.b ;
wire \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.cin ;
wire \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.b ;
wire \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.cin ;
wire \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.s ;
wire \add_32ns_32ns_32_2_1_U13.ce ;
wire \add_32ns_32ns_32_2_1_U13.clk ;
wire [31:0] \add_32ns_32ns_32_2_1_U13.din0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U13.din1 ;
wire [31:0] \add_32ns_32ns_32_2_1_U13.dout ;
wire \add_32ns_32ns_32_2_1_U13.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_5_U.a ;
wire [31:0] \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_5_U.ain_s0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_5_U.b ;
wire [31:0] \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_5_U.bin_s0 ;
wire \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_5_U.ce ;
wire \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_5_U.clk ;
wire \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_5_U.facout_s1 ;
wire \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_5_U.facout_s2 ;
wire [15:0] \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_5_U.fas_s1 ;
wire [15:0] \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_5_U.fas_s2 ;
wire \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_5_U.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_5_U.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.b ;
wire \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.cin ;
wire \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.b ;
wire \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.cin ;
wire \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.s ;
wire \add_33s_33s_33_2_1_U3.ce ;
wire \add_33s_33s_33_2_1_U3.clk ;
wire [32:0] \add_33s_33s_33_2_1_U3.din0 ;
wire [32:0] \add_33s_33s_33_2_1_U3.din1 ;
wire [32:0] \add_33s_33s_33_2_1_U3.dout ;
wire \add_33s_33s_33_2_1_U3.reset ;
wire [32:0] \add_33s_33s_33_2_1_U3.top_add_33s_33s_33_2_1_Adder_0_U.a ;
wire [32:0] \add_33s_33s_33_2_1_U3.top_add_33s_33s_33_2_1_Adder_0_U.ain_s0 ;
wire [32:0] \add_33s_33s_33_2_1_U3.top_add_33s_33s_33_2_1_Adder_0_U.b ;
wire [32:0] \add_33s_33s_33_2_1_U3.top_add_33s_33s_33_2_1_Adder_0_U.bin_s0 ;
wire \add_33s_33s_33_2_1_U3.top_add_33s_33s_33_2_1_Adder_0_U.ce ;
wire \add_33s_33s_33_2_1_U3.top_add_33s_33s_33_2_1_Adder_0_U.clk ;
wire \add_33s_33s_33_2_1_U3.top_add_33s_33s_33_2_1_Adder_0_U.facout_s1 ;
wire \add_33s_33s_33_2_1_U3.top_add_33s_33s_33_2_1_Adder_0_U.facout_s2 ;
wire [15:0] \add_33s_33s_33_2_1_U3.top_add_33s_33s_33_2_1_Adder_0_U.fas_s1 ;
wire [16:0] \add_33s_33s_33_2_1_U3.top_add_33s_33s_33_2_1_Adder_0_U.fas_s2 ;
wire \add_33s_33s_33_2_1_U3.top_add_33s_33s_33_2_1_Adder_0_U.reset ;
wire [32:0] \add_33s_33s_33_2_1_U3.top_add_33s_33s_33_2_1_Adder_0_U.s ;
wire [15:0] \add_33s_33s_33_2_1_U3.top_add_33s_33s_33_2_1_Adder_0_U.u1.a ;
wire [15:0] \add_33s_33s_33_2_1_U3.top_add_33s_33s_33_2_1_Adder_0_U.u1.b ;
wire \add_33s_33s_33_2_1_U3.top_add_33s_33s_33_2_1_Adder_0_U.u1.cin ;
wire \add_33s_33s_33_2_1_U3.top_add_33s_33s_33_2_1_Adder_0_U.u1.cout ;
wire [15:0] \add_33s_33s_33_2_1_U3.top_add_33s_33s_33_2_1_Adder_0_U.u1.s ;
wire [16:0] \add_33s_33s_33_2_1_U3.top_add_33s_33s_33_2_1_Adder_0_U.u2.a ;
wire [16:0] \add_33s_33s_33_2_1_U3.top_add_33s_33s_33_2_1_Adder_0_U.u2.b ;
wire \add_33s_33s_33_2_1_U3.top_add_33s_33s_33_2_1_Adder_0_U.u2.cin ;
wire \add_33s_33s_33_2_1_U3.top_add_33s_33s_33_2_1_Adder_0_U.u2.cout ;
wire [16:0] \add_33s_33s_33_2_1_U3.top_add_33s_33s_33_2_1_Adder_0_U.u2.s ;
wire \add_35s_35s_35_2_1_U11.ce ;
wire \add_35s_35s_35_2_1_U11.clk ;
wire [34:0] \add_35s_35s_35_2_1_U11.din0 ;
wire [34:0] \add_35s_35s_35_2_1_U11.din1 ;
wire [34:0] \add_35s_35s_35_2_1_U11.dout ;
wire \add_35s_35s_35_2_1_U11.reset ;
wire [34:0] \add_35s_35s_35_2_1_U11.top_add_35s_35s_35_2_1_Adder_6_U.a ;
wire [34:0] \add_35s_35s_35_2_1_U11.top_add_35s_35s_35_2_1_Adder_6_U.ain_s0 ;
wire [34:0] \add_35s_35s_35_2_1_U11.top_add_35s_35s_35_2_1_Adder_6_U.b ;
wire [34:0] \add_35s_35s_35_2_1_U11.top_add_35s_35s_35_2_1_Adder_6_U.bin_s0 ;
wire \add_35s_35s_35_2_1_U11.top_add_35s_35s_35_2_1_Adder_6_U.ce ;
wire \add_35s_35s_35_2_1_U11.top_add_35s_35s_35_2_1_Adder_6_U.clk ;
wire \add_35s_35s_35_2_1_U11.top_add_35s_35s_35_2_1_Adder_6_U.facout_s1 ;
wire \add_35s_35s_35_2_1_U11.top_add_35s_35s_35_2_1_Adder_6_U.facout_s2 ;
wire [16:0] \add_35s_35s_35_2_1_U11.top_add_35s_35s_35_2_1_Adder_6_U.fas_s1 ;
wire [17:0] \add_35s_35s_35_2_1_U11.top_add_35s_35s_35_2_1_Adder_6_U.fas_s2 ;
wire \add_35s_35s_35_2_1_U11.top_add_35s_35s_35_2_1_Adder_6_U.reset ;
wire [34:0] \add_35s_35s_35_2_1_U11.top_add_35s_35s_35_2_1_Adder_6_U.s ;
wire [16:0] \add_35s_35s_35_2_1_U11.top_add_35s_35s_35_2_1_Adder_6_U.u1.a ;
wire [16:0] \add_35s_35s_35_2_1_U11.top_add_35s_35s_35_2_1_Adder_6_U.u1.b ;
wire \add_35s_35s_35_2_1_U11.top_add_35s_35s_35_2_1_Adder_6_U.u1.cin ;
wire \add_35s_35s_35_2_1_U11.top_add_35s_35s_35_2_1_Adder_6_U.u1.cout ;
wire [16:0] \add_35s_35s_35_2_1_U11.top_add_35s_35s_35_2_1_Adder_6_U.u1.s ;
wire [17:0] \add_35s_35s_35_2_1_U11.top_add_35s_35s_35_2_1_Adder_6_U.u2.a ;
wire [17:0] \add_35s_35s_35_2_1_U11.top_add_35s_35s_35_2_1_Adder_6_U.u2.b ;
wire \add_35s_35s_35_2_1_U11.top_add_35s_35s_35_2_1_Adder_6_U.u2.cin ;
wire \add_35s_35s_35_2_1_U11.top_add_35s_35s_35_2_1_Adder_6_U.u2.cout ;
wire [17:0] \add_35s_35s_35_2_1_U11.top_add_35s_35s_35_2_1_Adder_6_U.u2.s ;
wire \add_43s_43s_43_2_1_U9.ce ;
wire \add_43s_43s_43_2_1_U9.clk ;
wire [42:0] \add_43s_43s_43_2_1_U9.din0 ;
wire [42:0] \add_43s_43s_43_2_1_U9.din1 ;
wire [42:0] \add_43s_43s_43_2_1_U9.dout ;
wire \add_43s_43s_43_2_1_U9.reset ;
wire [42:0] \add_43s_43s_43_2_1_U9.top_add_43s_43s_43_2_1_Adder_4_U.a ;
wire [42:0] \add_43s_43s_43_2_1_U9.top_add_43s_43s_43_2_1_Adder_4_U.ain_s0 ;
wire [42:0] \add_43s_43s_43_2_1_U9.top_add_43s_43s_43_2_1_Adder_4_U.b ;
wire [42:0] \add_43s_43s_43_2_1_U9.top_add_43s_43s_43_2_1_Adder_4_U.bin_s0 ;
wire \add_43s_43s_43_2_1_U9.top_add_43s_43s_43_2_1_Adder_4_U.ce ;
wire \add_43s_43s_43_2_1_U9.top_add_43s_43s_43_2_1_Adder_4_U.clk ;
wire \add_43s_43s_43_2_1_U9.top_add_43s_43s_43_2_1_Adder_4_U.facout_s1 ;
wire \add_43s_43s_43_2_1_U9.top_add_43s_43s_43_2_1_Adder_4_U.facout_s2 ;
wire [20:0] \add_43s_43s_43_2_1_U9.top_add_43s_43s_43_2_1_Adder_4_U.fas_s1 ;
wire [21:0] \add_43s_43s_43_2_1_U9.top_add_43s_43s_43_2_1_Adder_4_U.fas_s2 ;
wire \add_43s_43s_43_2_1_U9.top_add_43s_43s_43_2_1_Adder_4_U.reset ;
wire [42:0] \add_43s_43s_43_2_1_U9.top_add_43s_43s_43_2_1_Adder_4_U.s ;
wire [20:0] \add_43s_43s_43_2_1_U9.top_add_43s_43s_43_2_1_Adder_4_U.u1.a ;
wire [20:0] \add_43s_43s_43_2_1_U9.top_add_43s_43s_43_2_1_Adder_4_U.u1.b ;
wire \add_43s_43s_43_2_1_U9.top_add_43s_43s_43_2_1_Adder_4_U.u1.cin ;
wire \add_43s_43s_43_2_1_U9.top_add_43s_43s_43_2_1_Adder_4_U.u1.cout ;
wire [20:0] \add_43s_43s_43_2_1_U9.top_add_43s_43s_43_2_1_Adder_4_U.u1.s ;
wire [21:0] \add_43s_43s_43_2_1_U9.top_add_43s_43s_43_2_1_Adder_4_U.u2.a ;
wire [21:0] \add_43s_43s_43_2_1_U9.top_add_43s_43s_43_2_1_Adder_4_U.u2.b ;
wire \add_43s_43s_43_2_1_U9.top_add_43s_43s_43_2_1_Adder_4_U.u2.cin ;
wire \add_43s_43s_43_2_1_U9.top_add_43s_43s_43_2_1_Adder_4_U.u2.cout ;
wire [21:0] \add_43s_43s_43_2_1_U9.top_add_43s_43s_43_2_1_Adder_4_U.u2.s ;
wire [2:0] add_ln69_fu_232_p2;
wire and_ln785_1_fu_550_p2;
wire and_ln785_fu_545_p2;
wire and_ln786_fu_512_p2;
wire ap_CS_fsm_state1;
wire ap_CS_fsm_state10;
wire ap_CS_fsm_state11;
wire ap_CS_fsm_state12;
wire ap_CS_fsm_state13;
wire ap_CS_fsm_state14;
wire ap_CS_fsm_state15;
wire ap_CS_fsm_state16;
wire ap_CS_fsm_state17;
wire ap_CS_fsm_state18;
wire ap_CS_fsm_state19;
wire ap_CS_fsm_state2;
wire ap_CS_fsm_state20;
wire ap_CS_fsm_state21;
wire ap_CS_fsm_state22;
wire ap_CS_fsm_state23;
wire ap_CS_fsm_state24;
wire ap_CS_fsm_state25;
wire ap_CS_fsm_state26;
wire ap_CS_fsm_state27;
wire ap_CS_fsm_state28;
wire ap_CS_fsm_state29;
wire ap_CS_fsm_state30;
wire ap_CS_fsm_state4;
wire ap_CS_fsm_state5;
wire ap_CS_fsm_state6;
wire ap_CS_fsm_state7;
wire ap_CS_fsm_state8;
wire ap_CS_fsm_state9;
wire [29:0] ap_NS_fsm;
wire ap_clk;
wire ap_done;
wire ap_idle;
wire ap_ready;
wire ap_rst;
wire ap_start;
wire [3:0] grp_fu_189_p0;
wire [3:0] grp_fu_189_p1;
wire [7:0] grp_fu_189_p2;
wire [15:0] grp_fu_251_p1;
wire [15:0] grp_fu_251_p2;
wire [32:0] grp_fu_283_p0;
wire [32:0] grp_fu_283_p1;
wire [32:0] grp_fu_283_p2;
wire [28:0] grp_fu_312_p0;
wire [28:0] grp_fu_312_p2;
wire [28:0] grp_fu_345_p2;
wire [28:0] grp_fu_374_p2;
wire [28:0] grp_fu_391_p1;
wire [28:0] grp_fu_391_p2;
wire [28:0] grp_fu_400_p1;
wire [28:0] grp_fu_400_p2;
wire [42:0] grp_fu_420_p0;
wire [42:0] grp_fu_420_p1;
wire [42:0] grp_fu_420_p2;
wire [31:0] grp_fu_486_p2;
wire [34:0] grp_fu_600_p0;
wire [34:0] grp_fu_600_p1;
wire [34:0] grp_fu_600_p2;
wire [31:0] grp_fu_621_p2;
wire [31:0] grp_fu_645_p2;
wire icmp_ln851_1_fu_430_p2;
wire icmp_ln851_2_fu_606_p2;
wire icmp_ln851_fu_293_p2;
wire lhs_V_fu_382_p2;
wire \mul_4ns_4ns_8_4_1_U1.ce ;
wire \mul_4ns_4ns_8_4_1_U1.clk ;
wire [3:0] \mul_4ns_4ns_8_4_1_U1.din0 ;
wire [3:0] \mul_4ns_4ns_8_4_1_U1.din1 ;
wire [7:0] \mul_4ns_4ns_8_4_1_U1.dout ;
wire \mul_4ns_4ns_8_4_1_U1.reset ;
wire [3:0] \mul_4ns_4ns_8_4_1_U1.top_mul_4ns_4ns_8_4_1_Mul_DSP_0_U.a ;
wire [3:0] \mul_4ns_4ns_8_4_1_U1.top_mul_4ns_4ns_8_4_1_Mul_DSP_0_U.b ;
wire \mul_4ns_4ns_8_4_1_U1.top_mul_4ns_4ns_8_4_1_Mul_DSP_0_U.ce ;
wire \mul_4ns_4ns_8_4_1_U1.top_mul_4ns_4ns_8_4_1_Mul_DSP_0_U.clk ;
wire [7:0] \mul_4ns_4ns_8_4_1_U1.top_mul_4ns_4ns_8_4_1_Mul_DSP_0_U.p ;
wire [7:0] \mul_4ns_4ns_8_4_1_U1.top_mul_4ns_4ns_8_4_1_Mul_DSP_0_U.tmp_product ;
wire [31:0] op_0;
wire [1:0] op_10;
wire [31:0] op_11;
wire [31:0] op_12;
wire op_13;
wire [7:0] op_16;
wire [31:0] op_17;
wire [3:0] op_18_V_fu_555_p3;
wire [31:0] op_19;
wire [3:0] op_2;
wire [8:0] op_22_V_fu_262_p2;
wire [1:0] op_3;
wire [31:0] op_30;
wire op_30_ap_vld;
wire op_5;
wire [1:0] op_6_V_fu_203_p1;
wire [1:0] op_6_V_fu_203_p2;
wire op_8_V_fu_209_p2;
wire or_ln340_1_fu_521_p2;
wire or_ln340_fu_516_p2;
wire or_ln785_1_fu_540_p2;
wire or_ln785_fu_491_p2;
wire overflow_fu_507_p2;
wire p_Result_1_fu_563_p3;
wire p_Result_2_fu_626_p3;
wire [1:0] p_Result_3_fu_349_p1;
wire p_Result_3_fu_349_p3;
wire p_Result_s_fu_318_p3;
wire [3:0] p_Val2_1_fu_495_p3;
wire r_fu_356_p1;
wire [2:0] ret_1_fu_452_p2;
wire [28:0] ret_V_2_fu_330_p3;
wire [31:0] ret_V_7_fu_638_p3;
wire [2:0] ret_V_fu_226_p2;
wire [13:0] rhs_2_fu_272_p3;
wire [33:0] rhs_6_fu_589_p3;
wire [28:0] select_ln1192_fu_337_p3;
wire [3:0] select_ln340_fu_527_p3;
wire [31:0] select_ln353_fu_575_p3;
wire [15:0] select_ln546_fu_237_p3;
wire [28:0] select_ln69_1_fu_366_p3;
wire [2:0] select_ln69_fu_215_p3;
wire select_ln769_fu_359_p3;
wire [31:0] select_ln850_1_fu_570_p3;
wire [31:0] select_ln850_2_fu_633_p3;
wire [28:0] select_ln850_fu_325_p3;
wire [31:0] sext_ln1192_fu_268_p0;
wire [1:0] sext_ln1347_1_fu_449_p0;
wire [2:0] sext_ln1347_1_fu_449_p1;
wire [1:0] sext_ln1347_fu_446_p0;
wire [2:0] sext_ln1347_fu_446_p1;
wire [8:0] sext_ln69_1_fu_259_p1;
wire [8:0] sext_ln69_fu_256_p1;
wire [31:0] sext_ln703_1_fu_405_p0;
wire [2:0] sext_ln703_fu_223_p1;
wire [1:0] sext_ln781_fu_244_p0;
wire [3:0] sext_ln781_fu_244_p1;
wire [28:0] sext_ln850_fu_309_p1;
wire [1:0] sext_ln874_fu_378_p0;
wire [31:0] sext_ln874_fu_378_p1;
wire \shl_16ns_4ns_16_7_1_U2.ce ;
wire \shl_16ns_4ns_16_7_1_U2.clk ;
wire [15:0] \shl_16ns_4ns_16_7_1_U2.din0 ;
wire [15:0] \shl_16ns_4ns_16_7_1_U2.din1 ;
wire [3:0] \shl_16ns_4ns_16_7_1_U2.din1_cast ;
wire [3:0] \shl_16ns_4ns_16_7_1_U2.din1_mask ;
wire [15:0] \shl_16ns_4ns_16_7_1_U2.dout ;
wire \shl_16ns_4ns_16_7_1_U2.reset ;
wire [38:0] tmp_7_fu_409_p3;
wire [1:0] trunc_ln69_1_fu_199_p1;
wire trunc_ln69_fu_195_p1;
wire [1:0] trunc_ln731_fu_466_p1;
wire [31:0] trunc_ln851_1_fu_426_p0;
wire [9:0] trunc_ln851_1_fu_426_p1;
wire [1:0] trunc_ln851_2_fu_582_p1;
wire [31:0] trunc_ln851_fu_289_p0;
wire [4:0] trunc_ln851_fu_289_p1;
wire xor_ln785_1_fu_535_p2;
wire xor_ln785_fu_502_p2;
wire [7:0] zext_ln1345_fu_185_p1;


assign add_ln69_fu_232_p2 = ret_V_fu_226_p2 + select_ln69_reg_675;
assign op_22_V_fu_262_p2 = $signed(add_ln69_reg_680) + $signed(ret_reg_685);
assign ret_V_fu_226_p2 = $signed(op_6_V_reg_670) + $signed(2'h1);
assign _038_ = _043_ & ap_CS_fsm[0];
assign _039_ = ap_start & ap_CS_fsm[0];
assign and_ln785_1_fu_550_p2 = p_Result_5_reg_841 & and_ln785_fu_545_p2;
assign and_ln785_fu_545_p2 = tmp_5_reg_848 & or_ln785_1_fu_540_p2;
assign and_ln786_fu_512_p2 = tmp_5_reg_848 & p_Result_5_reg_841;
assign overflow_fu_507_p2 = xor_ln785_fu_502_p2 & or_ln785_reg_855;
assign _040_ = icmp_ln851_1_reg_812 & ap_CS_fsm[21];
assign _041_ = icmp_ln851_2_reg_891 & ap_CS_fsm[26];
assign _042_ = ap_CS_fsm[8] & icmp_ln851_reg_715;
assign xor_ln785_1_fu_535_p2 = ~ or_ln785_reg_855;
assign xor_ln785_fu_502_p2 = ~ p_Result_4_reg_829;
assign _043_ = ~ ap_start;
always @(posedge \add_29ns_29ns_29_2_1_U5.top_add_29ns_29ns_29_2_1_Adder_2_U.clk )
\add_29ns_29ns_29_2_1_U5.top_add_29ns_29ns_29_2_1_Adder_2_U.bin_s1  <= _045_;
always @(posedge \add_29ns_29ns_29_2_1_U5.top_add_29ns_29ns_29_2_1_Adder_2_U.clk )
\add_29ns_29ns_29_2_1_U5.top_add_29ns_29ns_29_2_1_Adder_2_U.ain_s1  <= _044_;
always @(posedge \add_29ns_29ns_29_2_1_U5.top_add_29ns_29ns_29_2_1_Adder_2_U.clk )
\add_29ns_29ns_29_2_1_U5.top_add_29ns_29ns_29_2_1_Adder_2_U.sum_s1  <= _047_;
always @(posedge \add_29ns_29ns_29_2_1_U5.top_add_29ns_29ns_29_2_1_Adder_2_U.clk )
\add_29ns_29ns_29_2_1_U5.top_add_29ns_29ns_29_2_1_Adder_2_U.carry_s1  <= _046_;
assign _045_ = \add_29ns_29ns_29_2_1_U5.top_add_29ns_29ns_29_2_1_Adder_2_U.ce  ? \add_29ns_29ns_29_2_1_U5.top_add_29ns_29ns_29_2_1_Adder_2_U.b [28:14] : \add_29ns_29ns_29_2_1_U5.top_add_29ns_29ns_29_2_1_Adder_2_U.bin_s1 ;
assign _044_ = \add_29ns_29ns_29_2_1_U5.top_add_29ns_29ns_29_2_1_Adder_2_U.ce  ? \add_29ns_29ns_29_2_1_U5.top_add_29ns_29ns_29_2_1_Adder_2_U.a [28:14] : \add_29ns_29ns_29_2_1_U5.top_add_29ns_29ns_29_2_1_Adder_2_U.ain_s1 ;
assign _046_ = \add_29ns_29ns_29_2_1_U5.top_add_29ns_29ns_29_2_1_Adder_2_U.ce  ? \add_29ns_29ns_29_2_1_U5.top_add_29ns_29ns_29_2_1_Adder_2_U.facout_s1  : \add_29ns_29ns_29_2_1_U5.top_add_29ns_29ns_29_2_1_Adder_2_U.carry_s1 ;
assign _047_ = \add_29ns_29ns_29_2_1_U5.top_add_29ns_29ns_29_2_1_Adder_2_U.ce  ? \add_29ns_29ns_29_2_1_U5.top_add_29ns_29ns_29_2_1_Adder_2_U.fas_s1  : \add_29ns_29ns_29_2_1_U5.top_add_29ns_29ns_29_2_1_Adder_2_U.sum_s1 ;
assign _048_ = \add_29ns_29ns_29_2_1_U5.top_add_29ns_29ns_29_2_1_Adder_2_U.u1.a  + \add_29ns_29ns_29_2_1_U5.top_add_29ns_29ns_29_2_1_Adder_2_U.u1.b ;
assign { \add_29ns_29ns_29_2_1_U5.top_add_29ns_29ns_29_2_1_Adder_2_U.u1.cout , \add_29ns_29ns_29_2_1_U5.top_add_29ns_29ns_29_2_1_Adder_2_U.u1.s  } = _048_ + \add_29ns_29ns_29_2_1_U5.top_add_29ns_29ns_29_2_1_Adder_2_U.u1.cin ;
assign _049_ = \add_29ns_29ns_29_2_1_U5.top_add_29ns_29ns_29_2_1_Adder_2_U.u2.a  + \add_29ns_29ns_29_2_1_U5.top_add_29ns_29ns_29_2_1_Adder_2_U.u2.b ;
assign { \add_29ns_29ns_29_2_1_U5.top_add_29ns_29ns_29_2_1_Adder_2_U.u2.cout , \add_29ns_29ns_29_2_1_U5.top_add_29ns_29ns_29_2_1_Adder_2_U.u2.s  } = _049_ + \add_29ns_29ns_29_2_1_U5.top_add_29ns_29ns_29_2_1_Adder_2_U.u2.cin ;
always @(posedge \add_29ns_29ns_29_2_1_U6.top_add_29ns_29ns_29_2_1_Adder_2_U.clk )
\add_29ns_29ns_29_2_1_U6.top_add_29ns_29ns_29_2_1_Adder_2_U.bin_s1  <= _051_;
always @(posedge \add_29ns_29ns_29_2_1_U6.top_add_29ns_29ns_29_2_1_Adder_2_U.clk )
\add_29ns_29ns_29_2_1_U6.top_add_29ns_29ns_29_2_1_Adder_2_U.ain_s1  <= _050_;
always @(posedge \add_29ns_29ns_29_2_1_U6.top_add_29ns_29ns_29_2_1_Adder_2_U.clk )
\add_29ns_29ns_29_2_1_U6.top_add_29ns_29ns_29_2_1_Adder_2_U.sum_s1  <= _053_;
always @(posedge \add_29ns_29ns_29_2_1_U6.top_add_29ns_29ns_29_2_1_Adder_2_U.clk )
\add_29ns_29ns_29_2_1_U6.top_add_29ns_29ns_29_2_1_Adder_2_U.carry_s1  <= _052_;
assign _051_ = \add_29ns_29ns_29_2_1_U6.top_add_29ns_29ns_29_2_1_Adder_2_U.ce  ? \add_29ns_29ns_29_2_1_U6.top_add_29ns_29ns_29_2_1_Adder_2_U.b [28:14] : \add_29ns_29ns_29_2_1_U6.top_add_29ns_29ns_29_2_1_Adder_2_U.bin_s1 ;
assign _050_ = \add_29ns_29ns_29_2_1_U6.top_add_29ns_29ns_29_2_1_Adder_2_U.ce  ? \add_29ns_29ns_29_2_1_U6.top_add_29ns_29ns_29_2_1_Adder_2_U.a [28:14] : \add_29ns_29ns_29_2_1_U6.top_add_29ns_29ns_29_2_1_Adder_2_U.ain_s1 ;
assign _052_ = \add_29ns_29ns_29_2_1_U6.top_add_29ns_29ns_29_2_1_Adder_2_U.ce  ? \add_29ns_29ns_29_2_1_U6.top_add_29ns_29ns_29_2_1_Adder_2_U.facout_s1  : \add_29ns_29ns_29_2_1_U6.top_add_29ns_29ns_29_2_1_Adder_2_U.carry_s1 ;
assign _053_ = \add_29ns_29ns_29_2_1_U6.top_add_29ns_29ns_29_2_1_Adder_2_U.ce  ? \add_29ns_29ns_29_2_1_U6.top_add_29ns_29ns_29_2_1_Adder_2_U.fas_s1  : \add_29ns_29ns_29_2_1_U6.top_add_29ns_29ns_29_2_1_Adder_2_U.sum_s1 ;
assign _054_ = \add_29ns_29ns_29_2_1_U6.top_add_29ns_29ns_29_2_1_Adder_2_U.u1.a  + \add_29ns_29ns_29_2_1_U6.top_add_29ns_29ns_29_2_1_Adder_2_U.u1.b ;
assign { \add_29ns_29ns_29_2_1_U6.top_add_29ns_29ns_29_2_1_Adder_2_U.u1.cout , \add_29ns_29ns_29_2_1_U6.top_add_29ns_29ns_29_2_1_Adder_2_U.u1.s  } = _054_ + \add_29ns_29ns_29_2_1_U6.top_add_29ns_29ns_29_2_1_Adder_2_U.u1.cin ;
assign _055_ = \add_29ns_29ns_29_2_1_U6.top_add_29ns_29ns_29_2_1_Adder_2_U.u2.a  + \add_29ns_29ns_29_2_1_U6.top_add_29ns_29ns_29_2_1_Adder_2_U.u2.b ;
assign { \add_29ns_29ns_29_2_1_U6.top_add_29ns_29ns_29_2_1_Adder_2_U.u2.cout , \add_29ns_29ns_29_2_1_U6.top_add_29ns_29ns_29_2_1_Adder_2_U.u2.s  } = _055_ + \add_29ns_29ns_29_2_1_U6.top_add_29ns_29ns_29_2_1_Adder_2_U.u2.cin ;
always @(posedge \add_29ns_29ns_29_2_1_U7.top_add_29ns_29ns_29_2_1_Adder_2_U.clk )
\add_29ns_29ns_29_2_1_U7.top_add_29ns_29ns_29_2_1_Adder_2_U.bin_s1  <= _057_;
always @(posedge \add_29ns_29ns_29_2_1_U7.top_add_29ns_29ns_29_2_1_Adder_2_U.clk )
\add_29ns_29ns_29_2_1_U7.top_add_29ns_29ns_29_2_1_Adder_2_U.ain_s1  <= _056_;
always @(posedge \add_29ns_29ns_29_2_1_U7.top_add_29ns_29ns_29_2_1_Adder_2_U.clk )
\add_29ns_29ns_29_2_1_U7.top_add_29ns_29ns_29_2_1_Adder_2_U.sum_s1  <= _059_;
always @(posedge \add_29ns_29ns_29_2_1_U7.top_add_29ns_29ns_29_2_1_Adder_2_U.clk )
\add_29ns_29ns_29_2_1_U7.top_add_29ns_29ns_29_2_1_Adder_2_U.carry_s1  <= _058_;
assign _057_ = \add_29ns_29ns_29_2_1_U7.top_add_29ns_29ns_29_2_1_Adder_2_U.ce  ? \add_29ns_29ns_29_2_1_U7.top_add_29ns_29ns_29_2_1_Adder_2_U.b [28:14] : \add_29ns_29ns_29_2_1_U7.top_add_29ns_29ns_29_2_1_Adder_2_U.bin_s1 ;
assign _056_ = \add_29ns_29ns_29_2_1_U7.top_add_29ns_29ns_29_2_1_Adder_2_U.ce  ? \add_29ns_29ns_29_2_1_U7.top_add_29ns_29ns_29_2_1_Adder_2_U.a [28:14] : \add_29ns_29ns_29_2_1_U7.top_add_29ns_29ns_29_2_1_Adder_2_U.ain_s1 ;
assign _058_ = \add_29ns_29ns_29_2_1_U7.top_add_29ns_29ns_29_2_1_Adder_2_U.ce  ? \add_29ns_29ns_29_2_1_U7.top_add_29ns_29ns_29_2_1_Adder_2_U.facout_s1  : \add_29ns_29ns_29_2_1_U7.top_add_29ns_29ns_29_2_1_Adder_2_U.carry_s1 ;
assign _059_ = \add_29ns_29ns_29_2_1_U7.top_add_29ns_29ns_29_2_1_Adder_2_U.ce  ? \add_29ns_29ns_29_2_1_U7.top_add_29ns_29ns_29_2_1_Adder_2_U.fas_s1  : \add_29ns_29ns_29_2_1_U7.top_add_29ns_29ns_29_2_1_Adder_2_U.sum_s1 ;
assign _060_ = \add_29ns_29ns_29_2_1_U7.top_add_29ns_29ns_29_2_1_Adder_2_U.u1.a  + \add_29ns_29ns_29_2_1_U7.top_add_29ns_29ns_29_2_1_Adder_2_U.u1.b ;
assign { \add_29ns_29ns_29_2_1_U7.top_add_29ns_29ns_29_2_1_Adder_2_U.u1.cout , \add_29ns_29ns_29_2_1_U7.top_add_29ns_29ns_29_2_1_Adder_2_U.u1.s  } = _060_ + \add_29ns_29ns_29_2_1_U7.top_add_29ns_29ns_29_2_1_Adder_2_U.u1.cin ;
assign _061_ = \add_29ns_29ns_29_2_1_U7.top_add_29ns_29ns_29_2_1_Adder_2_U.u2.a  + \add_29ns_29ns_29_2_1_U7.top_add_29ns_29ns_29_2_1_Adder_2_U.u2.b ;
assign { \add_29ns_29ns_29_2_1_U7.top_add_29ns_29ns_29_2_1_Adder_2_U.u2.cout , \add_29ns_29ns_29_2_1_U7.top_add_29ns_29ns_29_2_1_Adder_2_U.u2.s  } = _061_ + \add_29ns_29ns_29_2_1_U7.top_add_29ns_29ns_29_2_1_Adder_2_U.u2.cin ;
always @(posedge \add_29ns_29s_29_2_1_U8.top_add_29ns_29s_29_2_1_Adder_3_U.clk )
\add_29ns_29s_29_2_1_U8.top_add_29ns_29s_29_2_1_Adder_3_U.bin_s1  <= _063_;
always @(posedge \add_29ns_29s_29_2_1_U8.top_add_29ns_29s_29_2_1_Adder_3_U.clk )
\add_29ns_29s_29_2_1_U8.top_add_29ns_29s_29_2_1_Adder_3_U.ain_s1  <= _062_;
always @(posedge \add_29ns_29s_29_2_1_U8.top_add_29ns_29s_29_2_1_Adder_3_U.clk )
\add_29ns_29s_29_2_1_U8.top_add_29ns_29s_29_2_1_Adder_3_U.sum_s1  <= _065_;
always @(posedge \add_29ns_29s_29_2_1_U8.top_add_29ns_29s_29_2_1_Adder_3_U.clk )
\add_29ns_29s_29_2_1_U8.top_add_29ns_29s_29_2_1_Adder_3_U.carry_s1  <= _064_;
assign _063_ = \add_29ns_29s_29_2_1_U8.top_add_29ns_29s_29_2_1_Adder_3_U.ce  ? \add_29ns_29s_29_2_1_U8.top_add_29ns_29s_29_2_1_Adder_3_U.b [28:14] : \add_29ns_29s_29_2_1_U8.top_add_29ns_29s_29_2_1_Adder_3_U.bin_s1 ;
assign _062_ = \add_29ns_29s_29_2_1_U8.top_add_29ns_29s_29_2_1_Adder_3_U.ce  ? \add_29ns_29s_29_2_1_U8.top_add_29ns_29s_29_2_1_Adder_3_U.a [28:14] : \add_29ns_29s_29_2_1_U8.top_add_29ns_29s_29_2_1_Adder_3_U.ain_s1 ;
assign _064_ = \add_29ns_29s_29_2_1_U8.top_add_29ns_29s_29_2_1_Adder_3_U.ce  ? \add_29ns_29s_29_2_1_U8.top_add_29ns_29s_29_2_1_Adder_3_U.facout_s1  : \add_29ns_29s_29_2_1_U8.top_add_29ns_29s_29_2_1_Adder_3_U.carry_s1 ;
assign _065_ = \add_29ns_29s_29_2_1_U8.top_add_29ns_29s_29_2_1_Adder_3_U.ce  ? \add_29ns_29s_29_2_1_U8.top_add_29ns_29s_29_2_1_Adder_3_U.fas_s1  : \add_29ns_29s_29_2_1_U8.top_add_29ns_29s_29_2_1_Adder_3_U.sum_s1 ;
assign _066_ = \add_29ns_29s_29_2_1_U8.top_add_29ns_29s_29_2_1_Adder_3_U.u1.a  + \add_29ns_29s_29_2_1_U8.top_add_29ns_29s_29_2_1_Adder_3_U.u1.b ;
assign { \add_29ns_29s_29_2_1_U8.top_add_29ns_29s_29_2_1_Adder_3_U.u1.cout , \add_29ns_29s_29_2_1_U8.top_add_29ns_29s_29_2_1_Adder_3_U.u1.s  } = _066_ + \add_29ns_29s_29_2_1_U8.top_add_29ns_29s_29_2_1_Adder_3_U.u1.cin ;
assign _067_ = \add_29ns_29s_29_2_1_U8.top_add_29ns_29s_29_2_1_Adder_3_U.u2.a  + \add_29ns_29s_29_2_1_U8.top_add_29ns_29s_29_2_1_Adder_3_U.u2.b ;
assign { \add_29ns_29s_29_2_1_U8.top_add_29ns_29s_29_2_1_Adder_3_U.u2.cout , \add_29ns_29s_29_2_1_U8.top_add_29ns_29s_29_2_1_Adder_3_U.u2.s  } = _067_ + \add_29ns_29s_29_2_1_U8.top_add_29ns_29s_29_2_1_Adder_3_U.u2.cin ;
always @(posedge \add_29s_29ns_29_2_1_U4.top_add_29s_29ns_29_2_1_Adder_1_U.clk )
\add_29s_29ns_29_2_1_U4.top_add_29s_29ns_29_2_1_Adder_1_U.bin_s1  <= _069_;
always @(posedge \add_29s_29ns_29_2_1_U4.top_add_29s_29ns_29_2_1_Adder_1_U.clk )
\add_29s_29ns_29_2_1_U4.top_add_29s_29ns_29_2_1_Adder_1_U.ain_s1  <= _068_;
always @(posedge \add_29s_29ns_29_2_1_U4.top_add_29s_29ns_29_2_1_Adder_1_U.clk )
\add_29s_29ns_29_2_1_U4.top_add_29s_29ns_29_2_1_Adder_1_U.sum_s1  <= _071_;
always @(posedge \add_29s_29ns_29_2_1_U4.top_add_29s_29ns_29_2_1_Adder_1_U.clk )
\add_29s_29ns_29_2_1_U4.top_add_29s_29ns_29_2_1_Adder_1_U.carry_s1  <= _070_;
assign _069_ = \add_29s_29ns_29_2_1_U4.top_add_29s_29ns_29_2_1_Adder_1_U.ce  ? \add_29s_29ns_29_2_1_U4.top_add_29s_29ns_29_2_1_Adder_1_U.b [28:14] : \add_29s_29ns_29_2_1_U4.top_add_29s_29ns_29_2_1_Adder_1_U.bin_s1 ;
assign _068_ = \add_29s_29ns_29_2_1_U4.top_add_29s_29ns_29_2_1_Adder_1_U.ce  ? \add_29s_29ns_29_2_1_U4.top_add_29s_29ns_29_2_1_Adder_1_U.a [28:14] : \add_29s_29ns_29_2_1_U4.top_add_29s_29ns_29_2_1_Adder_1_U.ain_s1 ;
assign _070_ = \add_29s_29ns_29_2_1_U4.top_add_29s_29ns_29_2_1_Adder_1_U.ce  ? \add_29s_29ns_29_2_1_U4.top_add_29s_29ns_29_2_1_Adder_1_U.facout_s1  : \add_29s_29ns_29_2_1_U4.top_add_29s_29ns_29_2_1_Adder_1_U.carry_s1 ;
assign _071_ = \add_29s_29ns_29_2_1_U4.top_add_29s_29ns_29_2_1_Adder_1_U.ce  ? \add_29s_29ns_29_2_1_U4.top_add_29s_29ns_29_2_1_Adder_1_U.fas_s1  : \add_29s_29ns_29_2_1_U4.top_add_29s_29ns_29_2_1_Adder_1_U.sum_s1 ;
assign _072_ = \add_29s_29ns_29_2_1_U4.top_add_29s_29ns_29_2_1_Adder_1_U.u1.a  + \add_29s_29ns_29_2_1_U4.top_add_29s_29ns_29_2_1_Adder_1_U.u1.b ;
assign { \add_29s_29ns_29_2_1_U4.top_add_29s_29ns_29_2_1_Adder_1_U.u1.cout , \add_29s_29ns_29_2_1_U4.top_add_29s_29ns_29_2_1_Adder_1_U.u1.s  } = _072_ + \add_29s_29ns_29_2_1_U4.top_add_29s_29ns_29_2_1_Adder_1_U.u1.cin ;
assign _073_ = \add_29s_29ns_29_2_1_U4.top_add_29s_29ns_29_2_1_Adder_1_U.u2.a  + \add_29s_29ns_29_2_1_U4.top_add_29s_29ns_29_2_1_Adder_1_U.u2.b ;
assign { \add_29s_29ns_29_2_1_U4.top_add_29s_29ns_29_2_1_Adder_1_U.u2.cout , \add_29s_29ns_29_2_1_U4.top_add_29s_29ns_29_2_1_Adder_1_U.u2.s  } = _073_ + \add_29s_29ns_29_2_1_U4.top_add_29s_29ns_29_2_1_Adder_1_U.u2.cin ;
always @(posedge \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_5_U.clk )
\add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_5_U.bin_s1  <= _075_;
always @(posedge \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_5_U.clk )
\add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_5_U.ain_s1  <= _074_;
always @(posedge \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_5_U.clk )
\add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_5_U.sum_s1  <= _077_;
always @(posedge \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_5_U.clk )
\add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_5_U.carry_s1  <= _076_;
assign _075_ = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_5_U.ce  ? \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_5_U.b [31:16] : \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_5_U.bin_s1 ;
assign _074_ = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_5_U.ce  ? \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_5_U.a [31:16] : \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_5_U.ain_s1 ;
assign _076_ = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_5_U.ce  ? \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_5_U.facout_s1  : \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_5_U.carry_s1 ;
assign _077_ = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_5_U.ce  ? \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_5_U.fas_s1  : \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_5_U.sum_s1 ;
assign _078_ = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.a  + \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.b ;
assign { \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.cout , \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.s  } = _078_ + \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.cin ;
assign _079_ = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.a  + \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.b ;
assign { \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.cout , \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.s  } = _079_ + \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.cin ;
always @(posedge \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.clk )
\add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.bin_s1  <= _081_;
always @(posedge \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.clk )
\add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.ain_s1  <= _080_;
always @(posedge \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.clk )
\add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.sum_s1  <= _083_;
always @(posedge \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.clk )
\add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.carry_s1  <= _082_;
assign _081_ = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.ce  ? \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.b [31:16] : \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.bin_s1 ;
assign _080_ = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.ce  ? \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.a [31:16] : \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.ain_s1 ;
assign _082_ = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.ce  ? \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.facout_s1  : \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.carry_s1 ;
assign _083_ = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.ce  ? \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.fas_s1  : \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.sum_s1 ;
assign _084_ = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.a  + \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.b ;
assign { \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.cout , \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.s  } = _084_ + \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.cin ;
assign _085_ = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.a  + \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.b ;
assign { \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.cout , \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.s  } = _085_ + \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.cin ;
always @(posedge \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_5_U.clk )
\add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_5_U.bin_s1  <= _087_;
always @(posedge \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_5_U.clk )
\add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_5_U.ain_s1  <= _086_;
always @(posedge \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_5_U.clk )
\add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_5_U.sum_s1  <= _089_;
always @(posedge \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_5_U.clk )
\add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_5_U.carry_s1  <= _088_;
assign _087_ = \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_5_U.ce  ? \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_5_U.b [31:16] : \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_5_U.bin_s1 ;
assign _086_ = \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_5_U.ce  ? \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_5_U.a [31:16] : \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_5_U.ain_s1 ;
assign _088_ = \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_5_U.ce  ? \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_5_U.facout_s1  : \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_5_U.carry_s1 ;
assign _089_ = \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_5_U.ce  ? \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_5_U.fas_s1  : \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_5_U.sum_s1 ;
assign _090_ = \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.a  + \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.b ;
assign { \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.cout , \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.s  } = _090_ + \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.cin ;
assign _091_ = \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.a  + \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.b ;
assign { \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.cout , \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.s  } = _091_ + \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.cin ;
always @(posedge \add_33s_33s_33_2_1_U3.top_add_33s_33s_33_2_1_Adder_0_U.clk )
\add_33s_33s_33_2_1_U3.top_add_33s_33s_33_2_1_Adder_0_U.bin_s1  <= _093_;
always @(posedge \add_33s_33s_33_2_1_U3.top_add_33s_33s_33_2_1_Adder_0_U.clk )
\add_33s_33s_33_2_1_U3.top_add_33s_33s_33_2_1_Adder_0_U.ain_s1  <= _092_;
always @(posedge \add_33s_33s_33_2_1_U3.top_add_33s_33s_33_2_1_Adder_0_U.clk )
\add_33s_33s_33_2_1_U3.top_add_33s_33s_33_2_1_Adder_0_U.sum_s1  <= _095_;
always @(posedge \add_33s_33s_33_2_1_U3.top_add_33s_33s_33_2_1_Adder_0_U.clk )
\add_33s_33s_33_2_1_U3.top_add_33s_33s_33_2_1_Adder_0_U.carry_s1  <= _094_;
assign _093_ = \add_33s_33s_33_2_1_U3.top_add_33s_33s_33_2_1_Adder_0_U.ce  ? \add_33s_33s_33_2_1_U3.top_add_33s_33s_33_2_1_Adder_0_U.b [32:16] : \add_33s_33s_33_2_1_U3.top_add_33s_33s_33_2_1_Adder_0_U.bin_s1 ;
assign _092_ = \add_33s_33s_33_2_1_U3.top_add_33s_33s_33_2_1_Adder_0_U.ce  ? \add_33s_33s_33_2_1_U3.top_add_33s_33s_33_2_1_Adder_0_U.a [32:16] : \add_33s_33s_33_2_1_U3.top_add_33s_33s_33_2_1_Adder_0_U.ain_s1 ;
assign _094_ = \add_33s_33s_33_2_1_U3.top_add_33s_33s_33_2_1_Adder_0_U.ce  ? \add_33s_33s_33_2_1_U3.top_add_33s_33s_33_2_1_Adder_0_U.facout_s1  : \add_33s_33s_33_2_1_U3.top_add_33s_33s_33_2_1_Adder_0_U.carry_s1 ;
assign _095_ = \add_33s_33s_33_2_1_U3.top_add_33s_33s_33_2_1_Adder_0_U.ce  ? \add_33s_33s_33_2_1_U3.top_add_33s_33s_33_2_1_Adder_0_U.fas_s1  : \add_33s_33s_33_2_1_U3.top_add_33s_33s_33_2_1_Adder_0_U.sum_s1 ;
assign _096_ = \add_33s_33s_33_2_1_U3.top_add_33s_33s_33_2_1_Adder_0_U.u1.a  + \add_33s_33s_33_2_1_U3.top_add_33s_33s_33_2_1_Adder_0_U.u1.b ;
assign { \add_33s_33s_33_2_1_U3.top_add_33s_33s_33_2_1_Adder_0_U.u1.cout , \add_33s_33s_33_2_1_U3.top_add_33s_33s_33_2_1_Adder_0_U.u1.s  } = _096_ + \add_33s_33s_33_2_1_U3.top_add_33s_33s_33_2_1_Adder_0_U.u1.cin ;
assign _097_ = \add_33s_33s_33_2_1_U3.top_add_33s_33s_33_2_1_Adder_0_U.u2.a  + \add_33s_33s_33_2_1_U3.top_add_33s_33s_33_2_1_Adder_0_U.u2.b ;
assign { \add_33s_33s_33_2_1_U3.top_add_33s_33s_33_2_1_Adder_0_U.u2.cout , \add_33s_33s_33_2_1_U3.top_add_33s_33s_33_2_1_Adder_0_U.u2.s  } = _097_ + \add_33s_33s_33_2_1_U3.top_add_33s_33s_33_2_1_Adder_0_U.u2.cin ;
always @(posedge \add_35s_35s_35_2_1_U11.top_add_35s_35s_35_2_1_Adder_6_U.clk )
\add_35s_35s_35_2_1_U11.top_add_35s_35s_35_2_1_Adder_6_U.bin_s1  <= _099_;
always @(posedge \add_35s_35s_35_2_1_U11.top_add_35s_35s_35_2_1_Adder_6_U.clk )
\add_35s_35s_35_2_1_U11.top_add_35s_35s_35_2_1_Adder_6_U.ain_s1  <= _098_;
always @(posedge \add_35s_35s_35_2_1_U11.top_add_35s_35s_35_2_1_Adder_6_U.clk )
\add_35s_35s_35_2_1_U11.top_add_35s_35s_35_2_1_Adder_6_U.sum_s1  <= _101_;
always @(posedge \add_35s_35s_35_2_1_U11.top_add_35s_35s_35_2_1_Adder_6_U.clk )
\add_35s_35s_35_2_1_U11.top_add_35s_35s_35_2_1_Adder_6_U.carry_s1  <= _100_;
assign _099_ = \add_35s_35s_35_2_1_U11.top_add_35s_35s_35_2_1_Adder_6_U.ce  ? \add_35s_35s_35_2_1_U11.top_add_35s_35s_35_2_1_Adder_6_U.b [34:17] : \add_35s_35s_35_2_1_U11.top_add_35s_35s_35_2_1_Adder_6_U.bin_s1 ;
assign _098_ = \add_35s_35s_35_2_1_U11.top_add_35s_35s_35_2_1_Adder_6_U.ce  ? \add_35s_35s_35_2_1_U11.top_add_35s_35s_35_2_1_Adder_6_U.a [34:17] : \add_35s_35s_35_2_1_U11.top_add_35s_35s_35_2_1_Adder_6_U.ain_s1 ;
assign _100_ = \add_35s_35s_35_2_1_U11.top_add_35s_35s_35_2_1_Adder_6_U.ce  ? \add_35s_35s_35_2_1_U11.top_add_35s_35s_35_2_1_Adder_6_U.facout_s1  : \add_35s_35s_35_2_1_U11.top_add_35s_35s_35_2_1_Adder_6_U.carry_s1 ;
assign _101_ = \add_35s_35s_35_2_1_U11.top_add_35s_35s_35_2_1_Adder_6_U.ce  ? \add_35s_35s_35_2_1_U11.top_add_35s_35s_35_2_1_Adder_6_U.fas_s1  : \add_35s_35s_35_2_1_U11.top_add_35s_35s_35_2_1_Adder_6_U.sum_s1 ;
assign _102_ = \add_35s_35s_35_2_1_U11.top_add_35s_35s_35_2_1_Adder_6_U.u1.a  + \add_35s_35s_35_2_1_U11.top_add_35s_35s_35_2_1_Adder_6_U.u1.b ;
assign { \add_35s_35s_35_2_1_U11.top_add_35s_35s_35_2_1_Adder_6_U.u1.cout , \add_35s_35s_35_2_1_U11.top_add_35s_35s_35_2_1_Adder_6_U.u1.s  } = _102_ + \add_35s_35s_35_2_1_U11.top_add_35s_35s_35_2_1_Adder_6_U.u1.cin ;
assign _103_ = \add_35s_35s_35_2_1_U11.top_add_35s_35s_35_2_1_Adder_6_U.u2.a  + \add_35s_35s_35_2_1_U11.top_add_35s_35s_35_2_1_Adder_6_U.u2.b ;
assign { \add_35s_35s_35_2_1_U11.top_add_35s_35s_35_2_1_Adder_6_U.u2.cout , \add_35s_35s_35_2_1_U11.top_add_35s_35s_35_2_1_Adder_6_U.u2.s  } = _103_ + \add_35s_35s_35_2_1_U11.top_add_35s_35s_35_2_1_Adder_6_U.u2.cin ;
always @(posedge \add_43s_43s_43_2_1_U9.top_add_43s_43s_43_2_1_Adder_4_U.clk )
\add_43s_43s_43_2_1_U9.top_add_43s_43s_43_2_1_Adder_4_U.bin_s1  <= _105_;
always @(posedge \add_43s_43s_43_2_1_U9.top_add_43s_43s_43_2_1_Adder_4_U.clk )
\add_43s_43s_43_2_1_U9.top_add_43s_43s_43_2_1_Adder_4_U.ain_s1  <= _104_;
always @(posedge \add_43s_43s_43_2_1_U9.top_add_43s_43s_43_2_1_Adder_4_U.clk )
\add_43s_43s_43_2_1_U9.top_add_43s_43s_43_2_1_Adder_4_U.sum_s1  <= _107_;
always @(posedge \add_43s_43s_43_2_1_U9.top_add_43s_43s_43_2_1_Adder_4_U.clk )
\add_43s_43s_43_2_1_U9.top_add_43s_43s_43_2_1_Adder_4_U.carry_s1  <= _106_;
assign _105_ = \add_43s_43s_43_2_1_U9.top_add_43s_43s_43_2_1_Adder_4_U.ce  ? \add_43s_43s_43_2_1_U9.top_add_43s_43s_43_2_1_Adder_4_U.b [42:21] : \add_43s_43s_43_2_1_U9.top_add_43s_43s_43_2_1_Adder_4_U.bin_s1 ;
assign _104_ = \add_43s_43s_43_2_1_U9.top_add_43s_43s_43_2_1_Adder_4_U.ce  ? \add_43s_43s_43_2_1_U9.top_add_43s_43s_43_2_1_Adder_4_U.a [42:21] : \add_43s_43s_43_2_1_U9.top_add_43s_43s_43_2_1_Adder_4_U.ain_s1 ;
assign _106_ = \add_43s_43s_43_2_1_U9.top_add_43s_43s_43_2_1_Adder_4_U.ce  ? \add_43s_43s_43_2_1_U9.top_add_43s_43s_43_2_1_Adder_4_U.facout_s1  : \add_43s_43s_43_2_1_U9.top_add_43s_43s_43_2_1_Adder_4_U.carry_s1 ;
assign _107_ = \add_43s_43s_43_2_1_U9.top_add_43s_43s_43_2_1_Adder_4_U.ce  ? \add_43s_43s_43_2_1_U9.top_add_43s_43s_43_2_1_Adder_4_U.fas_s1  : \add_43s_43s_43_2_1_U9.top_add_43s_43s_43_2_1_Adder_4_U.sum_s1 ;
assign _108_ = \add_43s_43s_43_2_1_U9.top_add_43s_43s_43_2_1_Adder_4_U.u1.a  + \add_43s_43s_43_2_1_U9.top_add_43s_43s_43_2_1_Adder_4_U.u1.b ;
assign { \add_43s_43s_43_2_1_U9.top_add_43s_43s_43_2_1_Adder_4_U.u1.cout , \add_43s_43s_43_2_1_U9.top_add_43s_43s_43_2_1_Adder_4_U.u1.s  } = _108_ + \add_43s_43s_43_2_1_U9.top_add_43s_43s_43_2_1_Adder_4_U.u1.cin ;
assign _109_ = \add_43s_43s_43_2_1_U9.top_add_43s_43s_43_2_1_Adder_4_U.u2.a  + \add_43s_43s_43_2_1_U9.top_add_43s_43s_43_2_1_Adder_4_U.u2.b ;
assign { \add_43s_43s_43_2_1_U9.top_add_43s_43s_43_2_1_Adder_4_U.u2.cout , \add_43s_43s_43_2_1_U9.top_add_43s_43s_43_2_1_Adder_4_U.u2.s  } = _109_ + \add_43s_43s_43_2_1_U9.top_add_43s_43s_43_2_1_Adder_4_U.u2.cin ;
assign \mul_4ns_4ns_8_4_1_U1.top_mul_4ns_4ns_8_4_1_Mul_DSP_0_U.tmp_product  = \mul_4ns_4ns_8_4_1_U1.top_mul_4ns_4ns_8_4_1_Mul_DSP_0_U.a_reg0  * \mul_4ns_4ns_8_4_1_U1.top_mul_4ns_4ns_8_4_1_Mul_DSP_0_U.b_reg0 ;
always @(posedge \mul_4ns_4ns_8_4_1_U1.top_mul_4ns_4ns_8_4_1_Mul_DSP_0_U.clk )
\mul_4ns_4ns_8_4_1_U1.top_mul_4ns_4ns_8_4_1_Mul_DSP_0_U.a_reg0  <= _110_;
always @(posedge \mul_4ns_4ns_8_4_1_U1.top_mul_4ns_4ns_8_4_1_Mul_DSP_0_U.clk )
\mul_4ns_4ns_8_4_1_U1.top_mul_4ns_4ns_8_4_1_Mul_DSP_0_U.b_reg0  <= _111_;
always @(posedge \mul_4ns_4ns_8_4_1_U1.top_mul_4ns_4ns_8_4_1_Mul_DSP_0_U.clk )
\mul_4ns_4ns_8_4_1_U1.top_mul_4ns_4ns_8_4_1_Mul_DSP_0_U.buff0  <= _112_;
always @(posedge \mul_4ns_4ns_8_4_1_U1.top_mul_4ns_4ns_8_4_1_Mul_DSP_0_U.clk )
\mul_4ns_4ns_8_4_1_U1.top_mul_4ns_4ns_8_4_1_Mul_DSP_0_U.buff1  <= _113_;
assign _113_ = \mul_4ns_4ns_8_4_1_U1.top_mul_4ns_4ns_8_4_1_Mul_DSP_0_U.ce  ? \mul_4ns_4ns_8_4_1_U1.top_mul_4ns_4ns_8_4_1_Mul_DSP_0_U.buff0  : \mul_4ns_4ns_8_4_1_U1.top_mul_4ns_4ns_8_4_1_Mul_DSP_0_U.buff1 ;
assign _112_ = \mul_4ns_4ns_8_4_1_U1.top_mul_4ns_4ns_8_4_1_Mul_DSP_0_U.ce  ? \mul_4ns_4ns_8_4_1_U1.top_mul_4ns_4ns_8_4_1_Mul_DSP_0_U.tmp_product  : \mul_4ns_4ns_8_4_1_U1.top_mul_4ns_4ns_8_4_1_Mul_DSP_0_U.buff0 ;
assign _111_ = \mul_4ns_4ns_8_4_1_U1.top_mul_4ns_4ns_8_4_1_Mul_DSP_0_U.ce  ? \mul_4ns_4ns_8_4_1_U1.top_mul_4ns_4ns_8_4_1_Mul_DSP_0_U.b  : \mul_4ns_4ns_8_4_1_U1.top_mul_4ns_4ns_8_4_1_Mul_DSP_0_U.b_reg0 ;
assign _110_ = \mul_4ns_4ns_8_4_1_U1.top_mul_4ns_4ns_8_4_1_Mul_DSP_0_U.ce  ? \mul_4ns_4ns_8_4_1_U1.top_mul_4ns_4ns_8_4_1_Mul_DSP_0_U.a  : \mul_4ns_4ns_8_4_1_U1.top_mul_4ns_4ns_8_4_1_Mul_DSP_0_U.a_reg0 ;
always @(posedge \shl_16ns_4ns_16_7_1_U2.clk )
\shl_16ns_4ns_16_7_1_U2.dout_array[5]  <= _125_;
always @(posedge \shl_16ns_4ns_16_7_1_U2.clk )
\shl_16ns_4ns_16_7_1_U2.din1_cast_array[5]  <= _119_;
always @(posedge \shl_16ns_4ns_16_7_1_U2.clk )
\shl_16ns_4ns_16_7_1_U2.dout_array[4]  <= _124_;
always @(posedge \shl_16ns_4ns_16_7_1_U2.clk )
\shl_16ns_4ns_16_7_1_U2.din1_cast_array[4]  <= _118_;
always @(posedge \shl_16ns_4ns_16_7_1_U2.clk )
\shl_16ns_4ns_16_7_1_U2.dout_array[3]  <= _123_;
always @(posedge \shl_16ns_4ns_16_7_1_U2.clk )
\shl_16ns_4ns_16_7_1_U2.din1_cast_array[3]  <= _117_;
always @(posedge \shl_16ns_4ns_16_7_1_U2.clk )
\shl_16ns_4ns_16_7_1_U2.dout_array[2]  <= _122_;
always @(posedge \shl_16ns_4ns_16_7_1_U2.clk )
\shl_16ns_4ns_16_7_1_U2.din1_cast_array[2]  <= _116_;
always @(posedge \shl_16ns_4ns_16_7_1_U2.clk )
\shl_16ns_4ns_16_7_1_U2.dout_array[1]  <= _121_;
always @(posedge \shl_16ns_4ns_16_7_1_U2.clk )
\shl_16ns_4ns_16_7_1_U2.din1_cast_array[1]  <= _115_;
always @(posedge \shl_16ns_4ns_16_7_1_U2.clk )
\shl_16ns_4ns_16_7_1_U2.dout_array[0]  <= _120_;
always @(posedge \shl_16ns_4ns_16_7_1_U2.clk )
\shl_16ns_4ns_16_7_1_U2.din1_cast_array[0]  <= _114_;
assign _126_ = \shl_16ns_4ns_16_7_1_U2.ce  ? \shl_16ns_4ns_16_7_1_U2.din1_cast_array[4]  : \shl_16ns_4ns_16_7_1_U2.din1_cast_array[5] ;
assign _119_ = \shl_16ns_4ns_16_7_1_U2.reset  ? 4'h0 : _126_;
assign _127_ = \shl_16ns_4ns_16_7_1_U2.ce  ? _140_ : \shl_16ns_4ns_16_7_1_U2.dout_array[5] ;
assign _125_ = \shl_16ns_4ns_16_7_1_U2.reset  ? 16'h0000 : _127_;
assign _128_ = \shl_16ns_4ns_16_7_1_U2.ce  ? \shl_16ns_4ns_16_7_1_U2.din1_cast_array[3]  : \shl_16ns_4ns_16_7_1_U2.din1_cast_array[4] ;
assign _118_ = \shl_16ns_4ns_16_7_1_U2.reset  ? 4'h0 : _128_;
assign _129_ = \shl_16ns_4ns_16_7_1_U2.ce  ? _139_ : \shl_16ns_4ns_16_7_1_U2.dout_array[4] ;
assign _124_ = \shl_16ns_4ns_16_7_1_U2.reset  ? 16'h0000 : _129_;
assign _130_ = \shl_16ns_4ns_16_7_1_U2.ce  ? \shl_16ns_4ns_16_7_1_U2.din1_cast_array[2]  : \shl_16ns_4ns_16_7_1_U2.din1_cast_array[3] ;
assign _117_ = \shl_16ns_4ns_16_7_1_U2.reset  ? 4'h0 : _130_;
assign _131_ = \shl_16ns_4ns_16_7_1_U2.ce  ? _138_ : \shl_16ns_4ns_16_7_1_U2.dout_array[3] ;
assign _123_ = \shl_16ns_4ns_16_7_1_U2.reset  ? 16'h0000 : _131_;
assign _132_ = \shl_16ns_4ns_16_7_1_U2.ce  ? \shl_16ns_4ns_16_7_1_U2.din1_cast_array[1]  : \shl_16ns_4ns_16_7_1_U2.din1_cast_array[2] ;
assign _116_ = \shl_16ns_4ns_16_7_1_U2.reset  ? 4'h0 : _132_;
assign _133_ = \shl_16ns_4ns_16_7_1_U2.ce  ? \shl_16ns_4ns_16_7_1_U2.dout_array[1]  : \shl_16ns_4ns_16_7_1_U2.dout_array[2] ;
assign _122_ = \shl_16ns_4ns_16_7_1_U2.reset  ? 16'h0000 : _133_;
assign _134_ = \shl_16ns_4ns_16_7_1_U2.ce  ? \shl_16ns_4ns_16_7_1_U2.din1_cast_array[0]  : \shl_16ns_4ns_16_7_1_U2.din1_cast_array[1] ;
assign _115_ = \shl_16ns_4ns_16_7_1_U2.reset  ? 4'h0 : _134_;
assign _135_ = \shl_16ns_4ns_16_7_1_U2.ce  ? \shl_16ns_4ns_16_7_1_U2.dout_array[0]  : \shl_16ns_4ns_16_7_1_U2.dout_array[1] ;
assign _121_ = \shl_16ns_4ns_16_7_1_U2.reset  ? 16'h0000 : _135_;
assign _136_ = \shl_16ns_4ns_16_7_1_U2.ce  ? \shl_16ns_4ns_16_7_1_U2.din1 [3:0] : \shl_16ns_4ns_16_7_1_U2.din1_cast_array[0] ;
assign _114_ = \shl_16ns_4ns_16_7_1_U2.reset  ? 4'h0 : _136_;
assign _137_ = \shl_16ns_4ns_16_7_1_U2.ce  ? \shl_16ns_4ns_16_7_1_U2.din0  : \shl_16ns_4ns_16_7_1_U2.dout_array[0] ;
assign _120_ = \shl_16ns_4ns_16_7_1_U2.reset  ? 16'h0000 : _137_;
assign _138_ = \shl_16ns_4ns_16_7_1_U2.dout_array[2]  << { \shl_16ns_4ns_16_7_1_U2.din1_cast_array[2] [3], 3'h0 };
assign _139_ = \shl_16ns_4ns_16_7_1_U2.dout_array[3]  << { \shl_16ns_4ns_16_7_1_U2.din1_cast_array[3] [2], 2'h0 };
assign _140_ = \shl_16ns_4ns_16_7_1_U2.dout_array[4]  << { \shl_16ns_4ns_16_7_1_U2.din1_cast_array[4] [1], 1'h0 };
assign \shl_16ns_4ns_16_7_1_U2.dout  = \shl_16ns_4ns_16_7_1_U2.dout_array[5]  << \shl_16ns_4ns_16_7_1_U2.din1_cast_array[5] [0];
assign _141_ = | op_17[9:0];
assign _142_ = | trunc_ln851_2_reg_876;
assign _143_ = | op_12[4:0];
assign _144_ = { op_10[1], op_10[1], op_10[1], op_10[1], op_10[1], op_10[1], op_10[1], op_10[1], op_10[1], op_10[1], op_10[1], op_10[1], op_10[1], op_10[1], op_10[1], op_10[1], op_10[1], op_10[1], op_10[1], op_10[1], op_10[1], op_10[1], op_10[1], op_10[1], op_10[1], op_10[1], op_10[1], op_10[1], op_10[1], op_10[1], op_10 } != op_11;
assign or_ln340_1_fu_521_p2 = or_ln340_fu_516_p2 | and_ln786_fu_512_p2;
assign or_ln340_fu_516_p2 = p_Result_4_reg_829 | overflow_fu_507_p2;
assign or_ln785_1_fu_540_p2 = xor_ln785_1_fu_535_p2 | p_Result_4_reg_829;
assign or_ln785_fu_491_p2 = tmp_5_reg_848 | p_Result_5_reg_841;
always @(posedge ap_clk)
op_18_V_reg_866[1:0] <= 2'h0;
always @(posedge ap_clk)
trunc_ln851_2_reg_876 <= 2'h0;
always @(posedge ap_clk)
shl_ln781_reg_752 <= _033_;
always @(posedge ap_clk)
sext_ln850_reg_730 <= _032_;
always @(posedge ap_clk)
ret_reg_685 <= _026_;
always @(posedge ap_clk)
select_ln546_reg_690 <= _029_;
always @(posedge ap_clk)
ret_V_7_reg_913 <= _024_;
always @(posedge ap_clk)
ret_V_6_reg_896 <= _023_;
always @(posedge ap_clk)
ret_V_8_cast_reg_901 <= _025_;
always @(posedge ap_clk)
ret_V_5_reg_817 <= _022_;
always @(posedge ap_clk)
ret_V_5_cast_reg_822 <= _021_;
always @(posedge ap_clk)
ret_V_4_reg_787 <= _020_;
always @(posedge ap_clk)
ret_V_3_reg_757 <= _019_;
always @(posedge ap_clk)
select_ln69_1_reg_762 <= _030_;
always @(posedge ap_clk)
ret_V_2_reg_742 <= _018_;
always @(posedge ap_clk)
select_ln1192_reg_747 <= _027_;
always @(posedge ap_clk)
ret_V_1_reg_720 <= _017_;
always @(posedge ap_clk)
tmp_reg_725 <= _035_;
always @(posedge ap_clk)
p_Result_4_reg_829 <= _015_;
always @(posedge ap_clk)
trunc_ln731_reg_836 <= _036_;
always @(posedge ap_clk)
p_Result_5_reg_841 <= _016_;
always @(posedge ap_clk)
tmp_5_reg_848 <= _034_;
always @(posedge ap_clk)
or_ln785_reg_855 <= _014_;
always @(posedge ap_clk)
op_6_V_reg_670 <= _013_;
always @(posedge ap_clk)
select_ln69_reg_675 <= _031_;
always @(posedge ap_clk)
op_27_V_reg_797 <= _012_;
always @(posedge ap_clk)
op_22_V_reg_700 <= _010_;
always @(posedge ap_clk)
op_18_V_reg_866[3:2] <= _009_;
always @(posedge ap_clk)
select_ln353_reg_871 <= _028_;
always @(posedge ap_clk)
lhs_V_reg_772 <= _008_;
always @(posedge ap_clk)
op_25_V_reg_777 <= _011_;
always @(posedge ap_clk)
icmp_ln851_reg_715 <= _007_;
always @(posedge ap_clk)
icmp_ln851_2_reg_891 <= _006_;
always @(posedge ap_clk)
icmp_ln851_1_reg_812 <= _005_;
always @(posedge ap_clk)
add_ln69_reg_680 <= _003_;
always @(posedge ap_clk)
add_ln691_reg_737 <= _002_;
always @(posedge ap_clk)
add_ln691_2_reg_908 <= _001_;
always @(posedge ap_clk)
add_ln691_1_reg_861 <= _000_;
always @(posedge ap_clk)
ap_CS_fsm <= _004_;
assign _037_ = _039_ ? 2'h2 : 2'h1;
assign _145_ = ap_CS_fsm == 1'h1;
function [29:0] _420_;
input [29:0] a;
input [899:0] b;
input [29:0] s;
case (s)
30'b000000000000000000000000000001:
_420_ = b[29:0];
30'b000000000000000000000000000010:
_420_ = b[59:30];
30'b000000000000000000000000000100:
_420_ = b[89:60];
30'b000000000000000000000000001000:
_420_ = b[119:90];
30'b000000000000000000000000010000:
_420_ = b[149:120];
30'b000000000000000000000000100000:
_420_ = b[179:150];
30'b000000000000000000000001000000:
_420_ = b[209:180];
30'b000000000000000000000010000000:
_420_ = b[239:210];
30'b000000000000000000000100000000:
_420_ = b[269:240];
30'b000000000000000000001000000000:
_420_ = b[299:270];
30'b000000000000000000010000000000:
_420_ = b[329:300];
30'b000000000000000000100000000000:
_420_ = b[359:330];
30'b000000000000000001000000000000:
_420_ = b[389:360];
30'b000000000000000010000000000000:
_420_ = b[419:390];
30'b000000000000000100000000000000:
_420_ = b[449:420];
30'b000000000000001000000000000000:
_420_ = b[479:450];
30'b000000000000010000000000000000:
_420_ = b[509:480];
30'b000000000000100000000000000000:
_420_ = b[539:510];
30'b000000000001000000000000000000:
_420_ = b[569:540];
30'b000000000010000000000000000000:
_420_ = b[599:570];
30'b000000000100000000000000000000:
_420_ = b[629:600];
30'b000000001000000000000000000000:
_420_ = b[659:630];
30'b000000010000000000000000000000:
_420_ = b[689:660];
30'b000000100000000000000000000000:
_420_ = b[719:690];
30'b000001000000000000000000000000:
_420_ = b[749:720];
30'b000010000000000000000000000000:
_420_ = b[779:750];
30'b000100000000000000000000000000:
_420_ = b[809:780];
30'b001000000000000000000000000000:
_420_ = b[839:810];
30'b010000000000000000000000000000:
_420_ = b[869:840];
30'b100000000000000000000000000000:
_420_ = b[899:870];
30'b000000000000000000000000000000:
_420_ = a;
default:
_420_ = 30'bx;
endcase
endfunction
assign ap_NS_fsm = _420_(30'hxxxxxxxx, { 28'h0000000, _037_, 870'h00000004000000200000010000000800000040000002000000100000008000000400000020000001000000080000004000000200000010000000800000040000002000000100000008000000400000020000001000000080000004000000200000010000000800000000000001 }, { _145_, _174_, _173_, _172_, _171_, _170_, _169_, _168_, _167_, _166_, _165_, _164_, _163_, _162_, _161_, _160_, _159_, _158_, _157_, _156_, _155_, _154_, _153_, _152_, _151_, _150_, _149_, _148_, _147_, _146_ });
assign _146_ = ap_CS_fsm == 30'h20000000;
assign _147_ = ap_CS_fsm == 29'h10000000;
assign _148_ = ap_CS_fsm == 28'h8000000;
assign _149_ = ap_CS_fsm == 27'h4000000;
assign _150_ = ap_CS_fsm == 26'h2000000;
assign _151_ = ap_CS_fsm == 25'h1000000;
assign _152_ = ap_CS_fsm == 24'h800000;
assign _153_ = ap_CS_fsm == 23'h400000;
assign _154_ = ap_CS_fsm == 22'h200000;
assign _155_ = ap_CS_fsm == 21'h100000;
assign _156_ = ap_CS_fsm == 20'h80000;
assign _157_ = ap_CS_fsm == 19'h40000;
assign _158_ = ap_CS_fsm == 18'h20000;
assign _159_ = ap_CS_fsm == 17'h10000;
assign _160_ = ap_CS_fsm == 16'h8000;
assign _161_ = ap_CS_fsm == 15'h4000;
assign _162_ = ap_CS_fsm == 14'h2000;
assign _163_ = ap_CS_fsm == 13'h1000;
assign _164_ = ap_CS_fsm == 12'h800;
assign _165_ = ap_CS_fsm == 11'h400;
assign _166_ = ap_CS_fsm == 10'h200;
assign _167_ = ap_CS_fsm == 9'h100;
assign _168_ = ap_CS_fsm == 8'h80;
assign _169_ = ap_CS_fsm == 7'h40;
assign _170_ = ap_CS_fsm == 6'h20;
assign _171_ = ap_CS_fsm == 5'h10;
assign _172_ = ap_CS_fsm == 4'h8;
assign _173_ = ap_CS_fsm == 3'h4;
assign _174_ = ap_CS_fsm == 2'h2;
assign op_30_ap_vld = ap_CS_fsm[29] ? 1'h1 : 1'h0;
assign ap_idle = _038_ ? 1'h1 : 1'h0;
assign _033_ = ap_CS_fsm[10] ? grp_fu_251_p2 : shl_ln781_reg_752;
assign _032_ = ap_CS_fsm[7] ? { tmp_reg_725[27], tmp_reg_725 } : sext_ln850_reg_730;
assign _029_ = ap_CS_fsm[3] ? select_ln546_fu_237_p3 : select_ln546_reg_690;
assign _026_ = ap_CS_fsm[3] ? grp_fu_189_p2 : ret_reg_685;
assign _024_ = ap_CS_fsm[27] ? ret_V_7_fu_638_p3 : ret_V_7_reg_913;
assign _025_ = ap_CS_fsm[24] ? grp_fu_600_p2[33:2] : ret_V_8_cast_reg_901;
assign _023_ = ap_CS_fsm[24] ? grp_fu_600_p2 : ret_V_6_reg_896;
assign _021_ = ap_CS_fsm[19] ? grp_fu_420_p2[41:10] : ret_V_5_cast_reg_822;
assign _022_ = ap_CS_fsm[19] ? grp_fu_420_p2 : ret_V_5_reg_817;
assign _020_ = ap_CS_fsm[15] ? grp_fu_391_p2 : ret_V_4_reg_787;
assign _030_ = ap_CS_fsm[11] ? select_ln69_1_fu_366_p3 : select_ln69_1_reg_762;
assign _019_ = ap_CS_fsm[11] ? grp_fu_345_p2 : ret_V_3_reg_757;
assign _027_ = ap_CS_fsm[9] ? select_ln1192_fu_337_p3 : select_ln1192_reg_747;
assign _018_ = ap_CS_fsm[9] ? ret_V_2_fu_330_p3 : ret_V_2_reg_742;
assign _035_ = ap_CS_fsm[6] ? grp_fu_283_p2[32:5] : tmp_reg_725;
assign _017_ = ap_CS_fsm[6] ? grp_fu_283_p2 : ret_V_1_reg_720;
assign _034_ = ap_CS_fsm[20] ? ret_1_fu_452_p2[2] : tmp_5_reg_848;
assign _016_ = ap_CS_fsm[20] ? ret_1_fu_452_p2[1] : p_Result_5_reg_841;
assign _036_ = ap_CS_fsm[20] ? ret_1_fu_452_p2[1:0] : trunc_ln731_reg_836;
assign _015_ = ap_CS_fsm[20] ? ret_1_fu_452_p2[2] : p_Result_4_reg_829;
assign _014_ = ap_CS_fsm[21] ? or_ln785_fu_491_p2 : or_ln785_reg_855;
assign _031_ = ap_CS_fsm[0] ? select_ln69_fu_215_p3 : select_ln69_reg_675;
assign _013_ = ap_CS_fsm[0] ? op_6_V_fu_203_p2 : op_6_V_reg_670;
assign _012_ = ap_CS_fsm[17] ? grp_fu_400_p2 : op_27_V_reg_797;
assign _010_ = ap_CS_fsm[4] ? op_22_V_fu_262_p2 : op_22_V_reg_700;
assign _028_ = ap_CS_fsm[22] ? select_ln353_fu_575_p3 : select_ln353_reg_871;
assign _009_ = ap_CS_fsm[22] ? op_18_V_fu_555_p3[3:2] : op_18_V_reg_866[3:2];
assign _011_ = ap_CS_fsm[13] ? grp_fu_374_p2 : op_25_V_reg_777;
assign _008_ = ap_CS_fsm[13] ? lhs_V_fu_382_p2 : lhs_V_reg_772;
assign _007_ = ap_CS_fsm[5] ? icmp_ln851_fu_293_p2 : icmp_ln851_reg_715;
assign _006_ = ap_CS_fsm[23] ? icmp_ln851_2_fu_606_p2 : icmp_ln851_2_reg_891;
assign _005_ = ap_CS_fsm[18] ? icmp_ln851_1_fu_430_p2 : icmp_ln851_1_reg_812;
assign _003_ = ap_CS_fsm[1] ? add_ln69_fu_232_p2 : add_ln69_reg_680;
assign _002_ = _042_ ? grp_fu_312_p2 : add_ln691_reg_737;
assign _001_ = _041_ ? grp_fu_621_p2 : add_ln691_2_reg_908;
assign _000_ = _040_ ? grp_fu_486_p2 : add_ln691_1_reg_861;
assign _004_ = ap_rst ? 30'h00000001 : ap_NS_fsm;
assign op_6_V_fu_203_p2 = $signed(op_2[1:0]) - $signed(op_3);
assign ret_1_fu_452_p2 = $signed(op_3) - $signed(op_10);
assign icmp_ln851_1_fu_430_p2 = _141_ ? 1'h1 : 1'h0;
assign icmp_ln851_2_fu_606_p2 = _142_ ? 1'h1 : 1'h0;
assign icmp_ln851_fu_293_p2 = _143_ ? 1'h1 : 1'h0;
assign lhs_V_fu_382_p2 = _144_ ? 1'h1 : 1'h0;
assign op_18_V_fu_555_p3 = and_ln785_1_fu_550_p2 ? { trunc_ln731_reg_836, 2'h0 } : select_ln340_fu_527_p3;
assign ret_V_2_fu_330_p3 = ret_V_1_reg_720[32] ? select_ln850_fu_325_p3 : sext_ln850_reg_730;
assign ret_V_7_fu_638_p3 = ret_V_6_reg_896[34] ? select_ln850_2_fu_633_p3 : ret_V_8_cast_reg_901;
assign select_ln1192_fu_337_p3 = op_13 ? 29'h1fffffff : 29'h00000000;
assign select_ln340_fu_527_p3 = or_ln340_1_fu_521_p2 ? 4'h0 : { trunc_ln731_reg_836, 2'h0 };
assign select_ln353_fu_575_p3 = ret_V_5_reg_817[42] ? select_ln850_1_fu_570_p3 : ret_V_5_cast_reg_822;
assign select_ln546_fu_237_p3 = op_5 ? 16'hffff : 16'h0000;
assign select_ln69_1_fu_366_p3 = select_ln769_fu_359_p3 ? 29'h1fffffff : 29'h00000000;
assign select_ln69_fu_215_p3 = op_8_V_fu_209_p2 ? 3'h7 : 3'h0;
assign select_ln769_fu_359_p3 = op_3[1] ? op_5 : shl_ln781_reg_752[0];
assign select_ln850_1_fu_570_p3 = icmp_ln851_1_reg_812 ? add_ln691_1_reg_861 : ret_V_5_cast_reg_822;
assign select_ln850_2_fu_633_p3 = icmp_ln851_2_reg_891 ? add_ln691_2_reg_908 : ret_V_8_cast_reg_901;
assign select_ln850_fu_325_p3 = icmp_ln851_reg_715 ? add_ln691_reg_737 : sext_ln850_reg_730;
assign op_8_V_fu_209_p2 = op_2[0] ^ op_5;
assign ap_CS_fsm_state1 = ap_CS_fsm[0];
assign ap_CS_fsm_state10 = ap_CS_fsm[9];
assign ap_CS_fsm_state11 = ap_CS_fsm[10];
assign ap_CS_fsm_state12 = ap_CS_fsm[11];
assign ap_CS_fsm_state13 = ap_CS_fsm[12];
assign ap_CS_fsm_state14 = ap_CS_fsm[13];
assign ap_CS_fsm_state15 = ap_CS_fsm[14];
assign ap_CS_fsm_state16 = ap_CS_fsm[15];
assign ap_CS_fsm_state17 = ap_CS_fsm[16];
assign ap_CS_fsm_state18 = ap_CS_fsm[17];
assign ap_CS_fsm_state19 = ap_CS_fsm[18];
assign ap_CS_fsm_state2 = ap_CS_fsm[1];
assign ap_CS_fsm_state20 = ap_CS_fsm[19];
assign ap_CS_fsm_state21 = ap_CS_fsm[20];
assign ap_CS_fsm_state22 = ap_CS_fsm[21];
assign ap_CS_fsm_state23 = ap_CS_fsm[22];
assign ap_CS_fsm_state24 = ap_CS_fsm[23];
assign ap_CS_fsm_state25 = ap_CS_fsm[24];
assign ap_CS_fsm_state26 = ap_CS_fsm[25];
assign ap_CS_fsm_state27 = ap_CS_fsm[26];
assign ap_CS_fsm_state28 = ap_CS_fsm[27];
assign ap_CS_fsm_state29 = ap_CS_fsm[28];
assign ap_CS_fsm_state30 = ap_CS_fsm[29];
assign ap_CS_fsm_state4 = ap_CS_fsm[3];
assign ap_CS_fsm_state5 = ap_CS_fsm[4];
assign ap_CS_fsm_state6 = ap_CS_fsm[5];
assign ap_CS_fsm_state7 = ap_CS_fsm[6];
assign ap_CS_fsm_state8 = ap_CS_fsm[7];
assign ap_CS_fsm_state9 = ap_CS_fsm[8];
assign ap_done = op_30_ap_vld;
assign ap_ready = op_30_ap_vld;
assign grp_fu_189_p0 = op_2;
assign grp_fu_189_p1 = op_2;
assign grp_fu_251_p1 = { 12'h000, op_3[1], op_3[1], op_3 };
assign grp_fu_283_p0 = { op_22_V_reg_700[8], op_22_V_reg_700[8], op_22_V_reg_700[8], op_22_V_reg_700[8], op_22_V_reg_700[8], op_22_V_reg_700[8], op_22_V_reg_700[8], op_22_V_reg_700[8], op_22_V_reg_700[8], op_22_V_reg_700[8], op_22_V_reg_700[8], op_22_V_reg_700[8], op_22_V_reg_700[8], op_22_V_reg_700[8], op_22_V_reg_700[8], op_22_V_reg_700[8], op_22_V_reg_700[8], op_22_V_reg_700[8], op_22_V_reg_700[8], op_22_V_reg_700, 5'h00 };
assign grp_fu_283_p1 = { op_12[31], op_12 };
assign grp_fu_312_p0 = { tmp_reg_725[27], tmp_reg_725 };
assign grp_fu_391_p1 = { 28'h0000000, lhs_V_reg_772 };
assign grp_fu_400_p1 = { op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16 };
assign grp_fu_420_p0 = { op_27_V_reg_797[28], op_27_V_reg_797[28], op_27_V_reg_797[28], op_27_V_reg_797[28], op_27_V_reg_797, 10'h000 };
assign grp_fu_420_p1 = { op_17[31], op_17[31], op_17[31], op_17[31], op_17[31], op_17[31], op_17[31], op_17[31], op_17[31], op_17[31], op_17[31], op_17 };
assign grp_fu_600_p0 = { select_ln353_reg_871[31], select_ln353_reg_871, 2'h0 };
assign grp_fu_600_p1 = { op_18_V_reg_866[3], op_18_V_reg_866[3], op_18_V_reg_866[3], op_18_V_reg_866[3], op_18_V_reg_866[3], op_18_V_reg_866[3], op_18_V_reg_866[3], op_18_V_reg_866[3], op_18_V_reg_866[3], op_18_V_reg_866[3], op_18_V_reg_866[3], op_18_V_reg_866[3], op_18_V_reg_866[3], op_18_V_reg_866[3], op_18_V_reg_866[3], op_18_V_reg_866[3], op_18_V_reg_866[3], op_18_V_reg_866[3], op_18_V_reg_866[3], op_18_V_reg_866[3], op_18_V_reg_866[3], op_18_V_reg_866[3], op_18_V_reg_866[3], op_18_V_reg_866[3], op_18_V_reg_866[3], op_18_V_reg_866[3], op_18_V_reg_866[3], op_18_V_reg_866[3], op_18_V_reg_866[3], op_18_V_reg_866[3], op_18_V_reg_866[3], op_18_V_reg_866 };
assign op_30 = grp_fu_645_p2;
assign op_6_V_fu_203_p1 = op_3;
assign p_Result_1_fu_563_p3 = ret_V_5_reg_817[42];
assign p_Result_2_fu_626_p3 = ret_V_6_reg_896[34];
assign p_Result_3_fu_349_p1 = op_3;
assign p_Result_3_fu_349_p3 = op_3[1];
assign p_Result_s_fu_318_p3 = ret_V_1_reg_720[32];
assign p_Val2_1_fu_495_p3 = { trunc_ln731_reg_836, 2'h0 };
assign r_fu_356_p1 = shl_ln781_reg_752[0];
assign rhs_2_fu_272_p3 = { op_22_V_reg_700, 5'h00 };
assign rhs_6_fu_589_p3 = { select_ln353_reg_871, 2'h0 };
assign sext_ln1192_fu_268_p0 = op_12;
assign sext_ln1347_1_fu_449_p0 = op_10;
assign sext_ln1347_1_fu_449_p1 = { op_10[1], op_10 };
assign sext_ln1347_fu_446_p0 = op_3;
assign sext_ln1347_fu_446_p1 = { op_3[1], op_3 };
assign sext_ln69_1_fu_259_p1 = { add_ln69_reg_680[2], add_ln69_reg_680[2], add_ln69_reg_680[2], add_ln69_reg_680[2], add_ln69_reg_680[2], add_ln69_reg_680[2], add_ln69_reg_680 };
assign sext_ln69_fu_256_p1 = { ret_reg_685[7], ret_reg_685 };
assign sext_ln703_1_fu_405_p0 = op_17;
assign sext_ln703_fu_223_p1 = { op_6_V_reg_670[1], op_6_V_reg_670 };
assign sext_ln781_fu_244_p0 = op_3;
assign sext_ln781_fu_244_p1 = { op_3[1], op_3[1], op_3 };
assign sext_ln850_fu_309_p1 = { tmp_reg_725[27], tmp_reg_725 };
assign sext_ln874_fu_378_p0 = op_10;
assign sext_ln874_fu_378_p1 = { op_10[1], op_10[1], op_10[1], op_10[1], op_10[1], op_10[1], op_10[1], op_10[1], op_10[1], op_10[1], op_10[1], op_10[1], op_10[1], op_10[1], op_10[1], op_10[1], op_10[1], op_10[1], op_10[1], op_10[1], op_10[1], op_10[1], op_10[1], op_10[1], op_10[1], op_10[1], op_10[1], op_10[1], op_10[1], op_10[1], op_10 };
assign tmp_7_fu_409_p3 = { op_27_V_reg_797, 10'h000 };
assign trunc_ln69_1_fu_199_p1 = op_2[1:0];
assign trunc_ln69_fu_195_p1 = op_2[0];
assign trunc_ln731_fu_466_p1 = ret_1_fu_452_p2[1:0];
assign trunc_ln851_1_fu_426_p0 = op_17;
assign trunc_ln851_1_fu_426_p1 = op_17[9:0];
assign trunc_ln851_2_fu_582_p1 = op_18_V_fu_555_p3[1:0];
assign trunc_ln851_fu_289_p0 = op_12;
assign trunc_ln851_fu_289_p1 = op_12[4:0];
assign zext_ln1345_fu_185_p1 = { 4'h0, op_2 };
assign \shl_16ns_4ns_16_7_1_U2.din1_cast  = \shl_16ns_4ns_16_7_1_U2.din1 [3:0];
assign \shl_16ns_4ns_16_7_1_U2.din1_mask  = 4'h1;
assign \shl_16ns_4ns_16_7_1_U2.ce  = 1'h1;
assign \shl_16ns_4ns_16_7_1_U2.clk  = ap_clk;
assign \shl_16ns_4ns_16_7_1_U2.din0  = select_ln546_reg_690;
assign \shl_16ns_4ns_16_7_1_U2.din1  = { 12'h000, op_3[1], op_3[1], op_3 };
assign grp_fu_251_p2 = \shl_16ns_4ns_16_7_1_U2.dout ;
assign \shl_16ns_4ns_16_7_1_U2.reset  = ap_rst;
assign \mul_4ns_4ns_8_4_1_U1.top_mul_4ns_4ns_8_4_1_Mul_DSP_0_U.p  = \mul_4ns_4ns_8_4_1_U1.top_mul_4ns_4ns_8_4_1_Mul_DSP_0_U.buff1 ;
assign \mul_4ns_4ns_8_4_1_U1.top_mul_4ns_4ns_8_4_1_Mul_DSP_0_U.a  = \mul_4ns_4ns_8_4_1_U1.din0 ;
assign \mul_4ns_4ns_8_4_1_U1.top_mul_4ns_4ns_8_4_1_Mul_DSP_0_U.b  = \mul_4ns_4ns_8_4_1_U1.din1 ;
assign \mul_4ns_4ns_8_4_1_U1.top_mul_4ns_4ns_8_4_1_Mul_DSP_0_U.ce  = \mul_4ns_4ns_8_4_1_U1.ce ;
assign \mul_4ns_4ns_8_4_1_U1.top_mul_4ns_4ns_8_4_1_Mul_DSP_0_U.clk  = \mul_4ns_4ns_8_4_1_U1.clk ;
assign \mul_4ns_4ns_8_4_1_U1.dout  = \mul_4ns_4ns_8_4_1_U1.top_mul_4ns_4ns_8_4_1_Mul_DSP_0_U.p ;
assign \mul_4ns_4ns_8_4_1_U1.ce  = 1'h1;
assign \mul_4ns_4ns_8_4_1_U1.clk  = ap_clk;
assign \mul_4ns_4ns_8_4_1_U1.din0  = op_2;
assign \mul_4ns_4ns_8_4_1_U1.din1  = op_2;
assign grp_fu_189_p2 = \mul_4ns_4ns_8_4_1_U1.dout ;
assign \mul_4ns_4ns_8_4_1_U1.reset  = ap_rst;
assign \add_43s_43s_43_2_1_U9.top_add_43s_43s_43_2_1_Adder_4_U.ain_s0  = \add_43s_43s_43_2_1_U9.top_add_43s_43s_43_2_1_Adder_4_U.a ;
assign \add_43s_43s_43_2_1_U9.top_add_43s_43s_43_2_1_Adder_4_U.bin_s0  = \add_43s_43s_43_2_1_U9.top_add_43s_43s_43_2_1_Adder_4_U.b ;
assign \add_43s_43s_43_2_1_U9.top_add_43s_43s_43_2_1_Adder_4_U.s  = { \add_43s_43s_43_2_1_U9.top_add_43s_43s_43_2_1_Adder_4_U.fas_s2 , \add_43s_43s_43_2_1_U9.top_add_43s_43s_43_2_1_Adder_4_U.sum_s1  };
assign \add_43s_43s_43_2_1_U9.top_add_43s_43s_43_2_1_Adder_4_U.u2.a  = \add_43s_43s_43_2_1_U9.top_add_43s_43s_43_2_1_Adder_4_U.ain_s1 ;
assign \add_43s_43s_43_2_1_U9.top_add_43s_43s_43_2_1_Adder_4_U.u2.b  = \add_43s_43s_43_2_1_U9.top_add_43s_43s_43_2_1_Adder_4_U.bin_s1 ;
assign \add_43s_43s_43_2_1_U9.top_add_43s_43s_43_2_1_Adder_4_U.u2.cin  = \add_43s_43s_43_2_1_U9.top_add_43s_43s_43_2_1_Adder_4_U.carry_s1 ;
assign \add_43s_43s_43_2_1_U9.top_add_43s_43s_43_2_1_Adder_4_U.facout_s2  = \add_43s_43s_43_2_1_U9.top_add_43s_43s_43_2_1_Adder_4_U.u2.cout ;
assign \add_43s_43s_43_2_1_U9.top_add_43s_43s_43_2_1_Adder_4_U.fas_s2  = \add_43s_43s_43_2_1_U9.top_add_43s_43s_43_2_1_Adder_4_U.u2.s ;
assign \add_43s_43s_43_2_1_U9.top_add_43s_43s_43_2_1_Adder_4_U.u1.a  = \add_43s_43s_43_2_1_U9.top_add_43s_43s_43_2_1_Adder_4_U.a [20:0];
assign \add_43s_43s_43_2_1_U9.top_add_43s_43s_43_2_1_Adder_4_U.u1.b  = \add_43s_43s_43_2_1_U9.top_add_43s_43s_43_2_1_Adder_4_U.b [20:0];
assign \add_43s_43s_43_2_1_U9.top_add_43s_43s_43_2_1_Adder_4_U.u1.cin  = 1'h0;
assign \add_43s_43s_43_2_1_U9.top_add_43s_43s_43_2_1_Adder_4_U.facout_s1  = \add_43s_43s_43_2_1_U9.top_add_43s_43s_43_2_1_Adder_4_U.u1.cout ;
assign \add_43s_43s_43_2_1_U9.top_add_43s_43s_43_2_1_Adder_4_U.fas_s1  = \add_43s_43s_43_2_1_U9.top_add_43s_43s_43_2_1_Adder_4_U.u1.s ;
assign \add_43s_43s_43_2_1_U9.top_add_43s_43s_43_2_1_Adder_4_U.a  = \add_43s_43s_43_2_1_U9.din0 ;
assign \add_43s_43s_43_2_1_U9.top_add_43s_43s_43_2_1_Adder_4_U.b  = \add_43s_43s_43_2_1_U9.din1 ;
assign \add_43s_43s_43_2_1_U9.top_add_43s_43s_43_2_1_Adder_4_U.ce  = \add_43s_43s_43_2_1_U9.ce ;
assign \add_43s_43s_43_2_1_U9.top_add_43s_43s_43_2_1_Adder_4_U.clk  = \add_43s_43s_43_2_1_U9.clk ;
assign \add_43s_43s_43_2_1_U9.top_add_43s_43s_43_2_1_Adder_4_U.reset  = \add_43s_43s_43_2_1_U9.reset ;
assign \add_43s_43s_43_2_1_U9.dout  = \add_43s_43s_43_2_1_U9.top_add_43s_43s_43_2_1_Adder_4_U.s ;
assign \add_43s_43s_43_2_1_U9.ce  = 1'h1;
assign \add_43s_43s_43_2_1_U9.clk  = ap_clk;
assign \add_43s_43s_43_2_1_U9.din0  = { op_27_V_reg_797[28], op_27_V_reg_797[28], op_27_V_reg_797[28], op_27_V_reg_797[28], op_27_V_reg_797, 10'h000 };
assign \add_43s_43s_43_2_1_U9.din1  = { op_17[31], op_17[31], op_17[31], op_17[31], op_17[31], op_17[31], op_17[31], op_17[31], op_17[31], op_17[31], op_17[31], op_17 };
assign grp_fu_420_p2 = \add_43s_43s_43_2_1_U9.dout ;
assign \add_43s_43s_43_2_1_U9.reset  = ap_rst;
assign \add_35s_35s_35_2_1_U11.top_add_35s_35s_35_2_1_Adder_6_U.ain_s0  = \add_35s_35s_35_2_1_U11.top_add_35s_35s_35_2_1_Adder_6_U.a ;
assign \add_35s_35s_35_2_1_U11.top_add_35s_35s_35_2_1_Adder_6_U.bin_s0  = \add_35s_35s_35_2_1_U11.top_add_35s_35s_35_2_1_Adder_6_U.b ;
assign \add_35s_35s_35_2_1_U11.top_add_35s_35s_35_2_1_Adder_6_U.s  = { \add_35s_35s_35_2_1_U11.top_add_35s_35s_35_2_1_Adder_6_U.fas_s2 , \add_35s_35s_35_2_1_U11.top_add_35s_35s_35_2_1_Adder_6_U.sum_s1  };
assign \add_35s_35s_35_2_1_U11.top_add_35s_35s_35_2_1_Adder_6_U.u2.a  = \add_35s_35s_35_2_1_U11.top_add_35s_35s_35_2_1_Adder_6_U.ain_s1 ;
assign \add_35s_35s_35_2_1_U11.top_add_35s_35s_35_2_1_Adder_6_U.u2.b  = \add_35s_35s_35_2_1_U11.top_add_35s_35s_35_2_1_Adder_6_U.bin_s1 ;
assign \add_35s_35s_35_2_1_U11.top_add_35s_35s_35_2_1_Adder_6_U.u2.cin  = \add_35s_35s_35_2_1_U11.top_add_35s_35s_35_2_1_Adder_6_U.carry_s1 ;
assign \add_35s_35s_35_2_1_U11.top_add_35s_35s_35_2_1_Adder_6_U.facout_s2  = \add_35s_35s_35_2_1_U11.top_add_35s_35s_35_2_1_Adder_6_U.u2.cout ;
assign \add_35s_35s_35_2_1_U11.top_add_35s_35s_35_2_1_Adder_6_U.fas_s2  = \add_35s_35s_35_2_1_U11.top_add_35s_35s_35_2_1_Adder_6_U.u2.s ;
assign \add_35s_35s_35_2_1_U11.top_add_35s_35s_35_2_1_Adder_6_U.u1.a  = \add_35s_35s_35_2_1_U11.top_add_35s_35s_35_2_1_Adder_6_U.a [16:0];
assign \add_35s_35s_35_2_1_U11.top_add_35s_35s_35_2_1_Adder_6_U.u1.b  = \add_35s_35s_35_2_1_U11.top_add_35s_35s_35_2_1_Adder_6_U.b [16:0];
assign \add_35s_35s_35_2_1_U11.top_add_35s_35s_35_2_1_Adder_6_U.u1.cin  = 1'h0;
assign \add_35s_35s_35_2_1_U11.top_add_35s_35s_35_2_1_Adder_6_U.facout_s1  = \add_35s_35s_35_2_1_U11.top_add_35s_35s_35_2_1_Adder_6_U.u1.cout ;
assign \add_35s_35s_35_2_1_U11.top_add_35s_35s_35_2_1_Adder_6_U.fas_s1  = \add_35s_35s_35_2_1_U11.top_add_35s_35s_35_2_1_Adder_6_U.u1.s ;
assign \add_35s_35s_35_2_1_U11.top_add_35s_35s_35_2_1_Adder_6_U.a  = \add_35s_35s_35_2_1_U11.din0 ;
assign \add_35s_35s_35_2_1_U11.top_add_35s_35s_35_2_1_Adder_6_U.b  = \add_35s_35s_35_2_1_U11.din1 ;
assign \add_35s_35s_35_2_1_U11.top_add_35s_35s_35_2_1_Adder_6_U.ce  = \add_35s_35s_35_2_1_U11.ce ;
assign \add_35s_35s_35_2_1_U11.top_add_35s_35s_35_2_1_Adder_6_U.clk  = \add_35s_35s_35_2_1_U11.clk ;
assign \add_35s_35s_35_2_1_U11.top_add_35s_35s_35_2_1_Adder_6_U.reset  = \add_35s_35s_35_2_1_U11.reset ;
assign \add_35s_35s_35_2_1_U11.dout  = \add_35s_35s_35_2_1_U11.top_add_35s_35s_35_2_1_Adder_6_U.s ;
assign \add_35s_35s_35_2_1_U11.ce  = 1'h1;
assign \add_35s_35s_35_2_1_U11.clk  = ap_clk;
assign \add_35s_35s_35_2_1_U11.din0  = { select_ln353_reg_871[31], select_ln353_reg_871, 2'h0 };
assign \add_35s_35s_35_2_1_U11.din1  = { op_18_V_reg_866[3], op_18_V_reg_866[3], op_18_V_reg_866[3], op_18_V_reg_866[3], op_18_V_reg_866[3], op_18_V_reg_866[3], op_18_V_reg_866[3], op_18_V_reg_866[3], op_18_V_reg_866[3], op_18_V_reg_866[3], op_18_V_reg_866[3], op_18_V_reg_866[3], op_18_V_reg_866[3], op_18_V_reg_866[3], op_18_V_reg_866[3], op_18_V_reg_866[3], op_18_V_reg_866[3], op_18_V_reg_866[3], op_18_V_reg_866[3], op_18_V_reg_866[3], op_18_V_reg_866[3], op_18_V_reg_866[3], op_18_V_reg_866[3], op_18_V_reg_866[3], op_18_V_reg_866[3], op_18_V_reg_866[3], op_18_V_reg_866[3], op_18_V_reg_866[3], op_18_V_reg_866[3], op_18_V_reg_866[3], op_18_V_reg_866[3], op_18_V_reg_866 };
assign grp_fu_600_p2 = \add_35s_35s_35_2_1_U11.dout ;
assign \add_35s_35s_35_2_1_U11.reset  = ap_rst;
assign \add_33s_33s_33_2_1_U3.top_add_33s_33s_33_2_1_Adder_0_U.ain_s0  = \add_33s_33s_33_2_1_U3.top_add_33s_33s_33_2_1_Adder_0_U.a ;
assign \add_33s_33s_33_2_1_U3.top_add_33s_33s_33_2_1_Adder_0_U.bin_s0  = \add_33s_33s_33_2_1_U3.top_add_33s_33s_33_2_1_Adder_0_U.b ;
assign \add_33s_33s_33_2_1_U3.top_add_33s_33s_33_2_1_Adder_0_U.s  = { \add_33s_33s_33_2_1_U3.top_add_33s_33s_33_2_1_Adder_0_U.fas_s2 , \add_33s_33s_33_2_1_U3.top_add_33s_33s_33_2_1_Adder_0_U.sum_s1  };
assign \add_33s_33s_33_2_1_U3.top_add_33s_33s_33_2_1_Adder_0_U.u2.a  = \add_33s_33s_33_2_1_U3.top_add_33s_33s_33_2_1_Adder_0_U.ain_s1 ;
assign \add_33s_33s_33_2_1_U3.top_add_33s_33s_33_2_1_Adder_0_U.u2.b  = \add_33s_33s_33_2_1_U3.top_add_33s_33s_33_2_1_Adder_0_U.bin_s1 ;
assign \add_33s_33s_33_2_1_U3.top_add_33s_33s_33_2_1_Adder_0_U.u2.cin  = \add_33s_33s_33_2_1_U3.top_add_33s_33s_33_2_1_Adder_0_U.carry_s1 ;
assign \add_33s_33s_33_2_1_U3.top_add_33s_33s_33_2_1_Adder_0_U.facout_s2  = \add_33s_33s_33_2_1_U3.top_add_33s_33s_33_2_1_Adder_0_U.u2.cout ;
assign \add_33s_33s_33_2_1_U3.top_add_33s_33s_33_2_1_Adder_0_U.fas_s2  = \add_33s_33s_33_2_1_U3.top_add_33s_33s_33_2_1_Adder_0_U.u2.s ;
assign \add_33s_33s_33_2_1_U3.top_add_33s_33s_33_2_1_Adder_0_U.u1.a  = \add_33s_33s_33_2_1_U3.top_add_33s_33s_33_2_1_Adder_0_U.a [15:0];
assign \add_33s_33s_33_2_1_U3.top_add_33s_33s_33_2_1_Adder_0_U.u1.b  = \add_33s_33s_33_2_1_U3.top_add_33s_33s_33_2_1_Adder_0_U.b [15:0];
assign \add_33s_33s_33_2_1_U3.top_add_33s_33s_33_2_1_Adder_0_U.u1.cin  = 1'h0;
assign \add_33s_33s_33_2_1_U3.top_add_33s_33s_33_2_1_Adder_0_U.facout_s1  = \add_33s_33s_33_2_1_U3.top_add_33s_33s_33_2_1_Adder_0_U.u1.cout ;
assign \add_33s_33s_33_2_1_U3.top_add_33s_33s_33_2_1_Adder_0_U.fas_s1  = \add_33s_33s_33_2_1_U3.top_add_33s_33s_33_2_1_Adder_0_U.u1.s ;
assign \add_33s_33s_33_2_1_U3.top_add_33s_33s_33_2_1_Adder_0_U.a  = \add_33s_33s_33_2_1_U3.din0 ;
assign \add_33s_33s_33_2_1_U3.top_add_33s_33s_33_2_1_Adder_0_U.b  = \add_33s_33s_33_2_1_U3.din1 ;
assign \add_33s_33s_33_2_1_U3.top_add_33s_33s_33_2_1_Adder_0_U.ce  = \add_33s_33s_33_2_1_U3.ce ;
assign \add_33s_33s_33_2_1_U3.top_add_33s_33s_33_2_1_Adder_0_U.clk  = \add_33s_33s_33_2_1_U3.clk ;
assign \add_33s_33s_33_2_1_U3.top_add_33s_33s_33_2_1_Adder_0_U.reset  = \add_33s_33s_33_2_1_U3.reset ;
assign \add_33s_33s_33_2_1_U3.dout  = \add_33s_33s_33_2_1_U3.top_add_33s_33s_33_2_1_Adder_0_U.s ;
assign \add_33s_33s_33_2_1_U3.ce  = 1'h1;
assign \add_33s_33s_33_2_1_U3.clk  = ap_clk;
assign \add_33s_33s_33_2_1_U3.din0  = { op_22_V_reg_700[8], op_22_V_reg_700[8], op_22_V_reg_700[8], op_22_V_reg_700[8], op_22_V_reg_700[8], op_22_V_reg_700[8], op_22_V_reg_700[8], op_22_V_reg_700[8], op_22_V_reg_700[8], op_22_V_reg_700[8], op_22_V_reg_700[8], op_22_V_reg_700[8], op_22_V_reg_700[8], op_22_V_reg_700[8], op_22_V_reg_700[8], op_22_V_reg_700[8], op_22_V_reg_700[8], op_22_V_reg_700[8], op_22_V_reg_700[8], op_22_V_reg_700, 5'h00 };
assign \add_33s_33s_33_2_1_U3.din1  = { op_12[31], op_12 };
assign grp_fu_283_p2 = \add_33s_33s_33_2_1_U3.dout ;
assign \add_33s_33s_33_2_1_U3.reset  = ap_rst;
assign \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_5_U.ain_s0  = \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_5_U.a ;
assign \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_5_U.bin_s0  = \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_5_U.b ;
assign \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_5_U.s  = { \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_5_U.fas_s2 , \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_5_U.sum_s1  };
assign \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.a  = \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_5_U.ain_s1 ;
assign \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.b  = \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_5_U.bin_s1 ;
assign \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.cin  = \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_5_U.carry_s1 ;
assign \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_5_U.facout_s2  = \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.cout ;
assign \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_5_U.fas_s2  = \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.s ;
assign \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.a  = \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_5_U.a [15:0];
assign \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.b  = \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_5_U.b [15:0];
assign \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.cin  = 1'h0;
assign \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_5_U.facout_s1  = \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.cout ;
assign \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_5_U.fas_s1  = \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.s ;
assign \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_5_U.a  = \add_32ns_32ns_32_2_1_U13.din0 ;
assign \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_5_U.b  = \add_32ns_32ns_32_2_1_U13.din1 ;
assign \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_5_U.ce  = \add_32ns_32ns_32_2_1_U13.ce ;
assign \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_5_U.clk  = \add_32ns_32ns_32_2_1_U13.clk ;
assign \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_5_U.reset  = \add_32ns_32ns_32_2_1_U13.reset ;
assign \add_32ns_32ns_32_2_1_U13.dout  = \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_5_U.s ;
assign \add_32ns_32ns_32_2_1_U13.ce  = 1'h1;
assign \add_32ns_32ns_32_2_1_U13.clk  = ap_clk;
assign \add_32ns_32ns_32_2_1_U13.din0  = ret_V_7_reg_913;
assign \add_32ns_32ns_32_2_1_U13.din1  = op_19;
assign grp_fu_645_p2 = \add_32ns_32ns_32_2_1_U13.dout ;
assign \add_32ns_32ns_32_2_1_U13.reset  = ap_rst;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.ain_s0  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.a ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.bin_s0  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.b ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.s  = { \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.fas_s2 , \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.sum_s1  };
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.a  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.ain_s1 ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.b  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.bin_s1 ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.cin  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.carry_s1 ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.facout_s2  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.cout ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.fas_s2  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.s ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.a  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.a [15:0];
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.b  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.b [15:0];
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.cin  = 1'h0;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.facout_s1  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.cout ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.fas_s1  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.s ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.a  = \add_32ns_32ns_32_2_1_U12.din0 ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.b  = \add_32ns_32ns_32_2_1_U12.din1 ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.ce  = \add_32ns_32ns_32_2_1_U12.ce ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.clk  = \add_32ns_32ns_32_2_1_U12.clk ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.reset  = \add_32ns_32ns_32_2_1_U12.reset ;
assign \add_32ns_32ns_32_2_1_U12.dout  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.s ;
assign \add_32ns_32ns_32_2_1_U12.ce  = 1'h1;
assign \add_32ns_32ns_32_2_1_U12.clk  = ap_clk;
assign \add_32ns_32ns_32_2_1_U12.din0  = ret_V_8_cast_reg_901;
assign \add_32ns_32ns_32_2_1_U12.din1  = 32'd1;
assign grp_fu_621_p2 = \add_32ns_32ns_32_2_1_U12.dout ;
assign \add_32ns_32ns_32_2_1_U12.reset  = ap_rst;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_5_U.ain_s0  = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_5_U.a ;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_5_U.bin_s0  = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_5_U.b ;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_5_U.s  = { \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_5_U.fas_s2 , \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_5_U.sum_s1  };
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.a  = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_5_U.ain_s1 ;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.b  = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_5_U.bin_s1 ;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.cin  = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_5_U.carry_s1 ;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_5_U.facout_s2  = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.cout ;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_5_U.fas_s2  = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.s ;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.a  = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_5_U.a [15:0];
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.b  = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_5_U.b [15:0];
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.cin  = 1'h0;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_5_U.facout_s1  = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.cout ;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_5_U.fas_s1  = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.s ;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_5_U.a  = \add_32ns_32ns_32_2_1_U10.din0 ;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_5_U.b  = \add_32ns_32ns_32_2_1_U10.din1 ;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_5_U.ce  = \add_32ns_32ns_32_2_1_U10.ce ;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_5_U.clk  = \add_32ns_32ns_32_2_1_U10.clk ;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_5_U.reset  = \add_32ns_32ns_32_2_1_U10.reset ;
assign \add_32ns_32ns_32_2_1_U10.dout  = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_5_U.s ;
assign \add_32ns_32ns_32_2_1_U10.ce  = 1'h1;
assign \add_32ns_32ns_32_2_1_U10.clk  = ap_clk;
assign \add_32ns_32ns_32_2_1_U10.din0  = ret_V_5_cast_reg_822;
assign \add_32ns_32ns_32_2_1_U10.din1  = 32'd1;
assign grp_fu_486_p2 = \add_32ns_32ns_32_2_1_U10.dout ;
assign \add_32ns_32ns_32_2_1_U10.reset  = ap_rst;
assign \add_29s_29ns_29_2_1_U4.top_add_29s_29ns_29_2_1_Adder_1_U.ain_s0  = \add_29s_29ns_29_2_1_U4.top_add_29s_29ns_29_2_1_Adder_1_U.a ;
assign \add_29s_29ns_29_2_1_U4.top_add_29s_29ns_29_2_1_Adder_1_U.bin_s0  = \add_29s_29ns_29_2_1_U4.top_add_29s_29ns_29_2_1_Adder_1_U.b ;
assign \add_29s_29ns_29_2_1_U4.top_add_29s_29ns_29_2_1_Adder_1_U.s  = { \add_29s_29ns_29_2_1_U4.top_add_29s_29ns_29_2_1_Adder_1_U.fas_s2 , \add_29s_29ns_29_2_1_U4.top_add_29s_29ns_29_2_1_Adder_1_U.sum_s1  };
assign \add_29s_29ns_29_2_1_U4.top_add_29s_29ns_29_2_1_Adder_1_U.u2.a  = \add_29s_29ns_29_2_1_U4.top_add_29s_29ns_29_2_1_Adder_1_U.ain_s1 ;
assign \add_29s_29ns_29_2_1_U4.top_add_29s_29ns_29_2_1_Adder_1_U.u2.b  = \add_29s_29ns_29_2_1_U4.top_add_29s_29ns_29_2_1_Adder_1_U.bin_s1 ;
assign \add_29s_29ns_29_2_1_U4.top_add_29s_29ns_29_2_1_Adder_1_U.u2.cin  = \add_29s_29ns_29_2_1_U4.top_add_29s_29ns_29_2_1_Adder_1_U.carry_s1 ;
assign \add_29s_29ns_29_2_1_U4.top_add_29s_29ns_29_2_1_Adder_1_U.facout_s2  = \add_29s_29ns_29_2_1_U4.top_add_29s_29ns_29_2_1_Adder_1_U.u2.cout ;
assign \add_29s_29ns_29_2_1_U4.top_add_29s_29ns_29_2_1_Adder_1_U.fas_s2  = \add_29s_29ns_29_2_1_U4.top_add_29s_29ns_29_2_1_Adder_1_U.u2.s ;
assign \add_29s_29ns_29_2_1_U4.top_add_29s_29ns_29_2_1_Adder_1_U.u1.a  = \add_29s_29ns_29_2_1_U4.top_add_29s_29ns_29_2_1_Adder_1_U.a [13:0];
assign \add_29s_29ns_29_2_1_U4.top_add_29s_29ns_29_2_1_Adder_1_U.u1.b  = \add_29s_29ns_29_2_1_U4.top_add_29s_29ns_29_2_1_Adder_1_U.b [13:0];
assign \add_29s_29ns_29_2_1_U4.top_add_29s_29ns_29_2_1_Adder_1_U.u1.cin  = 1'h0;
assign \add_29s_29ns_29_2_1_U4.top_add_29s_29ns_29_2_1_Adder_1_U.facout_s1  = \add_29s_29ns_29_2_1_U4.top_add_29s_29ns_29_2_1_Adder_1_U.u1.cout ;
assign \add_29s_29ns_29_2_1_U4.top_add_29s_29ns_29_2_1_Adder_1_U.fas_s1  = \add_29s_29ns_29_2_1_U4.top_add_29s_29ns_29_2_1_Adder_1_U.u1.s ;
assign \add_29s_29ns_29_2_1_U4.top_add_29s_29ns_29_2_1_Adder_1_U.a  = \add_29s_29ns_29_2_1_U4.din0 ;
assign \add_29s_29ns_29_2_1_U4.top_add_29s_29ns_29_2_1_Adder_1_U.b  = \add_29s_29ns_29_2_1_U4.din1 ;
assign \add_29s_29ns_29_2_1_U4.top_add_29s_29ns_29_2_1_Adder_1_U.ce  = \add_29s_29ns_29_2_1_U4.ce ;
assign \add_29s_29ns_29_2_1_U4.top_add_29s_29ns_29_2_1_Adder_1_U.clk  = \add_29s_29ns_29_2_1_U4.clk ;
assign \add_29s_29ns_29_2_1_U4.top_add_29s_29ns_29_2_1_Adder_1_U.reset  = \add_29s_29ns_29_2_1_U4.reset ;
assign \add_29s_29ns_29_2_1_U4.dout  = \add_29s_29ns_29_2_1_U4.top_add_29s_29ns_29_2_1_Adder_1_U.s ;
assign \add_29s_29ns_29_2_1_U4.ce  = 1'h1;
assign \add_29s_29ns_29_2_1_U4.clk  = ap_clk;
assign \add_29s_29ns_29_2_1_U4.din0  = { tmp_reg_725[27], tmp_reg_725 };
assign \add_29s_29ns_29_2_1_U4.din1  = 29'h00000001;
assign grp_fu_312_p2 = \add_29s_29ns_29_2_1_U4.dout ;
assign \add_29s_29ns_29_2_1_U4.reset  = ap_rst;
assign \add_29ns_29s_29_2_1_U8.top_add_29ns_29s_29_2_1_Adder_3_U.ain_s0  = \add_29ns_29s_29_2_1_U8.top_add_29ns_29s_29_2_1_Adder_3_U.a ;
assign \add_29ns_29s_29_2_1_U8.top_add_29ns_29s_29_2_1_Adder_3_U.bin_s0  = \add_29ns_29s_29_2_1_U8.top_add_29ns_29s_29_2_1_Adder_3_U.b ;
assign \add_29ns_29s_29_2_1_U8.top_add_29ns_29s_29_2_1_Adder_3_U.s  = { \add_29ns_29s_29_2_1_U8.top_add_29ns_29s_29_2_1_Adder_3_U.fas_s2 , \add_29ns_29s_29_2_1_U8.top_add_29ns_29s_29_2_1_Adder_3_U.sum_s1  };
assign \add_29ns_29s_29_2_1_U8.top_add_29ns_29s_29_2_1_Adder_3_U.u2.a  = \add_29ns_29s_29_2_1_U8.top_add_29ns_29s_29_2_1_Adder_3_U.ain_s1 ;
assign \add_29ns_29s_29_2_1_U8.top_add_29ns_29s_29_2_1_Adder_3_U.u2.b  = \add_29ns_29s_29_2_1_U8.top_add_29ns_29s_29_2_1_Adder_3_U.bin_s1 ;
assign \add_29ns_29s_29_2_1_U8.top_add_29ns_29s_29_2_1_Adder_3_U.u2.cin  = \add_29ns_29s_29_2_1_U8.top_add_29ns_29s_29_2_1_Adder_3_U.carry_s1 ;
assign \add_29ns_29s_29_2_1_U8.top_add_29ns_29s_29_2_1_Adder_3_U.facout_s2  = \add_29ns_29s_29_2_1_U8.top_add_29ns_29s_29_2_1_Adder_3_U.u2.cout ;
assign \add_29ns_29s_29_2_1_U8.top_add_29ns_29s_29_2_1_Adder_3_U.fas_s2  = \add_29ns_29s_29_2_1_U8.top_add_29ns_29s_29_2_1_Adder_3_U.u2.s ;
assign \add_29ns_29s_29_2_1_U8.top_add_29ns_29s_29_2_1_Adder_3_U.u1.a  = \add_29ns_29s_29_2_1_U8.top_add_29ns_29s_29_2_1_Adder_3_U.a [13:0];
assign \add_29ns_29s_29_2_1_U8.top_add_29ns_29s_29_2_1_Adder_3_U.u1.b  = \add_29ns_29s_29_2_1_U8.top_add_29ns_29s_29_2_1_Adder_3_U.b [13:0];
assign \add_29ns_29s_29_2_1_U8.top_add_29ns_29s_29_2_1_Adder_3_U.u1.cin  = 1'h0;
assign \add_29ns_29s_29_2_1_U8.top_add_29ns_29s_29_2_1_Adder_3_U.facout_s1  = \add_29ns_29s_29_2_1_U8.top_add_29ns_29s_29_2_1_Adder_3_U.u1.cout ;
assign \add_29ns_29s_29_2_1_U8.top_add_29ns_29s_29_2_1_Adder_3_U.fas_s1  = \add_29ns_29s_29_2_1_U8.top_add_29ns_29s_29_2_1_Adder_3_U.u1.s ;
assign \add_29ns_29s_29_2_1_U8.top_add_29ns_29s_29_2_1_Adder_3_U.a  = \add_29ns_29s_29_2_1_U8.din0 ;
assign \add_29ns_29s_29_2_1_U8.top_add_29ns_29s_29_2_1_Adder_3_U.b  = \add_29ns_29s_29_2_1_U8.din1 ;
assign \add_29ns_29s_29_2_1_U8.top_add_29ns_29s_29_2_1_Adder_3_U.ce  = \add_29ns_29s_29_2_1_U8.ce ;
assign \add_29ns_29s_29_2_1_U8.top_add_29ns_29s_29_2_1_Adder_3_U.clk  = \add_29ns_29s_29_2_1_U8.clk ;
assign \add_29ns_29s_29_2_1_U8.top_add_29ns_29s_29_2_1_Adder_3_U.reset  = \add_29ns_29s_29_2_1_U8.reset ;
assign \add_29ns_29s_29_2_1_U8.dout  = \add_29ns_29s_29_2_1_U8.top_add_29ns_29s_29_2_1_Adder_3_U.s ;
assign \add_29ns_29s_29_2_1_U8.ce  = 1'h1;
assign \add_29ns_29s_29_2_1_U8.clk  = ap_clk;
assign \add_29ns_29s_29_2_1_U8.din0  = ret_V_4_reg_787;
assign \add_29ns_29s_29_2_1_U8.din1  = { op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16 };
assign grp_fu_400_p2 = \add_29ns_29s_29_2_1_U8.dout ;
assign \add_29ns_29s_29_2_1_U8.reset  = ap_rst;
assign \add_29ns_29ns_29_2_1_U7.top_add_29ns_29ns_29_2_1_Adder_2_U.ain_s0  = \add_29ns_29ns_29_2_1_U7.top_add_29ns_29ns_29_2_1_Adder_2_U.a ;
assign \add_29ns_29ns_29_2_1_U7.top_add_29ns_29ns_29_2_1_Adder_2_U.bin_s0  = \add_29ns_29ns_29_2_1_U7.top_add_29ns_29ns_29_2_1_Adder_2_U.b ;
assign \add_29ns_29ns_29_2_1_U7.top_add_29ns_29ns_29_2_1_Adder_2_U.s  = { \add_29ns_29ns_29_2_1_U7.top_add_29ns_29ns_29_2_1_Adder_2_U.fas_s2 , \add_29ns_29ns_29_2_1_U7.top_add_29ns_29ns_29_2_1_Adder_2_U.sum_s1  };
assign \add_29ns_29ns_29_2_1_U7.top_add_29ns_29ns_29_2_1_Adder_2_U.u2.a  = \add_29ns_29ns_29_2_1_U7.top_add_29ns_29ns_29_2_1_Adder_2_U.ain_s1 ;
assign \add_29ns_29ns_29_2_1_U7.top_add_29ns_29ns_29_2_1_Adder_2_U.u2.b  = \add_29ns_29ns_29_2_1_U7.top_add_29ns_29ns_29_2_1_Adder_2_U.bin_s1 ;
assign \add_29ns_29ns_29_2_1_U7.top_add_29ns_29ns_29_2_1_Adder_2_U.u2.cin  = \add_29ns_29ns_29_2_1_U7.top_add_29ns_29ns_29_2_1_Adder_2_U.carry_s1 ;
assign \add_29ns_29ns_29_2_1_U7.top_add_29ns_29ns_29_2_1_Adder_2_U.facout_s2  = \add_29ns_29ns_29_2_1_U7.top_add_29ns_29ns_29_2_1_Adder_2_U.u2.cout ;
assign \add_29ns_29ns_29_2_1_U7.top_add_29ns_29ns_29_2_1_Adder_2_U.fas_s2  = \add_29ns_29ns_29_2_1_U7.top_add_29ns_29ns_29_2_1_Adder_2_U.u2.s ;
assign \add_29ns_29ns_29_2_1_U7.top_add_29ns_29ns_29_2_1_Adder_2_U.u1.a  = \add_29ns_29ns_29_2_1_U7.top_add_29ns_29ns_29_2_1_Adder_2_U.a [13:0];
assign \add_29ns_29ns_29_2_1_U7.top_add_29ns_29ns_29_2_1_Adder_2_U.u1.b  = \add_29ns_29ns_29_2_1_U7.top_add_29ns_29ns_29_2_1_Adder_2_U.b [13:0];
assign \add_29ns_29ns_29_2_1_U7.top_add_29ns_29ns_29_2_1_Adder_2_U.u1.cin  = 1'h0;
assign \add_29ns_29ns_29_2_1_U7.top_add_29ns_29ns_29_2_1_Adder_2_U.facout_s1  = \add_29ns_29ns_29_2_1_U7.top_add_29ns_29ns_29_2_1_Adder_2_U.u1.cout ;
assign \add_29ns_29ns_29_2_1_U7.top_add_29ns_29ns_29_2_1_Adder_2_U.fas_s1  = \add_29ns_29ns_29_2_1_U7.top_add_29ns_29ns_29_2_1_Adder_2_U.u1.s ;
assign \add_29ns_29ns_29_2_1_U7.top_add_29ns_29ns_29_2_1_Adder_2_U.a  = \add_29ns_29ns_29_2_1_U7.din0 ;
assign \add_29ns_29ns_29_2_1_U7.top_add_29ns_29ns_29_2_1_Adder_2_U.b  = \add_29ns_29ns_29_2_1_U7.din1 ;
assign \add_29ns_29ns_29_2_1_U7.top_add_29ns_29ns_29_2_1_Adder_2_U.ce  = \add_29ns_29ns_29_2_1_U7.ce ;
assign \add_29ns_29ns_29_2_1_U7.top_add_29ns_29ns_29_2_1_Adder_2_U.clk  = \add_29ns_29ns_29_2_1_U7.clk ;
assign \add_29ns_29ns_29_2_1_U7.top_add_29ns_29ns_29_2_1_Adder_2_U.reset  = \add_29ns_29ns_29_2_1_U7.reset ;
assign \add_29ns_29ns_29_2_1_U7.dout  = \add_29ns_29ns_29_2_1_U7.top_add_29ns_29ns_29_2_1_Adder_2_U.s ;
assign \add_29ns_29ns_29_2_1_U7.ce  = 1'h1;
assign \add_29ns_29ns_29_2_1_U7.clk  = ap_clk;
assign \add_29ns_29ns_29_2_1_U7.din0  = op_25_V_reg_777;
assign \add_29ns_29ns_29_2_1_U7.din1  = { 28'h0000000, lhs_V_reg_772 };
assign grp_fu_391_p2 = \add_29ns_29ns_29_2_1_U7.dout ;
assign \add_29ns_29ns_29_2_1_U7.reset  = ap_rst;
assign \add_29ns_29ns_29_2_1_U6.top_add_29ns_29ns_29_2_1_Adder_2_U.ain_s0  = \add_29ns_29ns_29_2_1_U6.top_add_29ns_29ns_29_2_1_Adder_2_U.a ;
assign \add_29ns_29ns_29_2_1_U6.top_add_29ns_29ns_29_2_1_Adder_2_U.bin_s0  = \add_29ns_29ns_29_2_1_U6.top_add_29ns_29ns_29_2_1_Adder_2_U.b ;
assign \add_29ns_29ns_29_2_1_U6.top_add_29ns_29ns_29_2_1_Adder_2_U.s  = { \add_29ns_29ns_29_2_1_U6.top_add_29ns_29ns_29_2_1_Adder_2_U.fas_s2 , \add_29ns_29ns_29_2_1_U6.top_add_29ns_29ns_29_2_1_Adder_2_U.sum_s1  };
assign \add_29ns_29ns_29_2_1_U6.top_add_29ns_29ns_29_2_1_Adder_2_U.u2.a  = \add_29ns_29ns_29_2_1_U6.top_add_29ns_29ns_29_2_1_Adder_2_U.ain_s1 ;
assign \add_29ns_29ns_29_2_1_U6.top_add_29ns_29ns_29_2_1_Adder_2_U.u2.b  = \add_29ns_29ns_29_2_1_U6.top_add_29ns_29ns_29_2_1_Adder_2_U.bin_s1 ;
assign \add_29ns_29ns_29_2_1_U6.top_add_29ns_29ns_29_2_1_Adder_2_U.u2.cin  = \add_29ns_29ns_29_2_1_U6.top_add_29ns_29ns_29_2_1_Adder_2_U.carry_s1 ;
assign \add_29ns_29ns_29_2_1_U6.top_add_29ns_29ns_29_2_1_Adder_2_U.facout_s2  = \add_29ns_29ns_29_2_1_U6.top_add_29ns_29ns_29_2_1_Adder_2_U.u2.cout ;
assign \add_29ns_29ns_29_2_1_U6.top_add_29ns_29ns_29_2_1_Adder_2_U.fas_s2  = \add_29ns_29ns_29_2_1_U6.top_add_29ns_29ns_29_2_1_Adder_2_U.u2.s ;
assign \add_29ns_29ns_29_2_1_U6.top_add_29ns_29ns_29_2_1_Adder_2_U.u1.a  = \add_29ns_29ns_29_2_1_U6.top_add_29ns_29ns_29_2_1_Adder_2_U.a [13:0];
assign \add_29ns_29ns_29_2_1_U6.top_add_29ns_29ns_29_2_1_Adder_2_U.u1.b  = \add_29ns_29ns_29_2_1_U6.top_add_29ns_29ns_29_2_1_Adder_2_U.b [13:0];
assign \add_29ns_29ns_29_2_1_U6.top_add_29ns_29ns_29_2_1_Adder_2_U.u1.cin  = 1'h0;
assign \add_29ns_29ns_29_2_1_U6.top_add_29ns_29ns_29_2_1_Adder_2_U.facout_s1  = \add_29ns_29ns_29_2_1_U6.top_add_29ns_29ns_29_2_1_Adder_2_U.u1.cout ;
assign \add_29ns_29ns_29_2_1_U6.top_add_29ns_29ns_29_2_1_Adder_2_U.fas_s1  = \add_29ns_29ns_29_2_1_U6.top_add_29ns_29ns_29_2_1_Adder_2_U.u1.s ;
assign \add_29ns_29ns_29_2_1_U6.top_add_29ns_29ns_29_2_1_Adder_2_U.a  = \add_29ns_29ns_29_2_1_U6.din0 ;
assign \add_29ns_29ns_29_2_1_U6.top_add_29ns_29ns_29_2_1_Adder_2_U.b  = \add_29ns_29ns_29_2_1_U6.din1 ;
assign \add_29ns_29ns_29_2_1_U6.top_add_29ns_29ns_29_2_1_Adder_2_U.ce  = \add_29ns_29ns_29_2_1_U6.ce ;
assign \add_29ns_29ns_29_2_1_U6.top_add_29ns_29ns_29_2_1_Adder_2_U.clk  = \add_29ns_29ns_29_2_1_U6.clk ;
assign \add_29ns_29ns_29_2_1_U6.top_add_29ns_29ns_29_2_1_Adder_2_U.reset  = \add_29ns_29ns_29_2_1_U6.reset ;
assign \add_29ns_29ns_29_2_1_U6.dout  = \add_29ns_29ns_29_2_1_U6.top_add_29ns_29ns_29_2_1_Adder_2_U.s ;
assign \add_29ns_29ns_29_2_1_U6.ce  = 1'h1;
assign \add_29ns_29ns_29_2_1_U6.clk  = ap_clk;
assign \add_29ns_29ns_29_2_1_U6.din0  = ret_V_3_reg_757;
assign \add_29ns_29ns_29_2_1_U6.din1  = select_ln69_1_reg_762;
assign grp_fu_374_p2 = \add_29ns_29ns_29_2_1_U6.dout ;
assign \add_29ns_29ns_29_2_1_U6.reset  = ap_rst;
assign \add_29ns_29ns_29_2_1_U5.top_add_29ns_29ns_29_2_1_Adder_2_U.ain_s0  = \add_29ns_29ns_29_2_1_U5.top_add_29ns_29ns_29_2_1_Adder_2_U.a ;
assign \add_29ns_29ns_29_2_1_U5.top_add_29ns_29ns_29_2_1_Adder_2_U.bin_s0  = \add_29ns_29ns_29_2_1_U5.top_add_29ns_29ns_29_2_1_Adder_2_U.b ;
assign \add_29ns_29ns_29_2_1_U5.top_add_29ns_29ns_29_2_1_Adder_2_U.s  = { \add_29ns_29ns_29_2_1_U5.top_add_29ns_29ns_29_2_1_Adder_2_U.fas_s2 , \add_29ns_29ns_29_2_1_U5.top_add_29ns_29ns_29_2_1_Adder_2_U.sum_s1  };
assign \add_29ns_29ns_29_2_1_U5.top_add_29ns_29ns_29_2_1_Adder_2_U.u2.a  = \add_29ns_29ns_29_2_1_U5.top_add_29ns_29ns_29_2_1_Adder_2_U.ain_s1 ;
assign \add_29ns_29ns_29_2_1_U5.top_add_29ns_29ns_29_2_1_Adder_2_U.u2.b  = \add_29ns_29ns_29_2_1_U5.top_add_29ns_29ns_29_2_1_Adder_2_U.bin_s1 ;
assign \add_29ns_29ns_29_2_1_U5.top_add_29ns_29ns_29_2_1_Adder_2_U.u2.cin  = \add_29ns_29ns_29_2_1_U5.top_add_29ns_29ns_29_2_1_Adder_2_U.carry_s1 ;
assign \add_29ns_29ns_29_2_1_U5.top_add_29ns_29ns_29_2_1_Adder_2_U.facout_s2  = \add_29ns_29ns_29_2_1_U5.top_add_29ns_29ns_29_2_1_Adder_2_U.u2.cout ;
assign \add_29ns_29ns_29_2_1_U5.top_add_29ns_29ns_29_2_1_Adder_2_U.fas_s2  = \add_29ns_29ns_29_2_1_U5.top_add_29ns_29ns_29_2_1_Adder_2_U.u2.s ;
assign \add_29ns_29ns_29_2_1_U5.top_add_29ns_29ns_29_2_1_Adder_2_U.u1.a  = \add_29ns_29ns_29_2_1_U5.top_add_29ns_29ns_29_2_1_Adder_2_U.a [13:0];
assign \add_29ns_29ns_29_2_1_U5.top_add_29ns_29ns_29_2_1_Adder_2_U.u1.b  = \add_29ns_29ns_29_2_1_U5.top_add_29ns_29ns_29_2_1_Adder_2_U.b [13:0];
assign \add_29ns_29ns_29_2_1_U5.top_add_29ns_29ns_29_2_1_Adder_2_U.u1.cin  = 1'h0;
assign \add_29ns_29ns_29_2_1_U5.top_add_29ns_29ns_29_2_1_Adder_2_U.facout_s1  = \add_29ns_29ns_29_2_1_U5.top_add_29ns_29ns_29_2_1_Adder_2_U.u1.cout ;
assign \add_29ns_29ns_29_2_1_U5.top_add_29ns_29ns_29_2_1_Adder_2_U.fas_s1  = \add_29ns_29ns_29_2_1_U5.top_add_29ns_29ns_29_2_1_Adder_2_U.u1.s ;
assign \add_29ns_29ns_29_2_1_U5.top_add_29ns_29ns_29_2_1_Adder_2_U.a  = \add_29ns_29ns_29_2_1_U5.din0 ;
assign \add_29ns_29ns_29_2_1_U5.top_add_29ns_29ns_29_2_1_Adder_2_U.b  = \add_29ns_29ns_29_2_1_U5.din1 ;
assign \add_29ns_29ns_29_2_1_U5.top_add_29ns_29ns_29_2_1_Adder_2_U.ce  = \add_29ns_29ns_29_2_1_U5.ce ;
assign \add_29ns_29ns_29_2_1_U5.top_add_29ns_29ns_29_2_1_Adder_2_U.clk  = \add_29ns_29ns_29_2_1_U5.clk ;
assign \add_29ns_29ns_29_2_1_U5.top_add_29ns_29ns_29_2_1_Adder_2_U.reset  = \add_29ns_29ns_29_2_1_U5.reset ;
assign \add_29ns_29ns_29_2_1_U5.dout  = \add_29ns_29ns_29_2_1_U5.top_add_29ns_29ns_29_2_1_Adder_2_U.s ;
assign \add_29ns_29ns_29_2_1_U5.ce  = 1'h1;
assign \add_29ns_29ns_29_2_1_U5.clk  = ap_clk;
assign \add_29ns_29ns_29_2_1_U5.din0  = ret_V_2_reg_742;
assign \add_29ns_29ns_29_2_1_U5.din1  = select_ln1192_reg_747;
assign grp_fu_345_p2 = \add_29ns_29ns_29_2_1_U5.dout ;
assign \add_29ns_29ns_29_2_1_U5.reset  = ap_rst;
endmodule


// Machine B:
// Processed by function `add_clk_enable_signal` in `verilog_tricks.py`.
// Processed by function `remove_reset_signal` in `verilog_tricks.py`.
module top_B (
  ap_clk,
  ap_start,
  ap_done,
  ap_idle,
  ap_ready,
  op_0,
  op_2,
  op_3,
  op_5,
  op_10,
  op_11,
  op_12,
  op_13,
  op_16,
  op_17,
  op_19,
  op_30,
  op_30_ap_vld,
clk_enable
);
input clk_enable;


input ap_clk;
wire ap_rst;
assign ap_rst = op_30_ap_vld;
input ap_start;
input [31:0] op_0;
input [1:0] op_10;
input [31:0] op_11;
input [31:0] op_12;
input op_13;
input [7:0] op_16;
input [31:0] op_17;
input [31:0] op_19;
input [3:0] op_2;
input [1:0] op_3;
input op_5;
output ap_done;
output ap_idle;
output ap_ready;
output [31:0] op_30;
output op_30_ap_vld;


reg [31:0] add_ln691_1_reg_787;
reg [31:0] add_ln691_2_reg_809;
reg [2:0] add_ln69_reg_679;
reg [10:0] ap_CS_fsm = 11'h001;
reg icmp_ln851_1_reg_777;
reg icmp_ln851_2_reg_792;
reg icmp_ln851_reg_704;
reg lhs_V_reg_724;
reg [3:0] op_18_V_reg_782;
reg [8:0] op_22_V_reg_689;
reg [28:0] op_25_V_reg_729;
reg [28:0] op_27_V_reg_734;
reg p_Result_4_reg_739;
reg p_Result_5_reg_751;
reg [32:0] ret_V_1_reg_694;
reg [28:0] ret_V_2_reg_709;
reg [31:0] ret_V_5_cast_reg_770;
reg [42:0] ret_V_5_reg_765;
reg [31:0] ret_V_8_cast_reg_802;
reg [28:0] select_ln1192_reg_714;
reg [28:0] select_ln69_1_reg_684;
reg tmp_5_reg_758;
reg [27:0] tmp_reg_699;
reg [1:0] trunc_ln731_reg_746;
reg [32:0] _081_;
wire [31:0] _000_;
wire [31:0] _001_;
wire [2:0] _002_;
wire [10:0] _003_;
wire _004_;
wire _005_;
wire _006_;
wire _007_;
wire [1:0] _008_;
wire [8:0] _009_;
wire [28:0] _010_;
wire [28:0] _011_;
wire _012_;
wire _013_;
wire [32:0] _014_;
wire [28:0] _015_;
wire [31:0] _016_;
wire [42:0] _017_;
wire [32:0] _018_;
wire [31:0] _019_;
wire [28:0] _020_;
wire [28:0] _021_;
wire _022_;
wire [27:0] _023_;
wire [1:0] _024_;
wire [1:0] _025_;
wire _026_;
wire _027_;
wire _028_;
wire _029_;
wire _030_;
wire _031_;
wire _032_;
wire _033_;
wire _034_;
wire _035_;
wire _036_;
wire _037_;
wire _038_;
wire _039_;
wire _040_;
wire _041_;
wire _042_;
wire _043_;
wire _044_;
wire _045_;
wire [31:0] add_ln691_1_fu_573_p2;
wire [31:0] add_ln691_2_fu_638_p2;
wire [28:0] add_ln691_fu_352_p2;
wire [2:0] add_ln69_fu_265_p2;
wire and_ln785_1_fu_560_p2;
wire and_ln785_fu_555_p2;
wire and_ln786_fu_521_p2;
wire ap_CS_fsm_state1;
wire ap_CS_fsm_state10;
wire ap_CS_fsm_state11;
wire ap_CS_fsm_state2;
wire ap_CS_fsm_state3;
wire ap_CS_fsm_state4;
wire ap_CS_fsm_state5;
wire ap_CS_fsm_state6;
wire ap_CS_fsm_state7;
wire ap_CS_fsm_state8;
wire ap_CS_fsm_state9;
wire [10:0] ap_NS_fsm;
wire ap_clk;
wire ap_done;
wire ap_idle;
wire ap_ready;
wire ap_rst;
wire ap_start;
wire icmp_ln851_1_fu_493_p2;
wire icmp_ln851_2_fu_582_p2;
wire icmp_ln851_fu_336_p2;
wire lhs_V_fu_385_p2;
wire [3:0] \mul_4ns_4ns_8_1_1_U1.din0 ;
wire [3:0] \mul_4ns_4ns_8_1_1_U1.din1 ;
wire [7:0] \mul_4ns_4ns_8_1_1_U1.dout ;
wire [3:0] \mul_4ns_4ns_8_1_1_U1.top_mul_4ns_4ns_8_1_1_Multiplier_0_U.a ;
wire [3:0] \mul_4ns_4ns_8_1_1_U1.top_mul_4ns_4ns_8_1_1_Multiplier_0_U.b ;
wire [7:0] \mul_4ns_4ns_8_1_1_U1.top_mul_4ns_4ns_8_1_1_Multiplier_0_U.p ;
wire [31:0] op_0;
wire [1:0] op_10;
wire [31:0] op_11;
wire [31:0] op_12;
wire op_13;
wire [7:0] op_16;
wire [31:0] op_17;
wire [3:0] op_18_V_fu_565_p3;
wire [31:0] op_19;
wire [3:0] op_2;
wire [8:0] op_22_V_fu_295_p2;
wire [28:0] op_25_V_fu_395_p2;
wire [28:0] op_27_V_fu_412_p2;
wire [1:0] op_3;
wire [31:0] op_30;
wire op_30_ap_vld;
wire op_5;
wire [1:0] op_6_V_fu_193_p1;
wire [1:0] op_6_V_fu_193_p2;
wire op_8_V_fu_199_p2;
wire or_ln340_1_fu_530_p2;
wire or_ln340_fu_525_p2;
wire or_ln785_1_fu_550_p2;
wire or_ln785_fu_506_p2;
wire overflow_fu_515_p2;
wire p_Result_1_fu_588_p3;
wire p_Result_2_fu_643_p3;
wire [1:0] p_Result_3_fu_215_p1;
wire p_Result_3_fu_215_p3;
wire p_Result_s_fu_345_p3;
wire [3:0] p_Val2_1_fu_499_p3;
wire r_fu_245_p1;
wire [2:0] ret_1_fu_424_p2;
wire [32:0] ret_V_1_fu_316_p2;
wire [28:0] ret_V_2_fu_365_p3;
wire [28:0] ret_V_3_fu_391_p2;
wire [28:0] ret_V_4_fu_403_p2;
wire [42:0] ret_V_5_fu_473_p2;
wire [34:0] ret_V_6_fu_622_p2;
wire [34:0] ret_V_6_reg_797;
wire [31:0] ret_V_7_fu_655_p3;
wire [2:0] ret_V_fu_209_p2;
wire [3:0] ret_fu_282_p0;
wire [3:0] ret_fu_282_p1;
wire [7:0] ret_fu_282_p2;
wire [13:0] rhs_2_fu_305_p3;
wire [33:0] rhs_6_fu_610_p3;
wire [28:0] select_ln1192_fu_373_p3;
wire [3:0] select_ln340_fu_536_p3;
wire [31:0] select_ln353_fu_603_p3;
wire [15:0] select_ln546_fu_223_p3;
wire [28:0] select_ln69_1_fu_271_p3;
wire [2:0] select_ln69_fu_257_p3;
wire select_ln769_fu_249_p3;
wire [31:0] select_ln850_1_fu_598_p3;
wire [31:0] select_ln850_2_fu_650_p3;
wire [28:0] select_ln850_fu_358_p3;
wire [32:0] sext_ln1192_1_fu_312_p1;
wire [42:0] sext_ln1192_2_fu_469_p1;
wire [34:0] sext_ln1192_3_fu_618_p1;
wire [31:0] sext_ln1192_fu_301_p0;
wire [32:0] sext_ln1192_fu_301_p1;
wire [1:0] sext_ln1347_1_fu_421_p0;
wire [2:0] sext_ln1347_1_fu_421_p1;
wire [1:0] sext_ln1347_fu_418_p0;
wire [2:0] sext_ln1347_fu_418_p1;
wire [8:0] sext_ln69_1_fu_292_p1;
wire [28:0] sext_ln69_2_fu_408_p1;
wire [8:0] sext_ln69_fu_288_p1;
wire [31:0] sext_ln703_1_fu_458_p0;
wire [42:0] sext_ln703_1_fu_458_p1;
wire [34:0] sext_ln703_2_fu_595_p1;
wire [2:0] sext_ln703_fu_205_p1;
wire [1:0] sext_ln781_fu_231_p0;
wire [3:0] sext_ln781_fu_231_p1;
wire [28:0] sext_ln850_fu_342_p1;
wire [1:0] sext_ln874_fu_381_p0;
wire [31:0] sext_ln874_fu_381_p1;
wire [15:0] shl_ln781_fu_239_p2;
wire [38:0] tmp_7_fu_462_p3;
wire [1:0] trunc_ln69_1_fu_189_p1;
wire trunc_ln69_fu_185_p1;
wire [1:0] trunc_ln731_fu_438_p1;
wire [31:0] trunc_ln851_1_fu_489_p0;
wire [9:0] trunc_ln851_1_fu_489_p1;
wire [1:0] trunc_ln851_2_fu_578_p1;
wire [31:0] trunc_ln851_fu_332_p0;
wire [4:0] trunc_ln851_fu_332_p1;
wire xor_ln785_1_fu_544_p2;
wire xor_ln785_fu_510_p2;
wire [28:0] zext_ln1192_fu_400_p1;
wire [7:0] zext_ln1345_fu_279_p1;
wire [15:0] zext_ln781_fu_235_p1;


assign add_ln691_1_fu_573_p2 = ret_V_5_cast_reg_770 + 1'h1;
assign add_ln691_2_fu_638_p2 = ret_V_8_cast_reg_802 + 1'h1;
assign add_ln691_fu_352_p2 = $signed(tmp_reg_699) + $signed(2'h1);
assign add_ln69_fu_265_p2 = ret_V_fu_209_p2 + select_ln69_fu_257_p3;
assign op_22_V_fu_295_p2 = $signed(add_ln69_reg_679) + $signed(ret_fu_282_p2);
assign op_25_V_fu_395_p2 = ret_V_3_fu_391_p2 + select_ln69_1_reg_684;
assign op_27_V_fu_412_p2 = $signed(ret_V_4_fu_403_p2) + $signed(op_16);
assign op_30 = ret_V_7_fu_655_p3 + op_19;
assign ret_V_1_fu_316_p2 = $signed({ op_22_V_reg_689, 5'h00 }) + $signed(op_12);
assign ret_V_3_fu_391_p2 = ret_V_2_reg_709 + select_ln1192_reg_714;
assign ret_V_4_fu_403_p2 = op_25_V_reg_729 + lhs_V_reg_724;
assign { ret_V_5_fu_473_p2[42], ret_V_5_fu_473_p2[38:0] } = $signed({ op_27_V_reg_734, 10'h000 }) + $signed(op_17);
assign ret_V_6_fu_622_p2 = $signed({ select_ln353_fu_603_p3, 2'h0 }) + $signed(op_18_V_reg_782);
assign ret_V_fu_209_p2 = $signed(op_6_V_fu_193_p2) + $signed(2'h1);
assign _026_ = ap_CS_fsm[7] & icmp_ln851_1_reg_777;
assign _027_ = ap_CS_fsm[9] & icmp_ln851_2_reg_792;
assign _028_ = ap_CS_fsm[0] & _030_;
assign _029_ = ap_CS_fsm[0] & ap_start;
assign and_ln785_1_fu_560_p2 = p_Result_5_reg_751 & and_ln785_fu_555_p2;
assign and_ln785_fu_555_p2 = tmp_5_reg_758 & or_ln785_1_fu_550_p2;
assign and_ln786_fu_521_p2 = tmp_5_reg_758 & p_Result_5_reg_751;
assign overflow_fu_515_p2 = xor_ln785_fu_510_p2 & or_ln785_fu_506_p2;
assign xor_ln785_1_fu_544_p2 = ~ or_ln785_fu_506_p2;
assign xor_ln785_fu_510_p2 = ~ p_Result_4_reg_739;
assign _030_ = ~ ap_start;
assign \mul_4ns_4ns_8_1_1_U1.top_mul_4ns_4ns_8_1_1_Multiplier_0_U.p  = \mul_4ns_4ns_8_1_1_U1.top_mul_4ns_4ns_8_1_1_Multiplier_0_U.a  * \mul_4ns_4ns_8_1_1_U1.top_mul_4ns_4ns_8_1_1_Multiplier_0_U.b ;
assign _031_ = | op_17[9:0];
assign _032_ = | op_18_V_fu_565_p3[1:0];
assign _033_ = | op_12[4:0];
assign _034_ = { op_10[1], op_10[1], op_10[1], op_10[1], op_10[1], op_10[1], op_10[1], op_10[1], op_10[1], op_10[1], op_10[1], op_10[1], op_10[1], op_10[1], op_10[1], op_10[1], op_10[1], op_10[1], op_10[1], op_10[1], op_10[1], op_10[1], op_10[1], op_10[1], op_10[1], op_10[1], op_10[1], op_10[1], op_10[1], op_10[1], op_10 } != op_11;
assign or_ln340_1_fu_530_p2 = or_ln340_fu_525_p2 | and_ln786_fu_521_p2;
assign or_ln340_fu_525_p2 = p_Result_4_reg_739 | overflow_fu_515_p2;
assign or_ln785_1_fu_550_p2 = xor_ln785_1_fu_544_p2 | p_Result_4_reg_739;
assign or_ln785_fu_506_p2 = tmp_5_reg_758 | p_Result_5_reg_751;
always @(posedge ap_clk)
op_18_V_reg_782[1:0] <= 2'h0;
always @(posedge ap_clk)
_081_ <= _018_;
assign ret_V_6_reg_797[34:2] = _081_;
always @(posedge ap_clk)
ret_V_8_cast_reg_802 <= _019_;
always @(posedge ap_clk)
ret_V_2_reg_709 <= _015_;
always @(posedge ap_clk)
select_ln1192_reg_714 <= _020_;
always @(posedge ap_clk)
op_27_V_reg_734 <= _011_;
always @(posedge ap_clk)
op_22_V_reg_689 <= _009_;
always @(posedge ap_clk)
lhs_V_reg_724 <= _007_;
always @(posedge ap_clk)
op_25_V_reg_729 <= _010_;
always @(posedge ap_clk)
ret_V_1_reg_694 <= _014_;
always @(posedge ap_clk)
tmp_reg_699 <= _023_;
always @(posedge ap_clk)
icmp_ln851_reg_704 <= _006_;
always @(posedge ap_clk)
op_18_V_reg_782[3:2] <= _008_;
always @(posedge ap_clk)
icmp_ln851_2_reg_792 <= _005_;
always @(posedge ap_clk)
p_Result_4_reg_739 <= _012_;
always @(posedge ap_clk)
trunc_ln731_reg_746 <= _024_;
always @(posedge ap_clk)
p_Result_5_reg_751 <= _013_;
always @(posedge ap_clk)
tmp_5_reg_758 <= _022_;
always @(posedge ap_clk)
ret_V_5_reg_765 <= _017_;
always @(posedge ap_clk)
ret_V_5_cast_reg_770 <= _016_;
always @(posedge ap_clk)
icmp_ln851_1_reg_777 <= _004_;
always @(posedge ap_clk)
add_ln69_reg_679 <= _002_;
always @(posedge ap_clk)
select_ln69_1_reg_684 <= _021_;
always @(posedge ap_clk)
add_ln691_2_reg_809 <= _001_;
always @(posedge ap_clk)
add_ln691_1_reg_787 <= _000_;
always @(posedge ap_clk)
ap_CS_fsm <= _003_;
assign _025_ = _029_ ? 2'h2 : 2'h1;
assign _035_ = ap_CS_fsm == 1'h1;
function [10:0] _108_;
input [10:0] a;
input [120:0] b;
input [10:0] s;
case (s)
11'b00000000001:
_108_ = b[10:0];
11'b00000000010:
_108_ = b[21:11];
11'b00000000100:
_108_ = b[32:22];
11'b00000001000:
_108_ = b[43:33];
11'b00000010000:
_108_ = b[54:44];
11'b00000100000:
_108_ = b[65:55];
11'b00001000000:
_108_ = b[76:66];
11'b00010000000:
_108_ = b[87:77];
11'b00100000000:
_108_ = b[98:88];
11'b01000000000:
_108_ = b[109:99];
11'b10000000000:
_108_ = b[120:110];
11'b00000000000:
_108_ = a;
default:
_108_ = 11'bx;
endcase
endfunction
assign ap_NS_fsm = _108_(11'hxxx, { 9'h000, _025_, 110'h0020080200802008020080200001 }, { _035_, _045_, _044_, _043_, _042_, _041_, _040_, _039_, _038_, _037_, _036_ });
assign _036_ = ap_CS_fsm == 11'h400;
assign _037_ = ap_CS_fsm == 10'h200;
assign _038_ = ap_CS_fsm == 9'h100;
assign _039_ = ap_CS_fsm == 8'h80;
assign _040_ = ap_CS_fsm == 7'h40;
assign _041_ = ap_CS_fsm == 6'h20;
assign _042_ = ap_CS_fsm == 5'h10;
assign _043_ = ap_CS_fsm == 4'h8;
assign _044_ = ap_CS_fsm == 3'h4;
assign _045_ = ap_CS_fsm == 2'h2;
assign op_30_ap_vld = ap_CS_fsm[10] ? 1'h1 : 1'h0;
assign ap_idle = _028_ ? 1'h1 : 1'h0;
assign _019_ = ap_CS_fsm[8] ? ret_V_6_fu_622_p2[33:2] : ret_V_8_cast_reg_802;
assign _018_ = ap_CS_fsm[8] ? ret_V_6_fu_622_p2[34:2] : ret_V_6_reg_797[34:2];
assign _020_ = ap_CS_fsm[3] ? select_ln1192_fu_373_p3 : select_ln1192_reg_714;
assign _015_ = ap_CS_fsm[3] ? ret_V_2_fu_365_p3 : ret_V_2_reg_709;
assign _011_ = ap_CS_fsm[5] ? op_27_V_fu_412_p2 : op_27_V_reg_734;
assign _009_ = ap_CS_fsm[1] ? op_22_V_fu_295_p2 : op_22_V_reg_689;
assign _010_ = ap_CS_fsm[4] ? op_25_V_fu_395_p2 : op_25_V_reg_729;
assign _007_ = ap_CS_fsm[4] ? lhs_V_fu_385_p2 : lhs_V_reg_724;
assign _006_ = ap_CS_fsm[2] ? icmp_ln851_fu_336_p2 : icmp_ln851_reg_704;
assign _023_ = ap_CS_fsm[2] ? ret_V_1_fu_316_p2[32:5] : tmp_reg_699;
assign _014_ = ap_CS_fsm[2] ? ret_V_1_fu_316_p2 : ret_V_1_reg_694;
assign _005_ = ap_CS_fsm[7] ? icmp_ln851_2_fu_582_p2 : icmp_ln851_2_reg_792;
assign _008_ = ap_CS_fsm[7] ? op_18_V_fu_565_p3[3:2] : op_18_V_reg_782[3:2];
assign _004_ = ap_CS_fsm[6] ? icmp_ln851_1_fu_493_p2 : icmp_ln851_1_reg_777;
assign _016_ = ap_CS_fsm[6] ? { ret_V_5_fu_473_p2[42], ret_V_5_fu_473_p2[42], ret_V_5_fu_473_p2[42], ret_V_5_fu_473_p2[38:10] } : ret_V_5_cast_reg_770;
assign _017_ = ap_CS_fsm[6] ? { ret_V_5_fu_473_p2[42], ret_V_5_fu_473_p2[42], ret_V_5_fu_473_p2[42], ret_V_5_fu_473_p2[42], ret_V_5_fu_473_p2[38:0] } : ret_V_5_reg_765;
assign _022_ = ap_CS_fsm[6] ? ret_1_fu_424_p2[2] : tmp_5_reg_758;
assign _013_ = ap_CS_fsm[6] ? ret_1_fu_424_p2[1] : p_Result_5_reg_751;
assign _024_ = ap_CS_fsm[6] ? ret_1_fu_424_p2[1:0] : trunc_ln731_reg_746;
assign _012_ = ap_CS_fsm[6] ? ret_1_fu_424_p2[2] : p_Result_4_reg_739;
assign _021_ = ap_CS_fsm[0] ? select_ln69_1_fu_271_p3 : select_ln69_1_reg_684;
assign _002_ = ap_CS_fsm[0] ? add_ln69_fu_265_p2 : add_ln69_reg_679;
assign _001_ = _027_ ? add_ln691_2_fu_638_p2 : add_ln691_2_reg_809;
assign _000_ = _026_ ? add_ln691_1_fu_573_p2 : add_ln691_1_reg_787;
assign _003_ = ap_rst ? 11'h001 : ap_NS_fsm;
assign r_fu_245_p1 = select_ln546_fu_223_p3 << { op_3[1], op_3[1], op_3 };
assign op_6_V_fu_193_p2 = $signed(op_2[1:0]) - $signed(op_3);
assign ret_1_fu_424_p2 = $signed(op_3) - $signed(op_10);
assign icmp_ln851_1_fu_493_p2 = _031_ ? 1'h1 : 1'h0;
assign icmp_ln851_2_fu_582_p2 = _032_ ? 1'h1 : 1'h0;
assign icmp_ln851_fu_336_p2 = _033_ ? 1'h1 : 1'h0;
assign lhs_V_fu_385_p2 = _034_ ? 1'h1 : 1'h0;
assign op_18_V_fu_565_p3 = and_ln785_1_fu_560_p2 ? { trunc_ln731_reg_746, 2'h0 } : select_ln340_fu_536_p3;
assign ret_V_2_fu_365_p3 = ret_V_1_reg_694[32] ? select_ln850_fu_358_p3 : { tmp_reg_699[27], tmp_reg_699 };
assign ret_V_7_fu_655_p3 = ret_V_6_reg_797[34] ? select_ln850_2_fu_650_p3 : ret_V_8_cast_reg_802;
assign select_ln1192_fu_373_p3 = op_13 ? 29'h1fffffff : 29'h00000000;
assign select_ln340_fu_536_p3 = or_ln340_1_fu_530_p2 ? 4'h0 : { trunc_ln731_reg_746, 2'h0 };
assign select_ln353_fu_603_p3 = ret_V_5_reg_765[42] ? select_ln850_1_fu_598_p3 : ret_V_5_cast_reg_770;
assign select_ln546_fu_223_p3 = op_5 ? 16'hffff : 16'h0000;
assign select_ln69_1_fu_271_p3 = select_ln769_fu_249_p3 ? 29'h1fffffff : 29'h00000000;
assign select_ln69_fu_257_p3 = op_8_V_fu_199_p2 ? 3'h7 : 3'h0;
assign select_ln769_fu_249_p3 = op_3[1] ? op_5 : r_fu_245_p1;
assign select_ln850_1_fu_598_p3 = icmp_ln851_1_reg_777 ? add_ln691_1_reg_787 : ret_V_5_cast_reg_770;
assign select_ln850_2_fu_650_p3 = icmp_ln851_2_reg_792 ? add_ln691_2_reg_809 : ret_V_8_cast_reg_802;
assign select_ln850_fu_358_p3 = icmp_ln851_reg_704 ? add_ln691_fu_352_p2 : { tmp_reg_699[27], tmp_reg_699 };
assign op_8_V_fu_199_p2 = op_2[0] ^ op_5;
assign ap_CS_fsm_state1 = ap_CS_fsm[0];
assign ap_CS_fsm_state10 = ap_CS_fsm[9];
assign ap_CS_fsm_state11 = ap_CS_fsm[10];
assign ap_CS_fsm_state2 = ap_CS_fsm[1];
assign ap_CS_fsm_state3 = ap_CS_fsm[2];
assign ap_CS_fsm_state4 = ap_CS_fsm[3];
assign ap_CS_fsm_state5 = ap_CS_fsm[4];
assign ap_CS_fsm_state6 = ap_CS_fsm[5];
assign ap_CS_fsm_state7 = ap_CS_fsm[6];
assign ap_CS_fsm_state8 = ap_CS_fsm[7];
assign ap_CS_fsm_state9 = ap_CS_fsm[8];
assign ap_done = op_30_ap_vld;
assign ap_ready = op_30_ap_vld;
assign op_6_V_fu_193_p1 = op_3;
assign p_Result_1_fu_588_p3 = ret_V_5_reg_765[42];
assign p_Result_2_fu_643_p3 = ret_V_6_reg_797[34];
assign p_Result_3_fu_215_p1 = op_3;
assign p_Result_3_fu_215_p3 = op_3[1];
assign p_Result_s_fu_345_p3 = ret_V_1_reg_694[32];
assign p_Val2_1_fu_499_p3 = { trunc_ln731_reg_746, 2'h0 };
assign ret_V_5_fu_473_p2[41:39] = { ret_V_5_fu_473_p2[42], ret_V_5_fu_473_p2[42], ret_V_5_fu_473_p2[42] };
assign ret_fu_282_p0 = op_2;
assign ret_fu_282_p1 = op_2;
assign rhs_2_fu_305_p3 = { op_22_V_reg_689, 5'h00 };
assign rhs_6_fu_610_p3 = { select_ln353_fu_603_p3, 2'h0 };
assign sext_ln1192_1_fu_312_p1 = { op_22_V_reg_689[8], op_22_V_reg_689[8], op_22_V_reg_689[8], op_22_V_reg_689[8], op_22_V_reg_689[8], op_22_V_reg_689[8], op_22_V_reg_689[8], op_22_V_reg_689[8], op_22_V_reg_689[8], op_22_V_reg_689[8], op_22_V_reg_689[8], op_22_V_reg_689[8], op_22_V_reg_689[8], op_22_V_reg_689[8], op_22_V_reg_689[8], op_22_V_reg_689[8], op_22_V_reg_689[8], op_22_V_reg_689[8], op_22_V_reg_689[8], op_22_V_reg_689, 5'h00 };
assign sext_ln1192_2_fu_469_p1 = { op_27_V_reg_734[28], op_27_V_reg_734[28], op_27_V_reg_734[28], op_27_V_reg_734[28], op_27_V_reg_734, 10'h000 };
assign sext_ln1192_3_fu_618_p1 = { select_ln353_fu_603_p3[31], select_ln353_fu_603_p3, 2'h0 };
assign sext_ln1192_fu_301_p0 = op_12;
assign sext_ln1192_fu_301_p1 = { op_12[31], op_12 };
assign sext_ln1347_1_fu_421_p0 = op_10;
assign sext_ln1347_1_fu_421_p1 = { op_10[1], op_10 };
assign sext_ln1347_fu_418_p0 = op_3;
assign sext_ln1347_fu_418_p1 = { op_3[1], op_3 };
assign sext_ln69_1_fu_292_p1 = { add_ln69_reg_679[2], add_ln69_reg_679[2], add_ln69_reg_679[2], add_ln69_reg_679[2], add_ln69_reg_679[2], add_ln69_reg_679[2], add_ln69_reg_679 };
assign sext_ln69_2_fu_408_p1 = { op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16 };
assign sext_ln69_fu_288_p1 = { ret_fu_282_p2[7], ret_fu_282_p2 };
assign sext_ln703_1_fu_458_p0 = op_17;
assign sext_ln703_1_fu_458_p1 = { op_17[31], op_17[31], op_17[31], op_17[31], op_17[31], op_17[31], op_17[31], op_17[31], op_17[31], op_17[31], op_17[31], op_17 };
assign sext_ln703_2_fu_595_p1 = { op_18_V_reg_782[3], op_18_V_reg_782[3], op_18_V_reg_782[3], op_18_V_reg_782[3], op_18_V_reg_782[3], op_18_V_reg_782[3], op_18_V_reg_782[3], op_18_V_reg_782[3], op_18_V_reg_782[3], op_18_V_reg_782[3], op_18_V_reg_782[3], op_18_V_reg_782[3], op_18_V_reg_782[3], op_18_V_reg_782[3], op_18_V_reg_782[3], op_18_V_reg_782[3], op_18_V_reg_782[3], op_18_V_reg_782[3], op_18_V_reg_782[3], op_18_V_reg_782[3], op_18_V_reg_782[3], op_18_V_reg_782[3], op_18_V_reg_782[3], op_18_V_reg_782[3], op_18_V_reg_782[3], op_18_V_reg_782[3], op_18_V_reg_782[3], op_18_V_reg_782[3], op_18_V_reg_782[3], op_18_V_reg_782[3], op_18_V_reg_782[3], op_18_V_reg_782 };
assign sext_ln703_fu_205_p1 = { op_6_V_fu_193_p2[1], op_6_V_fu_193_p2 };
assign sext_ln781_fu_231_p0 = op_3;
assign sext_ln781_fu_231_p1 = { op_3[1], op_3[1], op_3 };
assign sext_ln850_fu_342_p1 = { tmp_reg_699[27], tmp_reg_699 };
assign sext_ln874_fu_381_p0 = op_10;
assign sext_ln874_fu_381_p1 = { op_10[1], op_10[1], op_10[1], op_10[1], op_10[1], op_10[1], op_10[1], op_10[1], op_10[1], op_10[1], op_10[1], op_10[1], op_10[1], op_10[1], op_10[1], op_10[1], op_10[1], op_10[1], op_10[1], op_10[1], op_10[1], op_10[1], op_10[1], op_10[1], op_10[1], op_10[1], op_10[1], op_10[1], op_10[1], op_10[1], op_10 };
assign shl_ln781_fu_239_p2[0] = r_fu_245_p1;
assign tmp_7_fu_462_p3 = { op_27_V_reg_734, 10'h000 };
assign trunc_ln69_1_fu_189_p1 = op_2[1:0];
assign trunc_ln69_fu_185_p1 = op_2[0];
assign trunc_ln731_fu_438_p1 = ret_1_fu_424_p2[1:0];
assign trunc_ln851_1_fu_489_p0 = op_17;
assign trunc_ln851_1_fu_489_p1 = op_17[9:0];
assign trunc_ln851_2_fu_578_p1 = op_18_V_fu_565_p3[1:0];
assign trunc_ln851_fu_332_p0 = op_12;
assign trunc_ln851_fu_332_p1 = op_12[4:0];
assign zext_ln1192_fu_400_p1 = { 28'h0000000, lhs_V_reg_724 };
assign zext_ln1345_fu_279_p1 = { 4'h0, op_2 };
assign zext_ln781_fu_235_p1 = { 12'h000, op_3[1], op_3[1], op_3 };
assign \mul_4ns_4ns_8_1_1_U1.top_mul_4ns_4ns_8_1_1_Multiplier_0_U.a  = \mul_4ns_4ns_8_1_1_U1.din0 ;
assign \mul_4ns_4ns_8_1_1_U1.top_mul_4ns_4ns_8_1_1_Multiplier_0_U.b  = \mul_4ns_4ns_8_1_1_U1.din1 ;
assign \mul_4ns_4ns_8_1_1_U1.dout  = \mul_4ns_4ns_8_1_1_U1.top_mul_4ns_4ns_8_1_1_Multiplier_0_U.p ;
assign \mul_4ns_4ns_8_1_1_U1.din0  = op_2;
assign \mul_4ns_4ns_8_1_1_U1.din1  = op_2;
assign ret_fu_282_p2 = \mul_4ns_4ns_8_1_1_U1.dout ;
endmodule


// Product machine:
module top_A_times_top_B (ap_start, op_0, op_10, op_11, op_12, op_13, op_16, op_17, op_19, op_2, op_3, op_5, ap_clk, unsafe_signal);
input ap_start;
input [31:0] op_0;
input [1:0] op_10;
input [31:0] op_11;
input [31:0] op_12;
input op_13;
input [7:0] op_16;
input [31:0] op_17;
input [31:0] op_19;
input [3:0] op_2;
input [1:0] op_3;
input op_5;
input ap_clk;
output unsafe_signal;
reg _setup;
initial _setup = 1'b0;
always @ (posedge ap_clk) _setup <= 1'b1;
reg ap_start_internal;
always @ (posedge ap_clk) if (!_setup) ap_start_internal <= ap_start;
reg [31:0] op_0_internal;
always @ (posedge ap_clk) if (!_setup) op_0_internal <= op_0;
reg [1:0] op_10_internal;
always @ (posedge ap_clk) if (!_setup) op_10_internal <= op_10;
reg [31:0] op_11_internal;
always @ (posedge ap_clk) if (!_setup) op_11_internal <= op_11;
reg [31:0] op_12_internal;
always @ (posedge ap_clk) if (!_setup) op_12_internal <= op_12;
reg op_13_internal;
always @ (posedge ap_clk) if (!_setup) op_13_internal <= op_13;
reg [7:0] op_16_internal;
always @ (posedge ap_clk) if (!_setup) op_16_internal <= op_16;
reg [31:0] op_17_internal;
always @ (posedge ap_clk) if (!_setup) op_17_internal <= op_17;
reg [31:0] op_19_internal;
always @ (posedge ap_clk) if (!_setup) op_19_internal <= op_19;
reg [3:0] op_2_internal;
always @ (posedge ap_clk) if (!_setup) op_2_internal <= op_2;
reg [1:0] op_3_internal;
always @ (posedge ap_clk) if (!_setup) op_3_internal <= op_3;
reg op_5_internal;
always @ (posedge ap_clk) if (!_setup) op_5_internal <= op_5;
wire ap_done_A;
wire ap_done_B;
wire ap_done_eq;
assign ap_done_eq = ap_done_A == ap_done_B;
wire ap_idle_A;
wire ap_idle_B;
wire ap_idle_eq;
assign ap_idle_eq = ap_idle_A == ap_idle_B;
wire ap_ready_A;
wire ap_ready_B;
wire ap_ready_eq;
assign ap_ready_eq = ap_ready_A == ap_ready_B;
wire [31:0] op_30_A;
wire [31:0] op_30_B;
wire op_30_eq;
assign op_30_eq = op_30_A == op_30_B;
wire op_30_ap_vld_A;
wire op_30_ap_vld_B;
wire clk_enable_A;
wire clk_enable_B;
assign clk_enable_A = _setup & (~op_30_ap_vld_A | op_30_ap_vld_B);
assign clk_enable_B = _setup;
wire divergent;
assign divergent = ~(ap_done_eq & ap_idle_eq & ap_ready_eq & op_30_eq);
assign unsafe_signal = op_30_ap_vld_A & op_30_ap_vld_B & divergent;
top_A instance_A (
    .ap_clk(ap_clk),
    .clk_enable(clk_enable_A),
    .ap_start(ap_start_internal),
    .op_0(op_0_internal),
    .op_10(op_10_internal),
    .op_11(op_11_internal),
    .op_12(op_12_internal),
    .op_13(op_13_internal),
    .op_16(op_16_internal),
    .op_17(op_17_internal),
    .op_19(op_19_internal),
    .op_2(op_2_internal),
    .op_3(op_3_internal),
    .op_5(op_5_internal),
    .ap_done(ap_done_A),
    .ap_idle(ap_idle_A),
    .ap_ready(ap_ready_A),
    .op_30(op_30_A),
    .op_30_ap_vld(op_30_ap_vld_A)
);
top_B instance_B (
    .ap_clk(ap_clk),
    .clk_enable(clk_enable_B),
    .ap_start(ap_start_internal),
    .op_0(op_0_internal),
    .op_10(op_10_internal),
    .op_11(op_11_internal),
    .op_12(op_12_internal),
    .op_13(op_13_internal),
    .op_16(op_16_internal),
    .op_17(op_17_internal),
    .op_19(op_19_internal),
    .op_2(op_2_internal),
    .op_3(op_3_internal),
    .op_5(op_5_internal),
    .ap_done(ap_done_B),
    .ap_idle(ap_idle_B),
    .ap_ready(ap_ready_B),
    .op_30(op_30_B),
    .op_30_ap_vld(op_30_ap_vld_B)
);
endmodule
