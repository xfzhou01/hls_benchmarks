// Processed by function `construct_kairos` in `verilog_tricks.py`.
// Machine A:
// Processed by function `add_clk_enable_signal` in `verilog_tricks.py`.
// Processed by function `remove_reset_signal` in `verilog_tricks.py`.
module top_A (
  ap_clk,
  ap_start,
  ap_done,
  ap_idle,
  ap_ready,
  op_0,
  op_3,
  op_4,
  op_6,
  op_7,
  op_12,
  op_15,
  op_16,
  op_17,
  op_18,
  op_29,
  op_29_ap_vld,
clk_enable
);
input clk_enable;


input ap_clk;
wire ap_rst;
assign ap_rst = op_29_ap_vld;
input ap_start;
input [1:0] op_0;
input [7:0] op_12;
input [7:0] op_15;
input [3:0] op_16;
input [7:0] op_17;
input [3:0] op_18;
input [3:0] op_3;
input op_4;
input [3:0] op_6;
input [15:0] op_7;
output ap_done;
output ap_idle;
output ap_ready;
output [31:0] op_29;
output op_29_ap_vld;


reg [8:0] add_ln69_reg_941;
reg [7:0] ap_CS_fsm = 8'h01;
reg icmp_ln786_reg_878;
reg icmp_ln851_1_reg_812;
reg icmp_ln851_2_reg_832;
reg icmp_ln851_reg_921;
reg [1:0] op_14_V_reg_893;
reg [5:0] op_20_V_reg_848;
reg or_ln785_reg_873;
reg p_Result_4_reg_858;
reg p_Result_5_reg_868;
reg [1:0] p_Val2_s_reg_863;
reg [1:0] ret_V_10_reg_827;
reg [31:0] ret_V_16_cast_reg_903;
reg [4:0] ret_V_21_reg_801;
reg [3:0] ret_V_23_reg_822;
reg [6:0] ret_V_25_reg_888;
reg [33:0] ret_V_26_reg_898;
reg [31:0] ret_V_27_reg_931;
reg [31:0] ret_V_28_reg_936;
reg [7:0] ret_V_2_reg_915;
reg [7:0] ret_V_3_reg_926;
reg [2:0] ret_V_6_reg_806;
reg [2:0] ret_V_7_reg_817;
reg [1:0] select_ln340_reg_883;
reg [4:0] sub_ln1497_reg_843;
reg tmp_6_reg_796;
reg [5:0] _082_;
reg [7:0] _088_;
wire [8:0] _000_;
wire [7:0] _001_;
wire _002_;
wire _003_;
wire _004_;
wire _005_;
wire [1:0] _006_;
wire [5:0] _007_;
wire _008_;
wire _009_;
wire _010_;
wire [5:0] _011_;
wire [1:0] _012_;
wire [1:0] _013_;
wire [31:0] _014_;
wire [7:0] _015_;
wire [4:0] _016_;
wire [3:0] _017_;
wire [6:0] _018_;
wire [33:0] _019_;
wire [31:0] _020_;
wire [31:0] _021_;
wire [7:0] _022_;
wire [7:0] _023_;
wire [2:0] _024_;
wire [2:0] _025_;
wire [1:0] _026_;
wire [4:0] _027_;
wire _028_;
wire [1:0] _029_;
wire _030_;
wire _031_;
wire _032_;
wire _033_;
wire _034_;
wire _035_;
wire _036_;
wire _037_;
wire _038_;
wire _039_;
wire _040_;
wire _041_;
wire _042_;
wire _043_;
wire _044_;
wire _045_;
wire [31:0] add_ln691_fu_701_p2;
wire [8:0] add_ln69_fu_766_p2;
wire and_ln340_fu_544_p2;
wire and_ln785_1_fu_606_p2;
wire and_ln785_fu_600_p2;
wire ap_CS_fsm_state1;
wire ap_CS_fsm_state2;
wire ap_CS_fsm_state3;
wire ap_CS_fsm_state4;
wire ap_CS_fsm_state5;
wire ap_CS_fsm_state6;
wire ap_CS_fsm_state7;
wire ap_CS_fsm_state8;
wire [7:0] ap_NS_fsm;
wire ap_clk;
wire ap_done;
wire ap_idle;
wire ap_ready;
wire ap_rst;
wire ap_start;
wire [31:0] conv_i2826_fu_365_p1;
wire [6:0] empty_fu_428_p1;
wire icmp_ln768_fu_490_p2;
wire icmp_ln786_fu_520_p2;
wire icmp_ln851_1_fu_231_p2;
wire icmp_ln851_2_fu_271_p2;
wire icmp_ln851_fu_679_p2;
wire lhs_fu_432_p0;
wire [6:0] lhs_fu_432_p3;
wire [31:0] lshr_ln1497_fu_368_p2;
wire [1:0] op_0;
wire [7:0] op_11_V_fu_403_p3;
wire [7:0] op_12;
wire op_13_V_fu_446_p3;
wire [1:0] op_14_V_fu_611_p3;
wire [7:0] op_15;
wire [3:0] op_16;
wire [7:0] op_17;
wire [3:0] op_18;
wire [5:0] op_20_V_fu_349_p2;
wire [5:0] op_22_V_fu_558_p4;
wire [31:0] op_25_V_fu_747_p2;
wire [31:0] op_29;
wire op_29_ap_vld;
wire [3:0] op_3;
wire op_4;
wire [3:0] op_6;
wire [15:0] op_7;
wire or_ln340_fu_532_p2;
wire or_ln785_1_fu_595_p2;
wire or_ln785_fu_496_p2;
wire or_ln786_fu_526_p2;
wire overflow_fu_508_p2;
wire p_Result_1_fu_277_p3;
wire p_Result_2_fu_303_p3;
wire p_Result_3_fu_691_p3;
wire p_Result_4_fu_454_p3;
wire p_Result_5_fu_472_p3;
wire p_Result_s_14_fu_720_p3;
wire [8:0] p_Result_s_fu_480_p4;
wire [9:0] p_Val2_5_fu_422_p2;
wire [9:0] p_Val2_5_reg_853;
wire [1:0] p_Val2_s_fu_462_p4;
wire [2:0] ret_V_11_fu_310_p2;
wire [9:0] ret_V_19_fu_659_p2;
wire [9:0] ret_V_19_reg_910;
wire [7:0] ret_V_20_fu_732_p3;
wire [4:0] ret_V_21_fu_211_p2;
wire [2:0] ret_V_22_fu_289_p3;
wire [3:0] ret_V_23_fu_251_p1;
wire [3:0] ret_V_23_fu_251_p2;
wire [2:0] ret_V_24_fu_323_p3;
wire [6:0] ret_V_25_fu_579_p2;
wire [33:0] ret_V_26_fu_632_p2;
wire [31:0] ret_V_27_fu_713_p3;
wire [31:0] ret_V_28_fu_756_p2;
wire [31:0] ret_V_29_fu_776_p2;
wire [7:0] ret_V_2_fu_665_p4;
wire [7:0] ret_V_3_fu_685_p2;
wire [2:0] ret_V_6_fu_217_p4;
wire [2:0] ret_V_7_fu_237_p2;
wire [6:0] ret_V_fu_440_p2;
wire [9:0] rhs_2_fu_415_p3;
wire [9:0] rhs_fu_651_p3;
wire [6:0] select_ln1192_fu_571_p3;
wire [2:0] select_ln1196_fu_243_p3;
wire [3:0] select_ln1497_fu_395_p3;
wire [1:0] select_ln340_fu_550_p3;
wire [2:0] select_ln850_1_fu_284_p3;
wire [2:0] select_ln850_2_fu_316_p3;
wire [31:0] select_ln850_3_fu_706_p3;
wire [7:0] select_ln850_fu_727_p3;
wire [33:0] sext_ln1192_1_fu_628_p1;
wire [31:0] sext_ln1192_2_fu_752_p1;
wire [31:0] sext_ln1192_3_fu_772_p1;
wire [9:0] sext_ln1192_fu_411_p1;
wire [31:0] sext_ln1497_1_fu_382_p1;
wire [3:0] sext_ln1497_fu_331_p0;
wire [4:0] sext_ln1497_fu_331_p1;
wire [5:0] sext_ln15_fu_296_p1;
wire [8:0] sext_ln21_fu_739_p1;
wire [6:0] sext_ln24_fu_567_p1;
wire [3:0] sext_ln545_fu_355_p0;
wire [31:0] sext_ln545_fu_355_p1;
wire [8:0] sext_ln69_1_fu_762_p1;
wire [31:0] sext_ln69_2_fu_781_p1;
wire [3:0] sext_ln69_3_fu_341_p1;
wire [31:0] sext_ln69_fu_743_p1;
wire [3:0] sext_ln703_1_fu_207_p0;
wire [4:0] sext_ln703_1_fu_207_p1;
wire [33:0] sext_ln703_2_fu_617_p1;
wire [3:0] sext_ln703_fu_648_p0;
wire [9:0] sext_ln703_fu_648_p1;
wire [2:0] sext_ln831_fu_300_p1;
wire [31:0] shl_ln1497_fu_385_p2;
wire [4:0] sub_ln1497_fu_335_p2;
wire tmp_6_fu_199_p3;
wire [7:0] tmp_8_fu_621_p3;
wire [3:0] tmp_fu_358_p1;
wire tmp_fu_358_p3;
wire trunc_ln1497_fu_374_p1;
wire [3:0] trunc_ln728_fu_391_p1;
wire [1:0] trunc_ln851_1_fu_227_p1;
wire [1:0] trunc_ln851_2_fu_267_p1;
wire trunc_ln851_3_fu_698_p1;
wire [1:0] trunc_ln851_fu_675_p1;
wire xor_ln340_fu_538_p2;
wire xor_ln785_1_fu_590_p2;
wire xor_ln785_fu_502_p2;
wire xor_ln786_1_fu_585_p2;
wire xor_ln786_fu_514_p2;
wire [3:0] zext_ln1497_fu_378_p1;
wire [5:0] zext_ln69_fu_345_p1;


assign add_ln691_fu_701_p2 = ret_V_16_cast_reg_903 + 1'h1;
assign add_ln69_fu_766_p2 = $signed(ret_V_20_fu_732_p3) + $signed(op_18);
assign op_20_V_fu_349_p2 = $signed({ 1'h0, ret_V_24_fu_323_p3[2], ret_V_24_fu_323_p3 }) + $signed(ret_V_22_fu_289_p3);
assign op_25_V_fu_747_p2 = $signed(ret_V_27_reg_931) + $signed(op_15);
assign op_29 = $signed(add_ln69_reg_941) + $signed(ret_V_29_fu_776_p2);
assign p_Val2_5_fu_422_p2 = $signed({ op_20_V_reg_848, 4'h0 }) + $signed({ select_ln1497_fu_395_p3, 4'h0 });
assign ret_V_11_fu_310_p2 = $signed(ret_V_10_reg_827) + $signed(2'h1);
assign ret_V_25_fu_579_p2 = $signed(p_Val2_5_reg_853[9:4]) + $signed(select_ln1192_fu_571_p3);
assign { ret_V_26_fu_632_p2[33], ret_V_26_fu_632_p2[7:0] } = $signed({ ret_V_25_reg_888, 1'h0 }) + $signed(op_14_V_fu_611_p3);
assign ret_V_28_fu_756_p2 = $signed(op_25_V_fu_747_p2) + $signed(op_16);
assign ret_V_29_fu_776_p2 = $signed(ret_V_28_reg_936) + $signed(op_17);
assign ret_V_3_fu_685_p2 = ret_V_19_fu_659_p2[9:2] + 1'h1;
assign ret_V_7_fu_237_p2 = ret_V_21_fu_211_p2[4:2] + 1'h1;
assign _030_ = ap_CS_fsm[0] & _032_;
assign _031_ = ap_CS_fsm[0] & ap_start;
assign and_ln340_fu_544_p2 = xor_ln340_fu_538_p2 & or_ln786_fu_526_p2;
assign and_ln785_1_fu_606_p2 = p_Result_5_reg_868 & and_ln785_fu_600_p2;
assign and_ln785_fu_600_p2 = xor_ln786_1_fu_585_p2 & or_ln785_1_fu_595_p2;
assign overflow_fu_508_p2 = xor_ln785_fu_502_p2 & or_ln785_fu_496_p2;
assign ret_V_19_fu_659_p2 = { op_3[3], op_3[3], op_3[3], op_3[3], op_3[3], op_3[3], op_3 } & { op_12, 2'h0 };
assign ret_V_fu_440_p2 = lhs_fu_432_p3 & op_7[6:0];
assign xor_ln786_fu_514_p2 = ~ op_7[6];
assign xor_ln785_fu_502_p2 = ~ op_7[15];
assign xor_ln340_fu_538_p2 = ~ or_ln340_fu_532_p2;
assign xor_ln785_1_fu_590_p2 = ~ or_ln785_reg_873;
assign xor_ln786_1_fu_585_p2 = ~ icmp_ln786_reg_878;
assign _032_ = ~ ap_start;
assign _033_ = ! ret_V_21_fu_211_p2[1:0];
assign _034_ = ! ret_V_23_fu_251_p2[1:0];
assign _035_ = ! ret_V_19_fu_659_p2[1:0];
assign _036_ = | op_7[15:7];
assign _037_ = op_7[15:7] != 9'h1ff;
assign or_ln340_fu_532_p2 = op_7[15] | overflow_fu_508_p2;
assign or_ln785_1_fu_595_p2 = xor_ln785_1_fu_590_p2 | p_Result_4_reg_858;
assign or_ln785_fu_496_p2 = op_7[6] | icmp_ln768_fu_490_p2;
assign or_ln786_fu_526_p2 = xor_ln786_fu_514_p2 | icmp_ln786_fu_520_p2;
always @(posedge ap_clk)
_082_ <= _011_;
assign p_Val2_5_reg_853[9:4] = _082_;
always @(posedge ap_clk)
sub_ln1497_reg_843 <= _027_;
always @(posedge ap_clk)
op_20_V_reg_848 <= _007_;
always @(posedge ap_clk)
op_14_V_reg_893 <= _006_;
always @(posedge ap_clk)
ret_V_26_reg_898 <= _019_;
always @(posedge ap_clk)
ret_V_16_cast_reg_903 <= _014_;
always @(posedge ap_clk)
_088_ <= _015_;
assign ret_V_19_reg_910[9:2] = _088_;
always @(posedge ap_clk)
ret_V_2_reg_915 <= _022_;
always @(posedge ap_clk)
icmp_ln851_reg_921 <= _005_;
always @(posedge ap_clk)
ret_V_3_reg_926 <= _023_;
always @(posedge ap_clk)
ret_V_27_reg_931 <= _020_;
always @(posedge ap_clk)
tmp_6_reg_796 <= _028_;
always @(posedge ap_clk)
ret_V_21_reg_801 <= _016_;
always @(posedge ap_clk)
ret_V_6_reg_806 <= _024_;
always @(posedge ap_clk)
icmp_ln851_1_reg_812 <= _003_;
always @(posedge ap_clk)
ret_V_7_reg_817 <= _025_;
always @(posedge ap_clk)
ret_V_23_reg_822 <= _017_;
always @(posedge ap_clk)
ret_V_10_reg_827 <= _013_;
always @(posedge ap_clk)
icmp_ln851_2_reg_832 <= _004_;
always @(posedge ap_clk)
p_Result_4_reg_858 <= _009_;
always @(posedge ap_clk)
p_Val2_s_reg_863 <= _012_;
always @(posedge ap_clk)
p_Result_5_reg_868 <= _010_;
always @(posedge ap_clk)
or_ln785_reg_873 <= _008_;
always @(posedge ap_clk)
icmp_ln786_reg_878 <= _002_;
always @(posedge ap_clk)
select_ln340_reg_883 <= _026_;
always @(posedge ap_clk)
ret_V_25_reg_888 <= _018_;
always @(posedge ap_clk)
ret_V_28_reg_936 <= _021_;
always @(posedge ap_clk)
add_ln69_reg_941 <= _000_;
always @(posedge ap_clk)
ap_CS_fsm <= _001_;
assign _029_ = _031_ ? 2'h2 : 2'h1;
assign _038_ = ap_CS_fsm == 1'h1;
function [7:0] _113_;
input [7:0] a;
input [63:0] b;
input [7:0] s;
case (s)
8'b00000001:
_113_ = b[7:0];
8'b00000010:
_113_ = b[15:8];
8'b00000100:
_113_ = b[23:16];
8'b00001000:
_113_ = b[31:24];
8'b00010000:
_113_ = b[39:32];
8'b00100000:
_113_ = b[47:40];
8'b01000000:
_113_ = b[55:48];
8'b10000000:
_113_ = b[63:56];
8'b00000000:
_113_ = a;
default:
_113_ = 8'bx;
endcase
endfunction
assign ap_NS_fsm = _113_(8'hxx, { 6'h00, _029_, 56'h04081020408001 }, { _038_, _045_, _044_, _043_, _042_, _041_, _040_, _039_ });
assign _039_ = ap_CS_fsm == 8'h80;
assign _040_ = ap_CS_fsm == 7'h40;
assign _041_ = ap_CS_fsm == 6'h20;
assign _042_ = ap_CS_fsm == 5'h10;
assign _043_ = ap_CS_fsm == 4'h8;
assign _044_ = ap_CS_fsm == 3'h4;
assign _045_ = ap_CS_fsm == 2'h2;
assign op_29_ap_vld = ap_CS_fsm[7] ? 1'h1 : 1'h0;
assign ap_idle = _030_ ? 1'h1 : 1'h0;
assign _011_ = ap_CS_fsm[2] ? p_Val2_5_fu_422_p2[9:4] : p_Val2_5_reg_853[9:4];
assign _007_ = ap_CS_fsm[1] ? op_20_V_fu_349_p2 : op_20_V_reg_848;
assign _027_ = ap_CS_fsm[1] ? sub_ln1497_fu_335_p2 : sub_ln1497_reg_843;
assign _014_ = ap_CS_fsm[4] ? { ret_V_26_fu_632_p2[33], ret_V_26_fu_632_p2[33], ret_V_26_fu_632_p2[33], ret_V_26_fu_632_p2[33], ret_V_26_fu_632_p2[33], ret_V_26_fu_632_p2[33], ret_V_26_fu_632_p2[33], ret_V_26_fu_632_p2[33], ret_V_26_fu_632_p2[33], ret_V_26_fu_632_p2[33], ret_V_26_fu_632_p2[33], ret_V_26_fu_632_p2[33], ret_V_26_fu_632_p2[33], ret_V_26_fu_632_p2[33], ret_V_26_fu_632_p2[33], ret_V_26_fu_632_p2[33], ret_V_26_fu_632_p2[33], ret_V_26_fu_632_p2[33], ret_V_26_fu_632_p2[33], ret_V_26_fu_632_p2[33], ret_V_26_fu_632_p2[33], ret_V_26_fu_632_p2[33], ret_V_26_fu_632_p2[33], ret_V_26_fu_632_p2[33], ret_V_26_fu_632_p2[33], ret_V_26_fu_632_p2[7:1] } : ret_V_16_cast_reg_903;
assign _019_ = ap_CS_fsm[4] ? { ret_V_26_fu_632_p2[33], ret_V_26_fu_632_p2[33], ret_V_26_fu_632_p2[33], ret_V_26_fu_632_p2[33], ret_V_26_fu_632_p2[33], ret_V_26_fu_632_p2[33], ret_V_26_fu_632_p2[33], ret_V_26_fu_632_p2[33], ret_V_26_fu_632_p2[33], ret_V_26_fu_632_p2[33], ret_V_26_fu_632_p2[33], ret_V_26_fu_632_p2[33], ret_V_26_fu_632_p2[33], ret_V_26_fu_632_p2[33], ret_V_26_fu_632_p2[33], ret_V_26_fu_632_p2[33], ret_V_26_fu_632_p2[33], ret_V_26_fu_632_p2[33], ret_V_26_fu_632_p2[33], ret_V_26_fu_632_p2[33], ret_V_26_fu_632_p2[33], ret_V_26_fu_632_p2[33], ret_V_26_fu_632_p2[33], ret_V_26_fu_632_p2[33], ret_V_26_fu_632_p2[33], ret_V_26_fu_632_p2[33], ret_V_26_fu_632_p2[7:0] } : ret_V_26_reg_898;
assign _006_ = ap_CS_fsm[4] ? op_14_V_fu_611_p3 : op_14_V_reg_893;
assign _020_ = ap_CS_fsm[5] ? ret_V_27_fu_713_p3 : ret_V_27_reg_931;
assign _023_ = ap_CS_fsm[5] ? ret_V_3_fu_685_p2 : ret_V_3_reg_926;
assign _005_ = ap_CS_fsm[5] ? icmp_ln851_fu_679_p2 : icmp_ln851_reg_921;
assign _022_ = ap_CS_fsm[5] ? ret_V_19_fu_659_p2[9:2] : ret_V_2_reg_915;
assign _015_ = ap_CS_fsm[5] ? ret_V_19_fu_659_p2[9:2] : ret_V_19_reg_910[9:2];
assign _004_ = ap_CS_fsm[0] ? icmp_ln851_2_fu_271_p2 : icmp_ln851_2_reg_832;
assign _013_ = ap_CS_fsm[0] ? ret_V_23_fu_251_p2[3:2] : ret_V_10_reg_827;
assign _017_ = ap_CS_fsm[0] ? ret_V_23_fu_251_p2 : ret_V_23_reg_822;
assign _025_ = ap_CS_fsm[0] ? ret_V_7_fu_237_p2 : ret_V_7_reg_817;
assign _003_ = ap_CS_fsm[0] ? icmp_ln851_1_fu_231_p2 : icmp_ln851_1_reg_812;
assign _024_ = ap_CS_fsm[0] ? ret_V_21_fu_211_p2[4:2] : ret_V_6_reg_806;
assign _016_ = ap_CS_fsm[0] ? ret_V_21_fu_211_p2 : ret_V_21_reg_801;
assign _028_ = ap_CS_fsm[0] ? op_0[1] : tmp_6_reg_796;
assign _018_ = ap_CS_fsm[3] ? ret_V_25_fu_579_p2 : ret_V_25_reg_888;
assign _026_ = ap_CS_fsm[3] ? select_ln340_fu_550_p3 : select_ln340_reg_883;
assign _002_ = ap_CS_fsm[3] ? icmp_ln786_fu_520_p2 : icmp_ln786_reg_878;
assign _008_ = ap_CS_fsm[3] ? or_ln785_fu_496_p2 : or_ln785_reg_873;
assign _010_ = ap_CS_fsm[3] ? op_7[6] : p_Result_5_reg_868;
assign _012_ = ap_CS_fsm[3] ? op_7[6:5] : p_Val2_s_reg_863;
assign _009_ = ap_CS_fsm[3] ? op_7[15] : p_Result_4_reg_858;
assign _000_ = ap_CS_fsm[6] ? add_ln69_fu_766_p2 : add_ln69_reg_941;
assign _021_ = ap_CS_fsm[6] ? ret_V_28_fu_756_p2 : ret_V_28_reg_936;
assign _001_ = ap_rst ? 8'h01 : ap_NS_fsm;
assign trunc_ln728_fu_391_p1 = tmp_6_reg_796 << { sub_ln1497_reg_843[4], sub_ln1497_reg_843[4], sub_ln1497_reg_843[4], sub_ln1497_reg_843[4], sub_ln1497_reg_843[4], sub_ln1497_reg_843[4], sub_ln1497_reg_843[4], sub_ln1497_reg_843[4], sub_ln1497_reg_843[4], sub_ln1497_reg_843[4], sub_ln1497_reg_843[4], sub_ln1497_reg_843[4], sub_ln1497_reg_843[4], sub_ln1497_reg_843[4], sub_ln1497_reg_843[4], sub_ln1497_reg_843[4], sub_ln1497_reg_843[4], sub_ln1497_reg_843[4], sub_ln1497_reg_843[4], sub_ln1497_reg_843[4], sub_ln1497_reg_843[4], sub_ln1497_reg_843[4], sub_ln1497_reg_843[4], sub_ln1497_reg_843[4], sub_ln1497_reg_843[4], sub_ln1497_reg_843[4], sub_ln1497_reg_843[4], sub_ln1497_reg_843 };
assign trunc_ln1497_fu_374_p1 = tmp_6_reg_796 >> { op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6 };
assign ret_V_21_fu_211_p2 = $signed(1'h0) - $signed(op_3);
assign sub_ln1497_fu_335_p2 = $signed(1'h0) - $signed(op_6);
assign icmp_ln768_fu_490_p2 = _036_ ? 1'h1 : 1'h0;
assign icmp_ln786_fu_520_p2 = _037_ ? 1'h1 : 1'h0;
assign icmp_ln851_1_fu_231_p2 = _033_ ? 1'h1 : 1'h0;
assign icmp_ln851_2_fu_271_p2 = _034_ ? 1'h1 : 1'h0;
assign icmp_ln851_fu_679_p2 = _035_ ? 1'h1 : 1'h0;
assign lhs_fu_432_p3 = op_4 ? 7'h40 : 7'h00;
assign op_14_V_fu_611_p3 = and_ln785_1_fu_606_p2 ? p_Val2_s_reg_863 : select_ln340_reg_883;
assign ret_V_20_fu_732_p3 = ret_V_19_reg_910[9] ? select_ln850_fu_727_p3 : ret_V_2_reg_915;
assign ret_V_22_fu_289_p3 = ret_V_21_reg_801[4] ? select_ln850_1_fu_284_p3 : ret_V_6_reg_806;
assign ret_V_24_fu_323_p3 = ret_V_23_reg_822[3] ? select_ln850_2_fu_316_p3 : { ret_V_10_reg_827[1], ret_V_10_reg_827 };
assign ret_V_27_fu_713_p3 = ret_V_26_reg_898[33] ? select_ln850_3_fu_706_p3 : ret_V_16_cast_reg_903;
assign select_ln1192_fu_571_p3 = ret_V_fu_440_p2[6] ? 7'h7f : 7'h00;
assign select_ln1196_fu_243_p3 = op_0[1] ? 3'h4 : 3'h0;
assign select_ln1497_fu_395_p3 = op_6[3] ? trunc_ln728_fu_391_p1 : { 3'h0, trunc_ln1497_fu_374_p1 };
assign select_ln340_fu_550_p3 = and_ln340_fu_544_p2 ? op_7[6:5] : 2'h0;
assign select_ln850_1_fu_284_p3 = icmp_ln851_1_reg_812 ? ret_V_6_reg_806 : ret_V_7_reg_817;
assign select_ln850_2_fu_316_p3 = icmp_ln851_2_reg_832 ? { ret_V_10_reg_827[1], ret_V_10_reg_827 } : ret_V_11_fu_310_p2;
assign select_ln850_3_fu_706_p3 = op_14_V_reg_893[0] ? add_ln691_fu_701_p2 : ret_V_16_cast_reg_903;
assign select_ln850_fu_727_p3 = icmp_ln851_reg_921 ? ret_V_2_reg_915 : ret_V_3_reg_926;
assign ret_V_23_fu_251_p2 = select_ln1196_fu_243_p3 ^ op_3;
assign ap_CS_fsm_state1 = ap_CS_fsm[0];
assign ap_CS_fsm_state2 = ap_CS_fsm[1];
assign ap_CS_fsm_state3 = ap_CS_fsm[2];
assign ap_CS_fsm_state4 = ap_CS_fsm[3];
assign ap_CS_fsm_state5 = ap_CS_fsm[4];
assign ap_CS_fsm_state6 = ap_CS_fsm[5];
assign ap_CS_fsm_state7 = ap_CS_fsm[6];
assign ap_CS_fsm_state8 = ap_CS_fsm[7];
assign ap_done = op_29_ap_vld;
assign ap_ready = op_29_ap_vld;
assign conv_i2826_fu_365_p1 = { 31'h00000000, tmp_6_reg_796 };
assign empty_fu_428_p1 = op_7[6:0];
assign lhs_fu_432_p0 = op_4;
assign lshr_ln1497_fu_368_p2[0] = trunc_ln1497_fu_374_p1;
assign op_11_V_fu_403_p3 = { select_ln1497_fu_395_p3, 4'h0 };
assign op_13_V_fu_446_p3 = ret_V_fu_440_p2[6];
assign op_22_V_fu_558_p4 = p_Val2_5_reg_853[9:4];
assign p_Result_1_fu_277_p3 = ret_V_21_reg_801[4];
assign p_Result_2_fu_303_p3 = ret_V_23_reg_822[3];
assign p_Result_3_fu_691_p3 = ret_V_26_reg_898[33];
assign p_Result_4_fu_454_p3 = op_7[15];
assign p_Result_5_fu_472_p3 = op_7[6];
assign p_Result_s_14_fu_720_p3 = ret_V_19_reg_910[9];
assign p_Result_s_fu_480_p4 = op_7[15:7];
assign p_Val2_s_fu_462_p4 = op_7[6:5];
assign ret_V_23_fu_251_p1 = op_3;
assign ret_V_26_fu_632_p2[32:8] = { ret_V_26_fu_632_p2[33], ret_V_26_fu_632_p2[33], ret_V_26_fu_632_p2[33], ret_V_26_fu_632_p2[33], ret_V_26_fu_632_p2[33], ret_V_26_fu_632_p2[33], ret_V_26_fu_632_p2[33], ret_V_26_fu_632_p2[33], ret_V_26_fu_632_p2[33], ret_V_26_fu_632_p2[33], ret_V_26_fu_632_p2[33], ret_V_26_fu_632_p2[33], ret_V_26_fu_632_p2[33], ret_V_26_fu_632_p2[33], ret_V_26_fu_632_p2[33], ret_V_26_fu_632_p2[33], ret_V_26_fu_632_p2[33], ret_V_26_fu_632_p2[33], ret_V_26_fu_632_p2[33], ret_V_26_fu_632_p2[33], ret_V_26_fu_632_p2[33], ret_V_26_fu_632_p2[33], ret_V_26_fu_632_p2[33], ret_V_26_fu_632_p2[33], ret_V_26_fu_632_p2[33] };
assign ret_V_2_fu_665_p4 = ret_V_19_fu_659_p2[9:2];
assign ret_V_6_fu_217_p4 = ret_V_21_fu_211_p2[4:2];
assign rhs_2_fu_415_p3 = { op_20_V_reg_848, 4'h0 };
assign rhs_fu_651_p3 = { op_12, 2'h0 };
assign sext_ln1192_1_fu_628_p1 = { ret_V_25_reg_888[6], ret_V_25_reg_888[6], ret_V_25_reg_888[6], ret_V_25_reg_888[6], ret_V_25_reg_888[6], ret_V_25_reg_888[6], ret_V_25_reg_888[6], ret_V_25_reg_888[6], ret_V_25_reg_888[6], ret_V_25_reg_888[6], ret_V_25_reg_888[6], ret_V_25_reg_888[6], ret_V_25_reg_888[6], ret_V_25_reg_888[6], ret_V_25_reg_888[6], ret_V_25_reg_888[6], ret_V_25_reg_888[6], ret_V_25_reg_888[6], ret_V_25_reg_888[6], ret_V_25_reg_888[6], ret_V_25_reg_888[6], ret_V_25_reg_888[6], ret_V_25_reg_888[6], ret_V_25_reg_888[6], ret_V_25_reg_888[6], ret_V_25_reg_888[6], ret_V_25_reg_888, 1'h0 };
assign sext_ln1192_2_fu_752_p1 = { op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16 };
assign sext_ln1192_3_fu_772_p1 = { op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17 };
assign sext_ln1192_fu_411_p1 = { select_ln1497_fu_395_p3[3], select_ln1497_fu_395_p3[3], select_ln1497_fu_395_p3, 4'h0 };
assign sext_ln1497_1_fu_382_p1 = { sub_ln1497_reg_843[4], sub_ln1497_reg_843[4], sub_ln1497_reg_843[4], sub_ln1497_reg_843[4], sub_ln1497_reg_843[4], sub_ln1497_reg_843[4], sub_ln1497_reg_843[4], sub_ln1497_reg_843[4], sub_ln1497_reg_843[4], sub_ln1497_reg_843[4], sub_ln1497_reg_843[4], sub_ln1497_reg_843[4], sub_ln1497_reg_843[4], sub_ln1497_reg_843[4], sub_ln1497_reg_843[4], sub_ln1497_reg_843[4], sub_ln1497_reg_843[4], sub_ln1497_reg_843[4], sub_ln1497_reg_843[4], sub_ln1497_reg_843[4], sub_ln1497_reg_843[4], sub_ln1497_reg_843[4], sub_ln1497_reg_843[4], sub_ln1497_reg_843[4], sub_ln1497_reg_843[4], sub_ln1497_reg_843[4], sub_ln1497_reg_843[4], sub_ln1497_reg_843 };
assign sext_ln1497_fu_331_p0 = op_6;
assign sext_ln1497_fu_331_p1 = { op_6[3], op_6 };
assign sext_ln15_fu_296_p1 = { ret_V_22_fu_289_p3[2], ret_V_22_fu_289_p3[2], ret_V_22_fu_289_p3[2], ret_V_22_fu_289_p3 };
assign sext_ln21_fu_739_p1 = { ret_V_20_fu_732_p3[7], ret_V_20_fu_732_p3 };
assign sext_ln24_fu_567_p1 = { p_Val2_5_reg_853[9], p_Val2_5_reg_853[9:4] };
assign sext_ln545_fu_355_p0 = op_6;
assign sext_ln545_fu_355_p1 = { op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6 };
assign sext_ln69_1_fu_762_p1 = { op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18 };
assign sext_ln69_2_fu_781_p1 = { add_ln69_reg_941[8], add_ln69_reg_941[8], add_ln69_reg_941[8], add_ln69_reg_941[8], add_ln69_reg_941[8], add_ln69_reg_941[8], add_ln69_reg_941[8], add_ln69_reg_941[8], add_ln69_reg_941[8], add_ln69_reg_941[8], add_ln69_reg_941[8], add_ln69_reg_941[8], add_ln69_reg_941[8], add_ln69_reg_941[8], add_ln69_reg_941[8], add_ln69_reg_941[8], add_ln69_reg_941[8], add_ln69_reg_941[8], add_ln69_reg_941[8], add_ln69_reg_941[8], add_ln69_reg_941[8], add_ln69_reg_941[8], add_ln69_reg_941[8], add_ln69_reg_941 };
assign sext_ln69_3_fu_341_p1 = { ret_V_24_fu_323_p3[2], ret_V_24_fu_323_p3 };
assign sext_ln69_fu_743_p1 = { op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15 };
assign sext_ln703_1_fu_207_p0 = op_3;
assign sext_ln703_1_fu_207_p1 = { op_3[3], op_3 };
assign sext_ln703_2_fu_617_p1 = { op_14_V_fu_611_p3[1], op_14_V_fu_611_p3[1], op_14_V_fu_611_p3[1], op_14_V_fu_611_p3[1], op_14_V_fu_611_p3[1], op_14_V_fu_611_p3[1], op_14_V_fu_611_p3[1], op_14_V_fu_611_p3[1], op_14_V_fu_611_p3[1], op_14_V_fu_611_p3[1], op_14_V_fu_611_p3[1], op_14_V_fu_611_p3[1], op_14_V_fu_611_p3[1], op_14_V_fu_611_p3[1], op_14_V_fu_611_p3[1], op_14_V_fu_611_p3[1], op_14_V_fu_611_p3[1], op_14_V_fu_611_p3[1], op_14_V_fu_611_p3[1], op_14_V_fu_611_p3[1], op_14_V_fu_611_p3[1], op_14_V_fu_611_p3[1], op_14_V_fu_611_p3[1], op_14_V_fu_611_p3[1], op_14_V_fu_611_p3[1], op_14_V_fu_611_p3[1], op_14_V_fu_611_p3[1], op_14_V_fu_611_p3[1], op_14_V_fu_611_p3[1], op_14_V_fu_611_p3[1], op_14_V_fu_611_p3[1], op_14_V_fu_611_p3[1], op_14_V_fu_611_p3 };
assign sext_ln703_fu_648_p0 = op_3;
assign sext_ln703_fu_648_p1 = { op_3[3], op_3[3], op_3[3], op_3[3], op_3[3], op_3[3], op_3 };
assign sext_ln831_fu_300_p1 = { ret_V_10_reg_827[1], ret_V_10_reg_827 };
assign shl_ln1497_fu_385_p2[3:0] = trunc_ln728_fu_391_p1;
assign tmp_6_fu_199_p3 = op_0[1];
assign tmp_8_fu_621_p3 = { ret_V_25_reg_888, 1'h0 };
assign tmp_fu_358_p1 = op_6;
assign tmp_fu_358_p3 = op_6[3];
assign trunc_ln851_1_fu_227_p1 = ret_V_21_fu_211_p2[1:0];
assign trunc_ln851_2_fu_267_p1 = ret_V_23_fu_251_p2[1:0];
assign trunc_ln851_3_fu_698_p1 = op_14_V_reg_893[0];
assign trunc_ln851_fu_675_p1 = ret_V_19_fu_659_p2[1:0];
assign zext_ln1497_fu_378_p1 = { 3'h0, trunc_ln1497_fu_374_p1 };
assign zext_ln69_fu_345_p1 = { 2'h0, ret_V_24_fu_323_p3[2], ret_V_24_fu_323_p3 };
endmodule


// Machine B:
// Processed by function `add_clk_enable_signal` in `verilog_tricks.py`.
// Processed by function `remove_reset_signal` in `verilog_tricks.py`.
module top_B (
  ap_clk,
  ap_start,
  ap_done,
  ap_idle,
  ap_ready,
  op_0,
  op_3,
  op_4,
  op_6,
  op_7,
  op_12,
  op_15,
  op_16,
  op_17,
  op_18,
  op_29,
  op_29_ap_vld,
clk_enable
);
input clk_enable;


input ap_clk;
wire ap_rst;
assign ap_rst = op_29_ap_vld;
input ap_start;
input [1:0] op_0;
input [7:0] op_12;
input [7:0] op_15;
input [3:0] op_16;
input [7:0] op_17;
input [3:0] op_18;
input [3:0] op_3;
input op_4;
input [3:0] op_6;
input [15:0] op_7;
output ap_done;
output ap_idle;
output ap_ready;
output [31:0] op_29;
output op_29_ap_vld;


reg [4:0] \add_10ns_10s_10_2_1_U8.top_add_10ns_10s_10_2_1_Adder_4_U.ain_s1 ;
reg [4:0] \add_10ns_10s_10_2_1_U8.top_add_10ns_10s_10_2_1_Adder_4_U.bin_s1 ;
reg \add_10ns_10s_10_2_1_U8.top_add_10ns_10s_10_2_1_Adder_4_U.carry_s1 ;
reg [4:0] \add_10ns_10s_10_2_1_U8.top_add_10ns_10s_10_2_1_Adder_4_U.sum_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s1 ;
reg \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.carry_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.sum_s1 ;
reg [15:0] \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.ain_s1 ;
reg [15:0] \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.bin_s1 ;
reg \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.carry_s1 ;
reg [15:0] \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.sum_s1 ;
reg [15:0] \add_32ns_32s_32_2_1_U14.top_add_32ns_32s_32_2_1_Adder_8_U.ain_s1 ;
reg [15:0] \add_32ns_32s_32_2_1_U14.top_add_32ns_32s_32_2_1_Adder_8_U.bin_s1 ;
reg \add_32ns_32s_32_2_1_U14.top_add_32ns_32s_32_2_1_Adder_8_U.carry_s1 ;
reg [15:0] \add_32ns_32s_32_2_1_U14.top_add_32ns_32s_32_2_1_Adder_8_U.sum_s1 ;
reg [15:0] \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_8_U.ain_s1 ;
reg [15:0] \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_8_U.bin_s1 ;
reg \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_8_U.carry_s1 ;
reg [15:0] \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_8_U.sum_s1 ;
reg [15:0] \add_32s_32ns_32_2_1_U17.top_add_32s_32ns_32_2_1_Adder_11_U.ain_s1 ;
reg [15:0] \add_32s_32ns_32_2_1_U17.top_add_32s_32ns_32_2_1_Adder_11_U.bin_s1 ;
reg \add_32s_32ns_32_2_1_U17.top_add_32s_32ns_32_2_1_Adder_11_U.carry_s1 ;
reg [15:0] \add_32s_32ns_32_2_1_U17.top_add_32s_32ns_32_2_1_Adder_11_U.sum_s1 ;
reg [16:0] \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_6_U.ain_s1 ;
reg [16:0] \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_6_U.bin_s1 ;
reg \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_6_U.carry_s1 ;
reg [16:0] \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_6_U.sum_s1 ;
reg [1:0] \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_1_U.ain_s1 ;
reg [1:0] \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_1_U.bin_s1 ;
reg \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_1_U.carry_s1 ;
reg \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_1_U.sum_s1 ;
reg [1:0] \add_3s_3ns_3_2_1_U6.top_add_3s_3ns_3_2_1_Adder_2_U.ain_s1 ;
reg [1:0] \add_3s_3ns_3_2_1_U6.top_add_3s_3ns_3_2_1_Adder_2_U.bin_s1 ;
reg \add_3s_3ns_3_2_1_U6.top_add_3s_3ns_3_2_1_Adder_2_U.carry_s1 ;
reg \add_3s_3ns_3_2_1_U6.top_add_3s_3ns_3_2_1_Adder_2_U.sum_s1 ;
reg [2:0] \add_6ns_6s_6_2_1_U7.top_add_6ns_6s_6_2_1_Adder_3_U.ain_s1 ;
reg [2:0] \add_6ns_6s_6_2_1_U7.top_add_6ns_6s_6_2_1_Adder_3_U.bin_s1 ;
reg \add_6ns_6s_6_2_1_U7.top_add_6ns_6s_6_2_1_Adder_3_U.carry_s1 ;
reg [2:0] \add_6ns_6s_6_2_1_U7.top_add_6ns_6s_6_2_1_Adder_3_U.sum_s1 ;
reg [3:0] \add_7s_7ns_7_2_1_U9.top_add_7s_7ns_7_2_1_Adder_5_U.ain_s1 ;
reg [3:0] \add_7s_7ns_7_2_1_U9.top_add_7s_7ns_7_2_1_Adder_5_U.bin_s1 ;
reg \add_7s_7ns_7_2_1_U9.top_add_7s_7ns_7_2_1_Adder_5_U.carry_s1 ;
reg [2:0] \add_7s_7ns_7_2_1_U9.top_add_7s_7ns_7_2_1_Adder_5_U.sum_s1 ;
reg [3:0] \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_9_U.ain_s1 ;
reg [3:0] \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_9_U.bin_s1 ;
reg \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_9_U.carry_s1 ;
reg [3:0] \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_9_U.sum_s1 ;
reg [4:0] \add_9s_9s_9_2_1_U16.top_add_9s_9s_9_2_1_Adder_10_U.ain_s1 ;
reg [4:0] \add_9s_9s_9_2_1_U16.top_add_9s_9s_9_2_1_Adder_10_U.bin_s1 ;
reg \add_9s_9s_9_2_1_U16.top_add_9s_9s_9_2_1_Adder_10_U.carry_s1 ;
reg [3:0] \add_9s_9s_9_2_1_U16.top_add_9s_9s_9_2_1_Adder_10_U.sum_s1 ;
reg [31:0] add_ln691_reg_1014;
reg [8:0] add_ln69_reg_1096;
reg [26:0] ap_CS_fsm = 27'h0000001;
reg icmp_ln768_reg_934;
reg icmp_ln786_reg_939;
reg icmp_ln851_1_reg_847;
reg icmp_ln851_2_reg_859;
reg icmp_ln851_reg_1046;
reg [31:0] \lshr_32ns_32s_32_7_1_U2.din1_cast_array[0] ;
reg [31:0] \lshr_32ns_32s_32_7_1_U2.din1_cast_array[1] ;
reg [31:0] \lshr_32ns_32s_32_7_1_U2.din1_cast_array[2] ;
reg [31:0] \lshr_32ns_32s_32_7_1_U2.din1_cast_array[3] ;
reg [31:0] \lshr_32ns_32s_32_7_1_U2.din1_cast_array[4] ;
reg [31:0] \lshr_32ns_32s_32_7_1_U2.din1_cast_array[5] ;
reg [31:0] \lshr_32ns_32s_32_7_1_U2.dout_array[0] ;
reg [31:0] \lshr_32ns_32s_32_7_1_U2.dout_array[1] ;
reg [31:0] \lshr_32ns_32s_32_7_1_U2.dout_array[2] ;
reg [31:0] \lshr_32ns_32s_32_7_1_U2.dout_array[3] ;
reg [31:0] \lshr_32ns_32s_32_7_1_U2.dout_array[4] ;
reg [31:0] \lshr_32ns_32s_32_7_1_U2.dout_array[5] ;
reg [1:0] op_14_V_reg_981;
reg [5:0] op_20_V_reg_909;
reg [5:0] op_22_V_reg_966;
reg [31:0] op_25_V_reg_1051;
reg or_ln785_reg_960;
reg p_Result_4_reg_914;
reg p_Result_5_reg_927;
reg [1:0] p_Val2_s_reg_921;
reg [1:0] ret_V_10_reg_837;
reg [2:0] ret_V_11_reg_869;
reg [31:0] ret_V_16_cast_reg_1007;
reg [7:0] ret_V_20_reg_1066;
reg [4:0] ret_V_21_reg_815;
reg [2:0] ret_V_22_reg_874;
reg [3:0] ret_V_23_reg_832;
reg [2:0] ret_V_24_reg_879;
reg [6:0] ret_V_25_reg_987;
reg [33:0] ret_V_26_reg_1002;
reg [31:0] ret_V_27_reg_1019;
reg [31:0] ret_V_28_reg_1071;
reg [31:0] ret_V_29_reg_1091;
reg [7:0] ret_V_2_reg_1029;
reg [7:0] ret_V_3_reg_1056;
reg [2:0] ret_V_6_reg_820;
reg [2:0] ret_V_7_reg_864;
reg [6:0] select_ln1192_reg_955;
reg [3:0] select_ln1497_reg_904;
reg [1:0] select_ln340_reg_971;
reg [2:0] sext_ln831_reg_852;
reg [31:0] \shl_32ns_32s_32_7_1_U3.din1_cast_array[0] ;
reg [31:0] \shl_32ns_32s_32_7_1_U3.din1_cast_array[1] ;
reg [31:0] \shl_32ns_32s_32_7_1_U3.din1_cast_array[2] ;
reg [31:0] \shl_32ns_32s_32_7_1_U3.din1_cast_array[3] ;
reg [31:0] \shl_32ns_32s_32_7_1_U3.din1_cast_array[4] ;
reg [31:0] \shl_32ns_32s_32_7_1_U3.din1_cast_array[5] ;
reg [31:0] \shl_32ns_32s_32_7_1_U3.dout_array[0] ;
reg [31:0] \shl_32ns_32s_32_7_1_U3.dout_array[1] ;
reg [31:0] \shl_32ns_32s_32_7_1_U3.dout_array[2] ;
reg [31:0] \shl_32ns_32s_32_7_1_U3.dout_array[3] ;
reg [31:0] \shl_32ns_32s_32_7_1_U3.dout_array[4] ;
reg [31:0] \shl_32ns_32s_32_7_1_U3.dout_array[5] ;
reg [2:0] \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.ain_s1 ;
reg [2:0] \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.bin_s1 ;
reg \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.carry_s1 ;
reg [1:0] \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.sum_s1 ;
reg [2:0] \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_0_U.ain_s1 ;
reg [2:0] \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_0_U.bin_s1 ;
reg \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_0_U.carry_s1 ;
reg [1:0] \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_0_U.sum_s1 ;
reg [4:0] sub_ln1497_reg_778;
reg tmp_6_reg_783;
reg tmp_reg_773;
reg trunc_ln1497_reg_889;
reg [3:0] trunc_ln728_reg_894;
reg [1:0] trunc_ln851_1_reg_827;
reg [1:0] trunc_ln851_2_reg_842;
reg [1:0] trunc_ln851_reg_1036;
reg [7:0] _541_;
wire [31:0] _000_;
wire [8:0] _001_;
wire [26:0] _002_;
wire _003_;
wire _004_;
wire _005_;
wire _006_;
wire _007_;
wire [1:0] _008_;
wire [5:0] _009_;
wire [5:0] _010_;
wire [31:0] _011_;
wire _012_;
wire _013_;
wire _014_;
wire [1:0] _015_;
wire [1:0] _016_;
wire [2:0] _017_;
wire [31:0] _018_;
wire [7:0] _019_;
wire [7:0] _020_;
wire [4:0] _021_;
wire [2:0] _022_;
wire [3:0] _023_;
wire [2:0] _024_;
wire [6:0] _025_;
wire [33:0] _026_;
wire [31:0] _027_;
wire [31:0] _028_;
wire [31:0] _029_;
wire [7:0] _030_;
wire [7:0] _031_;
wire [2:0] _032_;
wire [2:0] _033_;
wire [6:0] _034_;
wire [3:0] _035_;
wire [1:0] _036_;
wire [2:0] _037_;
wire [4:0] _038_;
wire _039_;
wire _040_;
wire _041_;
wire [3:0] _042_;
wire [1:0] _043_;
wire [1:0] _044_;
wire [1:0] _045_;
wire _046_;
wire _047_;
wire _048_;
wire _049_;
wire _050_;
wire _051_;
wire _052_;
wire _053_;
wire _054_;
wire [4:0] _055_;
wire [4:0] _056_;
wire _057_;
wire [4:0] _058_;
wire [5:0] _059_;
wire [5:0] _060_;
wire [15:0] _061_;
wire [15:0] _062_;
wire _063_;
wire [15:0] _064_;
wire [16:0] _065_;
wire [16:0] _066_;
wire [15:0] _067_;
wire [15:0] _068_;
wire _069_;
wire [15:0] _070_;
wire [16:0] _071_;
wire [16:0] _072_;
wire [15:0] _073_;
wire [15:0] _074_;
wire _075_;
wire [15:0] _076_;
wire [16:0] _077_;
wire [16:0] _078_;
wire [15:0] _079_;
wire [15:0] _080_;
wire _081_;
wire [15:0] _082_;
wire [16:0] _083_;
wire [16:0] _084_;
wire [15:0] _085_;
wire [15:0] _086_;
wire _087_;
wire [15:0] _088_;
wire [16:0] _089_;
wire [16:0] _090_;
wire [16:0] _091_;
wire [16:0] _092_;
wire _093_;
wire [16:0] _094_;
wire [17:0] _095_;
wire [17:0] _096_;
wire [1:0] _097_;
wire [1:0] _098_;
wire _099_;
wire _100_;
wire [1:0] _101_;
wire [2:0] _102_;
wire [1:0] _103_;
wire [1:0] _104_;
wire _105_;
wire _106_;
wire [1:0] _107_;
wire [2:0] _108_;
wire [2:0] _109_;
wire [2:0] _110_;
wire _111_;
wire [2:0] _112_;
wire [3:0] _113_;
wire [3:0] _114_;
wire [3:0] _115_;
wire [3:0] _116_;
wire _117_;
wire [2:0] _118_;
wire [3:0] _119_;
wire [4:0] _120_;
wire [3:0] _121_;
wire [3:0] _122_;
wire _123_;
wire [3:0] _124_;
wire [4:0] _125_;
wire [4:0] _126_;
wire [4:0] _127_;
wire [4:0] _128_;
wire _129_;
wire [3:0] _130_;
wire [4:0] _131_;
wire [5:0] _132_;
wire [31:0] _133_;
wire [31:0] _134_;
wire [31:0] _135_;
wire [31:0] _136_;
wire [31:0] _137_;
wire [31:0] _138_;
wire [31:0] _139_;
wire [31:0] _140_;
wire [31:0] _141_;
wire [31:0] _142_;
wire [31:0] _143_;
wire [31:0] _144_;
wire [31:0] _145_;
wire [31:0] _146_;
wire [31:0] _147_;
wire [31:0] _148_;
wire [31:0] _149_;
wire [31:0] _150_;
wire [31:0] _151_;
wire [31:0] _152_;
wire [31:0] _153_;
wire [31:0] _154_;
wire [31:0] _155_;
wire [31:0] _156_;
wire [31:0] _157_;
wire [31:0] _158_;
wire [31:0] _159_;
wire [31:0] _160_;
wire [31:0] _161_;
wire [31:0] _162_;
wire [31:0] _163_;
wire [31:0] _164_;
wire [31:0] _165_;
wire [31:0] _166_;
wire [31:0] _167_;
wire [31:0] _168_;
wire [31:0] _169_;
wire [31:0] _170_;
wire [31:0] _171_;
wire [31:0] _172_;
wire [31:0] _173_;
wire [31:0] _174_;
wire [31:0] _175_;
wire [31:0] _176_;
wire [31:0] _177_;
wire [31:0] _178_;
wire [31:0] _179_;
wire [31:0] _180_;
wire [31:0] _181_;
wire [31:0] _182_;
wire [31:0] _183_;
wire [31:0] _184_;
wire [31:0] _185_;
wire [31:0] _186_;
wire [31:0] _187_;
wire [31:0] _188_;
wire [31:0] _189_;
wire [31:0] _190_;
wire [31:0] _191_;
wire [31:0] _192_;
wire [2:0] _193_;
wire [2:0] _194_;
wire _195_;
wire [1:0] _196_;
wire [2:0] _197_;
wire [3:0] _198_;
wire [2:0] _199_;
wire [2:0] _200_;
wire _201_;
wire [1:0] _202_;
wire [2:0] _203_;
wire [3:0] _204_;
wire _205_;
wire _206_;
wire _207_;
wire _208_;
wire _209_;
wire _210_;
wire _211_;
wire _212_;
wire _213_;
wire _214_;
wire _215_;
wire _216_;
wire _217_;
wire _218_;
wire _219_;
wire _220_;
wire _221_;
wire _222_;
wire _223_;
wire _224_;
wire _225_;
wire _226_;
wire _227_;
wire _228_;
wire _229_;
wire _230_;
wire _231_;
wire _232_;
wire _233_;
wire \add_10ns_10s_10_2_1_U8.ce ;
wire \add_10ns_10s_10_2_1_U8.clk ;
wire [9:0] \add_10ns_10s_10_2_1_U8.din0 ;
wire [9:0] \add_10ns_10s_10_2_1_U8.din1 ;
wire [9:0] \add_10ns_10s_10_2_1_U8.dout ;
wire \add_10ns_10s_10_2_1_U8.reset ;
wire [9:0] \add_10ns_10s_10_2_1_U8.top_add_10ns_10s_10_2_1_Adder_4_U.a ;
wire [9:0] \add_10ns_10s_10_2_1_U8.top_add_10ns_10s_10_2_1_Adder_4_U.ain_s0 ;
wire [9:0] \add_10ns_10s_10_2_1_U8.top_add_10ns_10s_10_2_1_Adder_4_U.b ;
wire [9:0] \add_10ns_10s_10_2_1_U8.top_add_10ns_10s_10_2_1_Adder_4_U.bin_s0 ;
wire \add_10ns_10s_10_2_1_U8.top_add_10ns_10s_10_2_1_Adder_4_U.ce ;
wire \add_10ns_10s_10_2_1_U8.top_add_10ns_10s_10_2_1_Adder_4_U.clk ;
wire \add_10ns_10s_10_2_1_U8.top_add_10ns_10s_10_2_1_Adder_4_U.facout_s1 ;
wire \add_10ns_10s_10_2_1_U8.top_add_10ns_10s_10_2_1_Adder_4_U.facout_s2 ;
wire [4:0] \add_10ns_10s_10_2_1_U8.top_add_10ns_10s_10_2_1_Adder_4_U.fas_s1 ;
wire [4:0] \add_10ns_10s_10_2_1_U8.top_add_10ns_10s_10_2_1_Adder_4_U.fas_s2 ;
wire \add_10ns_10s_10_2_1_U8.top_add_10ns_10s_10_2_1_Adder_4_U.reset ;
wire [9:0] \add_10ns_10s_10_2_1_U8.top_add_10ns_10s_10_2_1_Adder_4_U.s ;
wire [4:0] \add_10ns_10s_10_2_1_U8.top_add_10ns_10s_10_2_1_Adder_4_U.u1.a ;
wire [4:0] \add_10ns_10s_10_2_1_U8.top_add_10ns_10s_10_2_1_Adder_4_U.u1.b ;
wire \add_10ns_10s_10_2_1_U8.top_add_10ns_10s_10_2_1_Adder_4_U.u1.cin ;
wire \add_10ns_10s_10_2_1_U8.top_add_10ns_10s_10_2_1_Adder_4_U.u1.cout ;
wire [4:0] \add_10ns_10s_10_2_1_U8.top_add_10ns_10s_10_2_1_Adder_4_U.u1.s ;
wire [4:0] \add_10ns_10s_10_2_1_U8.top_add_10ns_10s_10_2_1_Adder_4_U.u2.a ;
wire [4:0] \add_10ns_10s_10_2_1_U8.top_add_10ns_10s_10_2_1_Adder_4_U.u2.b ;
wire \add_10ns_10s_10_2_1_U8.top_add_10ns_10s_10_2_1_Adder_4_U.u2.cin ;
wire \add_10ns_10s_10_2_1_U8.top_add_10ns_10s_10_2_1_Adder_4_U.u2.cout ;
wire [4:0] \add_10ns_10s_10_2_1_U8.top_add_10ns_10s_10_2_1_Adder_4_U.u2.s ;
wire \add_32ns_32ns_32_2_1_U11.ce ;
wire \add_32ns_32ns_32_2_1_U11.clk ;
wire [31:0] \add_32ns_32ns_32_2_1_U11.din0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U11.din1 ;
wire [31:0] \add_32ns_32ns_32_2_1_U11.dout ;
wire \add_32ns_32ns_32_2_1_U11.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.a ;
wire [31:0] \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.b ;
wire [31:0] \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s0 ;
wire \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.ce ;
wire \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.clk ;
wire \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.facout_s1 ;
wire \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.facout_s2 ;
wire [15:0] \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s1 ;
wire [15:0] \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s2 ;
wire \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.b ;
wire \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cin ;
wire \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.b ;
wire \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cin ;
wire \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.s ;
wire \add_32ns_32s_32_2_1_U12.ce ;
wire \add_32ns_32s_32_2_1_U12.clk ;
wire [31:0] \add_32ns_32s_32_2_1_U12.din0 ;
wire [31:0] \add_32ns_32s_32_2_1_U12.din1 ;
wire [31:0] \add_32ns_32s_32_2_1_U12.dout ;
wire \add_32ns_32s_32_2_1_U12.reset ;
wire [31:0] \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.a ;
wire [31:0] \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.ain_s0 ;
wire [31:0] \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.b ;
wire [31:0] \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.bin_s0 ;
wire \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.ce ;
wire \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.clk ;
wire \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.facout_s1 ;
wire \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.facout_s2 ;
wire [15:0] \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.fas_s1 ;
wire [15:0] \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.fas_s2 ;
wire \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.reset ;
wire [31:0] \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.s ;
wire [15:0] \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.u1.a ;
wire [15:0] \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.u1.b ;
wire \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.u1.cin ;
wire \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.u1.cout ;
wire [15:0] \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.u1.s ;
wire [15:0] \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.u2.a ;
wire [15:0] \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.u2.b ;
wire \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.u2.cin ;
wire \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.u2.cout ;
wire [15:0] \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.u2.s ;
wire \add_32ns_32s_32_2_1_U14.ce ;
wire \add_32ns_32s_32_2_1_U14.clk ;
wire [31:0] \add_32ns_32s_32_2_1_U14.din0 ;
wire [31:0] \add_32ns_32s_32_2_1_U14.din1 ;
wire [31:0] \add_32ns_32s_32_2_1_U14.dout ;
wire \add_32ns_32s_32_2_1_U14.reset ;
wire [31:0] \add_32ns_32s_32_2_1_U14.top_add_32ns_32s_32_2_1_Adder_8_U.a ;
wire [31:0] \add_32ns_32s_32_2_1_U14.top_add_32ns_32s_32_2_1_Adder_8_U.ain_s0 ;
wire [31:0] \add_32ns_32s_32_2_1_U14.top_add_32ns_32s_32_2_1_Adder_8_U.b ;
wire [31:0] \add_32ns_32s_32_2_1_U14.top_add_32ns_32s_32_2_1_Adder_8_U.bin_s0 ;
wire \add_32ns_32s_32_2_1_U14.top_add_32ns_32s_32_2_1_Adder_8_U.ce ;
wire \add_32ns_32s_32_2_1_U14.top_add_32ns_32s_32_2_1_Adder_8_U.clk ;
wire \add_32ns_32s_32_2_1_U14.top_add_32ns_32s_32_2_1_Adder_8_U.facout_s1 ;
wire \add_32ns_32s_32_2_1_U14.top_add_32ns_32s_32_2_1_Adder_8_U.facout_s2 ;
wire [15:0] \add_32ns_32s_32_2_1_U14.top_add_32ns_32s_32_2_1_Adder_8_U.fas_s1 ;
wire [15:0] \add_32ns_32s_32_2_1_U14.top_add_32ns_32s_32_2_1_Adder_8_U.fas_s2 ;
wire \add_32ns_32s_32_2_1_U14.top_add_32ns_32s_32_2_1_Adder_8_U.reset ;
wire [31:0] \add_32ns_32s_32_2_1_U14.top_add_32ns_32s_32_2_1_Adder_8_U.s ;
wire [15:0] \add_32ns_32s_32_2_1_U14.top_add_32ns_32s_32_2_1_Adder_8_U.u1.a ;
wire [15:0] \add_32ns_32s_32_2_1_U14.top_add_32ns_32s_32_2_1_Adder_8_U.u1.b ;
wire \add_32ns_32s_32_2_1_U14.top_add_32ns_32s_32_2_1_Adder_8_U.u1.cin ;
wire \add_32ns_32s_32_2_1_U14.top_add_32ns_32s_32_2_1_Adder_8_U.u1.cout ;
wire [15:0] \add_32ns_32s_32_2_1_U14.top_add_32ns_32s_32_2_1_Adder_8_U.u1.s ;
wire [15:0] \add_32ns_32s_32_2_1_U14.top_add_32ns_32s_32_2_1_Adder_8_U.u2.a ;
wire [15:0] \add_32ns_32s_32_2_1_U14.top_add_32ns_32s_32_2_1_Adder_8_U.u2.b ;
wire \add_32ns_32s_32_2_1_U14.top_add_32ns_32s_32_2_1_Adder_8_U.u2.cin ;
wire \add_32ns_32s_32_2_1_U14.top_add_32ns_32s_32_2_1_Adder_8_U.u2.cout ;
wire [15:0] \add_32ns_32s_32_2_1_U14.top_add_32ns_32s_32_2_1_Adder_8_U.u2.s ;
wire \add_32ns_32s_32_2_1_U15.ce ;
wire \add_32ns_32s_32_2_1_U15.clk ;
wire [31:0] \add_32ns_32s_32_2_1_U15.din0 ;
wire [31:0] \add_32ns_32s_32_2_1_U15.din1 ;
wire [31:0] \add_32ns_32s_32_2_1_U15.dout ;
wire \add_32ns_32s_32_2_1_U15.reset ;
wire [31:0] \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_8_U.a ;
wire [31:0] \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_8_U.ain_s0 ;
wire [31:0] \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_8_U.b ;
wire [31:0] \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_8_U.bin_s0 ;
wire \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_8_U.ce ;
wire \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_8_U.clk ;
wire \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_8_U.facout_s1 ;
wire \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_8_U.facout_s2 ;
wire [15:0] \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_8_U.fas_s1 ;
wire [15:0] \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_8_U.fas_s2 ;
wire \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_8_U.reset ;
wire [31:0] \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_8_U.s ;
wire [15:0] \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_8_U.u1.a ;
wire [15:0] \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_8_U.u1.b ;
wire \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_8_U.u1.cin ;
wire \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_8_U.u1.cout ;
wire [15:0] \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_8_U.u1.s ;
wire [15:0] \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_8_U.u2.a ;
wire [15:0] \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_8_U.u2.b ;
wire \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_8_U.u2.cin ;
wire \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_8_U.u2.cout ;
wire [15:0] \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_8_U.u2.s ;
wire \add_32s_32ns_32_2_1_U17.ce ;
wire \add_32s_32ns_32_2_1_U17.clk ;
wire [31:0] \add_32s_32ns_32_2_1_U17.din0 ;
wire [31:0] \add_32s_32ns_32_2_1_U17.din1 ;
wire [31:0] \add_32s_32ns_32_2_1_U17.dout ;
wire \add_32s_32ns_32_2_1_U17.reset ;
wire [31:0] \add_32s_32ns_32_2_1_U17.top_add_32s_32ns_32_2_1_Adder_11_U.a ;
wire [31:0] \add_32s_32ns_32_2_1_U17.top_add_32s_32ns_32_2_1_Adder_11_U.ain_s0 ;
wire [31:0] \add_32s_32ns_32_2_1_U17.top_add_32s_32ns_32_2_1_Adder_11_U.b ;
wire [31:0] \add_32s_32ns_32_2_1_U17.top_add_32s_32ns_32_2_1_Adder_11_U.bin_s0 ;
wire \add_32s_32ns_32_2_1_U17.top_add_32s_32ns_32_2_1_Adder_11_U.ce ;
wire \add_32s_32ns_32_2_1_U17.top_add_32s_32ns_32_2_1_Adder_11_U.clk ;
wire \add_32s_32ns_32_2_1_U17.top_add_32s_32ns_32_2_1_Adder_11_U.facout_s1 ;
wire \add_32s_32ns_32_2_1_U17.top_add_32s_32ns_32_2_1_Adder_11_U.facout_s2 ;
wire [15:0] \add_32s_32ns_32_2_1_U17.top_add_32s_32ns_32_2_1_Adder_11_U.fas_s1 ;
wire [15:0] \add_32s_32ns_32_2_1_U17.top_add_32s_32ns_32_2_1_Adder_11_U.fas_s2 ;
wire \add_32s_32ns_32_2_1_U17.top_add_32s_32ns_32_2_1_Adder_11_U.reset ;
wire [31:0] \add_32s_32ns_32_2_1_U17.top_add_32s_32ns_32_2_1_Adder_11_U.s ;
wire [15:0] \add_32s_32ns_32_2_1_U17.top_add_32s_32ns_32_2_1_Adder_11_U.u1.a ;
wire [15:0] \add_32s_32ns_32_2_1_U17.top_add_32s_32ns_32_2_1_Adder_11_U.u1.b ;
wire \add_32s_32ns_32_2_1_U17.top_add_32s_32ns_32_2_1_Adder_11_U.u1.cin ;
wire \add_32s_32ns_32_2_1_U17.top_add_32s_32ns_32_2_1_Adder_11_U.u1.cout ;
wire [15:0] \add_32s_32ns_32_2_1_U17.top_add_32s_32ns_32_2_1_Adder_11_U.u1.s ;
wire [15:0] \add_32s_32ns_32_2_1_U17.top_add_32s_32ns_32_2_1_Adder_11_U.u2.a ;
wire [15:0] \add_32s_32ns_32_2_1_U17.top_add_32s_32ns_32_2_1_Adder_11_U.u2.b ;
wire \add_32s_32ns_32_2_1_U17.top_add_32s_32ns_32_2_1_Adder_11_U.u2.cin ;
wire \add_32s_32ns_32_2_1_U17.top_add_32s_32ns_32_2_1_Adder_11_U.u2.cout ;
wire [15:0] \add_32s_32ns_32_2_1_U17.top_add_32s_32ns_32_2_1_Adder_11_U.u2.s ;
wire \add_34s_34s_34_2_1_U10.ce ;
wire \add_34s_34s_34_2_1_U10.clk ;
wire [33:0] \add_34s_34s_34_2_1_U10.din0 ;
wire [33:0] \add_34s_34s_34_2_1_U10.din1 ;
wire [33:0] \add_34s_34s_34_2_1_U10.dout ;
wire \add_34s_34s_34_2_1_U10.reset ;
wire [33:0] \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_6_U.a ;
wire [33:0] \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_6_U.ain_s0 ;
wire [33:0] \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_6_U.b ;
wire [33:0] \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_6_U.bin_s0 ;
wire \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_6_U.ce ;
wire \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_6_U.clk ;
wire \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_6_U.facout_s1 ;
wire \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_6_U.facout_s2 ;
wire [16:0] \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_6_U.fas_s1 ;
wire [16:0] \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_6_U.fas_s2 ;
wire \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_6_U.reset ;
wire [33:0] \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_6_U.s ;
wire [16:0] \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_6_U.u1.a ;
wire [16:0] \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_6_U.u1.b ;
wire \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_6_U.u1.cin ;
wire \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_6_U.u1.cout ;
wire [16:0] \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_6_U.u1.s ;
wire [16:0] \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_6_U.u2.a ;
wire [16:0] \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_6_U.u2.b ;
wire \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_6_U.u2.cin ;
wire \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_6_U.u2.cout ;
wire [16:0] \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_6_U.u2.s ;
wire \add_3ns_3ns_3_2_1_U5.ce ;
wire \add_3ns_3ns_3_2_1_U5.clk ;
wire [2:0] \add_3ns_3ns_3_2_1_U5.din0 ;
wire [2:0] \add_3ns_3ns_3_2_1_U5.din1 ;
wire [2:0] \add_3ns_3ns_3_2_1_U5.dout ;
wire \add_3ns_3ns_3_2_1_U5.reset ;
wire [2:0] \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_1_U.a ;
wire [2:0] \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_1_U.ain_s0 ;
wire [2:0] \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_1_U.b ;
wire [2:0] \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_1_U.bin_s0 ;
wire \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_1_U.ce ;
wire \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_1_U.clk ;
wire \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_1_U.facout_s1 ;
wire \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_1_U.facout_s2 ;
wire \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_1_U.fas_s1 ;
wire [1:0] \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_1_U.fas_s2 ;
wire \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_1_U.reset ;
wire [2:0] \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_1_U.s ;
wire \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_1_U.u1.a ;
wire \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_1_U.u1.b ;
wire \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_1_U.u1.cin ;
wire \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_1_U.u1.cout ;
wire \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_1_U.u1.s ;
wire [1:0] \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_1_U.u2.a ;
wire [1:0] \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_1_U.u2.b ;
wire \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_1_U.u2.cin ;
wire \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_1_U.u2.cout ;
wire [1:0] \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_1_U.u2.s ;
wire \add_3s_3ns_3_2_1_U6.ce ;
wire \add_3s_3ns_3_2_1_U6.clk ;
wire [2:0] \add_3s_3ns_3_2_1_U6.din0 ;
wire [2:0] \add_3s_3ns_3_2_1_U6.din1 ;
wire [2:0] \add_3s_3ns_3_2_1_U6.dout ;
wire \add_3s_3ns_3_2_1_U6.reset ;
wire [2:0] \add_3s_3ns_3_2_1_U6.top_add_3s_3ns_3_2_1_Adder_2_U.a ;
wire [2:0] \add_3s_3ns_3_2_1_U6.top_add_3s_3ns_3_2_1_Adder_2_U.ain_s0 ;
wire [2:0] \add_3s_3ns_3_2_1_U6.top_add_3s_3ns_3_2_1_Adder_2_U.b ;
wire [2:0] \add_3s_3ns_3_2_1_U6.top_add_3s_3ns_3_2_1_Adder_2_U.bin_s0 ;
wire \add_3s_3ns_3_2_1_U6.top_add_3s_3ns_3_2_1_Adder_2_U.ce ;
wire \add_3s_3ns_3_2_1_U6.top_add_3s_3ns_3_2_1_Adder_2_U.clk ;
wire \add_3s_3ns_3_2_1_U6.top_add_3s_3ns_3_2_1_Adder_2_U.facout_s1 ;
wire \add_3s_3ns_3_2_1_U6.top_add_3s_3ns_3_2_1_Adder_2_U.facout_s2 ;
wire \add_3s_3ns_3_2_1_U6.top_add_3s_3ns_3_2_1_Adder_2_U.fas_s1 ;
wire [1:0] \add_3s_3ns_3_2_1_U6.top_add_3s_3ns_3_2_1_Adder_2_U.fas_s2 ;
wire \add_3s_3ns_3_2_1_U6.top_add_3s_3ns_3_2_1_Adder_2_U.reset ;
wire [2:0] \add_3s_3ns_3_2_1_U6.top_add_3s_3ns_3_2_1_Adder_2_U.s ;
wire \add_3s_3ns_3_2_1_U6.top_add_3s_3ns_3_2_1_Adder_2_U.u1.a ;
wire \add_3s_3ns_3_2_1_U6.top_add_3s_3ns_3_2_1_Adder_2_U.u1.b ;
wire \add_3s_3ns_3_2_1_U6.top_add_3s_3ns_3_2_1_Adder_2_U.u1.cin ;
wire \add_3s_3ns_3_2_1_U6.top_add_3s_3ns_3_2_1_Adder_2_U.u1.cout ;
wire \add_3s_3ns_3_2_1_U6.top_add_3s_3ns_3_2_1_Adder_2_U.u1.s ;
wire [1:0] \add_3s_3ns_3_2_1_U6.top_add_3s_3ns_3_2_1_Adder_2_U.u2.a ;
wire [1:0] \add_3s_3ns_3_2_1_U6.top_add_3s_3ns_3_2_1_Adder_2_U.u2.b ;
wire \add_3s_3ns_3_2_1_U6.top_add_3s_3ns_3_2_1_Adder_2_U.u2.cin ;
wire \add_3s_3ns_3_2_1_U6.top_add_3s_3ns_3_2_1_Adder_2_U.u2.cout ;
wire [1:0] \add_3s_3ns_3_2_1_U6.top_add_3s_3ns_3_2_1_Adder_2_U.u2.s ;
wire \add_6ns_6s_6_2_1_U7.ce ;
wire \add_6ns_6s_6_2_1_U7.clk ;
wire [5:0] \add_6ns_6s_6_2_1_U7.din0 ;
wire [5:0] \add_6ns_6s_6_2_1_U7.din1 ;
wire [5:0] \add_6ns_6s_6_2_1_U7.dout ;
wire \add_6ns_6s_6_2_1_U7.reset ;
wire [5:0] \add_6ns_6s_6_2_1_U7.top_add_6ns_6s_6_2_1_Adder_3_U.a ;
wire [5:0] \add_6ns_6s_6_2_1_U7.top_add_6ns_6s_6_2_1_Adder_3_U.ain_s0 ;
wire [5:0] \add_6ns_6s_6_2_1_U7.top_add_6ns_6s_6_2_1_Adder_3_U.b ;
wire [5:0] \add_6ns_6s_6_2_1_U7.top_add_6ns_6s_6_2_1_Adder_3_U.bin_s0 ;
wire \add_6ns_6s_6_2_1_U7.top_add_6ns_6s_6_2_1_Adder_3_U.ce ;
wire \add_6ns_6s_6_2_1_U7.top_add_6ns_6s_6_2_1_Adder_3_U.clk ;
wire \add_6ns_6s_6_2_1_U7.top_add_6ns_6s_6_2_1_Adder_3_U.facout_s1 ;
wire \add_6ns_6s_6_2_1_U7.top_add_6ns_6s_6_2_1_Adder_3_U.facout_s2 ;
wire [2:0] \add_6ns_6s_6_2_1_U7.top_add_6ns_6s_6_2_1_Adder_3_U.fas_s1 ;
wire [2:0] \add_6ns_6s_6_2_1_U7.top_add_6ns_6s_6_2_1_Adder_3_U.fas_s2 ;
wire \add_6ns_6s_6_2_1_U7.top_add_6ns_6s_6_2_1_Adder_3_U.reset ;
wire [5:0] \add_6ns_6s_6_2_1_U7.top_add_6ns_6s_6_2_1_Adder_3_U.s ;
wire [2:0] \add_6ns_6s_6_2_1_U7.top_add_6ns_6s_6_2_1_Adder_3_U.u1.a ;
wire [2:0] \add_6ns_6s_6_2_1_U7.top_add_6ns_6s_6_2_1_Adder_3_U.u1.b ;
wire \add_6ns_6s_6_2_1_U7.top_add_6ns_6s_6_2_1_Adder_3_U.u1.cin ;
wire \add_6ns_6s_6_2_1_U7.top_add_6ns_6s_6_2_1_Adder_3_U.u1.cout ;
wire [2:0] \add_6ns_6s_6_2_1_U7.top_add_6ns_6s_6_2_1_Adder_3_U.u1.s ;
wire [2:0] \add_6ns_6s_6_2_1_U7.top_add_6ns_6s_6_2_1_Adder_3_U.u2.a ;
wire [2:0] \add_6ns_6s_6_2_1_U7.top_add_6ns_6s_6_2_1_Adder_3_U.u2.b ;
wire \add_6ns_6s_6_2_1_U7.top_add_6ns_6s_6_2_1_Adder_3_U.u2.cin ;
wire \add_6ns_6s_6_2_1_U7.top_add_6ns_6s_6_2_1_Adder_3_U.u2.cout ;
wire [2:0] \add_6ns_6s_6_2_1_U7.top_add_6ns_6s_6_2_1_Adder_3_U.u2.s ;
wire \add_7s_7ns_7_2_1_U9.ce ;
wire \add_7s_7ns_7_2_1_U9.clk ;
wire [6:0] \add_7s_7ns_7_2_1_U9.din0 ;
wire [6:0] \add_7s_7ns_7_2_1_U9.din1 ;
wire [6:0] \add_7s_7ns_7_2_1_U9.dout ;
wire \add_7s_7ns_7_2_1_U9.reset ;
wire [6:0] \add_7s_7ns_7_2_1_U9.top_add_7s_7ns_7_2_1_Adder_5_U.a ;
wire [6:0] \add_7s_7ns_7_2_1_U9.top_add_7s_7ns_7_2_1_Adder_5_U.ain_s0 ;
wire [6:0] \add_7s_7ns_7_2_1_U9.top_add_7s_7ns_7_2_1_Adder_5_U.b ;
wire [6:0] \add_7s_7ns_7_2_1_U9.top_add_7s_7ns_7_2_1_Adder_5_U.bin_s0 ;
wire \add_7s_7ns_7_2_1_U9.top_add_7s_7ns_7_2_1_Adder_5_U.ce ;
wire \add_7s_7ns_7_2_1_U9.top_add_7s_7ns_7_2_1_Adder_5_U.clk ;
wire \add_7s_7ns_7_2_1_U9.top_add_7s_7ns_7_2_1_Adder_5_U.facout_s1 ;
wire \add_7s_7ns_7_2_1_U9.top_add_7s_7ns_7_2_1_Adder_5_U.facout_s2 ;
wire [2:0] \add_7s_7ns_7_2_1_U9.top_add_7s_7ns_7_2_1_Adder_5_U.fas_s1 ;
wire [3:0] \add_7s_7ns_7_2_1_U9.top_add_7s_7ns_7_2_1_Adder_5_U.fas_s2 ;
wire \add_7s_7ns_7_2_1_U9.top_add_7s_7ns_7_2_1_Adder_5_U.reset ;
wire [6:0] \add_7s_7ns_7_2_1_U9.top_add_7s_7ns_7_2_1_Adder_5_U.s ;
wire [2:0] \add_7s_7ns_7_2_1_U9.top_add_7s_7ns_7_2_1_Adder_5_U.u1.a ;
wire [2:0] \add_7s_7ns_7_2_1_U9.top_add_7s_7ns_7_2_1_Adder_5_U.u1.b ;
wire \add_7s_7ns_7_2_1_U9.top_add_7s_7ns_7_2_1_Adder_5_U.u1.cin ;
wire \add_7s_7ns_7_2_1_U9.top_add_7s_7ns_7_2_1_Adder_5_U.u1.cout ;
wire [2:0] \add_7s_7ns_7_2_1_U9.top_add_7s_7ns_7_2_1_Adder_5_U.u1.s ;
wire [3:0] \add_7s_7ns_7_2_1_U9.top_add_7s_7ns_7_2_1_Adder_5_U.u2.a ;
wire [3:0] \add_7s_7ns_7_2_1_U9.top_add_7s_7ns_7_2_1_Adder_5_U.u2.b ;
wire \add_7s_7ns_7_2_1_U9.top_add_7s_7ns_7_2_1_Adder_5_U.u2.cin ;
wire \add_7s_7ns_7_2_1_U9.top_add_7s_7ns_7_2_1_Adder_5_U.u2.cout ;
wire [3:0] \add_7s_7ns_7_2_1_U9.top_add_7s_7ns_7_2_1_Adder_5_U.u2.s ;
wire \add_8ns_8ns_8_2_1_U13.ce ;
wire \add_8ns_8ns_8_2_1_U13.clk ;
wire [7:0] \add_8ns_8ns_8_2_1_U13.din0 ;
wire [7:0] \add_8ns_8ns_8_2_1_U13.din1 ;
wire [7:0] \add_8ns_8ns_8_2_1_U13.dout ;
wire \add_8ns_8ns_8_2_1_U13.reset ;
wire [7:0] \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_9_U.a ;
wire [7:0] \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_9_U.ain_s0 ;
wire [7:0] \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_9_U.b ;
wire [7:0] \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_9_U.bin_s0 ;
wire \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_9_U.ce ;
wire \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_9_U.clk ;
wire \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_9_U.facout_s1 ;
wire \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_9_U.facout_s2 ;
wire [3:0] \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_9_U.fas_s1 ;
wire [3:0] \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_9_U.fas_s2 ;
wire \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_9_U.reset ;
wire [7:0] \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_9_U.s ;
wire [3:0] \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_9_U.u1.a ;
wire [3:0] \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_9_U.u1.b ;
wire \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_9_U.u1.cin ;
wire \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_9_U.u1.cout ;
wire [3:0] \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_9_U.u1.s ;
wire [3:0] \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_9_U.u2.a ;
wire [3:0] \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_9_U.u2.b ;
wire \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_9_U.u2.cin ;
wire \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_9_U.u2.cout ;
wire [3:0] \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_9_U.u2.s ;
wire \add_9s_9s_9_2_1_U16.ce ;
wire \add_9s_9s_9_2_1_U16.clk ;
wire [8:0] \add_9s_9s_9_2_1_U16.din0 ;
wire [8:0] \add_9s_9s_9_2_1_U16.din1 ;
wire [8:0] \add_9s_9s_9_2_1_U16.dout ;
wire \add_9s_9s_9_2_1_U16.reset ;
wire [8:0] \add_9s_9s_9_2_1_U16.top_add_9s_9s_9_2_1_Adder_10_U.a ;
wire [8:0] \add_9s_9s_9_2_1_U16.top_add_9s_9s_9_2_1_Adder_10_U.ain_s0 ;
wire [8:0] \add_9s_9s_9_2_1_U16.top_add_9s_9s_9_2_1_Adder_10_U.b ;
wire [8:0] \add_9s_9s_9_2_1_U16.top_add_9s_9s_9_2_1_Adder_10_U.bin_s0 ;
wire \add_9s_9s_9_2_1_U16.top_add_9s_9s_9_2_1_Adder_10_U.ce ;
wire \add_9s_9s_9_2_1_U16.top_add_9s_9s_9_2_1_Adder_10_U.clk ;
wire \add_9s_9s_9_2_1_U16.top_add_9s_9s_9_2_1_Adder_10_U.facout_s1 ;
wire \add_9s_9s_9_2_1_U16.top_add_9s_9s_9_2_1_Adder_10_U.facout_s2 ;
wire [3:0] \add_9s_9s_9_2_1_U16.top_add_9s_9s_9_2_1_Adder_10_U.fas_s1 ;
wire [4:0] \add_9s_9s_9_2_1_U16.top_add_9s_9s_9_2_1_Adder_10_U.fas_s2 ;
wire \add_9s_9s_9_2_1_U16.top_add_9s_9s_9_2_1_Adder_10_U.reset ;
wire [8:0] \add_9s_9s_9_2_1_U16.top_add_9s_9s_9_2_1_Adder_10_U.s ;
wire [3:0] \add_9s_9s_9_2_1_U16.top_add_9s_9s_9_2_1_Adder_10_U.u1.a ;
wire [3:0] \add_9s_9s_9_2_1_U16.top_add_9s_9s_9_2_1_Adder_10_U.u1.b ;
wire \add_9s_9s_9_2_1_U16.top_add_9s_9s_9_2_1_Adder_10_U.u1.cin ;
wire \add_9s_9s_9_2_1_U16.top_add_9s_9s_9_2_1_Adder_10_U.u1.cout ;
wire [3:0] \add_9s_9s_9_2_1_U16.top_add_9s_9s_9_2_1_Adder_10_U.u1.s ;
wire [4:0] \add_9s_9s_9_2_1_U16.top_add_9s_9s_9_2_1_Adder_10_U.u2.a ;
wire [4:0] \add_9s_9s_9_2_1_U16.top_add_9s_9s_9_2_1_Adder_10_U.u2.b ;
wire \add_9s_9s_9_2_1_U16.top_add_9s_9s_9_2_1_Adder_10_U.u2.cin ;
wire \add_9s_9s_9_2_1_U16.top_add_9s_9s_9_2_1_Adder_10_U.u2.cout ;
wire [4:0] \add_9s_9s_9_2_1_U16.top_add_9s_9s_9_2_1_Adder_10_U.u2.s ;
wire and_ln340_fu_543_p2;
wire and_ln785_1_fu_585_p2;
wire and_ln785_fu_579_p2;
wire ap_CS_fsm_state1;
wire ap_CS_fsm_state10;
wire ap_CS_fsm_state11;
wire ap_CS_fsm_state12;
wire ap_CS_fsm_state13;
wire ap_CS_fsm_state14;
wire ap_CS_fsm_state15;
wire ap_CS_fsm_state16;
wire ap_CS_fsm_state17;
wire ap_CS_fsm_state18;
wire ap_CS_fsm_state19;
wire ap_CS_fsm_state2;
wire ap_CS_fsm_state20;
wire ap_CS_fsm_state21;
wire ap_CS_fsm_state22;
wire ap_CS_fsm_state23;
wire ap_CS_fsm_state24;
wire ap_CS_fsm_state25;
wire ap_CS_fsm_state26;
wire ap_CS_fsm_state27;
wire ap_CS_fsm_state3;
wire ap_CS_fsm_state4;
wire ap_CS_fsm_state5;
wire ap_CS_fsm_state6;
wire ap_CS_fsm_state7;
wire ap_CS_fsm_state8;
wire ap_CS_fsm_state9;
wire [26:0] ap_NS_fsm;
wire ap_clk;
wire ap_done;
wire ap_idle;
wire ap_ready;
wire ap_rst;
wire ap_start;
wire [31:0] conv_i2826_fu_228_p1;
wire [6:0] empty_fu_392_p1;
wire [4:0] grp_fu_211_p1;
wire [4:0] grp_fu_211_p2;
wire [31:0] grp_fu_232_p1;
wire [31:0] grp_fu_232_p2;
wire [31:0] grp_fu_241_p1;
wire [31:0] grp_fu_241_p2;
wire [4:0] grp_fu_251_p1;
wire [4:0] grp_fu_251_p2;
wire [2:0] grp_fu_302_p2;
wire [2:0] grp_fu_315_p0;
wire [2:0] grp_fu_315_p2;
wire [5:0] grp_fu_377_p0;
wire [5:0] grp_fu_377_p1;
wire [5:0] grp_fu_377_p2;
wire [9:0] grp_fu_484_p0;
wire [9:0] grp_fu_484_p1;
wire [9:0] grp_fu_484_p2;
wire [6:0] grp_fu_559_p0;
wire [6:0] grp_fu_559_p2;
wire [33:0] grp_fu_610_p0;
wire [33:0] grp_fu_610_p1;
wire [33:0] grp_fu_610_p2;
wire [31:0] grp_fu_626_p2;
wire [31:0] grp_fu_689_p1;
wire [31:0] grp_fu_689_p2;
wire [7:0] grp_fu_699_p2;
wire [31:0] grp_fu_708_p1;
wire [31:0] grp_fu_708_p2;
wire [31:0] grp_fu_739_p1;
wire [31:0] grp_fu_739_p2;
wire [8:0] grp_fu_748_p0;
wire [8:0] grp_fu_748_p1;
wire [8:0] grp_fu_748_p2;
wire [31:0] grp_fu_757_p0;
wire [31:0] grp_fu_757_p2;
wire icmp_ln768_fu_454_p2;
wire icmp_ln786_fu_460_p2;
wire icmp_ln851_1_fu_297_p2;
wire icmp_ln851_2_fu_310_p2;
wire icmp_ln851_fu_694_p2;
wire lhs_fu_396_p0;
wire [6:0] lhs_fu_396_p3;
wire \lshr_32ns_32s_32_7_1_U2.ce ;
wire \lshr_32ns_32s_32_7_1_U2.clk ;
wire [31:0] \lshr_32ns_32s_32_7_1_U2.din0 ;
wire [31:0] \lshr_32ns_32s_32_7_1_U2.din1 ;
wire [31:0] \lshr_32ns_32s_32_7_1_U2.din1_cast ;
wire [31:0] \lshr_32ns_32s_32_7_1_U2.din1_mask ;
wire [31:0] \lshr_32ns_32s_32_7_1_U2.dout ;
wire \lshr_32ns_32s_32_7_1_U2.reset ;
wire [1:0] op_0;
wire [7:0] op_11_V_fu_466_p3;
wire [7:0] op_12;
wire op_13_V_fu_410_p3;
wire [1:0] op_14_V_fu_590_p3;
wire [7:0] op_15;
wire [3:0] op_16;
wire [7:0] op_17;
wire [3:0] op_18;
wire [31:0] op_29;
wire op_29_ap_vld;
wire [3:0] op_3;
wire op_4;
wire [3:0] op_6;
wire [15:0] op_7;
wire or_ln340_fu_532_p2;
wire or_ln785_1_fu_574_p2;
wire or_ln785_fu_498_p2;
wire or_ln786_fu_527_p2;
wire overflow_fu_517_p2;
wire p_Result_1_fu_321_p3;
wire p_Result_2_fu_340_p3;
wire p_Result_3_fu_631_p3;
wire p_Result_s_14_fu_713_p3;
wire [8:0] p_Result_s_fu_444_p4;
wire [9:0] ret_V_19_fu_665_p2;
wire [9:0] ret_V_19_reg_1024;
wire [7:0] ret_V_20_fu_725_p3;
wire [2:0] ret_V_22_fu_333_p3;
wire [3:0] ret_V_23_fu_278_p1;
wire [3:0] ret_V_23_fu_278_p2;
wire [2:0] ret_V_24_fu_352_p3;
wire [31:0] ret_V_27_fu_647_p3;
wire [6:0] ret_V_fu_404_p2;
wire [9:0] rhs_fu_657_p3;
wire [6:0] select_ln1192_fu_490_p3;
wire [2:0] select_ln1196_fu_271_p3;
wire [3:0] select_ln1497_fu_386_p3;
wire [1:0] select_ln340_fu_549_p3;
wire [2:0] select_ln850_1_fu_328_p3;
wire [2:0] select_ln850_2_fu_347_p3;
wire [31:0] select_ln850_3_fu_641_p3;
wire [7:0] select_ln850_fu_720_p3;
wire [3:0] sext_ln1497_fu_199_p0;
wire [3:0] sext_ln545_fu_225_p0;
wire [3:0] sext_ln69_3_fu_370_p1;
wire [3:0] sext_ln703_1_fu_247_p0;
wire [3:0] sext_ln703_fu_654_p0;
wire [9:0] sext_ln703_fu_654_p1;
wire [2:0] sext_ln831_fu_307_p1;
wire \shl_32ns_32s_32_7_1_U3.ce ;
wire \shl_32ns_32s_32_7_1_U3.clk ;
wire [31:0] \shl_32ns_32s_32_7_1_U3.din0 ;
wire [31:0] \shl_32ns_32s_32_7_1_U3.din1 ;
wire [31:0] \shl_32ns_32s_32_7_1_U3.din1_cast ;
wire [31:0] \shl_32ns_32s_32_7_1_U3.din1_mask ;
wire [31:0] \shl_32ns_32s_32_7_1_U3.dout ;
wire \shl_32ns_32s_32_7_1_U3.reset ;
wire \sub_5ns_5s_5_2_1_U1.ce ;
wire \sub_5ns_5s_5_2_1_U1.clk ;
wire [4:0] \sub_5ns_5s_5_2_1_U1.din0 ;
wire [4:0] \sub_5ns_5s_5_2_1_U1.din1 ;
wire [4:0] \sub_5ns_5s_5_2_1_U1.dout ;
wire \sub_5ns_5s_5_2_1_U1.reset ;
wire [4:0] \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.a ;
wire [4:0] \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.ain_s0 ;
wire [4:0] \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.b ;
wire [4:0] \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.bin_s0 ;
wire \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.ce ;
wire \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.clk ;
wire \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.facout_s1 ;
wire \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.facout_s2 ;
wire [1:0] \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.fas_s1 ;
wire [2:0] \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.fas_s2 ;
wire \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.reset ;
wire [4:0] \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.s ;
wire [1:0] \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.u1.a ;
wire [1:0] \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.u1.b ;
wire \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.u1.cin ;
wire \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.u1.cout ;
wire [1:0] \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.u1.s ;
wire [2:0] \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.u2.a ;
wire [2:0] \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.u2.b ;
wire \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.u2.cin ;
wire \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.u2.cout ;
wire [2:0] \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.u2.s ;
wire \sub_5ns_5s_5_2_1_U4.ce ;
wire \sub_5ns_5s_5_2_1_U4.clk ;
wire [4:0] \sub_5ns_5s_5_2_1_U4.din0 ;
wire [4:0] \sub_5ns_5s_5_2_1_U4.din1 ;
wire [4:0] \sub_5ns_5s_5_2_1_U4.dout ;
wire \sub_5ns_5s_5_2_1_U4.reset ;
wire [4:0] \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_0_U.a ;
wire [4:0] \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_0_U.ain_s0 ;
wire [4:0] \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_0_U.b ;
wire [4:0] \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_0_U.bin_s0 ;
wire \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_0_U.ce ;
wire \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_0_U.clk ;
wire \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_0_U.facout_s1 ;
wire \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_0_U.facout_s2 ;
wire [1:0] \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_0_U.fas_s1 ;
wire [2:0] \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_0_U.fas_s2 ;
wire \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_0_U.reset ;
wire [4:0] \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_0_U.s ;
wire [1:0] \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_0_U.u1.a ;
wire [1:0] \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_0_U.u1.b ;
wire \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_0_U.u1.cin ;
wire \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_0_U.u1.cout ;
wire [1:0] \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_0_U.u1.s ;
wire [2:0] \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_0_U.u2.a ;
wire [2:0] \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_0_U.u2.b ;
wire \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_0_U.u2.cin ;
wire \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_0_U.u2.cout ;
wire [2:0] \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_0_U.u2.s ;
wire tmp_6_fu_217_p3;
wire [7:0] tmp_8_fu_599_p3;
wire [3:0] tmp_fu_203_p1;
wire trunc_ln1497_fu_362_p1;
wire [3:0] trunc_ln728_fu_366_p1;
wire [1:0] trunc_ln851_1_fu_267_p1;
wire [1:0] trunc_ln851_2_fu_293_p1;
wire trunc_ln851_3_fu_638_p1;
wire [1:0] trunc_ln851_fu_681_p1;
wire xor_ln340_fu_537_p2;
wire xor_ln785_1_fu_569_p2;
wire xor_ln785_fu_512_p2;
wire xor_ln786_1_fu_564_p2;
wire xor_ln786_fu_522_p2;
wire [3:0] zext_ln1497_fu_383_p1;


assign _046_ = _050_ & ap_CS_fsm[8];
assign _047_ = tmp_reg_773 & ap_CS_fsm[8];
assign _048_ = _051_ & ap_CS_fsm[0];
assign _049_ = ap_start & ap_CS_fsm[0];
assign and_ln340_fu_543_p2 = xor_ln340_fu_537_p2 & or_ln786_fu_527_p2;
assign and_ln785_1_fu_585_p2 = p_Result_5_reg_927 & and_ln785_fu_579_p2;
assign and_ln785_fu_579_p2 = xor_ln786_1_fu_564_p2 & or_ln785_1_fu_574_p2;
assign overflow_fu_517_p2 = xor_ln785_fu_512_p2 & or_ln785_reg_960;
assign ret_V_19_fu_665_p2 = { op_3[3], op_3[3], op_3[3], op_3[3], op_3[3], op_3[3], op_3 } & { op_12, 2'h0 };
assign ret_V_fu_404_p2 = lhs_fu_396_p3 & op_7[6:0];
assign xor_ln786_fu_522_p2 = ~ p_Result_5_reg_927;
assign xor_ln785_fu_512_p2 = ~ p_Result_4_reg_914;
assign xor_ln340_fu_537_p2 = ~ or_ln340_fu_532_p2;
assign xor_ln785_1_fu_569_p2 = ~ or_ln785_reg_960;
assign xor_ln786_1_fu_564_p2 = ~ icmp_ln786_reg_939;
assign _050_ = ~ tmp_reg_773;
assign _051_ = ~ ap_start;
assign _052_ = ! trunc_ln851_1_reg_827;
assign _053_ = ! trunc_ln851_2_reg_842;
assign _054_ = ! trunc_ln851_reg_1036;
always @(posedge \add_10ns_10s_10_2_1_U8.top_add_10ns_10s_10_2_1_Adder_4_U.clk )
\add_10ns_10s_10_2_1_U8.top_add_10ns_10s_10_2_1_Adder_4_U.bin_s1  <= _056_;
always @(posedge \add_10ns_10s_10_2_1_U8.top_add_10ns_10s_10_2_1_Adder_4_U.clk )
\add_10ns_10s_10_2_1_U8.top_add_10ns_10s_10_2_1_Adder_4_U.ain_s1  <= _055_;
always @(posedge \add_10ns_10s_10_2_1_U8.top_add_10ns_10s_10_2_1_Adder_4_U.clk )
\add_10ns_10s_10_2_1_U8.top_add_10ns_10s_10_2_1_Adder_4_U.sum_s1  <= _058_;
always @(posedge \add_10ns_10s_10_2_1_U8.top_add_10ns_10s_10_2_1_Adder_4_U.clk )
\add_10ns_10s_10_2_1_U8.top_add_10ns_10s_10_2_1_Adder_4_U.carry_s1  <= _057_;
assign _056_ = \add_10ns_10s_10_2_1_U8.top_add_10ns_10s_10_2_1_Adder_4_U.ce  ? \add_10ns_10s_10_2_1_U8.top_add_10ns_10s_10_2_1_Adder_4_U.b [9:5] : \add_10ns_10s_10_2_1_U8.top_add_10ns_10s_10_2_1_Adder_4_U.bin_s1 ;
assign _055_ = \add_10ns_10s_10_2_1_U8.top_add_10ns_10s_10_2_1_Adder_4_U.ce  ? \add_10ns_10s_10_2_1_U8.top_add_10ns_10s_10_2_1_Adder_4_U.a [9:5] : \add_10ns_10s_10_2_1_U8.top_add_10ns_10s_10_2_1_Adder_4_U.ain_s1 ;
assign _057_ = \add_10ns_10s_10_2_1_U8.top_add_10ns_10s_10_2_1_Adder_4_U.ce  ? \add_10ns_10s_10_2_1_U8.top_add_10ns_10s_10_2_1_Adder_4_U.facout_s1  : \add_10ns_10s_10_2_1_U8.top_add_10ns_10s_10_2_1_Adder_4_U.carry_s1 ;
assign _058_ = \add_10ns_10s_10_2_1_U8.top_add_10ns_10s_10_2_1_Adder_4_U.ce  ? \add_10ns_10s_10_2_1_U8.top_add_10ns_10s_10_2_1_Adder_4_U.fas_s1  : \add_10ns_10s_10_2_1_U8.top_add_10ns_10s_10_2_1_Adder_4_U.sum_s1 ;
assign _059_ = \add_10ns_10s_10_2_1_U8.top_add_10ns_10s_10_2_1_Adder_4_U.u1.a  + \add_10ns_10s_10_2_1_U8.top_add_10ns_10s_10_2_1_Adder_4_U.u1.b ;
assign { \add_10ns_10s_10_2_1_U8.top_add_10ns_10s_10_2_1_Adder_4_U.u1.cout , \add_10ns_10s_10_2_1_U8.top_add_10ns_10s_10_2_1_Adder_4_U.u1.s  } = _059_ + \add_10ns_10s_10_2_1_U8.top_add_10ns_10s_10_2_1_Adder_4_U.u1.cin ;
assign _060_ = \add_10ns_10s_10_2_1_U8.top_add_10ns_10s_10_2_1_Adder_4_U.u2.a  + \add_10ns_10s_10_2_1_U8.top_add_10ns_10s_10_2_1_Adder_4_U.u2.b ;
assign { \add_10ns_10s_10_2_1_U8.top_add_10ns_10s_10_2_1_Adder_4_U.u2.cout , \add_10ns_10s_10_2_1_U8.top_add_10ns_10s_10_2_1_Adder_4_U.u2.s  } = _060_ + \add_10ns_10s_10_2_1_U8.top_add_10ns_10s_10_2_1_Adder_4_U.u2.cin ;
always @(posedge \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.clk )
\add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s1  <= _062_;
always @(posedge \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.clk )
\add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s1  <= _061_;
always @(posedge \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.clk )
\add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.sum_s1  <= _064_;
always @(posedge \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.clk )
\add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.carry_s1  <= _063_;
assign _062_ = \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.ce  ? \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.b [31:16] : \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s1 ;
assign _061_ = \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.ce  ? \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.a [31:16] : \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s1 ;
assign _063_ = \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.ce  ? \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.facout_s1  : \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.carry_s1 ;
assign _064_ = \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.ce  ? \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s1  : \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.sum_s1 ;
assign _065_ = \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.a  + \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.b ;
assign { \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cout , \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.s  } = _065_ + \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cin ;
assign _066_ = \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.a  + \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.b ;
assign { \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cout , \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.s  } = _066_ + \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cin ;
always @(posedge \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.clk )
\add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.bin_s1  <= _068_;
always @(posedge \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.clk )
\add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.ain_s1  <= _067_;
always @(posedge \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.clk )
\add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.sum_s1  <= _070_;
always @(posedge \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.clk )
\add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.carry_s1  <= _069_;
assign _068_ = \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.ce  ? \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.b [31:16] : \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.bin_s1 ;
assign _067_ = \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.ce  ? \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.a [31:16] : \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.ain_s1 ;
assign _069_ = \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.ce  ? \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.facout_s1  : \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.carry_s1 ;
assign _070_ = \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.ce  ? \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.fas_s1  : \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.sum_s1 ;
assign _071_ = \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.u1.a  + \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.u1.b ;
assign { \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.u1.cout , \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.u1.s  } = _071_ + \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.u1.cin ;
assign _072_ = \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.u2.a  + \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.u2.b ;
assign { \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.u2.cout , \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.u2.s  } = _072_ + \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.u2.cin ;
always @(posedge \add_32ns_32s_32_2_1_U14.top_add_32ns_32s_32_2_1_Adder_8_U.clk )
\add_32ns_32s_32_2_1_U14.top_add_32ns_32s_32_2_1_Adder_8_U.bin_s1  <= _074_;
always @(posedge \add_32ns_32s_32_2_1_U14.top_add_32ns_32s_32_2_1_Adder_8_U.clk )
\add_32ns_32s_32_2_1_U14.top_add_32ns_32s_32_2_1_Adder_8_U.ain_s1  <= _073_;
always @(posedge \add_32ns_32s_32_2_1_U14.top_add_32ns_32s_32_2_1_Adder_8_U.clk )
\add_32ns_32s_32_2_1_U14.top_add_32ns_32s_32_2_1_Adder_8_U.sum_s1  <= _076_;
always @(posedge \add_32ns_32s_32_2_1_U14.top_add_32ns_32s_32_2_1_Adder_8_U.clk )
\add_32ns_32s_32_2_1_U14.top_add_32ns_32s_32_2_1_Adder_8_U.carry_s1  <= _075_;
assign _074_ = \add_32ns_32s_32_2_1_U14.top_add_32ns_32s_32_2_1_Adder_8_U.ce  ? \add_32ns_32s_32_2_1_U14.top_add_32ns_32s_32_2_1_Adder_8_U.b [31:16] : \add_32ns_32s_32_2_1_U14.top_add_32ns_32s_32_2_1_Adder_8_U.bin_s1 ;
assign _073_ = \add_32ns_32s_32_2_1_U14.top_add_32ns_32s_32_2_1_Adder_8_U.ce  ? \add_32ns_32s_32_2_1_U14.top_add_32ns_32s_32_2_1_Adder_8_U.a [31:16] : \add_32ns_32s_32_2_1_U14.top_add_32ns_32s_32_2_1_Adder_8_U.ain_s1 ;
assign _075_ = \add_32ns_32s_32_2_1_U14.top_add_32ns_32s_32_2_1_Adder_8_U.ce  ? \add_32ns_32s_32_2_1_U14.top_add_32ns_32s_32_2_1_Adder_8_U.facout_s1  : \add_32ns_32s_32_2_1_U14.top_add_32ns_32s_32_2_1_Adder_8_U.carry_s1 ;
assign _076_ = \add_32ns_32s_32_2_1_U14.top_add_32ns_32s_32_2_1_Adder_8_U.ce  ? \add_32ns_32s_32_2_1_U14.top_add_32ns_32s_32_2_1_Adder_8_U.fas_s1  : \add_32ns_32s_32_2_1_U14.top_add_32ns_32s_32_2_1_Adder_8_U.sum_s1 ;
assign _077_ = \add_32ns_32s_32_2_1_U14.top_add_32ns_32s_32_2_1_Adder_8_U.u1.a  + \add_32ns_32s_32_2_1_U14.top_add_32ns_32s_32_2_1_Adder_8_U.u1.b ;
assign { \add_32ns_32s_32_2_1_U14.top_add_32ns_32s_32_2_1_Adder_8_U.u1.cout , \add_32ns_32s_32_2_1_U14.top_add_32ns_32s_32_2_1_Adder_8_U.u1.s  } = _077_ + \add_32ns_32s_32_2_1_U14.top_add_32ns_32s_32_2_1_Adder_8_U.u1.cin ;
assign _078_ = \add_32ns_32s_32_2_1_U14.top_add_32ns_32s_32_2_1_Adder_8_U.u2.a  + \add_32ns_32s_32_2_1_U14.top_add_32ns_32s_32_2_1_Adder_8_U.u2.b ;
assign { \add_32ns_32s_32_2_1_U14.top_add_32ns_32s_32_2_1_Adder_8_U.u2.cout , \add_32ns_32s_32_2_1_U14.top_add_32ns_32s_32_2_1_Adder_8_U.u2.s  } = _078_ + \add_32ns_32s_32_2_1_U14.top_add_32ns_32s_32_2_1_Adder_8_U.u2.cin ;
always @(posedge \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_8_U.clk )
\add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_8_U.bin_s1  <= _080_;
always @(posedge \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_8_U.clk )
\add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_8_U.ain_s1  <= _079_;
always @(posedge \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_8_U.clk )
\add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_8_U.sum_s1  <= _082_;
always @(posedge \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_8_U.clk )
\add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_8_U.carry_s1  <= _081_;
assign _080_ = \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_8_U.ce  ? \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_8_U.b [31:16] : \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_8_U.bin_s1 ;
assign _079_ = \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_8_U.ce  ? \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_8_U.a [31:16] : \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_8_U.ain_s1 ;
assign _081_ = \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_8_U.ce  ? \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_8_U.facout_s1  : \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_8_U.carry_s1 ;
assign _082_ = \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_8_U.ce  ? \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_8_U.fas_s1  : \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_8_U.sum_s1 ;
assign _083_ = \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_8_U.u1.a  + \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_8_U.u1.b ;
assign { \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_8_U.u1.cout , \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_8_U.u1.s  } = _083_ + \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_8_U.u1.cin ;
assign _084_ = \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_8_U.u2.a  + \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_8_U.u2.b ;
assign { \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_8_U.u2.cout , \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_8_U.u2.s  } = _084_ + \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_8_U.u2.cin ;
always @(posedge \add_32s_32ns_32_2_1_U17.top_add_32s_32ns_32_2_1_Adder_11_U.clk )
\add_32s_32ns_32_2_1_U17.top_add_32s_32ns_32_2_1_Adder_11_U.bin_s1  <= _086_;
always @(posedge \add_32s_32ns_32_2_1_U17.top_add_32s_32ns_32_2_1_Adder_11_U.clk )
\add_32s_32ns_32_2_1_U17.top_add_32s_32ns_32_2_1_Adder_11_U.ain_s1  <= _085_;
always @(posedge \add_32s_32ns_32_2_1_U17.top_add_32s_32ns_32_2_1_Adder_11_U.clk )
\add_32s_32ns_32_2_1_U17.top_add_32s_32ns_32_2_1_Adder_11_U.sum_s1  <= _088_;
always @(posedge \add_32s_32ns_32_2_1_U17.top_add_32s_32ns_32_2_1_Adder_11_U.clk )
\add_32s_32ns_32_2_1_U17.top_add_32s_32ns_32_2_1_Adder_11_U.carry_s1  <= _087_;
assign _086_ = \add_32s_32ns_32_2_1_U17.top_add_32s_32ns_32_2_1_Adder_11_U.ce  ? \add_32s_32ns_32_2_1_U17.top_add_32s_32ns_32_2_1_Adder_11_U.b [31:16] : \add_32s_32ns_32_2_1_U17.top_add_32s_32ns_32_2_1_Adder_11_U.bin_s1 ;
assign _085_ = \add_32s_32ns_32_2_1_U17.top_add_32s_32ns_32_2_1_Adder_11_U.ce  ? \add_32s_32ns_32_2_1_U17.top_add_32s_32ns_32_2_1_Adder_11_U.a [31:16] : \add_32s_32ns_32_2_1_U17.top_add_32s_32ns_32_2_1_Adder_11_U.ain_s1 ;
assign _087_ = \add_32s_32ns_32_2_1_U17.top_add_32s_32ns_32_2_1_Adder_11_U.ce  ? \add_32s_32ns_32_2_1_U17.top_add_32s_32ns_32_2_1_Adder_11_U.facout_s1  : \add_32s_32ns_32_2_1_U17.top_add_32s_32ns_32_2_1_Adder_11_U.carry_s1 ;
assign _088_ = \add_32s_32ns_32_2_1_U17.top_add_32s_32ns_32_2_1_Adder_11_U.ce  ? \add_32s_32ns_32_2_1_U17.top_add_32s_32ns_32_2_1_Adder_11_U.fas_s1  : \add_32s_32ns_32_2_1_U17.top_add_32s_32ns_32_2_1_Adder_11_U.sum_s1 ;
assign _089_ = \add_32s_32ns_32_2_1_U17.top_add_32s_32ns_32_2_1_Adder_11_U.u1.a  + \add_32s_32ns_32_2_1_U17.top_add_32s_32ns_32_2_1_Adder_11_U.u1.b ;
assign { \add_32s_32ns_32_2_1_U17.top_add_32s_32ns_32_2_1_Adder_11_U.u1.cout , \add_32s_32ns_32_2_1_U17.top_add_32s_32ns_32_2_1_Adder_11_U.u1.s  } = _089_ + \add_32s_32ns_32_2_1_U17.top_add_32s_32ns_32_2_1_Adder_11_U.u1.cin ;
assign _090_ = \add_32s_32ns_32_2_1_U17.top_add_32s_32ns_32_2_1_Adder_11_U.u2.a  + \add_32s_32ns_32_2_1_U17.top_add_32s_32ns_32_2_1_Adder_11_U.u2.b ;
assign { \add_32s_32ns_32_2_1_U17.top_add_32s_32ns_32_2_1_Adder_11_U.u2.cout , \add_32s_32ns_32_2_1_U17.top_add_32s_32ns_32_2_1_Adder_11_U.u2.s  } = _090_ + \add_32s_32ns_32_2_1_U17.top_add_32s_32ns_32_2_1_Adder_11_U.u2.cin ;
always @(posedge \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_6_U.clk )
\add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_6_U.bin_s1  <= _092_;
always @(posedge \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_6_U.clk )
\add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_6_U.ain_s1  <= _091_;
always @(posedge \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_6_U.clk )
\add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_6_U.sum_s1  <= _094_;
always @(posedge \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_6_U.clk )
\add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_6_U.carry_s1  <= _093_;
assign _092_ = \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_6_U.ce  ? \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_6_U.b [33:17] : \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_6_U.bin_s1 ;
assign _091_ = \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_6_U.ce  ? \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_6_U.a [33:17] : \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_6_U.ain_s1 ;
assign _093_ = \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_6_U.ce  ? \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_6_U.facout_s1  : \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_6_U.carry_s1 ;
assign _094_ = \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_6_U.ce  ? \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_6_U.fas_s1  : \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_6_U.sum_s1 ;
assign _095_ = \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_6_U.u1.a  + \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_6_U.u1.b ;
assign { \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_6_U.u1.cout , \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_6_U.u1.s  } = _095_ + \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_6_U.u1.cin ;
assign _096_ = \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_6_U.u2.a  + \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_6_U.u2.b ;
assign { \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_6_U.u2.cout , \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_6_U.u2.s  } = _096_ + \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_6_U.u2.cin ;
always @(posedge \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_1_U.clk )
\add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_1_U.bin_s1  <= _098_;
always @(posedge \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_1_U.clk )
\add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_1_U.ain_s1  <= _097_;
always @(posedge \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_1_U.clk )
\add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_1_U.sum_s1  <= _100_;
always @(posedge \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_1_U.clk )
\add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_1_U.carry_s1  <= _099_;
assign _098_ = \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_1_U.ce  ? \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_1_U.b [2:1] : \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_1_U.bin_s1 ;
assign _097_ = \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_1_U.ce  ? \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_1_U.a [2:1] : \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_1_U.ain_s1 ;
assign _099_ = \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_1_U.ce  ? \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_1_U.facout_s1  : \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_1_U.carry_s1 ;
assign _100_ = \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_1_U.ce  ? \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_1_U.fas_s1  : \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_1_U.sum_s1 ;
assign _101_ = \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_1_U.u1.a  + \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_1_U.u1.b ;
assign { \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_1_U.u1.cout , \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_1_U.u1.s  } = _101_ + \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_1_U.u1.cin ;
assign _102_ = \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_1_U.u2.a  + \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_1_U.u2.b ;
assign { \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_1_U.u2.cout , \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_1_U.u2.s  } = _102_ + \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_1_U.u2.cin ;
always @(posedge \add_3s_3ns_3_2_1_U6.top_add_3s_3ns_3_2_1_Adder_2_U.clk )
\add_3s_3ns_3_2_1_U6.top_add_3s_3ns_3_2_1_Adder_2_U.bin_s1  <= _104_;
always @(posedge \add_3s_3ns_3_2_1_U6.top_add_3s_3ns_3_2_1_Adder_2_U.clk )
\add_3s_3ns_3_2_1_U6.top_add_3s_3ns_3_2_1_Adder_2_U.ain_s1  <= _103_;
always @(posedge \add_3s_3ns_3_2_1_U6.top_add_3s_3ns_3_2_1_Adder_2_U.clk )
\add_3s_3ns_3_2_1_U6.top_add_3s_3ns_3_2_1_Adder_2_U.sum_s1  <= _106_;
always @(posedge \add_3s_3ns_3_2_1_U6.top_add_3s_3ns_3_2_1_Adder_2_U.clk )
\add_3s_3ns_3_2_1_U6.top_add_3s_3ns_3_2_1_Adder_2_U.carry_s1  <= _105_;
assign _104_ = \add_3s_3ns_3_2_1_U6.top_add_3s_3ns_3_2_1_Adder_2_U.ce  ? \add_3s_3ns_3_2_1_U6.top_add_3s_3ns_3_2_1_Adder_2_U.b [2:1] : \add_3s_3ns_3_2_1_U6.top_add_3s_3ns_3_2_1_Adder_2_U.bin_s1 ;
assign _103_ = \add_3s_3ns_3_2_1_U6.top_add_3s_3ns_3_2_1_Adder_2_U.ce  ? \add_3s_3ns_3_2_1_U6.top_add_3s_3ns_3_2_1_Adder_2_U.a [2:1] : \add_3s_3ns_3_2_1_U6.top_add_3s_3ns_3_2_1_Adder_2_U.ain_s1 ;
assign _105_ = \add_3s_3ns_3_2_1_U6.top_add_3s_3ns_3_2_1_Adder_2_U.ce  ? \add_3s_3ns_3_2_1_U6.top_add_3s_3ns_3_2_1_Adder_2_U.facout_s1  : \add_3s_3ns_3_2_1_U6.top_add_3s_3ns_3_2_1_Adder_2_U.carry_s1 ;
assign _106_ = \add_3s_3ns_3_2_1_U6.top_add_3s_3ns_3_2_1_Adder_2_U.ce  ? \add_3s_3ns_3_2_1_U6.top_add_3s_3ns_3_2_1_Adder_2_U.fas_s1  : \add_3s_3ns_3_2_1_U6.top_add_3s_3ns_3_2_1_Adder_2_U.sum_s1 ;
assign _107_ = \add_3s_3ns_3_2_1_U6.top_add_3s_3ns_3_2_1_Adder_2_U.u1.a  + \add_3s_3ns_3_2_1_U6.top_add_3s_3ns_3_2_1_Adder_2_U.u1.b ;
assign { \add_3s_3ns_3_2_1_U6.top_add_3s_3ns_3_2_1_Adder_2_U.u1.cout , \add_3s_3ns_3_2_1_U6.top_add_3s_3ns_3_2_1_Adder_2_U.u1.s  } = _107_ + \add_3s_3ns_3_2_1_U6.top_add_3s_3ns_3_2_1_Adder_2_U.u1.cin ;
assign _108_ = \add_3s_3ns_3_2_1_U6.top_add_3s_3ns_3_2_1_Adder_2_U.u2.a  + \add_3s_3ns_3_2_1_U6.top_add_3s_3ns_3_2_1_Adder_2_U.u2.b ;
assign { \add_3s_3ns_3_2_1_U6.top_add_3s_3ns_3_2_1_Adder_2_U.u2.cout , \add_3s_3ns_3_2_1_U6.top_add_3s_3ns_3_2_1_Adder_2_U.u2.s  } = _108_ + \add_3s_3ns_3_2_1_U6.top_add_3s_3ns_3_2_1_Adder_2_U.u2.cin ;
always @(posedge \add_6ns_6s_6_2_1_U7.top_add_6ns_6s_6_2_1_Adder_3_U.clk )
\add_6ns_6s_6_2_1_U7.top_add_6ns_6s_6_2_1_Adder_3_U.bin_s1  <= _110_;
always @(posedge \add_6ns_6s_6_2_1_U7.top_add_6ns_6s_6_2_1_Adder_3_U.clk )
\add_6ns_6s_6_2_1_U7.top_add_6ns_6s_6_2_1_Adder_3_U.ain_s1  <= _109_;
always @(posedge \add_6ns_6s_6_2_1_U7.top_add_6ns_6s_6_2_1_Adder_3_U.clk )
\add_6ns_6s_6_2_1_U7.top_add_6ns_6s_6_2_1_Adder_3_U.sum_s1  <= _112_;
always @(posedge \add_6ns_6s_6_2_1_U7.top_add_6ns_6s_6_2_1_Adder_3_U.clk )
\add_6ns_6s_6_2_1_U7.top_add_6ns_6s_6_2_1_Adder_3_U.carry_s1  <= _111_;
assign _110_ = \add_6ns_6s_6_2_1_U7.top_add_6ns_6s_6_2_1_Adder_3_U.ce  ? \add_6ns_6s_6_2_1_U7.top_add_6ns_6s_6_2_1_Adder_3_U.b [5:3] : \add_6ns_6s_6_2_1_U7.top_add_6ns_6s_6_2_1_Adder_3_U.bin_s1 ;
assign _109_ = \add_6ns_6s_6_2_1_U7.top_add_6ns_6s_6_2_1_Adder_3_U.ce  ? \add_6ns_6s_6_2_1_U7.top_add_6ns_6s_6_2_1_Adder_3_U.a [5:3] : \add_6ns_6s_6_2_1_U7.top_add_6ns_6s_6_2_1_Adder_3_U.ain_s1 ;
assign _111_ = \add_6ns_6s_6_2_1_U7.top_add_6ns_6s_6_2_1_Adder_3_U.ce  ? \add_6ns_6s_6_2_1_U7.top_add_6ns_6s_6_2_1_Adder_3_U.facout_s1  : \add_6ns_6s_6_2_1_U7.top_add_6ns_6s_6_2_1_Adder_3_U.carry_s1 ;
assign _112_ = \add_6ns_6s_6_2_1_U7.top_add_6ns_6s_6_2_1_Adder_3_U.ce  ? \add_6ns_6s_6_2_1_U7.top_add_6ns_6s_6_2_1_Adder_3_U.fas_s1  : \add_6ns_6s_6_2_1_U7.top_add_6ns_6s_6_2_1_Adder_3_U.sum_s1 ;
assign _113_ = \add_6ns_6s_6_2_1_U7.top_add_6ns_6s_6_2_1_Adder_3_U.u1.a  + \add_6ns_6s_6_2_1_U7.top_add_6ns_6s_6_2_1_Adder_3_U.u1.b ;
assign { \add_6ns_6s_6_2_1_U7.top_add_6ns_6s_6_2_1_Adder_3_U.u1.cout , \add_6ns_6s_6_2_1_U7.top_add_6ns_6s_6_2_1_Adder_3_U.u1.s  } = _113_ + \add_6ns_6s_6_2_1_U7.top_add_6ns_6s_6_2_1_Adder_3_U.u1.cin ;
assign _114_ = \add_6ns_6s_6_2_1_U7.top_add_6ns_6s_6_2_1_Adder_3_U.u2.a  + \add_6ns_6s_6_2_1_U7.top_add_6ns_6s_6_2_1_Adder_3_U.u2.b ;
assign { \add_6ns_6s_6_2_1_U7.top_add_6ns_6s_6_2_1_Adder_3_U.u2.cout , \add_6ns_6s_6_2_1_U7.top_add_6ns_6s_6_2_1_Adder_3_U.u2.s  } = _114_ + \add_6ns_6s_6_2_1_U7.top_add_6ns_6s_6_2_1_Adder_3_U.u2.cin ;
always @(posedge \add_7s_7ns_7_2_1_U9.top_add_7s_7ns_7_2_1_Adder_5_U.clk )
\add_7s_7ns_7_2_1_U9.top_add_7s_7ns_7_2_1_Adder_5_U.bin_s1  <= _116_;
always @(posedge \add_7s_7ns_7_2_1_U9.top_add_7s_7ns_7_2_1_Adder_5_U.clk )
\add_7s_7ns_7_2_1_U9.top_add_7s_7ns_7_2_1_Adder_5_U.ain_s1  <= _115_;
always @(posedge \add_7s_7ns_7_2_1_U9.top_add_7s_7ns_7_2_1_Adder_5_U.clk )
\add_7s_7ns_7_2_1_U9.top_add_7s_7ns_7_2_1_Adder_5_U.sum_s1  <= _118_;
always @(posedge \add_7s_7ns_7_2_1_U9.top_add_7s_7ns_7_2_1_Adder_5_U.clk )
\add_7s_7ns_7_2_1_U9.top_add_7s_7ns_7_2_1_Adder_5_U.carry_s1  <= _117_;
assign _116_ = \add_7s_7ns_7_2_1_U9.top_add_7s_7ns_7_2_1_Adder_5_U.ce  ? \add_7s_7ns_7_2_1_U9.top_add_7s_7ns_7_2_1_Adder_5_U.b [6:3] : \add_7s_7ns_7_2_1_U9.top_add_7s_7ns_7_2_1_Adder_5_U.bin_s1 ;
assign _115_ = \add_7s_7ns_7_2_1_U9.top_add_7s_7ns_7_2_1_Adder_5_U.ce  ? \add_7s_7ns_7_2_1_U9.top_add_7s_7ns_7_2_1_Adder_5_U.a [6:3] : \add_7s_7ns_7_2_1_U9.top_add_7s_7ns_7_2_1_Adder_5_U.ain_s1 ;
assign _117_ = \add_7s_7ns_7_2_1_U9.top_add_7s_7ns_7_2_1_Adder_5_U.ce  ? \add_7s_7ns_7_2_1_U9.top_add_7s_7ns_7_2_1_Adder_5_U.facout_s1  : \add_7s_7ns_7_2_1_U9.top_add_7s_7ns_7_2_1_Adder_5_U.carry_s1 ;
assign _118_ = \add_7s_7ns_7_2_1_U9.top_add_7s_7ns_7_2_1_Adder_5_U.ce  ? \add_7s_7ns_7_2_1_U9.top_add_7s_7ns_7_2_1_Adder_5_U.fas_s1  : \add_7s_7ns_7_2_1_U9.top_add_7s_7ns_7_2_1_Adder_5_U.sum_s1 ;
assign _119_ = \add_7s_7ns_7_2_1_U9.top_add_7s_7ns_7_2_1_Adder_5_U.u1.a  + \add_7s_7ns_7_2_1_U9.top_add_7s_7ns_7_2_1_Adder_5_U.u1.b ;
assign { \add_7s_7ns_7_2_1_U9.top_add_7s_7ns_7_2_1_Adder_5_U.u1.cout , \add_7s_7ns_7_2_1_U9.top_add_7s_7ns_7_2_1_Adder_5_U.u1.s  } = _119_ + \add_7s_7ns_7_2_1_U9.top_add_7s_7ns_7_2_1_Adder_5_U.u1.cin ;
assign _120_ = \add_7s_7ns_7_2_1_U9.top_add_7s_7ns_7_2_1_Adder_5_U.u2.a  + \add_7s_7ns_7_2_1_U9.top_add_7s_7ns_7_2_1_Adder_5_U.u2.b ;
assign { \add_7s_7ns_7_2_1_U9.top_add_7s_7ns_7_2_1_Adder_5_U.u2.cout , \add_7s_7ns_7_2_1_U9.top_add_7s_7ns_7_2_1_Adder_5_U.u2.s  } = _120_ + \add_7s_7ns_7_2_1_U9.top_add_7s_7ns_7_2_1_Adder_5_U.u2.cin ;
always @(posedge \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_9_U.clk )
\add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_9_U.bin_s1  <= _122_;
always @(posedge \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_9_U.clk )
\add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_9_U.ain_s1  <= _121_;
always @(posedge \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_9_U.clk )
\add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_9_U.sum_s1  <= _124_;
always @(posedge \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_9_U.clk )
\add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_9_U.carry_s1  <= _123_;
assign _122_ = \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_9_U.ce  ? \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_9_U.b [7:4] : \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_9_U.bin_s1 ;
assign _121_ = \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_9_U.ce  ? \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_9_U.a [7:4] : \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_9_U.ain_s1 ;
assign _123_ = \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_9_U.ce  ? \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_9_U.facout_s1  : \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_9_U.carry_s1 ;
assign _124_ = \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_9_U.ce  ? \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_9_U.fas_s1  : \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_9_U.sum_s1 ;
assign _125_ = \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_9_U.u1.a  + \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_9_U.u1.b ;
assign { \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_9_U.u1.cout , \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_9_U.u1.s  } = _125_ + \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_9_U.u1.cin ;
assign _126_ = \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_9_U.u2.a  + \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_9_U.u2.b ;
assign { \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_9_U.u2.cout , \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_9_U.u2.s  } = _126_ + \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_9_U.u2.cin ;
always @(posedge \add_9s_9s_9_2_1_U16.top_add_9s_9s_9_2_1_Adder_10_U.clk )
\add_9s_9s_9_2_1_U16.top_add_9s_9s_9_2_1_Adder_10_U.bin_s1  <= _128_;
always @(posedge \add_9s_9s_9_2_1_U16.top_add_9s_9s_9_2_1_Adder_10_U.clk )
\add_9s_9s_9_2_1_U16.top_add_9s_9s_9_2_1_Adder_10_U.ain_s1  <= _127_;
always @(posedge \add_9s_9s_9_2_1_U16.top_add_9s_9s_9_2_1_Adder_10_U.clk )
\add_9s_9s_9_2_1_U16.top_add_9s_9s_9_2_1_Adder_10_U.sum_s1  <= _130_;
always @(posedge \add_9s_9s_9_2_1_U16.top_add_9s_9s_9_2_1_Adder_10_U.clk )
\add_9s_9s_9_2_1_U16.top_add_9s_9s_9_2_1_Adder_10_U.carry_s1  <= _129_;
assign _128_ = \add_9s_9s_9_2_1_U16.top_add_9s_9s_9_2_1_Adder_10_U.ce  ? \add_9s_9s_9_2_1_U16.top_add_9s_9s_9_2_1_Adder_10_U.b [8:4] : \add_9s_9s_9_2_1_U16.top_add_9s_9s_9_2_1_Adder_10_U.bin_s1 ;
assign _127_ = \add_9s_9s_9_2_1_U16.top_add_9s_9s_9_2_1_Adder_10_U.ce  ? \add_9s_9s_9_2_1_U16.top_add_9s_9s_9_2_1_Adder_10_U.a [8:4] : \add_9s_9s_9_2_1_U16.top_add_9s_9s_9_2_1_Adder_10_U.ain_s1 ;
assign _129_ = \add_9s_9s_9_2_1_U16.top_add_9s_9s_9_2_1_Adder_10_U.ce  ? \add_9s_9s_9_2_1_U16.top_add_9s_9s_9_2_1_Adder_10_U.facout_s1  : \add_9s_9s_9_2_1_U16.top_add_9s_9s_9_2_1_Adder_10_U.carry_s1 ;
assign _130_ = \add_9s_9s_9_2_1_U16.top_add_9s_9s_9_2_1_Adder_10_U.ce  ? \add_9s_9s_9_2_1_U16.top_add_9s_9s_9_2_1_Adder_10_U.fas_s1  : \add_9s_9s_9_2_1_U16.top_add_9s_9s_9_2_1_Adder_10_U.sum_s1 ;
assign _131_ = \add_9s_9s_9_2_1_U16.top_add_9s_9s_9_2_1_Adder_10_U.u1.a  + \add_9s_9s_9_2_1_U16.top_add_9s_9s_9_2_1_Adder_10_U.u1.b ;
assign { \add_9s_9s_9_2_1_U16.top_add_9s_9s_9_2_1_Adder_10_U.u1.cout , \add_9s_9s_9_2_1_U16.top_add_9s_9s_9_2_1_Adder_10_U.u1.s  } = _131_ + \add_9s_9s_9_2_1_U16.top_add_9s_9s_9_2_1_Adder_10_U.u1.cin ;
assign _132_ = \add_9s_9s_9_2_1_U16.top_add_9s_9s_9_2_1_Adder_10_U.u2.a  + \add_9s_9s_9_2_1_U16.top_add_9s_9s_9_2_1_Adder_10_U.u2.b ;
assign { \add_9s_9s_9_2_1_U16.top_add_9s_9s_9_2_1_Adder_10_U.u2.cout , \add_9s_9s_9_2_1_U16.top_add_9s_9s_9_2_1_Adder_10_U.u2.s  } = _132_ + \add_9s_9s_9_2_1_U16.top_add_9s_9s_9_2_1_Adder_10_U.u2.cin ;
always @(posedge \lshr_32ns_32s_32_7_1_U2.clk )
\lshr_32ns_32s_32_7_1_U2.dout_array[5]  <= _144_;
always @(posedge \lshr_32ns_32s_32_7_1_U2.clk )
\lshr_32ns_32s_32_7_1_U2.din1_cast_array[5]  <= _138_;
always @(posedge \lshr_32ns_32s_32_7_1_U2.clk )
\lshr_32ns_32s_32_7_1_U2.dout_array[4]  <= _143_;
always @(posedge \lshr_32ns_32s_32_7_1_U2.clk )
\lshr_32ns_32s_32_7_1_U2.din1_cast_array[4]  <= _137_;
always @(posedge \lshr_32ns_32s_32_7_1_U2.clk )
\lshr_32ns_32s_32_7_1_U2.dout_array[3]  <= _142_;
always @(posedge \lshr_32ns_32s_32_7_1_U2.clk )
\lshr_32ns_32s_32_7_1_U2.din1_cast_array[3]  <= _136_;
always @(posedge \lshr_32ns_32s_32_7_1_U2.clk )
\lshr_32ns_32s_32_7_1_U2.dout_array[2]  <= _141_;
always @(posedge \lshr_32ns_32s_32_7_1_U2.clk )
\lshr_32ns_32s_32_7_1_U2.din1_cast_array[2]  <= _135_;
always @(posedge \lshr_32ns_32s_32_7_1_U2.clk )
\lshr_32ns_32s_32_7_1_U2.dout_array[1]  <= _140_;
always @(posedge \lshr_32ns_32s_32_7_1_U2.clk )
\lshr_32ns_32s_32_7_1_U2.din1_cast_array[1]  <= _134_;
always @(posedge \lshr_32ns_32s_32_7_1_U2.clk )
\lshr_32ns_32s_32_7_1_U2.dout_array[0]  <= _139_;
always @(posedge \lshr_32ns_32s_32_7_1_U2.clk )
\lshr_32ns_32s_32_7_1_U2.din1_cast_array[0]  <= _133_;
assign _145_ = \lshr_32ns_32s_32_7_1_U2.ce  ? \lshr_32ns_32s_32_7_1_U2.din1_cast_array[4]  : \lshr_32ns_32s_32_7_1_U2.din1_cast_array[5] ;
assign _138_ = \lshr_32ns_32s_32_7_1_U2.reset  ? 32'd0 : _145_;
assign _146_ = \lshr_32ns_32s_32_7_1_U2.ce  ? _162_ : \lshr_32ns_32s_32_7_1_U2.dout_array[5] ;
assign _144_ = \lshr_32ns_32s_32_7_1_U2.reset  ? 32'd0 : _146_;
assign _147_ = \lshr_32ns_32s_32_7_1_U2.ce  ? \lshr_32ns_32s_32_7_1_U2.din1_cast_array[3]  : \lshr_32ns_32s_32_7_1_U2.din1_cast_array[4] ;
assign _137_ = \lshr_32ns_32s_32_7_1_U2.reset  ? 32'd0 : _147_;
assign _148_ = \lshr_32ns_32s_32_7_1_U2.ce  ? _161_ : \lshr_32ns_32s_32_7_1_U2.dout_array[4] ;
assign _143_ = \lshr_32ns_32s_32_7_1_U2.reset  ? 32'd0 : _148_;
assign _149_ = \lshr_32ns_32s_32_7_1_U2.ce  ? \lshr_32ns_32s_32_7_1_U2.din1_cast_array[2]  : \lshr_32ns_32s_32_7_1_U2.din1_cast_array[3] ;
assign _136_ = \lshr_32ns_32s_32_7_1_U2.reset  ? 32'd0 : _149_;
assign _150_ = \lshr_32ns_32s_32_7_1_U2.ce  ? _160_ : \lshr_32ns_32s_32_7_1_U2.dout_array[3] ;
assign _142_ = \lshr_32ns_32s_32_7_1_U2.reset  ? 32'd0 : _150_;
assign _151_ = \lshr_32ns_32s_32_7_1_U2.ce  ? \lshr_32ns_32s_32_7_1_U2.din1_cast_array[1]  : \lshr_32ns_32s_32_7_1_U2.din1_cast_array[2] ;
assign _135_ = \lshr_32ns_32s_32_7_1_U2.reset  ? 32'd0 : _151_;
assign _152_ = \lshr_32ns_32s_32_7_1_U2.ce  ? _159_ : \lshr_32ns_32s_32_7_1_U2.dout_array[2] ;
assign _141_ = \lshr_32ns_32s_32_7_1_U2.reset  ? 32'd0 : _152_;
assign _153_ = \lshr_32ns_32s_32_7_1_U2.ce  ? \lshr_32ns_32s_32_7_1_U2.din1_cast_array[0]  : \lshr_32ns_32s_32_7_1_U2.din1_cast_array[1] ;
assign _134_ = \lshr_32ns_32s_32_7_1_U2.reset  ? 32'd0 : _153_;
assign _154_ = \lshr_32ns_32s_32_7_1_U2.ce  ? _158_ : \lshr_32ns_32s_32_7_1_U2.dout_array[1] ;
assign _140_ = \lshr_32ns_32s_32_7_1_U2.reset  ? 32'd0 : _154_;
assign _155_ = \lshr_32ns_32s_32_7_1_U2.ce  ? \lshr_32ns_32s_32_7_1_U2.din1  : \lshr_32ns_32s_32_7_1_U2.din1_cast_array[0] ;
assign _133_ = \lshr_32ns_32s_32_7_1_U2.reset  ? 32'd0 : _155_;
assign _156_ = \lshr_32ns_32s_32_7_1_U2.ce  ? _157_ : \lshr_32ns_32s_32_7_1_U2.dout_array[0] ;
assign _139_ = \lshr_32ns_32s_32_7_1_U2.reset  ? 32'd0 : _156_;
assign _157_ = \lshr_32ns_32s_32_7_1_U2.din0  >> { \lshr_32ns_32s_32_7_1_U2.din1 [31:30], 30'h00000000 };
assign _158_ = \lshr_32ns_32s_32_7_1_U2.dout_array[0]  >> { \lshr_32ns_32s_32_7_1_U2.din1_cast_array[0] [29:25], 25'h0000000 };
assign _159_ = \lshr_32ns_32s_32_7_1_U2.dout_array[1]  >> { \lshr_32ns_32s_32_7_1_U2.din1_cast_array[1] [24:20], 20'h00000 };
assign _160_ = \lshr_32ns_32s_32_7_1_U2.dout_array[2]  >> { \lshr_32ns_32s_32_7_1_U2.din1_cast_array[2] [19:15], 15'h0000 };
assign _161_ = \lshr_32ns_32s_32_7_1_U2.dout_array[3]  >> { \lshr_32ns_32s_32_7_1_U2.din1_cast_array[3] [14:10], 10'h000 };
assign _162_ = \lshr_32ns_32s_32_7_1_U2.dout_array[4]  >> { \lshr_32ns_32s_32_7_1_U2.din1_cast_array[4] [9:5], 5'h00 };
assign \lshr_32ns_32s_32_7_1_U2.dout  = \lshr_32ns_32s_32_7_1_U2.dout_array[5]  >> \lshr_32ns_32s_32_7_1_U2.din1_cast_array[5] [4:0];
always @(posedge \shl_32ns_32s_32_7_1_U3.clk )
\shl_32ns_32s_32_7_1_U3.dout_array[5]  <= _174_;
always @(posedge \shl_32ns_32s_32_7_1_U3.clk )
\shl_32ns_32s_32_7_1_U3.din1_cast_array[5]  <= _168_;
always @(posedge \shl_32ns_32s_32_7_1_U3.clk )
\shl_32ns_32s_32_7_1_U3.dout_array[4]  <= _173_;
always @(posedge \shl_32ns_32s_32_7_1_U3.clk )
\shl_32ns_32s_32_7_1_U3.din1_cast_array[4]  <= _167_;
always @(posedge \shl_32ns_32s_32_7_1_U3.clk )
\shl_32ns_32s_32_7_1_U3.dout_array[3]  <= _172_;
always @(posedge \shl_32ns_32s_32_7_1_U3.clk )
\shl_32ns_32s_32_7_1_U3.din1_cast_array[3]  <= _166_;
always @(posedge \shl_32ns_32s_32_7_1_U3.clk )
\shl_32ns_32s_32_7_1_U3.dout_array[2]  <= _171_;
always @(posedge \shl_32ns_32s_32_7_1_U3.clk )
\shl_32ns_32s_32_7_1_U3.din1_cast_array[2]  <= _165_;
always @(posedge \shl_32ns_32s_32_7_1_U3.clk )
\shl_32ns_32s_32_7_1_U3.dout_array[1]  <= _170_;
always @(posedge \shl_32ns_32s_32_7_1_U3.clk )
\shl_32ns_32s_32_7_1_U3.din1_cast_array[1]  <= _164_;
always @(posedge \shl_32ns_32s_32_7_1_U3.clk )
\shl_32ns_32s_32_7_1_U3.dout_array[0]  <= _169_;
always @(posedge \shl_32ns_32s_32_7_1_U3.clk )
\shl_32ns_32s_32_7_1_U3.din1_cast_array[0]  <= _163_;
assign _175_ = \shl_32ns_32s_32_7_1_U3.ce  ? \shl_32ns_32s_32_7_1_U3.din1_cast_array[4]  : \shl_32ns_32s_32_7_1_U3.din1_cast_array[5] ;
assign _168_ = \shl_32ns_32s_32_7_1_U3.reset  ? 32'd0 : _175_;
assign _176_ = \shl_32ns_32s_32_7_1_U3.ce  ? _192_ : \shl_32ns_32s_32_7_1_U3.dout_array[5] ;
assign _174_ = \shl_32ns_32s_32_7_1_U3.reset  ? 32'd0 : _176_;
assign _177_ = \shl_32ns_32s_32_7_1_U3.ce  ? \shl_32ns_32s_32_7_1_U3.din1_cast_array[3]  : \shl_32ns_32s_32_7_1_U3.din1_cast_array[4] ;
assign _167_ = \shl_32ns_32s_32_7_1_U3.reset  ? 32'd0 : _177_;
assign _178_ = \shl_32ns_32s_32_7_1_U3.ce  ? _191_ : \shl_32ns_32s_32_7_1_U3.dout_array[4] ;
assign _173_ = \shl_32ns_32s_32_7_1_U3.reset  ? 32'd0 : _178_;
assign _179_ = \shl_32ns_32s_32_7_1_U3.ce  ? \shl_32ns_32s_32_7_1_U3.din1_cast_array[2]  : \shl_32ns_32s_32_7_1_U3.din1_cast_array[3] ;
assign _166_ = \shl_32ns_32s_32_7_1_U3.reset  ? 32'd0 : _179_;
assign _180_ = \shl_32ns_32s_32_7_1_U3.ce  ? _190_ : \shl_32ns_32s_32_7_1_U3.dout_array[3] ;
assign _172_ = \shl_32ns_32s_32_7_1_U3.reset  ? 32'd0 : _180_;
assign _181_ = \shl_32ns_32s_32_7_1_U3.ce  ? \shl_32ns_32s_32_7_1_U3.din1_cast_array[1]  : \shl_32ns_32s_32_7_1_U3.din1_cast_array[2] ;
assign _165_ = \shl_32ns_32s_32_7_1_U3.reset  ? 32'd0 : _181_;
assign _182_ = \shl_32ns_32s_32_7_1_U3.ce  ? _189_ : \shl_32ns_32s_32_7_1_U3.dout_array[2] ;
assign _171_ = \shl_32ns_32s_32_7_1_U3.reset  ? 32'd0 : _182_;
assign _183_ = \shl_32ns_32s_32_7_1_U3.ce  ? \shl_32ns_32s_32_7_1_U3.din1_cast_array[0]  : \shl_32ns_32s_32_7_1_U3.din1_cast_array[1] ;
assign _164_ = \shl_32ns_32s_32_7_1_U3.reset  ? 32'd0 : _183_;
assign _184_ = \shl_32ns_32s_32_7_1_U3.ce  ? _188_ : \shl_32ns_32s_32_7_1_U3.dout_array[1] ;
assign _170_ = \shl_32ns_32s_32_7_1_U3.reset  ? 32'd0 : _184_;
assign _185_ = \shl_32ns_32s_32_7_1_U3.ce  ? \shl_32ns_32s_32_7_1_U3.din1  : \shl_32ns_32s_32_7_1_U3.din1_cast_array[0] ;
assign _163_ = \shl_32ns_32s_32_7_1_U3.reset  ? 32'd0 : _185_;
assign _186_ = \shl_32ns_32s_32_7_1_U3.ce  ? _187_ : \shl_32ns_32s_32_7_1_U3.dout_array[0] ;
assign _169_ = \shl_32ns_32s_32_7_1_U3.reset  ? 32'd0 : _186_;
assign _187_ = \shl_32ns_32s_32_7_1_U3.din0  << { \shl_32ns_32s_32_7_1_U3.din1 [31:30], 30'h00000000 };
assign _188_ = \shl_32ns_32s_32_7_1_U3.dout_array[0]  << { \shl_32ns_32s_32_7_1_U3.din1_cast_array[0] [29:25], 25'h0000000 };
assign _189_ = \shl_32ns_32s_32_7_1_U3.dout_array[1]  << { \shl_32ns_32s_32_7_1_U3.din1_cast_array[1] [24:20], 20'h00000 };
assign _190_ = \shl_32ns_32s_32_7_1_U3.dout_array[2]  << { \shl_32ns_32s_32_7_1_U3.din1_cast_array[2] [19:15], 15'h0000 };
assign _191_ = \shl_32ns_32s_32_7_1_U3.dout_array[3]  << { \shl_32ns_32s_32_7_1_U3.din1_cast_array[3] [14:10], 10'h000 };
assign _192_ = \shl_32ns_32s_32_7_1_U3.dout_array[4]  << { \shl_32ns_32s_32_7_1_U3.din1_cast_array[4] [9:5], 5'h00 };
assign \shl_32ns_32s_32_7_1_U3.dout  = \shl_32ns_32s_32_7_1_U3.dout_array[5]  << \shl_32ns_32s_32_7_1_U3.din1_cast_array[5] [4:0];
assign \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.bin_s0  = ~ \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.b ;
always @(posedge \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.clk )
\sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.bin_s1  <= _194_;
always @(posedge \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.clk )
\sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.ain_s1  <= _193_;
always @(posedge \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.clk )
\sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.sum_s1  <= _196_;
always @(posedge \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.clk )
\sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.carry_s1  <= _195_;
assign _194_ = \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.ce  ? \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.bin_s0 [4:2] : \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.bin_s1 ;
assign _193_ = \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.ce  ? \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.a [4:2] : \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.ain_s1 ;
assign _195_ = \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.ce  ? \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.facout_s1  : \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.carry_s1 ;
assign _196_ = \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.ce  ? \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.fas_s1  : \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.sum_s1 ;
assign _197_ = \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.u1.a  + \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.u1.b ;
assign { \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.u1.cout , \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.u1.s  } = _197_ + \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.u1.cin ;
assign _198_ = \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.u2.a  + \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.u2.b ;
assign { \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.u2.cout , \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.u2.s  } = _198_ + \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.u2.cin ;
assign \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_0_U.bin_s0  = ~ \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_0_U.b ;
always @(posedge \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_0_U.clk )
\sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_0_U.bin_s1  <= _200_;
always @(posedge \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_0_U.clk )
\sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_0_U.ain_s1  <= _199_;
always @(posedge \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_0_U.clk )
\sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_0_U.sum_s1  <= _202_;
always @(posedge \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_0_U.clk )
\sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_0_U.carry_s1  <= _201_;
assign _200_ = \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_0_U.ce  ? \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_0_U.bin_s0 [4:2] : \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_0_U.bin_s1 ;
assign _199_ = \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_0_U.ce  ? \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_0_U.a [4:2] : \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_0_U.ain_s1 ;
assign _201_ = \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_0_U.ce  ? \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_0_U.facout_s1  : \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_0_U.carry_s1 ;
assign _202_ = \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_0_U.ce  ? \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_0_U.fas_s1  : \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_0_U.sum_s1 ;
assign _203_ = \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_0_U.u1.a  + \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_0_U.u1.b ;
assign { \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_0_U.u1.cout , \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_0_U.u1.s  } = _203_ + \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_0_U.u1.cin ;
assign _204_ = \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_0_U.u2.a  + \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_0_U.u2.b ;
assign { \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_0_U.u2.cout , \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_0_U.u2.s  } = _204_ + \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_0_U.u2.cin ;
assign _205_ = | op_7[15:7];
assign _206_ = op_7[15:7] != 9'h1ff;
assign or_ln340_fu_532_p2 = p_Result_4_reg_914 | overflow_fu_517_p2;
assign or_ln785_1_fu_574_p2 = xor_ln785_1_fu_569_p2 | p_Result_4_reg_914;
assign or_ln785_fu_498_p2 = p_Result_5_reg_927 | icmp_ln768_reg_934;
assign or_ln786_fu_527_p2 = xor_ln786_fu_522_p2 | icmp_ln786_reg_939;
always @(posedge ap_clk)
trunc_ln851_reg_1036 <= 2'h0;
always @(posedge ap_clk)
trunc_ln728_reg_894 <= _042_;
always @(posedge ap_clk)
trunc_ln1497_reg_889 <= _041_;
always @(posedge ap_clk)
tmp_reg_773 <= _040_;
always @(posedge ap_clk)
tmp_6_reg_783 <= _039_;
always @(posedge ap_clk)
sub_ln1497_reg_778 <= _038_;
always @(posedge ap_clk)
select_ln340_reg_971 <= _036_;
always @(posedge ap_clk)
ret_V_3_reg_1056 <= _031_;
always @(posedge ap_clk)
ret_V_27_reg_1019 <= _027_;
always @(posedge ap_clk)
ret_V_22_reg_874 <= _022_;
always @(posedge ap_clk)
ret_V_24_reg_879 <= _024_;
always @(posedge ap_clk)
ret_V_20_reg_1066 <= _020_;
always @(posedge ap_clk)
ret_V_28_reg_1071 <= _028_;
always @(posedge ap_clk)
_541_ <= _019_;
assign ret_V_19_reg_1024[9:2] = _541_;
always @(posedge ap_clk)
ret_V_2_reg_1029 <= _030_;
always @(posedge ap_clk)
ret_V_26_reg_1002 <= _026_;
always @(posedge ap_clk)
ret_V_16_cast_reg_1007 <= _018_;
always @(posedge ap_clk)
ret_V_7_reg_864 <= _033_;
always @(posedge ap_clk)
ret_V_11_reg_869 <= _017_;
always @(posedge ap_clk)
ret_V_21_reg_815 <= _021_;
always @(posedge ap_clk)
ret_V_6_reg_820 <= _032_;
always @(posedge ap_clk)
trunc_ln851_1_reg_827 <= _043_;
always @(posedge ap_clk)
ret_V_23_reg_832 <= _023_;
always @(posedge ap_clk)
ret_V_10_reg_837 <= _016_;
always @(posedge ap_clk)
trunc_ln851_2_reg_842 <= _044_;
always @(posedge ap_clk)
or_ln785_reg_960 <= _012_;
always @(posedge ap_clk)
op_22_V_reg_966 <= _010_;
always @(posedge ap_clk)
select_ln1497_reg_904 <= _035_;
always @(posedge ap_clk)
op_20_V_reg_909 <= _009_;
always @(posedge ap_clk)
op_14_V_reg_981 <= _008_;
always @(posedge ap_clk)
ret_V_25_reg_987 <= _025_;
always @(posedge ap_clk)
icmp_ln851_reg_1046 <= _007_;
always @(posedge ap_clk)
op_25_V_reg_1051 <= _011_;
always @(posedge ap_clk)
icmp_ln851_1_reg_847 <= _005_;
always @(posedge ap_clk)
sext_ln831_reg_852 <= _037_;
always @(posedge ap_clk)
icmp_ln851_2_reg_859 <= _006_;
always @(posedge ap_clk)
p_Result_4_reg_914 <= _013_;
always @(posedge ap_clk)
p_Val2_s_reg_921 <= _015_;
always @(posedge ap_clk)
p_Result_5_reg_927 <= _014_;
always @(posedge ap_clk)
icmp_ln768_reg_934 <= _003_;
always @(posedge ap_clk)
icmp_ln786_reg_939 <= _004_;
always @(posedge ap_clk)
select_ln1192_reg_955 <= _034_;
always @(posedge ap_clk)
ret_V_29_reg_1091 <= _029_;
always @(posedge ap_clk)
add_ln69_reg_1096 <= _001_;
always @(posedge ap_clk)
add_ln691_reg_1014 <= _000_;
always @(posedge ap_clk)
ap_CS_fsm <= _002_;
assign _045_ = _049_ ? 2'h2 : 2'h1;
assign _207_ = ap_CS_fsm == 1'h1;
function [26:0] _576_;
input [26:0] a;
input [728:0] b;
input [26:0] s;
case (s)
27'b000000000000000000000000001:
_576_ = b[26:0];
27'b000000000000000000000000010:
_576_ = b[53:27];
27'b000000000000000000000000100:
_576_ = b[80:54];
27'b000000000000000000000001000:
_576_ = b[107:81];
27'b000000000000000000000010000:
_576_ = b[134:108];
27'b000000000000000000000100000:
_576_ = b[161:135];
27'b000000000000000000001000000:
_576_ = b[188:162];
27'b000000000000000000010000000:
_576_ = b[215:189];
27'b000000000000000000100000000:
_576_ = b[242:216];
27'b000000000000000001000000000:
_576_ = b[269:243];
27'b000000000000000010000000000:
_576_ = b[296:270];
27'b000000000000000100000000000:
_576_ = b[323:297];
27'b000000000000001000000000000:
_576_ = b[350:324];
27'b000000000000010000000000000:
_576_ = b[377:351];
27'b000000000000100000000000000:
_576_ = b[404:378];
27'b000000000001000000000000000:
_576_ = b[431:405];
27'b000000000010000000000000000:
_576_ = b[458:432];
27'b000000000100000000000000000:
_576_ = b[485:459];
27'b000000001000000000000000000:
_576_ = b[512:486];
27'b000000010000000000000000000:
_576_ = b[539:513];
27'b000000100000000000000000000:
_576_ = b[566:540];
27'b000001000000000000000000000:
_576_ = b[593:567];
27'b000010000000000000000000000:
_576_ = b[620:594];
27'b000100000000000000000000000:
_576_ = b[647:621];
27'b001000000000000000000000000:
_576_ = b[674:648];
27'b010000000000000000000000000:
_576_ = b[701:675];
27'b100000000000000000000000000:
_576_ = b[728:702];
27'b000000000000000000000000000:
_576_ = a;
default:
_576_ = 27'bx;
endcase
endfunction
assign ap_NS_fsm = _576_(27'hxxxxxxx, { 25'h0000000, _045_, 702'h00000020000008000002000000800000200000080000020000008000002000000800000200000080000020000008000002000000800000200000080000020000008000002000000800000200000080000020000000000001 }, { _207_, _233_, _232_, _231_, _230_, _229_, _228_, _227_, _226_, _225_, _224_, _223_, _222_, _221_, _220_, _219_, _218_, _217_, _216_, _215_, _214_, _213_, _212_, _211_, _210_, _209_, _208_ });
assign _208_ = ap_CS_fsm == 27'h4000000;
assign _209_ = ap_CS_fsm == 26'h2000000;
assign _210_ = ap_CS_fsm == 25'h1000000;
assign _211_ = ap_CS_fsm == 24'h800000;
assign _212_ = ap_CS_fsm == 23'h400000;
assign _213_ = ap_CS_fsm == 22'h200000;
assign _214_ = ap_CS_fsm == 21'h100000;
assign _215_ = ap_CS_fsm == 20'h80000;
assign _216_ = ap_CS_fsm == 19'h40000;
assign _217_ = ap_CS_fsm == 18'h20000;
assign _218_ = ap_CS_fsm == 17'h10000;
assign _219_ = ap_CS_fsm == 16'h8000;
assign _220_ = ap_CS_fsm == 15'h4000;
assign _221_ = ap_CS_fsm == 14'h2000;
assign _222_ = ap_CS_fsm == 13'h1000;
assign _223_ = ap_CS_fsm == 12'h800;
assign _224_ = ap_CS_fsm == 11'h400;
assign _225_ = ap_CS_fsm == 10'h200;
assign _226_ = ap_CS_fsm == 9'h100;
assign _227_ = ap_CS_fsm == 8'h80;
assign _228_ = ap_CS_fsm == 7'h40;
assign _229_ = ap_CS_fsm == 6'h20;
assign _230_ = ap_CS_fsm == 5'h10;
assign _231_ = ap_CS_fsm == 4'h8;
assign _232_ = ap_CS_fsm == 3'h4;
assign _233_ = ap_CS_fsm == 2'h2;
assign op_29_ap_vld = ap_CS_fsm[26] ? 1'h1 : 1'h0;
assign ap_idle = _048_ ? 1'h1 : 1'h0;
assign _042_ = _047_ ? grp_fu_241_p2[3:0] : trunc_ln728_reg_894;
assign _041_ = _046_ ? grp_fu_232_p2[0] : trunc_ln1497_reg_889;
assign _040_ = ap_CS_fsm[0] ? op_6[3] : tmp_reg_773;
assign _039_ = ap_CS_fsm[2] ? op_0[1] : tmp_6_reg_783;
assign _038_ = ap_CS_fsm[1] ? grp_fu_211_p2 : sub_ln1497_reg_778;
assign _036_ = ap_CS_fsm[12] ? select_ln340_fu_549_p3 : select_ln340_reg_971;
assign _031_ = ap_CS_fsm[21] ? grp_fu_699_p2 : ret_V_3_reg_1056;
assign _027_ = ap_CS_fsm[18] ? ret_V_27_fu_647_p3 : ret_V_27_reg_1019;
assign _024_ = ap_CS_fsm[7] ? ret_V_24_fu_352_p3 : ret_V_24_reg_879;
assign _022_ = ap_CS_fsm[7] ? ret_V_22_fu_333_p3 : ret_V_22_reg_874;
assign _028_ = ap_CS_fsm[22] ? grp_fu_708_p2 : ret_V_28_reg_1071;
assign _020_ = ap_CS_fsm[22] ? ret_V_20_fu_725_p3 : ret_V_20_reg_1066;
assign _030_ = ap_CS_fsm[19] ? ret_V_19_fu_665_p2[9:2] : ret_V_2_reg_1029;
assign _019_ = ap_CS_fsm[19] ? ret_V_19_fu_665_p2[9:2] : ret_V_19_reg_1024[9:2];
assign _018_ = ap_CS_fsm[15] ? grp_fu_610_p2[32:1] : ret_V_16_cast_reg_1007;
assign _026_ = ap_CS_fsm[15] ? grp_fu_610_p2 : ret_V_26_reg_1002;
assign _017_ = ap_CS_fsm[6] ? grp_fu_315_p2 : ret_V_11_reg_869;
assign _033_ = ap_CS_fsm[6] ? grp_fu_302_p2 : ret_V_7_reg_864;
assign _044_ = ap_CS_fsm[4] ? ret_V_23_fu_278_p2[1:0] : trunc_ln851_2_reg_842;
assign _016_ = ap_CS_fsm[4] ? ret_V_23_fu_278_p2[3:2] : ret_V_10_reg_837;
assign _023_ = ap_CS_fsm[4] ? ret_V_23_fu_278_p2 : ret_V_23_reg_832;
assign _043_ = ap_CS_fsm[4] ? grp_fu_251_p2[1:0] : trunc_ln851_1_reg_827;
assign _032_ = ap_CS_fsm[4] ? grp_fu_251_p2[4:2] : ret_V_6_reg_820;
assign _021_ = ap_CS_fsm[4] ? grp_fu_251_p2 : ret_V_21_reg_815;
assign _010_ = ap_CS_fsm[11] ? grp_fu_484_p2[9:4] : op_22_V_reg_966;
assign _012_ = ap_CS_fsm[11] ? or_ln785_fu_498_p2 : or_ln785_reg_960;
assign _009_ = ap_CS_fsm[9] ? grp_fu_377_p2 : op_20_V_reg_909;
assign _035_ = ap_CS_fsm[9] ? select_ln1497_fu_386_p3 : select_ln1497_reg_904;
assign _025_ = ap_CS_fsm[13] ? grp_fu_559_p2 : ret_V_25_reg_987;
assign _008_ = ap_CS_fsm[13] ? op_14_V_fu_590_p3 : op_14_V_reg_981;
assign _011_ = ap_CS_fsm[20] ? grp_fu_689_p2 : op_25_V_reg_1051;
assign _007_ = ap_CS_fsm[20] ? icmp_ln851_fu_694_p2 : icmp_ln851_reg_1046;
assign _006_ = ap_CS_fsm[5] ? icmp_ln851_2_fu_310_p2 : icmp_ln851_2_reg_859;
assign _037_ = ap_CS_fsm[5] ? { ret_V_10_reg_837[1], ret_V_10_reg_837 } : sext_ln831_reg_852;
assign _005_ = ap_CS_fsm[5] ? icmp_ln851_1_fu_297_p2 : icmp_ln851_1_reg_847;
assign _034_ = ap_CS_fsm[10] ? select_ln1192_fu_490_p3 : select_ln1192_reg_955;
assign _004_ = ap_CS_fsm[10] ? icmp_ln786_fu_460_p2 : icmp_ln786_reg_939;
assign _003_ = ap_CS_fsm[10] ? icmp_ln768_fu_454_p2 : icmp_ln768_reg_934;
assign _014_ = ap_CS_fsm[10] ? op_7[6] : p_Result_5_reg_927;
assign _015_ = ap_CS_fsm[10] ? op_7[6:5] : p_Val2_s_reg_921;
assign _013_ = ap_CS_fsm[10] ? op_7[15] : p_Result_4_reg_914;
assign _001_ = ap_CS_fsm[24] ? grp_fu_748_p2 : add_ln69_reg_1096;
assign _029_ = ap_CS_fsm[24] ? grp_fu_739_p2 : ret_V_29_reg_1091;
assign _000_ = ap_CS_fsm[17] ? grp_fu_626_p2 : add_ln691_reg_1014;
assign _002_ = ap_rst ? 27'h0000001 : ap_NS_fsm;
assign icmp_ln768_fu_454_p2 = _205_ ? 1'h1 : 1'h0;
assign icmp_ln786_fu_460_p2 = _206_ ? 1'h1 : 1'h0;
assign icmp_ln851_1_fu_297_p2 = _052_ ? 1'h1 : 1'h0;
assign icmp_ln851_2_fu_310_p2 = _053_ ? 1'h1 : 1'h0;
assign icmp_ln851_fu_694_p2 = _054_ ? 1'h1 : 1'h0;
assign lhs_fu_396_p3 = op_4 ? 7'h40 : 7'h00;
assign op_14_V_fu_590_p3 = and_ln785_1_fu_585_p2 ? p_Val2_s_reg_921 : select_ln340_reg_971;
assign ret_V_20_fu_725_p3 = ret_V_19_reg_1024[9] ? select_ln850_fu_720_p3 : ret_V_2_reg_1029;
assign ret_V_22_fu_333_p3 = ret_V_21_reg_815[4] ? select_ln850_1_fu_328_p3 : ret_V_6_reg_820;
assign ret_V_24_fu_352_p3 = ret_V_23_reg_832[3] ? select_ln850_2_fu_347_p3 : sext_ln831_reg_852;
assign ret_V_27_fu_647_p3 = ret_V_26_reg_1002[33] ? select_ln850_3_fu_641_p3 : ret_V_16_cast_reg_1007;
assign select_ln1192_fu_490_p3 = ret_V_fu_404_p2[6] ? 7'h7f : 7'h00;
assign select_ln1196_fu_271_p3 = tmp_6_reg_783 ? 3'h4 : 3'h0;
assign select_ln1497_fu_386_p3 = tmp_reg_773 ? trunc_ln728_reg_894 : { 3'h0, trunc_ln1497_reg_889 };
assign select_ln340_fu_549_p3 = and_ln340_fu_543_p2 ? p_Val2_s_reg_921 : 2'h0;
assign select_ln850_1_fu_328_p3 = icmp_ln851_1_reg_847 ? ret_V_6_reg_820 : ret_V_7_reg_864;
assign select_ln850_2_fu_347_p3 = icmp_ln851_2_reg_859 ? sext_ln831_reg_852 : ret_V_11_reg_869;
assign select_ln850_3_fu_641_p3 = op_14_V_reg_981[0] ? add_ln691_reg_1014 : ret_V_16_cast_reg_1007;
assign select_ln850_fu_720_p3 = icmp_ln851_reg_1046 ? ret_V_2_reg_1029 : ret_V_3_reg_1056;
assign ret_V_23_fu_278_p2 = { 1'h0, select_ln1196_fu_271_p3 } ^ op_3;
assign ap_CS_fsm_state1 = ap_CS_fsm[0];
assign ap_CS_fsm_state10 = ap_CS_fsm[9];
assign ap_CS_fsm_state11 = ap_CS_fsm[10];
assign ap_CS_fsm_state12 = ap_CS_fsm[11];
assign ap_CS_fsm_state13 = ap_CS_fsm[12];
assign ap_CS_fsm_state14 = ap_CS_fsm[13];
assign ap_CS_fsm_state15 = ap_CS_fsm[14];
assign ap_CS_fsm_state16 = ap_CS_fsm[15];
assign ap_CS_fsm_state17 = ap_CS_fsm[16];
assign ap_CS_fsm_state18 = ap_CS_fsm[17];
assign ap_CS_fsm_state19 = ap_CS_fsm[18];
assign ap_CS_fsm_state2 = ap_CS_fsm[1];
assign ap_CS_fsm_state20 = ap_CS_fsm[19];
assign ap_CS_fsm_state21 = ap_CS_fsm[20];
assign ap_CS_fsm_state22 = ap_CS_fsm[21];
assign ap_CS_fsm_state23 = ap_CS_fsm[22];
assign ap_CS_fsm_state24 = ap_CS_fsm[23];
assign ap_CS_fsm_state25 = ap_CS_fsm[24];
assign ap_CS_fsm_state26 = ap_CS_fsm[25];
assign ap_CS_fsm_state27 = ap_CS_fsm[26];
assign ap_CS_fsm_state3 = ap_CS_fsm[2];
assign ap_CS_fsm_state4 = ap_CS_fsm[3];
assign ap_CS_fsm_state5 = ap_CS_fsm[4];
assign ap_CS_fsm_state6 = ap_CS_fsm[5];
assign ap_CS_fsm_state7 = ap_CS_fsm[6];
assign ap_CS_fsm_state8 = ap_CS_fsm[7];
assign ap_CS_fsm_state9 = ap_CS_fsm[8];
assign ap_done = op_29_ap_vld;
assign ap_ready = op_29_ap_vld;
assign conv_i2826_fu_228_p1 = { 31'h00000000, op_0[1] };
assign empty_fu_392_p1 = op_7[6:0];
assign grp_fu_211_p1 = { op_6[3], op_6 };
assign grp_fu_232_p1 = { op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6 };
assign grp_fu_241_p1 = { sub_ln1497_reg_778[4], sub_ln1497_reg_778[4], sub_ln1497_reg_778[4], sub_ln1497_reg_778[4], sub_ln1497_reg_778[4], sub_ln1497_reg_778[4], sub_ln1497_reg_778[4], sub_ln1497_reg_778[4], sub_ln1497_reg_778[4], sub_ln1497_reg_778[4], sub_ln1497_reg_778[4], sub_ln1497_reg_778[4], sub_ln1497_reg_778[4], sub_ln1497_reg_778[4], sub_ln1497_reg_778[4], sub_ln1497_reg_778[4], sub_ln1497_reg_778[4], sub_ln1497_reg_778[4], sub_ln1497_reg_778[4], sub_ln1497_reg_778[4], sub_ln1497_reg_778[4], sub_ln1497_reg_778[4], sub_ln1497_reg_778[4], sub_ln1497_reg_778[4], sub_ln1497_reg_778[4], sub_ln1497_reg_778[4], sub_ln1497_reg_778[4], sub_ln1497_reg_778 };
assign grp_fu_251_p1 = { op_3[3], op_3 };
assign grp_fu_315_p0 = { ret_V_10_reg_837[1], ret_V_10_reg_837 };
assign grp_fu_377_p0 = { 2'h0, ret_V_24_reg_879[2], ret_V_24_reg_879 };
assign grp_fu_377_p1 = { ret_V_22_reg_874[2], ret_V_22_reg_874[2], ret_V_22_reg_874[2], ret_V_22_reg_874 };
assign grp_fu_484_p0 = { op_20_V_reg_909, 4'h0 };
assign grp_fu_484_p1 = { select_ln1497_reg_904[3], select_ln1497_reg_904[3], select_ln1497_reg_904, 4'h0 };
assign grp_fu_559_p0 = { op_22_V_reg_966[5], op_22_V_reg_966 };
assign grp_fu_610_p0 = { ret_V_25_reg_987[6], ret_V_25_reg_987[6], ret_V_25_reg_987[6], ret_V_25_reg_987[6], ret_V_25_reg_987[6], ret_V_25_reg_987[6], ret_V_25_reg_987[6], ret_V_25_reg_987[6], ret_V_25_reg_987[6], ret_V_25_reg_987[6], ret_V_25_reg_987[6], ret_V_25_reg_987[6], ret_V_25_reg_987[6], ret_V_25_reg_987[6], ret_V_25_reg_987[6], ret_V_25_reg_987[6], ret_V_25_reg_987[6], ret_V_25_reg_987[6], ret_V_25_reg_987[6], ret_V_25_reg_987[6], ret_V_25_reg_987[6], ret_V_25_reg_987[6], ret_V_25_reg_987[6], ret_V_25_reg_987[6], ret_V_25_reg_987[6], ret_V_25_reg_987[6], ret_V_25_reg_987, 1'h0 };
assign grp_fu_610_p1 = { op_14_V_reg_981[1], op_14_V_reg_981[1], op_14_V_reg_981[1], op_14_V_reg_981[1], op_14_V_reg_981[1], op_14_V_reg_981[1], op_14_V_reg_981[1], op_14_V_reg_981[1], op_14_V_reg_981[1], op_14_V_reg_981[1], op_14_V_reg_981[1], op_14_V_reg_981[1], op_14_V_reg_981[1], op_14_V_reg_981[1], op_14_V_reg_981[1], op_14_V_reg_981[1], op_14_V_reg_981[1], op_14_V_reg_981[1], op_14_V_reg_981[1], op_14_V_reg_981[1], op_14_V_reg_981[1], op_14_V_reg_981[1], op_14_V_reg_981[1], op_14_V_reg_981[1], op_14_V_reg_981[1], op_14_V_reg_981[1], op_14_V_reg_981[1], op_14_V_reg_981[1], op_14_V_reg_981[1], op_14_V_reg_981[1], op_14_V_reg_981[1], op_14_V_reg_981[1], op_14_V_reg_981 };
assign grp_fu_689_p1 = { op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15 };
assign grp_fu_708_p1 = { op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16 };
assign grp_fu_739_p1 = { op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17 };
assign grp_fu_748_p0 = { ret_V_20_reg_1066[7], ret_V_20_reg_1066 };
assign grp_fu_748_p1 = { op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18 };
assign grp_fu_757_p0 = { add_ln69_reg_1096[8], add_ln69_reg_1096[8], add_ln69_reg_1096[8], add_ln69_reg_1096[8], add_ln69_reg_1096[8], add_ln69_reg_1096[8], add_ln69_reg_1096[8], add_ln69_reg_1096[8], add_ln69_reg_1096[8], add_ln69_reg_1096[8], add_ln69_reg_1096[8], add_ln69_reg_1096[8], add_ln69_reg_1096[8], add_ln69_reg_1096[8], add_ln69_reg_1096[8], add_ln69_reg_1096[8], add_ln69_reg_1096[8], add_ln69_reg_1096[8], add_ln69_reg_1096[8], add_ln69_reg_1096[8], add_ln69_reg_1096[8], add_ln69_reg_1096[8], add_ln69_reg_1096[8], add_ln69_reg_1096 };
assign lhs_fu_396_p0 = op_4;
assign op_11_V_fu_466_p3 = { select_ln1497_reg_904, 4'h0 };
assign op_13_V_fu_410_p3 = ret_V_fu_404_p2[6];
assign op_29 = grp_fu_757_p2;
assign p_Result_1_fu_321_p3 = ret_V_21_reg_815[4];
assign p_Result_2_fu_340_p3 = ret_V_23_reg_832[3];
assign p_Result_3_fu_631_p3 = ret_V_26_reg_1002[33];
assign p_Result_s_14_fu_713_p3 = ret_V_19_reg_1024[9];
assign p_Result_s_fu_444_p4 = op_7[15:7];
assign ret_V_23_fu_278_p1 = op_3;
assign rhs_fu_657_p3 = { op_12, 2'h0 };
assign sext_ln1497_fu_199_p0 = op_6;
assign sext_ln545_fu_225_p0 = op_6;
assign sext_ln69_3_fu_370_p1 = { ret_V_24_reg_879[2], ret_V_24_reg_879 };
assign sext_ln703_1_fu_247_p0 = op_3;
assign sext_ln703_fu_654_p0 = op_3;
assign sext_ln703_fu_654_p1 = { op_3[3], op_3[3], op_3[3], op_3[3], op_3[3], op_3[3], op_3 };
assign sext_ln831_fu_307_p1 = { ret_V_10_reg_837[1], ret_V_10_reg_837 };
assign tmp_6_fu_217_p3 = op_0[1];
assign tmp_8_fu_599_p3 = { ret_V_25_reg_987, 1'h0 };
assign tmp_fu_203_p1 = op_6;
assign trunc_ln1497_fu_362_p1 = grp_fu_232_p2[0];
assign trunc_ln728_fu_366_p1 = grp_fu_241_p2[3:0];
assign trunc_ln851_1_fu_267_p1 = grp_fu_251_p2[1:0];
assign trunc_ln851_2_fu_293_p1 = ret_V_23_fu_278_p2[1:0];
assign trunc_ln851_3_fu_638_p1 = op_14_V_reg_981[0];
assign trunc_ln851_fu_681_p1 = ret_V_19_fu_665_p2[1:0];
assign zext_ln1497_fu_383_p1 = { 3'h0, trunc_ln1497_reg_889 };
assign \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_0_U.ain_s0  = \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_0_U.a ;
assign \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_0_U.s  = { \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_0_U.fas_s2 , \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_0_U.sum_s1  };
assign \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_0_U.u2.a  = \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_0_U.ain_s1 ;
assign \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_0_U.u2.b  = \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_0_U.bin_s1 ;
assign \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_0_U.u2.cin  = \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_0_U.carry_s1 ;
assign \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_0_U.facout_s2  = \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_0_U.u2.cout ;
assign \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_0_U.fas_s2  = \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_0_U.u2.s ;
assign \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_0_U.u1.a  = \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_0_U.a [1:0];
assign \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_0_U.u1.b  = \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_0_U.bin_s0 [1:0];
assign \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_0_U.u1.cin  = 1'h1;
assign \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_0_U.facout_s1  = \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_0_U.u1.cout ;
assign \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_0_U.fas_s1  = \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_0_U.u1.s ;
assign \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_0_U.a  = \sub_5ns_5s_5_2_1_U4.din0 ;
assign \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_0_U.b  = \sub_5ns_5s_5_2_1_U4.din1 ;
assign \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_0_U.ce  = \sub_5ns_5s_5_2_1_U4.ce ;
assign \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_0_U.clk  = \sub_5ns_5s_5_2_1_U4.clk ;
assign \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_0_U.reset  = \sub_5ns_5s_5_2_1_U4.reset ;
assign \sub_5ns_5s_5_2_1_U4.dout  = \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_0_U.s ;
assign \sub_5ns_5s_5_2_1_U4.ce  = 1'h1;
assign \sub_5ns_5s_5_2_1_U4.clk  = ap_clk;
assign \sub_5ns_5s_5_2_1_U4.din0  = 5'h00;
assign \sub_5ns_5s_5_2_1_U4.din1  = { op_3[3], op_3 };
assign grp_fu_251_p2 = \sub_5ns_5s_5_2_1_U4.dout ;
assign \sub_5ns_5s_5_2_1_U4.reset  = ap_rst;
assign \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.ain_s0  = \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.a ;
assign \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.s  = { \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.fas_s2 , \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.sum_s1  };
assign \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.u2.a  = \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.ain_s1 ;
assign \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.u2.b  = \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.bin_s1 ;
assign \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.u2.cin  = \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.carry_s1 ;
assign \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.facout_s2  = \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.u2.cout ;
assign \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.fas_s2  = \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.u2.s ;
assign \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.u1.a  = \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.a [1:0];
assign \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.u1.b  = \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.bin_s0 [1:0];
assign \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.u1.cin  = 1'h1;
assign \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.facout_s1  = \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.u1.cout ;
assign \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.fas_s1  = \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.u1.s ;
assign \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.a  = \sub_5ns_5s_5_2_1_U1.din0 ;
assign \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.b  = \sub_5ns_5s_5_2_1_U1.din1 ;
assign \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.ce  = \sub_5ns_5s_5_2_1_U1.ce ;
assign \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.clk  = \sub_5ns_5s_5_2_1_U1.clk ;
assign \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.reset  = \sub_5ns_5s_5_2_1_U1.reset ;
assign \sub_5ns_5s_5_2_1_U1.dout  = \sub_5ns_5s_5_2_1_U1.top_sub_5ns_5s_5_2_1_Adder_0_U.s ;
assign \sub_5ns_5s_5_2_1_U1.ce  = 1'h1;
assign \sub_5ns_5s_5_2_1_U1.clk  = ap_clk;
assign \sub_5ns_5s_5_2_1_U1.din0  = 5'h00;
assign \sub_5ns_5s_5_2_1_U1.din1  = { op_6[3], op_6 };
assign grp_fu_211_p2 = \sub_5ns_5s_5_2_1_U1.dout ;
assign \sub_5ns_5s_5_2_1_U1.reset  = ap_rst;
assign \shl_32ns_32s_32_7_1_U3.din1_cast  = \shl_32ns_32s_32_7_1_U3.din1 ;
assign \shl_32ns_32s_32_7_1_U3.din1_mask  = 32'd31;
assign \shl_32ns_32s_32_7_1_U3.ce  = 1'h1;
assign \shl_32ns_32s_32_7_1_U3.clk  = ap_clk;
assign \shl_32ns_32s_32_7_1_U3.din0  = { 31'h00000000, op_0[1] };
assign \shl_32ns_32s_32_7_1_U3.din1  = { sub_ln1497_reg_778[4], sub_ln1497_reg_778[4], sub_ln1497_reg_778[4], sub_ln1497_reg_778[4], sub_ln1497_reg_778[4], sub_ln1497_reg_778[4], sub_ln1497_reg_778[4], sub_ln1497_reg_778[4], sub_ln1497_reg_778[4], sub_ln1497_reg_778[4], sub_ln1497_reg_778[4], sub_ln1497_reg_778[4], sub_ln1497_reg_778[4], sub_ln1497_reg_778[4], sub_ln1497_reg_778[4], sub_ln1497_reg_778[4], sub_ln1497_reg_778[4], sub_ln1497_reg_778[4], sub_ln1497_reg_778[4], sub_ln1497_reg_778[4], sub_ln1497_reg_778[4], sub_ln1497_reg_778[4], sub_ln1497_reg_778[4], sub_ln1497_reg_778[4], sub_ln1497_reg_778[4], sub_ln1497_reg_778[4], sub_ln1497_reg_778[4], sub_ln1497_reg_778 };
assign grp_fu_241_p2 = \shl_32ns_32s_32_7_1_U3.dout ;
assign \shl_32ns_32s_32_7_1_U3.reset  = ap_rst;
assign \lshr_32ns_32s_32_7_1_U2.din1_cast  = \lshr_32ns_32s_32_7_1_U2.din1 ;
assign \lshr_32ns_32s_32_7_1_U2.din1_mask  = 32'd31;
assign \lshr_32ns_32s_32_7_1_U2.ce  = 1'h1;
assign \lshr_32ns_32s_32_7_1_U2.clk  = ap_clk;
assign \lshr_32ns_32s_32_7_1_U2.din0  = { 31'h00000000, op_0[1] };
assign \lshr_32ns_32s_32_7_1_U2.din1  = { op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6[3], op_6 };
assign grp_fu_232_p2 = \lshr_32ns_32s_32_7_1_U2.dout ;
assign \lshr_32ns_32s_32_7_1_U2.reset  = ap_rst;
assign \add_9s_9s_9_2_1_U16.top_add_9s_9s_9_2_1_Adder_10_U.ain_s0  = \add_9s_9s_9_2_1_U16.top_add_9s_9s_9_2_1_Adder_10_U.a ;
assign \add_9s_9s_9_2_1_U16.top_add_9s_9s_9_2_1_Adder_10_U.bin_s0  = \add_9s_9s_9_2_1_U16.top_add_9s_9s_9_2_1_Adder_10_U.b ;
assign \add_9s_9s_9_2_1_U16.top_add_9s_9s_9_2_1_Adder_10_U.s  = { \add_9s_9s_9_2_1_U16.top_add_9s_9s_9_2_1_Adder_10_U.fas_s2 , \add_9s_9s_9_2_1_U16.top_add_9s_9s_9_2_1_Adder_10_U.sum_s1  };
assign \add_9s_9s_9_2_1_U16.top_add_9s_9s_9_2_1_Adder_10_U.u2.a  = \add_9s_9s_9_2_1_U16.top_add_9s_9s_9_2_1_Adder_10_U.ain_s1 ;
assign \add_9s_9s_9_2_1_U16.top_add_9s_9s_9_2_1_Adder_10_U.u2.b  = \add_9s_9s_9_2_1_U16.top_add_9s_9s_9_2_1_Adder_10_U.bin_s1 ;
assign \add_9s_9s_9_2_1_U16.top_add_9s_9s_9_2_1_Adder_10_U.u2.cin  = \add_9s_9s_9_2_1_U16.top_add_9s_9s_9_2_1_Adder_10_U.carry_s1 ;
assign \add_9s_9s_9_2_1_U16.top_add_9s_9s_9_2_1_Adder_10_U.facout_s2  = \add_9s_9s_9_2_1_U16.top_add_9s_9s_9_2_1_Adder_10_U.u2.cout ;
assign \add_9s_9s_9_2_1_U16.top_add_9s_9s_9_2_1_Adder_10_U.fas_s2  = \add_9s_9s_9_2_1_U16.top_add_9s_9s_9_2_1_Adder_10_U.u2.s ;
assign \add_9s_9s_9_2_1_U16.top_add_9s_9s_9_2_1_Adder_10_U.u1.a  = \add_9s_9s_9_2_1_U16.top_add_9s_9s_9_2_1_Adder_10_U.a [3:0];
assign \add_9s_9s_9_2_1_U16.top_add_9s_9s_9_2_1_Adder_10_U.u1.b  = \add_9s_9s_9_2_1_U16.top_add_9s_9s_9_2_1_Adder_10_U.b [3:0];
assign \add_9s_9s_9_2_1_U16.top_add_9s_9s_9_2_1_Adder_10_U.u1.cin  = 1'h0;
assign \add_9s_9s_9_2_1_U16.top_add_9s_9s_9_2_1_Adder_10_U.facout_s1  = \add_9s_9s_9_2_1_U16.top_add_9s_9s_9_2_1_Adder_10_U.u1.cout ;
assign \add_9s_9s_9_2_1_U16.top_add_9s_9s_9_2_1_Adder_10_U.fas_s1  = \add_9s_9s_9_2_1_U16.top_add_9s_9s_9_2_1_Adder_10_U.u1.s ;
assign \add_9s_9s_9_2_1_U16.top_add_9s_9s_9_2_1_Adder_10_U.a  = \add_9s_9s_9_2_1_U16.din0 ;
assign \add_9s_9s_9_2_1_U16.top_add_9s_9s_9_2_1_Adder_10_U.b  = \add_9s_9s_9_2_1_U16.din1 ;
assign \add_9s_9s_9_2_1_U16.top_add_9s_9s_9_2_1_Adder_10_U.ce  = \add_9s_9s_9_2_1_U16.ce ;
assign \add_9s_9s_9_2_1_U16.top_add_9s_9s_9_2_1_Adder_10_U.clk  = \add_9s_9s_9_2_1_U16.clk ;
assign \add_9s_9s_9_2_1_U16.top_add_9s_9s_9_2_1_Adder_10_U.reset  = \add_9s_9s_9_2_1_U16.reset ;
assign \add_9s_9s_9_2_1_U16.dout  = \add_9s_9s_9_2_1_U16.top_add_9s_9s_9_2_1_Adder_10_U.s ;
assign \add_9s_9s_9_2_1_U16.ce  = 1'h1;
assign \add_9s_9s_9_2_1_U16.clk  = ap_clk;
assign \add_9s_9s_9_2_1_U16.din0  = { ret_V_20_reg_1066[7], ret_V_20_reg_1066 };
assign \add_9s_9s_9_2_1_U16.din1  = { op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18 };
assign grp_fu_748_p2 = \add_9s_9s_9_2_1_U16.dout ;
assign \add_9s_9s_9_2_1_U16.reset  = ap_rst;
assign \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_9_U.ain_s0  = \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_9_U.a ;
assign \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_9_U.bin_s0  = \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_9_U.b ;
assign \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_9_U.s  = { \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_9_U.fas_s2 , \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_9_U.sum_s1  };
assign \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_9_U.u2.a  = \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_9_U.ain_s1 ;
assign \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_9_U.u2.b  = \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_9_U.bin_s1 ;
assign \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_9_U.u2.cin  = \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_9_U.carry_s1 ;
assign \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_9_U.facout_s2  = \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_9_U.u2.cout ;
assign \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_9_U.fas_s2  = \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_9_U.u2.s ;
assign \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_9_U.u1.a  = \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_9_U.a [3:0];
assign \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_9_U.u1.b  = \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_9_U.b [3:0];
assign \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_9_U.u1.cin  = 1'h0;
assign \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_9_U.facout_s1  = \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_9_U.u1.cout ;
assign \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_9_U.fas_s1  = \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_9_U.u1.s ;
assign \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_9_U.a  = \add_8ns_8ns_8_2_1_U13.din0 ;
assign \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_9_U.b  = \add_8ns_8ns_8_2_1_U13.din1 ;
assign \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_9_U.ce  = \add_8ns_8ns_8_2_1_U13.ce ;
assign \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_9_U.clk  = \add_8ns_8ns_8_2_1_U13.clk ;
assign \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_9_U.reset  = \add_8ns_8ns_8_2_1_U13.reset ;
assign \add_8ns_8ns_8_2_1_U13.dout  = \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_9_U.s ;
assign \add_8ns_8ns_8_2_1_U13.ce  = 1'h1;
assign \add_8ns_8ns_8_2_1_U13.clk  = ap_clk;
assign \add_8ns_8ns_8_2_1_U13.din0  = ret_V_2_reg_1029;
assign \add_8ns_8ns_8_2_1_U13.din1  = 8'h01;
assign grp_fu_699_p2 = \add_8ns_8ns_8_2_1_U13.dout ;
assign \add_8ns_8ns_8_2_1_U13.reset  = ap_rst;
assign \add_7s_7ns_7_2_1_U9.top_add_7s_7ns_7_2_1_Adder_5_U.ain_s0  = \add_7s_7ns_7_2_1_U9.top_add_7s_7ns_7_2_1_Adder_5_U.a ;
assign \add_7s_7ns_7_2_1_U9.top_add_7s_7ns_7_2_1_Adder_5_U.bin_s0  = \add_7s_7ns_7_2_1_U9.top_add_7s_7ns_7_2_1_Adder_5_U.b ;
assign \add_7s_7ns_7_2_1_U9.top_add_7s_7ns_7_2_1_Adder_5_U.s  = { \add_7s_7ns_7_2_1_U9.top_add_7s_7ns_7_2_1_Adder_5_U.fas_s2 , \add_7s_7ns_7_2_1_U9.top_add_7s_7ns_7_2_1_Adder_5_U.sum_s1  };
assign \add_7s_7ns_7_2_1_U9.top_add_7s_7ns_7_2_1_Adder_5_U.u2.a  = \add_7s_7ns_7_2_1_U9.top_add_7s_7ns_7_2_1_Adder_5_U.ain_s1 ;
assign \add_7s_7ns_7_2_1_U9.top_add_7s_7ns_7_2_1_Adder_5_U.u2.b  = \add_7s_7ns_7_2_1_U9.top_add_7s_7ns_7_2_1_Adder_5_U.bin_s1 ;
assign \add_7s_7ns_7_2_1_U9.top_add_7s_7ns_7_2_1_Adder_5_U.u2.cin  = \add_7s_7ns_7_2_1_U9.top_add_7s_7ns_7_2_1_Adder_5_U.carry_s1 ;
assign \add_7s_7ns_7_2_1_U9.top_add_7s_7ns_7_2_1_Adder_5_U.facout_s2  = \add_7s_7ns_7_2_1_U9.top_add_7s_7ns_7_2_1_Adder_5_U.u2.cout ;
assign \add_7s_7ns_7_2_1_U9.top_add_7s_7ns_7_2_1_Adder_5_U.fas_s2  = \add_7s_7ns_7_2_1_U9.top_add_7s_7ns_7_2_1_Adder_5_U.u2.s ;
assign \add_7s_7ns_7_2_1_U9.top_add_7s_7ns_7_2_1_Adder_5_U.u1.a  = \add_7s_7ns_7_2_1_U9.top_add_7s_7ns_7_2_1_Adder_5_U.a [2:0];
assign \add_7s_7ns_7_2_1_U9.top_add_7s_7ns_7_2_1_Adder_5_U.u1.b  = \add_7s_7ns_7_2_1_U9.top_add_7s_7ns_7_2_1_Adder_5_U.b [2:0];
assign \add_7s_7ns_7_2_1_U9.top_add_7s_7ns_7_2_1_Adder_5_U.u1.cin  = 1'h0;
assign \add_7s_7ns_7_2_1_U9.top_add_7s_7ns_7_2_1_Adder_5_U.facout_s1  = \add_7s_7ns_7_2_1_U9.top_add_7s_7ns_7_2_1_Adder_5_U.u1.cout ;
assign \add_7s_7ns_7_2_1_U9.top_add_7s_7ns_7_2_1_Adder_5_U.fas_s1  = \add_7s_7ns_7_2_1_U9.top_add_7s_7ns_7_2_1_Adder_5_U.u1.s ;
assign \add_7s_7ns_7_2_1_U9.top_add_7s_7ns_7_2_1_Adder_5_U.a  = \add_7s_7ns_7_2_1_U9.din0 ;
assign \add_7s_7ns_7_2_1_U9.top_add_7s_7ns_7_2_1_Adder_5_U.b  = \add_7s_7ns_7_2_1_U9.din1 ;
assign \add_7s_7ns_7_2_1_U9.top_add_7s_7ns_7_2_1_Adder_5_U.ce  = \add_7s_7ns_7_2_1_U9.ce ;
assign \add_7s_7ns_7_2_1_U9.top_add_7s_7ns_7_2_1_Adder_5_U.clk  = \add_7s_7ns_7_2_1_U9.clk ;
assign \add_7s_7ns_7_2_1_U9.top_add_7s_7ns_7_2_1_Adder_5_U.reset  = \add_7s_7ns_7_2_1_U9.reset ;
assign \add_7s_7ns_7_2_1_U9.dout  = \add_7s_7ns_7_2_1_U9.top_add_7s_7ns_7_2_1_Adder_5_U.s ;
assign \add_7s_7ns_7_2_1_U9.ce  = 1'h1;
assign \add_7s_7ns_7_2_1_U9.clk  = ap_clk;
assign \add_7s_7ns_7_2_1_U9.din0  = { op_22_V_reg_966[5], op_22_V_reg_966 };
assign \add_7s_7ns_7_2_1_U9.din1  = select_ln1192_reg_955;
assign grp_fu_559_p2 = \add_7s_7ns_7_2_1_U9.dout ;
assign \add_7s_7ns_7_2_1_U9.reset  = ap_rst;
assign \add_6ns_6s_6_2_1_U7.top_add_6ns_6s_6_2_1_Adder_3_U.ain_s0  = \add_6ns_6s_6_2_1_U7.top_add_6ns_6s_6_2_1_Adder_3_U.a ;
assign \add_6ns_6s_6_2_1_U7.top_add_6ns_6s_6_2_1_Adder_3_U.bin_s0  = \add_6ns_6s_6_2_1_U7.top_add_6ns_6s_6_2_1_Adder_3_U.b ;
assign \add_6ns_6s_6_2_1_U7.top_add_6ns_6s_6_2_1_Adder_3_U.s  = { \add_6ns_6s_6_2_1_U7.top_add_6ns_6s_6_2_1_Adder_3_U.fas_s2 , \add_6ns_6s_6_2_1_U7.top_add_6ns_6s_6_2_1_Adder_3_U.sum_s1  };
assign \add_6ns_6s_6_2_1_U7.top_add_6ns_6s_6_2_1_Adder_3_U.u2.a  = \add_6ns_6s_6_2_1_U7.top_add_6ns_6s_6_2_1_Adder_3_U.ain_s1 ;
assign \add_6ns_6s_6_2_1_U7.top_add_6ns_6s_6_2_1_Adder_3_U.u2.b  = \add_6ns_6s_6_2_1_U7.top_add_6ns_6s_6_2_1_Adder_3_U.bin_s1 ;
assign \add_6ns_6s_6_2_1_U7.top_add_6ns_6s_6_2_1_Adder_3_U.u2.cin  = \add_6ns_6s_6_2_1_U7.top_add_6ns_6s_6_2_1_Adder_3_U.carry_s1 ;
assign \add_6ns_6s_6_2_1_U7.top_add_6ns_6s_6_2_1_Adder_3_U.facout_s2  = \add_6ns_6s_6_2_1_U7.top_add_6ns_6s_6_2_1_Adder_3_U.u2.cout ;
assign \add_6ns_6s_6_2_1_U7.top_add_6ns_6s_6_2_1_Adder_3_U.fas_s2  = \add_6ns_6s_6_2_1_U7.top_add_6ns_6s_6_2_1_Adder_3_U.u2.s ;
assign \add_6ns_6s_6_2_1_U7.top_add_6ns_6s_6_2_1_Adder_3_U.u1.a  = \add_6ns_6s_6_2_1_U7.top_add_6ns_6s_6_2_1_Adder_3_U.a [2:0];
assign \add_6ns_6s_6_2_1_U7.top_add_6ns_6s_6_2_1_Adder_3_U.u1.b  = \add_6ns_6s_6_2_1_U7.top_add_6ns_6s_6_2_1_Adder_3_U.b [2:0];
assign \add_6ns_6s_6_2_1_U7.top_add_6ns_6s_6_2_1_Adder_3_U.u1.cin  = 1'h0;
assign \add_6ns_6s_6_2_1_U7.top_add_6ns_6s_6_2_1_Adder_3_U.facout_s1  = \add_6ns_6s_6_2_1_U7.top_add_6ns_6s_6_2_1_Adder_3_U.u1.cout ;
assign \add_6ns_6s_6_2_1_U7.top_add_6ns_6s_6_2_1_Adder_3_U.fas_s1  = \add_6ns_6s_6_2_1_U7.top_add_6ns_6s_6_2_1_Adder_3_U.u1.s ;
assign \add_6ns_6s_6_2_1_U7.top_add_6ns_6s_6_2_1_Adder_3_U.a  = \add_6ns_6s_6_2_1_U7.din0 ;
assign \add_6ns_6s_6_2_1_U7.top_add_6ns_6s_6_2_1_Adder_3_U.b  = \add_6ns_6s_6_2_1_U7.din1 ;
assign \add_6ns_6s_6_2_1_U7.top_add_6ns_6s_6_2_1_Adder_3_U.ce  = \add_6ns_6s_6_2_1_U7.ce ;
assign \add_6ns_6s_6_2_1_U7.top_add_6ns_6s_6_2_1_Adder_3_U.clk  = \add_6ns_6s_6_2_1_U7.clk ;
assign \add_6ns_6s_6_2_1_U7.top_add_6ns_6s_6_2_1_Adder_3_U.reset  = \add_6ns_6s_6_2_1_U7.reset ;
assign \add_6ns_6s_6_2_1_U7.dout  = \add_6ns_6s_6_2_1_U7.top_add_6ns_6s_6_2_1_Adder_3_U.s ;
assign \add_6ns_6s_6_2_1_U7.ce  = 1'h1;
assign \add_6ns_6s_6_2_1_U7.clk  = ap_clk;
assign \add_6ns_6s_6_2_1_U7.din0  = { 2'h0, ret_V_24_reg_879[2], ret_V_24_reg_879 };
assign \add_6ns_6s_6_2_1_U7.din1  = { ret_V_22_reg_874[2], ret_V_22_reg_874[2], ret_V_22_reg_874[2], ret_V_22_reg_874 };
assign grp_fu_377_p2 = \add_6ns_6s_6_2_1_U7.dout ;
assign \add_6ns_6s_6_2_1_U7.reset  = ap_rst;
assign \add_3s_3ns_3_2_1_U6.top_add_3s_3ns_3_2_1_Adder_2_U.ain_s0  = \add_3s_3ns_3_2_1_U6.top_add_3s_3ns_3_2_1_Adder_2_U.a ;
assign \add_3s_3ns_3_2_1_U6.top_add_3s_3ns_3_2_1_Adder_2_U.bin_s0  = \add_3s_3ns_3_2_1_U6.top_add_3s_3ns_3_2_1_Adder_2_U.b ;
assign \add_3s_3ns_3_2_1_U6.top_add_3s_3ns_3_2_1_Adder_2_U.s  = { \add_3s_3ns_3_2_1_U6.top_add_3s_3ns_3_2_1_Adder_2_U.fas_s2 , \add_3s_3ns_3_2_1_U6.top_add_3s_3ns_3_2_1_Adder_2_U.sum_s1  };
assign \add_3s_3ns_3_2_1_U6.top_add_3s_3ns_3_2_1_Adder_2_U.u2.a  = \add_3s_3ns_3_2_1_U6.top_add_3s_3ns_3_2_1_Adder_2_U.ain_s1 ;
assign \add_3s_3ns_3_2_1_U6.top_add_3s_3ns_3_2_1_Adder_2_U.u2.b  = \add_3s_3ns_3_2_1_U6.top_add_3s_3ns_3_2_1_Adder_2_U.bin_s1 ;
assign \add_3s_3ns_3_2_1_U6.top_add_3s_3ns_3_2_1_Adder_2_U.u2.cin  = \add_3s_3ns_3_2_1_U6.top_add_3s_3ns_3_2_1_Adder_2_U.carry_s1 ;
assign \add_3s_3ns_3_2_1_U6.top_add_3s_3ns_3_2_1_Adder_2_U.facout_s2  = \add_3s_3ns_3_2_1_U6.top_add_3s_3ns_3_2_1_Adder_2_U.u2.cout ;
assign \add_3s_3ns_3_2_1_U6.top_add_3s_3ns_3_2_1_Adder_2_U.fas_s2  = \add_3s_3ns_3_2_1_U6.top_add_3s_3ns_3_2_1_Adder_2_U.u2.s ;
assign \add_3s_3ns_3_2_1_U6.top_add_3s_3ns_3_2_1_Adder_2_U.u1.a  = \add_3s_3ns_3_2_1_U6.top_add_3s_3ns_3_2_1_Adder_2_U.a [0];
assign \add_3s_3ns_3_2_1_U6.top_add_3s_3ns_3_2_1_Adder_2_U.u1.b  = \add_3s_3ns_3_2_1_U6.top_add_3s_3ns_3_2_1_Adder_2_U.b [0];
assign \add_3s_3ns_3_2_1_U6.top_add_3s_3ns_3_2_1_Adder_2_U.u1.cin  = 1'h0;
assign \add_3s_3ns_3_2_1_U6.top_add_3s_3ns_3_2_1_Adder_2_U.facout_s1  = \add_3s_3ns_3_2_1_U6.top_add_3s_3ns_3_2_1_Adder_2_U.u1.cout ;
assign \add_3s_3ns_3_2_1_U6.top_add_3s_3ns_3_2_1_Adder_2_U.fas_s1  = \add_3s_3ns_3_2_1_U6.top_add_3s_3ns_3_2_1_Adder_2_U.u1.s ;
assign \add_3s_3ns_3_2_1_U6.top_add_3s_3ns_3_2_1_Adder_2_U.a  = \add_3s_3ns_3_2_1_U6.din0 ;
assign \add_3s_3ns_3_2_1_U6.top_add_3s_3ns_3_2_1_Adder_2_U.b  = \add_3s_3ns_3_2_1_U6.din1 ;
assign \add_3s_3ns_3_2_1_U6.top_add_3s_3ns_3_2_1_Adder_2_U.ce  = \add_3s_3ns_3_2_1_U6.ce ;
assign \add_3s_3ns_3_2_1_U6.top_add_3s_3ns_3_2_1_Adder_2_U.clk  = \add_3s_3ns_3_2_1_U6.clk ;
assign \add_3s_3ns_3_2_1_U6.top_add_3s_3ns_3_2_1_Adder_2_U.reset  = \add_3s_3ns_3_2_1_U6.reset ;
assign \add_3s_3ns_3_2_1_U6.dout  = \add_3s_3ns_3_2_1_U6.top_add_3s_3ns_3_2_1_Adder_2_U.s ;
assign \add_3s_3ns_3_2_1_U6.ce  = 1'h1;
assign \add_3s_3ns_3_2_1_U6.clk  = ap_clk;
assign \add_3s_3ns_3_2_1_U6.din0  = { ret_V_10_reg_837[1], ret_V_10_reg_837 };
assign \add_3s_3ns_3_2_1_U6.din1  = 3'h1;
assign grp_fu_315_p2 = \add_3s_3ns_3_2_1_U6.dout ;
assign \add_3s_3ns_3_2_1_U6.reset  = ap_rst;
assign \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_1_U.ain_s0  = \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_1_U.a ;
assign \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_1_U.bin_s0  = \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_1_U.b ;
assign \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_1_U.s  = { \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_1_U.fas_s2 , \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_1_U.sum_s1  };
assign \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_1_U.u2.a  = \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_1_U.ain_s1 ;
assign \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_1_U.u2.b  = \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_1_U.bin_s1 ;
assign \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_1_U.u2.cin  = \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_1_U.carry_s1 ;
assign \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_1_U.facout_s2  = \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_1_U.u2.cout ;
assign \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_1_U.fas_s2  = \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_1_U.u2.s ;
assign \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_1_U.u1.a  = \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_1_U.a [0];
assign \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_1_U.u1.b  = \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_1_U.b [0];
assign \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_1_U.u1.cin  = 1'h0;
assign \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_1_U.facout_s1  = \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_1_U.u1.cout ;
assign \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_1_U.fas_s1  = \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_1_U.u1.s ;
assign \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_1_U.a  = \add_3ns_3ns_3_2_1_U5.din0 ;
assign \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_1_U.b  = \add_3ns_3ns_3_2_1_U5.din1 ;
assign \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_1_U.ce  = \add_3ns_3ns_3_2_1_U5.ce ;
assign \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_1_U.clk  = \add_3ns_3ns_3_2_1_U5.clk ;
assign \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_1_U.reset  = \add_3ns_3ns_3_2_1_U5.reset ;
assign \add_3ns_3ns_3_2_1_U5.dout  = \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_1_U.s ;
assign \add_3ns_3ns_3_2_1_U5.ce  = 1'h1;
assign \add_3ns_3ns_3_2_1_U5.clk  = ap_clk;
assign \add_3ns_3ns_3_2_1_U5.din0  = ret_V_6_reg_820;
assign \add_3ns_3ns_3_2_1_U5.din1  = 3'h1;
assign grp_fu_302_p2 = \add_3ns_3ns_3_2_1_U5.dout ;
assign \add_3ns_3ns_3_2_1_U5.reset  = ap_rst;
assign \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_6_U.ain_s0  = \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_6_U.a ;
assign \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_6_U.bin_s0  = \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_6_U.b ;
assign \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_6_U.s  = { \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_6_U.fas_s2 , \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_6_U.sum_s1  };
assign \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_6_U.u2.a  = \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_6_U.ain_s1 ;
assign \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_6_U.u2.b  = \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_6_U.bin_s1 ;
assign \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_6_U.u2.cin  = \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_6_U.carry_s1 ;
assign \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_6_U.facout_s2  = \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_6_U.u2.cout ;
assign \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_6_U.fas_s2  = \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_6_U.u2.s ;
assign \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_6_U.u1.a  = \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_6_U.a [16:0];
assign \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_6_U.u1.b  = \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_6_U.b [16:0];
assign \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_6_U.u1.cin  = 1'h0;
assign \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_6_U.facout_s1  = \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_6_U.u1.cout ;
assign \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_6_U.fas_s1  = \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_6_U.u1.s ;
assign \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_6_U.a  = \add_34s_34s_34_2_1_U10.din0 ;
assign \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_6_U.b  = \add_34s_34s_34_2_1_U10.din1 ;
assign \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_6_U.ce  = \add_34s_34s_34_2_1_U10.ce ;
assign \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_6_U.clk  = \add_34s_34s_34_2_1_U10.clk ;
assign \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_6_U.reset  = \add_34s_34s_34_2_1_U10.reset ;
assign \add_34s_34s_34_2_1_U10.dout  = \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_6_U.s ;
assign \add_34s_34s_34_2_1_U10.ce  = 1'h1;
assign \add_34s_34s_34_2_1_U10.clk  = ap_clk;
assign \add_34s_34s_34_2_1_U10.din0  = { ret_V_25_reg_987[6], ret_V_25_reg_987[6], ret_V_25_reg_987[6], ret_V_25_reg_987[6], ret_V_25_reg_987[6], ret_V_25_reg_987[6], ret_V_25_reg_987[6], ret_V_25_reg_987[6], ret_V_25_reg_987[6], ret_V_25_reg_987[6], ret_V_25_reg_987[6], ret_V_25_reg_987[6], ret_V_25_reg_987[6], ret_V_25_reg_987[6], ret_V_25_reg_987[6], ret_V_25_reg_987[6], ret_V_25_reg_987[6], ret_V_25_reg_987[6], ret_V_25_reg_987[6], ret_V_25_reg_987[6], ret_V_25_reg_987[6], ret_V_25_reg_987[6], ret_V_25_reg_987[6], ret_V_25_reg_987[6], ret_V_25_reg_987[6], ret_V_25_reg_987[6], ret_V_25_reg_987, 1'h0 };
assign \add_34s_34s_34_2_1_U10.din1  = { op_14_V_reg_981[1], op_14_V_reg_981[1], op_14_V_reg_981[1], op_14_V_reg_981[1], op_14_V_reg_981[1], op_14_V_reg_981[1], op_14_V_reg_981[1], op_14_V_reg_981[1], op_14_V_reg_981[1], op_14_V_reg_981[1], op_14_V_reg_981[1], op_14_V_reg_981[1], op_14_V_reg_981[1], op_14_V_reg_981[1], op_14_V_reg_981[1], op_14_V_reg_981[1], op_14_V_reg_981[1], op_14_V_reg_981[1], op_14_V_reg_981[1], op_14_V_reg_981[1], op_14_V_reg_981[1], op_14_V_reg_981[1], op_14_V_reg_981[1], op_14_V_reg_981[1], op_14_V_reg_981[1], op_14_V_reg_981[1], op_14_V_reg_981[1], op_14_V_reg_981[1], op_14_V_reg_981[1], op_14_V_reg_981[1], op_14_V_reg_981[1], op_14_V_reg_981[1], op_14_V_reg_981 };
assign grp_fu_610_p2 = \add_34s_34s_34_2_1_U10.dout ;
assign \add_34s_34s_34_2_1_U10.reset  = ap_rst;
assign \add_32s_32ns_32_2_1_U17.top_add_32s_32ns_32_2_1_Adder_11_U.ain_s0  = \add_32s_32ns_32_2_1_U17.top_add_32s_32ns_32_2_1_Adder_11_U.a ;
assign \add_32s_32ns_32_2_1_U17.top_add_32s_32ns_32_2_1_Adder_11_U.bin_s0  = \add_32s_32ns_32_2_1_U17.top_add_32s_32ns_32_2_1_Adder_11_U.b ;
assign \add_32s_32ns_32_2_1_U17.top_add_32s_32ns_32_2_1_Adder_11_U.s  = { \add_32s_32ns_32_2_1_U17.top_add_32s_32ns_32_2_1_Adder_11_U.fas_s2 , \add_32s_32ns_32_2_1_U17.top_add_32s_32ns_32_2_1_Adder_11_U.sum_s1  };
assign \add_32s_32ns_32_2_1_U17.top_add_32s_32ns_32_2_1_Adder_11_U.u2.a  = \add_32s_32ns_32_2_1_U17.top_add_32s_32ns_32_2_1_Adder_11_U.ain_s1 ;
assign \add_32s_32ns_32_2_1_U17.top_add_32s_32ns_32_2_1_Adder_11_U.u2.b  = \add_32s_32ns_32_2_1_U17.top_add_32s_32ns_32_2_1_Adder_11_U.bin_s1 ;
assign \add_32s_32ns_32_2_1_U17.top_add_32s_32ns_32_2_1_Adder_11_U.u2.cin  = \add_32s_32ns_32_2_1_U17.top_add_32s_32ns_32_2_1_Adder_11_U.carry_s1 ;
assign \add_32s_32ns_32_2_1_U17.top_add_32s_32ns_32_2_1_Adder_11_U.facout_s2  = \add_32s_32ns_32_2_1_U17.top_add_32s_32ns_32_2_1_Adder_11_U.u2.cout ;
assign \add_32s_32ns_32_2_1_U17.top_add_32s_32ns_32_2_1_Adder_11_U.fas_s2  = \add_32s_32ns_32_2_1_U17.top_add_32s_32ns_32_2_1_Adder_11_U.u2.s ;
assign \add_32s_32ns_32_2_1_U17.top_add_32s_32ns_32_2_1_Adder_11_U.u1.a  = \add_32s_32ns_32_2_1_U17.top_add_32s_32ns_32_2_1_Adder_11_U.a [15:0];
assign \add_32s_32ns_32_2_1_U17.top_add_32s_32ns_32_2_1_Adder_11_U.u1.b  = \add_32s_32ns_32_2_1_U17.top_add_32s_32ns_32_2_1_Adder_11_U.b [15:0];
assign \add_32s_32ns_32_2_1_U17.top_add_32s_32ns_32_2_1_Adder_11_U.u1.cin  = 1'h0;
assign \add_32s_32ns_32_2_1_U17.top_add_32s_32ns_32_2_1_Adder_11_U.facout_s1  = \add_32s_32ns_32_2_1_U17.top_add_32s_32ns_32_2_1_Adder_11_U.u1.cout ;
assign \add_32s_32ns_32_2_1_U17.top_add_32s_32ns_32_2_1_Adder_11_U.fas_s1  = \add_32s_32ns_32_2_1_U17.top_add_32s_32ns_32_2_1_Adder_11_U.u1.s ;
assign \add_32s_32ns_32_2_1_U17.top_add_32s_32ns_32_2_1_Adder_11_U.a  = \add_32s_32ns_32_2_1_U17.din0 ;
assign \add_32s_32ns_32_2_1_U17.top_add_32s_32ns_32_2_1_Adder_11_U.b  = \add_32s_32ns_32_2_1_U17.din1 ;
assign \add_32s_32ns_32_2_1_U17.top_add_32s_32ns_32_2_1_Adder_11_U.ce  = \add_32s_32ns_32_2_1_U17.ce ;
assign \add_32s_32ns_32_2_1_U17.top_add_32s_32ns_32_2_1_Adder_11_U.clk  = \add_32s_32ns_32_2_1_U17.clk ;
assign \add_32s_32ns_32_2_1_U17.top_add_32s_32ns_32_2_1_Adder_11_U.reset  = \add_32s_32ns_32_2_1_U17.reset ;
assign \add_32s_32ns_32_2_1_U17.dout  = \add_32s_32ns_32_2_1_U17.top_add_32s_32ns_32_2_1_Adder_11_U.s ;
assign \add_32s_32ns_32_2_1_U17.ce  = 1'h1;
assign \add_32s_32ns_32_2_1_U17.clk  = ap_clk;
assign \add_32s_32ns_32_2_1_U17.din0  = { add_ln69_reg_1096[8], add_ln69_reg_1096[8], add_ln69_reg_1096[8], add_ln69_reg_1096[8], add_ln69_reg_1096[8], add_ln69_reg_1096[8], add_ln69_reg_1096[8], add_ln69_reg_1096[8], add_ln69_reg_1096[8], add_ln69_reg_1096[8], add_ln69_reg_1096[8], add_ln69_reg_1096[8], add_ln69_reg_1096[8], add_ln69_reg_1096[8], add_ln69_reg_1096[8], add_ln69_reg_1096[8], add_ln69_reg_1096[8], add_ln69_reg_1096[8], add_ln69_reg_1096[8], add_ln69_reg_1096[8], add_ln69_reg_1096[8], add_ln69_reg_1096[8], add_ln69_reg_1096[8], add_ln69_reg_1096 };
assign \add_32s_32ns_32_2_1_U17.din1  = ret_V_29_reg_1091;
assign grp_fu_757_p2 = \add_32s_32ns_32_2_1_U17.dout ;
assign \add_32s_32ns_32_2_1_U17.reset  = ap_rst;
assign \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_8_U.ain_s0  = \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_8_U.a ;
assign \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_8_U.bin_s0  = \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_8_U.b ;
assign \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_8_U.s  = { \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_8_U.fas_s2 , \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_8_U.sum_s1  };
assign \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_8_U.u2.a  = \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_8_U.ain_s1 ;
assign \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_8_U.u2.b  = \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_8_U.bin_s1 ;
assign \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_8_U.u2.cin  = \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_8_U.carry_s1 ;
assign \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_8_U.facout_s2  = \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_8_U.u2.cout ;
assign \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_8_U.fas_s2  = \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_8_U.u2.s ;
assign \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_8_U.u1.a  = \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_8_U.a [15:0];
assign \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_8_U.u1.b  = \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_8_U.b [15:0];
assign \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_8_U.u1.cin  = 1'h0;
assign \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_8_U.facout_s1  = \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_8_U.u1.cout ;
assign \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_8_U.fas_s1  = \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_8_U.u1.s ;
assign \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_8_U.a  = \add_32ns_32s_32_2_1_U15.din0 ;
assign \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_8_U.b  = \add_32ns_32s_32_2_1_U15.din1 ;
assign \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_8_U.ce  = \add_32ns_32s_32_2_1_U15.ce ;
assign \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_8_U.clk  = \add_32ns_32s_32_2_1_U15.clk ;
assign \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_8_U.reset  = \add_32ns_32s_32_2_1_U15.reset ;
assign \add_32ns_32s_32_2_1_U15.dout  = \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_8_U.s ;
assign \add_32ns_32s_32_2_1_U15.ce  = 1'h1;
assign \add_32ns_32s_32_2_1_U15.clk  = ap_clk;
assign \add_32ns_32s_32_2_1_U15.din0  = ret_V_28_reg_1071;
assign \add_32ns_32s_32_2_1_U15.din1  = { op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17 };
assign grp_fu_739_p2 = \add_32ns_32s_32_2_1_U15.dout ;
assign \add_32ns_32s_32_2_1_U15.reset  = ap_rst;
assign \add_32ns_32s_32_2_1_U14.top_add_32ns_32s_32_2_1_Adder_8_U.ain_s0  = \add_32ns_32s_32_2_1_U14.top_add_32ns_32s_32_2_1_Adder_8_U.a ;
assign \add_32ns_32s_32_2_1_U14.top_add_32ns_32s_32_2_1_Adder_8_U.bin_s0  = \add_32ns_32s_32_2_1_U14.top_add_32ns_32s_32_2_1_Adder_8_U.b ;
assign \add_32ns_32s_32_2_1_U14.top_add_32ns_32s_32_2_1_Adder_8_U.s  = { \add_32ns_32s_32_2_1_U14.top_add_32ns_32s_32_2_1_Adder_8_U.fas_s2 , \add_32ns_32s_32_2_1_U14.top_add_32ns_32s_32_2_1_Adder_8_U.sum_s1  };
assign \add_32ns_32s_32_2_1_U14.top_add_32ns_32s_32_2_1_Adder_8_U.u2.a  = \add_32ns_32s_32_2_1_U14.top_add_32ns_32s_32_2_1_Adder_8_U.ain_s1 ;
assign \add_32ns_32s_32_2_1_U14.top_add_32ns_32s_32_2_1_Adder_8_U.u2.b  = \add_32ns_32s_32_2_1_U14.top_add_32ns_32s_32_2_1_Adder_8_U.bin_s1 ;
assign \add_32ns_32s_32_2_1_U14.top_add_32ns_32s_32_2_1_Adder_8_U.u2.cin  = \add_32ns_32s_32_2_1_U14.top_add_32ns_32s_32_2_1_Adder_8_U.carry_s1 ;
assign \add_32ns_32s_32_2_1_U14.top_add_32ns_32s_32_2_1_Adder_8_U.facout_s2  = \add_32ns_32s_32_2_1_U14.top_add_32ns_32s_32_2_1_Adder_8_U.u2.cout ;
assign \add_32ns_32s_32_2_1_U14.top_add_32ns_32s_32_2_1_Adder_8_U.fas_s2  = \add_32ns_32s_32_2_1_U14.top_add_32ns_32s_32_2_1_Adder_8_U.u2.s ;
assign \add_32ns_32s_32_2_1_U14.top_add_32ns_32s_32_2_1_Adder_8_U.u1.a  = \add_32ns_32s_32_2_1_U14.top_add_32ns_32s_32_2_1_Adder_8_U.a [15:0];
assign \add_32ns_32s_32_2_1_U14.top_add_32ns_32s_32_2_1_Adder_8_U.u1.b  = \add_32ns_32s_32_2_1_U14.top_add_32ns_32s_32_2_1_Adder_8_U.b [15:0];
assign \add_32ns_32s_32_2_1_U14.top_add_32ns_32s_32_2_1_Adder_8_U.u1.cin  = 1'h0;
assign \add_32ns_32s_32_2_1_U14.top_add_32ns_32s_32_2_1_Adder_8_U.facout_s1  = \add_32ns_32s_32_2_1_U14.top_add_32ns_32s_32_2_1_Adder_8_U.u1.cout ;
assign \add_32ns_32s_32_2_1_U14.top_add_32ns_32s_32_2_1_Adder_8_U.fas_s1  = \add_32ns_32s_32_2_1_U14.top_add_32ns_32s_32_2_1_Adder_8_U.u1.s ;
assign \add_32ns_32s_32_2_1_U14.top_add_32ns_32s_32_2_1_Adder_8_U.a  = \add_32ns_32s_32_2_1_U14.din0 ;
assign \add_32ns_32s_32_2_1_U14.top_add_32ns_32s_32_2_1_Adder_8_U.b  = \add_32ns_32s_32_2_1_U14.din1 ;
assign \add_32ns_32s_32_2_1_U14.top_add_32ns_32s_32_2_1_Adder_8_U.ce  = \add_32ns_32s_32_2_1_U14.ce ;
assign \add_32ns_32s_32_2_1_U14.top_add_32ns_32s_32_2_1_Adder_8_U.clk  = \add_32ns_32s_32_2_1_U14.clk ;
assign \add_32ns_32s_32_2_1_U14.top_add_32ns_32s_32_2_1_Adder_8_U.reset  = \add_32ns_32s_32_2_1_U14.reset ;
assign \add_32ns_32s_32_2_1_U14.dout  = \add_32ns_32s_32_2_1_U14.top_add_32ns_32s_32_2_1_Adder_8_U.s ;
assign \add_32ns_32s_32_2_1_U14.ce  = 1'h1;
assign \add_32ns_32s_32_2_1_U14.clk  = ap_clk;
assign \add_32ns_32s_32_2_1_U14.din0  = op_25_V_reg_1051;
assign \add_32ns_32s_32_2_1_U14.din1  = { op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16 };
assign grp_fu_708_p2 = \add_32ns_32s_32_2_1_U14.dout ;
assign \add_32ns_32s_32_2_1_U14.reset  = ap_rst;
assign \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.ain_s0  = \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.a ;
assign \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.bin_s0  = \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.b ;
assign \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.s  = { \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.fas_s2 , \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.sum_s1  };
assign \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.u2.a  = \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.ain_s1 ;
assign \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.u2.b  = \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.bin_s1 ;
assign \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.u2.cin  = \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.carry_s1 ;
assign \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.facout_s2  = \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.u2.cout ;
assign \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.fas_s2  = \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.u2.s ;
assign \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.u1.a  = \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.a [15:0];
assign \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.u1.b  = \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.b [15:0];
assign \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.u1.cin  = 1'h0;
assign \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.facout_s1  = \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.u1.cout ;
assign \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.fas_s1  = \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.u1.s ;
assign \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.a  = \add_32ns_32s_32_2_1_U12.din0 ;
assign \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.b  = \add_32ns_32s_32_2_1_U12.din1 ;
assign \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.ce  = \add_32ns_32s_32_2_1_U12.ce ;
assign \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.clk  = \add_32ns_32s_32_2_1_U12.clk ;
assign \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.reset  = \add_32ns_32s_32_2_1_U12.reset ;
assign \add_32ns_32s_32_2_1_U12.dout  = \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_8_U.s ;
assign \add_32ns_32s_32_2_1_U12.ce  = 1'h1;
assign \add_32ns_32s_32_2_1_U12.clk  = ap_clk;
assign \add_32ns_32s_32_2_1_U12.din0  = ret_V_27_reg_1019;
assign \add_32ns_32s_32_2_1_U12.din1  = { op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15 };
assign grp_fu_689_p2 = \add_32ns_32s_32_2_1_U12.dout ;
assign \add_32ns_32s_32_2_1_U12.reset  = ap_rst;
assign \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s0  = \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.a ;
assign \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s0  = \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.b ;
assign \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.s  = { \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s2 , \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.sum_s1  };
assign \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.a  = \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s1 ;
assign \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.b  = \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s1 ;
assign \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cin  = \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.carry_s1 ;
assign \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.facout_s2  = \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cout ;
assign \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s2  = \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.s ;
assign \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.a  = \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.a [15:0];
assign \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.b  = \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.b [15:0];
assign \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cin  = 1'h0;
assign \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.facout_s1  = \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cout ;
assign \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s1  = \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.s ;
assign \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.a  = \add_32ns_32ns_32_2_1_U11.din0 ;
assign \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.b  = \add_32ns_32ns_32_2_1_U11.din1 ;
assign \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.ce  = \add_32ns_32ns_32_2_1_U11.ce ;
assign \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.clk  = \add_32ns_32ns_32_2_1_U11.clk ;
assign \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.reset  = \add_32ns_32ns_32_2_1_U11.reset ;
assign \add_32ns_32ns_32_2_1_U11.dout  = \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.s ;
assign \add_32ns_32ns_32_2_1_U11.ce  = 1'h1;
assign \add_32ns_32ns_32_2_1_U11.clk  = ap_clk;
assign \add_32ns_32ns_32_2_1_U11.din0  = ret_V_16_cast_reg_1007;
assign \add_32ns_32ns_32_2_1_U11.din1  = 32'd1;
assign grp_fu_626_p2 = \add_32ns_32ns_32_2_1_U11.dout ;
assign \add_32ns_32ns_32_2_1_U11.reset  = ap_rst;
assign \add_10ns_10s_10_2_1_U8.top_add_10ns_10s_10_2_1_Adder_4_U.ain_s0  = \add_10ns_10s_10_2_1_U8.top_add_10ns_10s_10_2_1_Adder_4_U.a ;
assign \add_10ns_10s_10_2_1_U8.top_add_10ns_10s_10_2_1_Adder_4_U.bin_s0  = \add_10ns_10s_10_2_1_U8.top_add_10ns_10s_10_2_1_Adder_4_U.b ;
assign \add_10ns_10s_10_2_1_U8.top_add_10ns_10s_10_2_1_Adder_4_U.s  = { \add_10ns_10s_10_2_1_U8.top_add_10ns_10s_10_2_1_Adder_4_U.fas_s2 , \add_10ns_10s_10_2_1_U8.top_add_10ns_10s_10_2_1_Adder_4_U.sum_s1  };
assign \add_10ns_10s_10_2_1_U8.top_add_10ns_10s_10_2_1_Adder_4_U.u2.a  = \add_10ns_10s_10_2_1_U8.top_add_10ns_10s_10_2_1_Adder_4_U.ain_s1 ;
assign \add_10ns_10s_10_2_1_U8.top_add_10ns_10s_10_2_1_Adder_4_U.u2.b  = \add_10ns_10s_10_2_1_U8.top_add_10ns_10s_10_2_1_Adder_4_U.bin_s1 ;
assign \add_10ns_10s_10_2_1_U8.top_add_10ns_10s_10_2_1_Adder_4_U.u2.cin  = \add_10ns_10s_10_2_1_U8.top_add_10ns_10s_10_2_1_Adder_4_U.carry_s1 ;
assign \add_10ns_10s_10_2_1_U8.top_add_10ns_10s_10_2_1_Adder_4_U.facout_s2  = \add_10ns_10s_10_2_1_U8.top_add_10ns_10s_10_2_1_Adder_4_U.u2.cout ;
assign \add_10ns_10s_10_2_1_U8.top_add_10ns_10s_10_2_1_Adder_4_U.fas_s2  = \add_10ns_10s_10_2_1_U8.top_add_10ns_10s_10_2_1_Adder_4_U.u2.s ;
assign \add_10ns_10s_10_2_1_U8.top_add_10ns_10s_10_2_1_Adder_4_U.u1.a  = \add_10ns_10s_10_2_1_U8.top_add_10ns_10s_10_2_1_Adder_4_U.a [4:0];
assign \add_10ns_10s_10_2_1_U8.top_add_10ns_10s_10_2_1_Adder_4_U.u1.b  = \add_10ns_10s_10_2_1_U8.top_add_10ns_10s_10_2_1_Adder_4_U.b [4:0];
assign \add_10ns_10s_10_2_1_U8.top_add_10ns_10s_10_2_1_Adder_4_U.u1.cin  = 1'h0;
assign \add_10ns_10s_10_2_1_U8.top_add_10ns_10s_10_2_1_Adder_4_U.facout_s1  = \add_10ns_10s_10_2_1_U8.top_add_10ns_10s_10_2_1_Adder_4_U.u1.cout ;
assign \add_10ns_10s_10_2_1_U8.top_add_10ns_10s_10_2_1_Adder_4_U.fas_s1  = \add_10ns_10s_10_2_1_U8.top_add_10ns_10s_10_2_1_Adder_4_U.u1.s ;
assign \add_10ns_10s_10_2_1_U8.top_add_10ns_10s_10_2_1_Adder_4_U.a  = \add_10ns_10s_10_2_1_U8.din0 ;
assign \add_10ns_10s_10_2_1_U8.top_add_10ns_10s_10_2_1_Adder_4_U.b  = \add_10ns_10s_10_2_1_U8.din1 ;
assign \add_10ns_10s_10_2_1_U8.top_add_10ns_10s_10_2_1_Adder_4_U.ce  = \add_10ns_10s_10_2_1_U8.ce ;
assign \add_10ns_10s_10_2_1_U8.top_add_10ns_10s_10_2_1_Adder_4_U.clk  = \add_10ns_10s_10_2_1_U8.clk ;
assign \add_10ns_10s_10_2_1_U8.top_add_10ns_10s_10_2_1_Adder_4_U.reset  = \add_10ns_10s_10_2_1_U8.reset ;
assign \add_10ns_10s_10_2_1_U8.dout  = \add_10ns_10s_10_2_1_U8.top_add_10ns_10s_10_2_1_Adder_4_U.s ;
assign \add_10ns_10s_10_2_1_U8.ce  = 1'h1;
assign \add_10ns_10s_10_2_1_U8.clk  = ap_clk;
assign \add_10ns_10s_10_2_1_U8.din0  = { op_20_V_reg_909, 4'h0 };
assign \add_10ns_10s_10_2_1_U8.din1  = { select_ln1497_reg_904[3], select_ln1497_reg_904[3], select_ln1497_reg_904, 4'h0 };
assign grp_fu_484_p2 = \add_10ns_10s_10_2_1_U8.dout ;
assign \add_10ns_10s_10_2_1_U8.reset  = ap_rst;
endmodule


// Product machine:
module top_A_times_top_B (ap_start, op_0, op_12, op_15, op_16, op_17, op_18, op_3, op_4, op_6, op_7, ap_clk, unsafe_signal);
input ap_start;
input [1:0] op_0;
input [7:0] op_12;
input [7:0] op_15;
input [3:0] op_16;
input [7:0] op_17;
input [3:0] op_18;
input [3:0] op_3;
input op_4;
input [3:0] op_6;
input [15:0] op_7;
input ap_clk;
output unsafe_signal;
reg _setup;
initial _setup = 1'b0;
always @ (posedge ap_clk) _setup <= 1'b1;
reg ap_start_internal;
always @ (posedge ap_clk) if (!_setup) ap_start_internal <= ap_start;
reg [1:0] op_0_internal;
always @ (posedge ap_clk) if (!_setup) op_0_internal <= op_0;
reg [7:0] op_12_internal;
always @ (posedge ap_clk) if (!_setup) op_12_internal <= op_12;
reg [7:0] op_15_internal;
always @ (posedge ap_clk) if (!_setup) op_15_internal <= op_15;
reg [3:0] op_16_internal;
always @ (posedge ap_clk) if (!_setup) op_16_internal <= op_16;
reg [7:0] op_17_internal;
always @ (posedge ap_clk) if (!_setup) op_17_internal <= op_17;
reg [3:0] op_18_internal;
always @ (posedge ap_clk) if (!_setup) op_18_internal <= op_18;
reg [3:0] op_3_internal;
always @ (posedge ap_clk) if (!_setup) op_3_internal <= op_3;
reg op_4_internal;
always @ (posedge ap_clk) if (!_setup) op_4_internal <= op_4;
reg [3:0] op_6_internal;
always @ (posedge ap_clk) if (!_setup) op_6_internal <= op_6;
reg [15:0] op_7_internal;
always @ (posedge ap_clk) if (!_setup) op_7_internal <= op_7;
wire ap_done_A;
wire ap_done_B;
wire ap_done_eq;
assign ap_done_eq = ap_done_A == ap_done_B;
wire ap_idle_A;
wire ap_idle_B;
wire ap_idle_eq;
assign ap_idle_eq = ap_idle_A == ap_idle_B;
wire ap_ready_A;
wire ap_ready_B;
wire ap_ready_eq;
assign ap_ready_eq = ap_ready_A == ap_ready_B;
wire [31:0] op_29_A;
wire [31:0] op_29_B;
wire op_29_eq;
assign op_29_eq = op_29_A == op_29_B;
wire op_29_ap_vld_A;
wire op_29_ap_vld_B;
wire clk_enable_A;
wire clk_enable_B;
assign clk_enable_A = _setup & (~op_29_ap_vld_A | op_29_ap_vld_B);
assign clk_enable_B = _setup;
wire divergent;
assign divergent = ~(ap_done_eq & ap_idle_eq & ap_ready_eq & op_29_eq);
assign unsafe_signal = op_29_ap_vld_A & op_29_ap_vld_B & divergent;
top_A instance_A (
    .ap_clk(ap_clk),
    .clk_enable(clk_enable_A),
    .ap_start(ap_start_internal),
    .op_0(op_0_internal),
    .op_12(op_12_internal),
    .op_15(op_15_internal),
    .op_16(op_16_internal),
    .op_17(op_17_internal),
    .op_18(op_18_internal),
    .op_3(op_3_internal),
    .op_4(op_4_internal),
    .op_6(op_6_internal),
    .op_7(op_7_internal),
    .ap_done(ap_done_A),
    .ap_idle(ap_idle_A),
    .ap_ready(ap_ready_A),
    .op_29(op_29_A),
    .op_29_ap_vld(op_29_ap_vld_A)
);
top_B instance_B (
    .ap_clk(ap_clk),
    .clk_enable(clk_enable_B),
    .ap_start(ap_start_internal),
    .op_0(op_0_internal),
    .op_12(op_12_internal),
    .op_15(op_15_internal),
    .op_16(op_16_internal),
    .op_17(op_17_internal),
    .op_18(op_18_internal),
    .op_3(op_3_internal),
    .op_4(op_4_internal),
    .op_6(op_6_internal),
    .op_7(op_7_internal),
    .ap_done(ap_done_B),
    .ap_idle(ap_idle_B),
    .ap_ready(ap_ready_B),
    .op_29(op_29_B),
    .op_29_ap_vld(op_29_ap_vld_B)
);
endmodule
