// Processed by function `construct_kairos` in `verilog_tricks.py`.
// Machine A:
// Processed by function `add_clk_enable_signal` in `verilog_tricks.py`.
// Processed by function `remove_reset_signal` in `verilog_tricks.py`.
module top_A (
  ap_clk,
  ap_start,
  ap_done,
  ap_idle,
  ap_ready,
  op_0,
  op_1,
  op_2,
  op_3,
  op_4,
  op_7,
  op_8,
  op_10,
  op_14,
  op_15,
  op_16,
  op_29,
  op_29_ap_vld,
clk_enable
);
input clk_enable;


input ap_clk;
wire ap_rst;
assign ap_rst = op_29_ap_vld;
input ap_start;
input [3:0] op_0;
input [7:0] op_1;
input [1:0] op_10;
input [7:0] op_14;
input [3:0] op_15;
input [7:0] op_16;
input [1:0] op_2;
input op_3;
input [31:0] op_4;
input [1:0] op_7;
input op_8;
output ap_done;
output ap_idle;
output ap_ready;
output [31:0] op_29;
output op_29_ap_vld;


reg \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_11_U.ain_s1 ;
reg \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_11_U.bin_s1 ;
reg \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_11_U.carry_s1 ;
reg \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_11_U.sum_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.ain_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.bin_s1 ;
reg \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.carry_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.sum_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_8_U.ain_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_8_U.bin_s1 ;
reg \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_8_U.carry_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_8_U.sum_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_8_U.ain_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_8_U.bin_s1 ;
reg \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_8_U.carry_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_8_U.sum_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.ain_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.bin_s1 ;
reg \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.carry_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.sum_s1 ;
reg [15:0] \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_9_U.ain_s1 ;
reg [15:0] \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_9_U.bin_s1 ;
reg \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_9_U.carry_s1 ;
reg [15:0] \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_9_U.sum_s1 ;
reg [16:0] \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_7_U.ain_s1 ;
reg [16:0] \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_7_U.bin_s1 ;
reg \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_7_U.carry_s1 ;
reg [16:0] \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_7_U.sum_s1 ;
reg [17:0] \add_35s_35s_35_2_1_U13.top_add_35s_35s_35_2_1_Adder_10_U.ain_s1 ;
reg [17:0] \add_35s_35s_35_2_1_U13.top_add_35s_35s_35_2_1_Adder_10_U.bin_s1 ;
reg \add_35s_35s_35_2_1_U13.top_add_35s_35s_35_2_1_Adder_10_U.carry_s1 ;
reg [16:0] \add_35s_35s_35_2_1_U13.top_add_35s_35s_35_2_1_Adder_10_U.sum_s1 ;
reg [1:0] \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_2_U.ain_s1 ;
reg [1:0] \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_2_U.bin_s1 ;
reg \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_2_U.carry_s1 ;
reg \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_2_U.sum_s1 ;
reg [1:0] \add_3s_3ns_3_2_1_U2.top_add_3s_3ns_3_2_1_Adder_1_U.ain_s1 ;
reg [1:0] \add_3s_3ns_3_2_1_U2.top_add_3s_3ns_3_2_1_Adder_1_U.bin_s1 ;
reg \add_3s_3ns_3_2_1_U2.top_add_3s_3ns_3_2_1_Adder_1_U.carry_s1 ;
reg \add_3s_3ns_3_2_1_U2.top_add_3s_3ns_3_2_1_Adder_1_U.sum_s1 ;
reg [2:0] \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_6_U.ain_s1 ;
reg [2:0] \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_6_U.bin_s1 ;
reg \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_6_U.carry_s1 ;
reg [1:0] \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_6_U.sum_s1 ;
reg [2:0] \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.ain_s1 ;
reg [2:0] \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.bin_s1 ;
reg \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.carry_s1 ;
reg [1:0] \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.sum_s1 ;
reg [2:0] \add_5s_5ns_5_2_1_U5.top_add_5s_5ns_5_2_1_Adder_4_U.ain_s1 ;
reg [2:0] \add_5s_5ns_5_2_1_U5.top_add_5s_5ns_5_2_1_Adder_4_U.bin_s1 ;
reg \add_5s_5ns_5_2_1_U5.top_add_5s_5ns_5_2_1_Adder_4_U.carry_s1 ;
reg [1:0] \add_5s_5ns_5_2_1_U5.top_add_5s_5ns_5_2_1_Adder_4_U.sum_s1 ;
reg [2:0] \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_3_U.ain_s1 ;
reg [2:0] \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_3_U.bin_s1 ;
reg \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_3_U.carry_s1 ;
reg [1:0] \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_3_U.sum_s1 ;
reg [31:0] add_ln691_1_reg_808;
reg [31:0] add_ln691_2_reg_880;
reg [4:0] add_ln691_reg_708;
reg [1:0] add_ln69_1_reg_875;
reg [31:0] add_ln69_reg_900;
reg [29:0] ap_CS_fsm = 30'h00000001;
reg icmp_ln1495_reg_771;
reg icmp_ln1498_1_reg_729;
reg icmp_ln1498_reg_739;
reg icmp_ln851_1_reg_853;
reg icmp_ln851_reg_628;
reg [31:0] \lshr_32ns_32s_32_7_1_U9.din1_cast_array[0] ;
reg [31:0] \lshr_32ns_32s_32_7_1_U9.din1_cast_array[1] ;
reg [31:0] \lshr_32ns_32s_32_7_1_U9.din1_cast_array[2] ;
reg [31:0] \lshr_32ns_32s_32_7_1_U9.din1_cast_array[3] ;
reg [31:0] \lshr_32ns_32s_32_7_1_U9.din1_cast_array[4] ;
reg [31:0] \lshr_32ns_32s_32_7_1_U9.din1_cast_array[5] ;
reg [31:0] \lshr_32ns_32s_32_7_1_U9.dout_array[0] ;
reg [31:0] \lshr_32ns_32s_32_7_1_U9.dout_array[1] ;
reg [31:0] \lshr_32ns_32s_32_7_1_U9.dout_array[2] ;
reg [31:0] \lshr_32ns_32s_32_7_1_U9.dout_array[3] ;
reg [31:0] \lshr_32ns_32s_32_7_1_U9.dout_array[4] ;
reg [31:0] \lshr_32ns_32s_32_7_1_U9.dout_array[5] ;
reg [1:0] op_17_V_reg_833;
reg [2:0] op_21_V_reg_660;
reg [4:0] op_23_V_reg_776;
reg [31:0] op_25_V_reg_838;
reg op_6_V_reg_703;
reg [1:0] ret_V_11_reg_885;
reg [4:0] ret_V_12_reg_633;
reg [2:0] ret_V_13_reg_655;
reg [4:0] ret_V_14_reg_680;
reg [31:0] ret_V_15_cast_reg_868;
reg [4:0] ret_V_15_reg_734;
reg [33:0] ret_V_16_reg_796;
reg [31:0] ret_V_17_reg_813;
reg [34:0] ret_V_18_reg_863;
reg [31:0] ret_V_19_reg_890;
reg [2:0] ret_V_3_reg_650;
reg [31:0] ret_V_7_cast_reg_801;
reg [1:0] ret_V_reg_638;
reg [2:0] sext_ln835_reg_643;
reg [4:0] sext_ln850_reg_690;
reg [31:0] \shl_32ns_32s_32_7_1_U8.din1_cast_array[0] ;
reg [31:0] \shl_32ns_32s_32_7_1_U8.din1_cast_array[1] ;
reg [31:0] \shl_32ns_32s_32_7_1_U8.din1_cast_array[2] ;
reg [31:0] \shl_32ns_32s_32_7_1_U8.din1_cast_array[3] ;
reg [31:0] \shl_32ns_32s_32_7_1_U8.din1_cast_array[4] ;
reg [31:0] \shl_32ns_32s_32_7_1_U8.din1_cast_array[5] ;
reg [31:0] \shl_32ns_32s_32_7_1_U8.dout_array[0] ;
reg [31:0] \shl_32ns_32s_32_7_1_U8.dout_array[1] ;
reg [31:0] \shl_32ns_32s_32_7_1_U8.dout_array[2] ;
reg [31:0] \shl_32ns_32s_32_7_1_U8.dout_array[3] ;
reg [31:0] \shl_32ns_32s_32_7_1_U8.dout_array[4] ;
reg [31:0] \shl_32ns_32s_32_7_1_U8.dout_array[5] ;
reg [1:0] \sub_3ns_3s_3_2_1_U6.top_sub_3ns_3s_3_2_1_Adder_5_U.ain_s1 ;
reg [1:0] \sub_3ns_3s_3_2_1_U6.top_sub_3ns_3s_3_2_1_Adder_5_U.bin_s1 ;
reg \sub_3ns_3s_3_2_1_U6.top_sub_3ns_3s_3_2_1_Adder_5_U.carry_s1 ;
reg \sub_3ns_3s_3_2_1_U6.top_sub_3ns_3s_3_2_1_Adder_5_U.sum_s1 ;
reg [2:0] sub_ln1497_reg_745;
reg [3:0] tmp_2_reg_685;
reg tmp_reg_724;
reg trunc_ln1497_1_reg_823;
reg [1:0] trunc_ln1497_reg_818;
wire [31:0] _000_;
wire [31:0] _001_;
wire [4:0] _002_;
wire [1:0] _003_;
wire [31:0] _004_;
wire [29:0] _005_;
wire _006_;
wire _007_;
wire _008_;
wire _009_;
wire _010_;
wire [1:0] _011_;
wire [2:0] _012_;
wire [4:0] _013_;
wire [31:0] _014_;
wire _015_;
wire [1:0] _016_;
wire [4:0] _017_;
wire [2:0] _018_;
wire [4:0] _019_;
wire [31:0] _020_;
wire [4:0] _021_;
wire [33:0] _022_;
wire [31:0] _023_;
wire [34:0] _024_;
wire [31:0] _025_;
wire [2:0] _026_;
wire [31:0] _027_;
wire [1:0] _028_;
wire [2:0] _029_;
wire [4:0] _030_;
wire [2:0] _031_;
wire [3:0] _032_;
wire _033_;
wire _034_;
wire [1:0] _035_;
wire [1:0] _036_;
wire _037_;
wire _038_;
wire _039_;
wire _040_;
wire _041_;
wire _042_;
wire _043_;
wire _044_;
wire _045_;
wire _046_;
wire _047_;
wire _048_;
wire _049_;
wire _050_;
wire _051_;
wire _052_;
wire [1:0] _053_;
wire [1:0] _054_;
wire [15:0] _055_;
wire [15:0] _056_;
wire _057_;
wire [15:0] _058_;
wire [16:0] _059_;
wire [16:0] _060_;
wire [15:0] _061_;
wire [15:0] _062_;
wire _063_;
wire [15:0] _064_;
wire [16:0] _065_;
wire [16:0] _066_;
wire [15:0] _067_;
wire [15:0] _068_;
wire _069_;
wire [15:0] _070_;
wire [16:0] _071_;
wire [16:0] _072_;
wire [15:0] _073_;
wire [15:0] _074_;
wire _075_;
wire [15:0] _076_;
wire [16:0] _077_;
wire [16:0] _078_;
wire [15:0] _079_;
wire [15:0] _080_;
wire _081_;
wire [15:0] _082_;
wire [16:0] _083_;
wire [16:0] _084_;
wire [16:0] _085_;
wire [16:0] _086_;
wire _087_;
wire [16:0] _088_;
wire [17:0] _089_;
wire [17:0] _090_;
wire [17:0] _091_;
wire [17:0] _092_;
wire _093_;
wire [16:0] _094_;
wire [17:0] _095_;
wire [18:0] _096_;
wire [1:0] _097_;
wire [1:0] _098_;
wire _099_;
wire _100_;
wire [1:0] _101_;
wire [2:0] _102_;
wire [1:0] _103_;
wire [1:0] _104_;
wire _105_;
wire _106_;
wire [1:0] _107_;
wire [2:0] _108_;
wire [2:0] _109_;
wire [2:0] _110_;
wire _111_;
wire [1:0] _112_;
wire [2:0] _113_;
wire [3:0] _114_;
wire [2:0] _115_;
wire [2:0] _116_;
wire _117_;
wire [1:0] _118_;
wire [2:0] _119_;
wire [3:0] _120_;
wire [2:0] _121_;
wire [2:0] _122_;
wire _123_;
wire [1:0] _124_;
wire [2:0] _125_;
wire [3:0] _126_;
wire [2:0] _127_;
wire [2:0] _128_;
wire _129_;
wire [1:0] _130_;
wire [2:0] _131_;
wire [3:0] _132_;
wire [31:0] _133_;
wire [31:0] _134_;
wire [31:0] _135_;
wire [31:0] _136_;
wire [31:0] _137_;
wire [31:0] _138_;
wire [31:0] _139_;
wire [31:0] _140_;
wire [31:0] _141_;
wire [31:0] _142_;
wire [31:0] _143_;
wire [31:0] _144_;
wire [31:0] _145_;
wire [31:0] _146_;
wire [31:0] _147_;
wire [31:0] _148_;
wire [31:0] _149_;
wire [31:0] _150_;
wire [31:0] _151_;
wire [31:0] _152_;
wire [31:0] _153_;
wire [31:0] _154_;
wire [31:0] _155_;
wire [31:0] _156_;
wire [31:0] _157_;
wire [31:0] _158_;
wire [31:0] _159_;
wire [31:0] _160_;
wire [31:0] _161_;
wire [31:0] _162_;
wire [31:0] _163_;
wire [31:0] _164_;
wire [31:0] _165_;
wire [31:0] _166_;
wire [31:0] _167_;
wire [31:0] _168_;
wire [31:0] _169_;
wire [31:0] _170_;
wire [31:0] _171_;
wire [31:0] _172_;
wire [31:0] _173_;
wire [31:0] _174_;
wire [31:0] _175_;
wire [31:0] _176_;
wire [31:0] _177_;
wire [31:0] _178_;
wire [31:0] _179_;
wire [31:0] _180_;
wire [31:0] _181_;
wire [31:0] _182_;
wire [31:0] _183_;
wire [31:0] _184_;
wire [31:0] _185_;
wire [31:0] _186_;
wire [31:0] _187_;
wire [31:0] _188_;
wire [31:0] _189_;
wire [31:0] _190_;
wire [31:0] _191_;
wire [31:0] _192_;
wire [1:0] _193_;
wire [1:0] _194_;
wire _195_;
wire _196_;
wire [1:0] _197_;
wire [2:0] _198_;
wire _199_;
wire _200_;
wire _201_;
wire _202_;
wire _203_;
wire _204_;
wire _205_;
wire _206_;
wire _207_;
wire _208_;
wire _209_;
wire _210_;
wire _211_;
wire _212_;
wire _213_;
wire _214_;
wire _215_;
wire _216_;
wire _217_;
wire _218_;
wire _219_;
wire _220_;
wire _221_;
wire _222_;
wire _223_;
wire _224_;
wire _225_;
wire _226_;
wire _227_;
wire _228_;
wire _229_;
wire _230_;
wire _231_;
wire \add_2ns_2ns_2_2_1_U14.ce ;
wire \add_2ns_2ns_2_2_1_U14.clk ;
wire [1:0] \add_2ns_2ns_2_2_1_U14.din0 ;
wire [1:0] \add_2ns_2ns_2_2_1_U14.din1 ;
wire [1:0] \add_2ns_2ns_2_2_1_U14.dout ;
wire \add_2ns_2ns_2_2_1_U14.reset ;
wire [1:0] \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_11_U.a ;
wire [1:0] \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_11_U.ain_s0 ;
wire [1:0] \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_11_U.b ;
wire [1:0] \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_11_U.bin_s0 ;
wire \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_11_U.ce ;
wire \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_11_U.clk ;
wire \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_11_U.facout_s1 ;
wire \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_11_U.facout_s2 ;
wire \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_11_U.fas_s1 ;
wire \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_11_U.fas_s2 ;
wire \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_11_U.reset ;
wire [1:0] \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_11_U.s ;
wire \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_11_U.u1.a ;
wire \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_11_U.u1.b ;
wire \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_11_U.u1.cin ;
wire \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_11_U.u1.cout ;
wire \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_11_U.u1.s ;
wire \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_11_U.u2.a ;
wire \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_11_U.u2.b ;
wire \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_11_U.u2.cin ;
wire \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_11_U.u2.cout ;
wire \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_11_U.u2.s ;
wire \add_32ns_32ns_32_2_1_U11.ce ;
wire \add_32ns_32ns_32_2_1_U11.clk ;
wire [31:0] \add_32ns_32ns_32_2_1_U11.din0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U11.din1 ;
wire [31:0] \add_32ns_32ns_32_2_1_U11.dout ;
wire \add_32ns_32ns_32_2_1_U11.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.a ;
wire [31:0] \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.ain_s0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.b ;
wire [31:0] \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.bin_s0 ;
wire \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.ce ;
wire \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.clk ;
wire \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.facout_s1 ;
wire \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.facout_s2 ;
wire [15:0] \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.fas_s1 ;
wire [15:0] \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.fas_s2 ;
wire \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.u1.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.u1.b ;
wire \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.u1.cin ;
wire \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.u1.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.u1.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.u2.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.u2.b ;
wire \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.u2.cin ;
wire \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.u2.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.u2.s ;
wire \add_32ns_32ns_32_2_1_U15.ce ;
wire \add_32ns_32ns_32_2_1_U15.clk ;
wire [31:0] \add_32ns_32ns_32_2_1_U15.din0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U15.din1 ;
wire [31:0] \add_32ns_32ns_32_2_1_U15.dout ;
wire \add_32ns_32ns_32_2_1_U15.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_8_U.a ;
wire [31:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_8_U.ain_s0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_8_U.b ;
wire [31:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_8_U.bin_s0 ;
wire \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_8_U.ce ;
wire \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_8_U.clk ;
wire \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_8_U.facout_s1 ;
wire \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_8_U.facout_s2 ;
wire [15:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_8_U.fas_s1 ;
wire [15:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_8_U.fas_s2 ;
wire \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_8_U.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_8_U.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_8_U.u1.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_8_U.u1.b ;
wire \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_8_U.u1.cin ;
wire \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_8_U.u1.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_8_U.u1.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_8_U.u2.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_8_U.u2.b ;
wire \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_8_U.u2.cin ;
wire \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_8_U.u2.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_8_U.u2.s ;
wire \add_32ns_32ns_32_2_1_U16.ce ;
wire \add_32ns_32ns_32_2_1_U16.clk ;
wire [31:0] \add_32ns_32ns_32_2_1_U16.din0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U16.din1 ;
wire [31:0] \add_32ns_32ns_32_2_1_U16.dout ;
wire \add_32ns_32ns_32_2_1_U16.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_8_U.a ;
wire [31:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_8_U.ain_s0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_8_U.b ;
wire [31:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_8_U.bin_s0 ;
wire \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_8_U.ce ;
wire \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_8_U.clk ;
wire \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_8_U.facout_s1 ;
wire \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_8_U.facout_s2 ;
wire [15:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_8_U.fas_s1 ;
wire [15:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_8_U.fas_s2 ;
wire \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_8_U.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_8_U.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_8_U.u1.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_8_U.u1.b ;
wire \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_8_U.u1.cin ;
wire \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_8_U.u1.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_8_U.u1.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_8_U.u2.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_8_U.u2.b ;
wire \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_8_U.u2.cin ;
wire \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_8_U.u2.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_8_U.u2.s ;
wire \add_32ns_32ns_32_2_1_U17.ce ;
wire \add_32ns_32ns_32_2_1_U17.clk ;
wire [31:0] \add_32ns_32ns_32_2_1_U17.din0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U17.din1 ;
wire [31:0] \add_32ns_32ns_32_2_1_U17.dout ;
wire \add_32ns_32ns_32_2_1_U17.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.a ;
wire [31:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.ain_s0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.b ;
wire [31:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.bin_s0 ;
wire \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.ce ;
wire \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.clk ;
wire \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.facout_s1 ;
wire \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.facout_s2 ;
wire [15:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.fas_s1 ;
wire [15:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.fas_s2 ;
wire \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.u1.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.u1.b ;
wire \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.u1.cin ;
wire \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.u1.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.u1.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.u2.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.u2.b ;
wire \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.u2.cin ;
wire \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.u2.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.u2.s ;
wire \add_32ns_32s_32_2_1_U12.ce ;
wire \add_32ns_32s_32_2_1_U12.clk ;
wire [31:0] \add_32ns_32s_32_2_1_U12.din0 ;
wire [31:0] \add_32ns_32s_32_2_1_U12.din1 ;
wire [31:0] \add_32ns_32s_32_2_1_U12.dout ;
wire \add_32ns_32s_32_2_1_U12.reset ;
wire [31:0] \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_9_U.a ;
wire [31:0] \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_9_U.ain_s0 ;
wire [31:0] \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_9_U.b ;
wire [31:0] \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_9_U.bin_s0 ;
wire \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_9_U.ce ;
wire \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_9_U.clk ;
wire \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_9_U.facout_s1 ;
wire \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_9_U.facout_s2 ;
wire [15:0] \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_9_U.fas_s1 ;
wire [15:0] \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_9_U.fas_s2 ;
wire \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_9_U.reset ;
wire [31:0] \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_9_U.s ;
wire [15:0] \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_9_U.u1.a ;
wire [15:0] \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_9_U.u1.b ;
wire \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_9_U.u1.cin ;
wire \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_9_U.u1.cout ;
wire [15:0] \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_9_U.u1.s ;
wire [15:0] \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_9_U.u2.a ;
wire [15:0] \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_9_U.u2.b ;
wire \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_9_U.u2.cin ;
wire \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_9_U.u2.cout ;
wire [15:0] \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_9_U.u2.s ;
wire \add_34s_34s_34_2_1_U10.ce ;
wire \add_34s_34s_34_2_1_U10.clk ;
wire [33:0] \add_34s_34s_34_2_1_U10.din0 ;
wire [33:0] \add_34s_34s_34_2_1_U10.din1 ;
wire [33:0] \add_34s_34s_34_2_1_U10.dout ;
wire \add_34s_34s_34_2_1_U10.reset ;
wire [33:0] \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_7_U.a ;
wire [33:0] \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_7_U.ain_s0 ;
wire [33:0] \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_7_U.b ;
wire [33:0] \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_7_U.bin_s0 ;
wire \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_7_U.ce ;
wire \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_7_U.clk ;
wire \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_7_U.facout_s1 ;
wire \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_7_U.facout_s2 ;
wire [16:0] \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_7_U.fas_s1 ;
wire [16:0] \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_7_U.fas_s2 ;
wire \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_7_U.reset ;
wire [33:0] \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_7_U.s ;
wire [16:0] \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_7_U.u1.a ;
wire [16:0] \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_7_U.u1.b ;
wire \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_7_U.u1.cin ;
wire \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_7_U.u1.cout ;
wire [16:0] \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_7_U.u1.s ;
wire [16:0] \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_7_U.u2.a ;
wire [16:0] \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_7_U.u2.b ;
wire \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_7_U.u2.cin ;
wire \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_7_U.u2.cout ;
wire [16:0] \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_7_U.u2.s ;
wire \add_35s_35s_35_2_1_U13.ce ;
wire \add_35s_35s_35_2_1_U13.clk ;
wire [34:0] \add_35s_35s_35_2_1_U13.din0 ;
wire [34:0] \add_35s_35s_35_2_1_U13.din1 ;
wire [34:0] \add_35s_35s_35_2_1_U13.dout ;
wire \add_35s_35s_35_2_1_U13.reset ;
wire [34:0] \add_35s_35s_35_2_1_U13.top_add_35s_35s_35_2_1_Adder_10_U.a ;
wire [34:0] \add_35s_35s_35_2_1_U13.top_add_35s_35s_35_2_1_Adder_10_U.ain_s0 ;
wire [34:0] \add_35s_35s_35_2_1_U13.top_add_35s_35s_35_2_1_Adder_10_U.b ;
wire [34:0] \add_35s_35s_35_2_1_U13.top_add_35s_35s_35_2_1_Adder_10_U.bin_s0 ;
wire \add_35s_35s_35_2_1_U13.top_add_35s_35s_35_2_1_Adder_10_U.ce ;
wire \add_35s_35s_35_2_1_U13.top_add_35s_35s_35_2_1_Adder_10_U.clk ;
wire \add_35s_35s_35_2_1_U13.top_add_35s_35s_35_2_1_Adder_10_U.facout_s1 ;
wire \add_35s_35s_35_2_1_U13.top_add_35s_35s_35_2_1_Adder_10_U.facout_s2 ;
wire [16:0] \add_35s_35s_35_2_1_U13.top_add_35s_35s_35_2_1_Adder_10_U.fas_s1 ;
wire [17:0] \add_35s_35s_35_2_1_U13.top_add_35s_35s_35_2_1_Adder_10_U.fas_s2 ;
wire \add_35s_35s_35_2_1_U13.top_add_35s_35s_35_2_1_Adder_10_U.reset ;
wire [34:0] \add_35s_35s_35_2_1_U13.top_add_35s_35s_35_2_1_Adder_10_U.s ;
wire [16:0] \add_35s_35s_35_2_1_U13.top_add_35s_35s_35_2_1_Adder_10_U.u1.a ;
wire [16:0] \add_35s_35s_35_2_1_U13.top_add_35s_35s_35_2_1_Adder_10_U.u1.b ;
wire \add_35s_35s_35_2_1_U13.top_add_35s_35s_35_2_1_Adder_10_U.u1.cin ;
wire \add_35s_35s_35_2_1_U13.top_add_35s_35s_35_2_1_Adder_10_U.u1.cout ;
wire [16:0] \add_35s_35s_35_2_1_U13.top_add_35s_35s_35_2_1_Adder_10_U.u1.s ;
wire [17:0] \add_35s_35s_35_2_1_U13.top_add_35s_35s_35_2_1_Adder_10_U.u2.a ;
wire [17:0] \add_35s_35s_35_2_1_U13.top_add_35s_35s_35_2_1_Adder_10_U.u2.b ;
wire \add_35s_35s_35_2_1_U13.top_add_35s_35s_35_2_1_Adder_10_U.u2.cin ;
wire \add_35s_35s_35_2_1_U13.top_add_35s_35s_35_2_1_Adder_10_U.u2.cout ;
wire [17:0] \add_35s_35s_35_2_1_U13.top_add_35s_35s_35_2_1_Adder_10_U.u2.s ;
wire \add_3ns_3ns_3_2_1_U3.ce ;
wire \add_3ns_3ns_3_2_1_U3.clk ;
wire [2:0] \add_3ns_3ns_3_2_1_U3.din0 ;
wire [2:0] \add_3ns_3ns_3_2_1_U3.din1 ;
wire [2:0] \add_3ns_3ns_3_2_1_U3.dout ;
wire \add_3ns_3ns_3_2_1_U3.reset ;
wire [2:0] \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_2_U.a ;
wire [2:0] \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_2_U.ain_s0 ;
wire [2:0] \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_2_U.b ;
wire [2:0] \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_2_U.bin_s0 ;
wire \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_2_U.ce ;
wire \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_2_U.clk ;
wire \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_2_U.facout_s1 ;
wire \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_2_U.facout_s2 ;
wire \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_2_U.fas_s1 ;
wire [1:0] \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_2_U.fas_s2 ;
wire \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_2_U.reset ;
wire [2:0] \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_2_U.s ;
wire \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_2_U.u1.a ;
wire \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_2_U.u1.b ;
wire \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_2_U.u1.cin ;
wire \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_2_U.u1.cout ;
wire \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_2_U.u1.s ;
wire [1:0] \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_2_U.u2.a ;
wire [1:0] \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_2_U.u2.b ;
wire \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_2_U.u2.cin ;
wire \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_2_U.u2.cout ;
wire [1:0] \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_2_U.u2.s ;
wire \add_3s_3ns_3_2_1_U2.ce ;
wire \add_3s_3ns_3_2_1_U2.clk ;
wire [2:0] \add_3s_3ns_3_2_1_U2.din0 ;
wire [2:0] \add_3s_3ns_3_2_1_U2.din1 ;
wire [2:0] \add_3s_3ns_3_2_1_U2.dout ;
wire \add_3s_3ns_3_2_1_U2.reset ;
wire [2:0] \add_3s_3ns_3_2_1_U2.top_add_3s_3ns_3_2_1_Adder_1_U.a ;
wire [2:0] \add_3s_3ns_3_2_1_U2.top_add_3s_3ns_3_2_1_Adder_1_U.ain_s0 ;
wire [2:0] \add_3s_3ns_3_2_1_U2.top_add_3s_3ns_3_2_1_Adder_1_U.b ;
wire [2:0] \add_3s_3ns_3_2_1_U2.top_add_3s_3ns_3_2_1_Adder_1_U.bin_s0 ;
wire \add_3s_3ns_3_2_1_U2.top_add_3s_3ns_3_2_1_Adder_1_U.ce ;
wire \add_3s_3ns_3_2_1_U2.top_add_3s_3ns_3_2_1_Adder_1_U.clk ;
wire \add_3s_3ns_3_2_1_U2.top_add_3s_3ns_3_2_1_Adder_1_U.facout_s1 ;
wire \add_3s_3ns_3_2_1_U2.top_add_3s_3ns_3_2_1_Adder_1_U.facout_s2 ;
wire \add_3s_3ns_3_2_1_U2.top_add_3s_3ns_3_2_1_Adder_1_U.fas_s1 ;
wire [1:0] \add_3s_3ns_3_2_1_U2.top_add_3s_3ns_3_2_1_Adder_1_U.fas_s2 ;
wire \add_3s_3ns_3_2_1_U2.top_add_3s_3ns_3_2_1_Adder_1_U.reset ;
wire [2:0] \add_3s_3ns_3_2_1_U2.top_add_3s_3ns_3_2_1_Adder_1_U.s ;
wire \add_3s_3ns_3_2_1_U2.top_add_3s_3ns_3_2_1_Adder_1_U.u1.a ;
wire \add_3s_3ns_3_2_1_U2.top_add_3s_3ns_3_2_1_Adder_1_U.u1.b ;
wire \add_3s_3ns_3_2_1_U2.top_add_3s_3ns_3_2_1_Adder_1_U.u1.cin ;
wire \add_3s_3ns_3_2_1_U2.top_add_3s_3ns_3_2_1_Adder_1_U.u1.cout ;
wire \add_3s_3ns_3_2_1_U2.top_add_3s_3ns_3_2_1_Adder_1_U.u1.s ;
wire [1:0] \add_3s_3ns_3_2_1_U2.top_add_3s_3ns_3_2_1_Adder_1_U.u2.a ;
wire [1:0] \add_3s_3ns_3_2_1_U2.top_add_3s_3ns_3_2_1_Adder_1_U.u2.b ;
wire \add_3s_3ns_3_2_1_U2.top_add_3s_3ns_3_2_1_Adder_1_U.u2.cin ;
wire \add_3s_3ns_3_2_1_U2.top_add_3s_3ns_3_2_1_Adder_1_U.u2.cout ;
wire [1:0] \add_3s_3ns_3_2_1_U2.top_add_3s_3ns_3_2_1_Adder_1_U.u2.s ;
wire \add_5ns_5ns_5_2_1_U7.ce ;
wire \add_5ns_5ns_5_2_1_U7.clk ;
wire [4:0] \add_5ns_5ns_5_2_1_U7.din0 ;
wire [4:0] \add_5ns_5ns_5_2_1_U7.din1 ;
wire [4:0] \add_5ns_5ns_5_2_1_U7.dout ;
wire \add_5ns_5ns_5_2_1_U7.reset ;
wire [4:0] \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_6_U.a ;
wire [4:0] \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_6_U.ain_s0 ;
wire [4:0] \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_6_U.b ;
wire [4:0] \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_6_U.bin_s0 ;
wire \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_6_U.ce ;
wire \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_6_U.clk ;
wire \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_6_U.facout_s1 ;
wire \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_6_U.facout_s2 ;
wire [1:0] \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_6_U.fas_s1 ;
wire [2:0] \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_6_U.fas_s2 ;
wire \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_6_U.reset ;
wire [4:0] \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_6_U.s ;
wire [1:0] \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_6_U.u1.a ;
wire [1:0] \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_6_U.u1.b ;
wire \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_6_U.u1.cin ;
wire \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_6_U.u1.cout ;
wire [1:0] \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_6_U.u1.s ;
wire [2:0] \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_6_U.u2.a ;
wire [2:0] \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_6_U.u2.b ;
wire \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_6_U.u2.cin ;
wire \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_6_U.u2.cout ;
wire [2:0] \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_6_U.u2.s ;
wire \add_5ns_5s_5_2_1_U1.ce ;
wire \add_5ns_5s_5_2_1_U1.clk ;
wire [4:0] \add_5ns_5s_5_2_1_U1.din0 ;
wire [4:0] \add_5ns_5s_5_2_1_U1.din1 ;
wire [4:0] \add_5ns_5s_5_2_1_U1.dout ;
wire \add_5ns_5s_5_2_1_U1.reset ;
wire [4:0] \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.a ;
wire [4:0] \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.ain_s0 ;
wire [4:0] \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.b ;
wire [4:0] \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.bin_s0 ;
wire \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.ce ;
wire \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.clk ;
wire \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.facout_s1 ;
wire \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.facout_s2 ;
wire [1:0] \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.fas_s1 ;
wire [2:0] \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.fas_s2 ;
wire \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.reset ;
wire [4:0] \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.s ;
wire [1:0] \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.u1.a ;
wire [1:0] \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.u1.b ;
wire \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.u1.cin ;
wire \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.u1.cout ;
wire [1:0] \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.u1.s ;
wire [2:0] \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.u2.a ;
wire [2:0] \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.u2.b ;
wire \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.u2.cin ;
wire \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.u2.cout ;
wire [2:0] \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.u2.s ;
wire \add_5s_5ns_5_2_1_U5.ce ;
wire \add_5s_5ns_5_2_1_U5.clk ;
wire [4:0] \add_5s_5ns_5_2_1_U5.din0 ;
wire [4:0] \add_5s_5ns_5_2_1_U5.din1 ;
wire [4:0] \add_5s_5ns_5_2_1_U5.dout ;
wire \add_5s_5ns_5_2_1_U5.reset ;
wire [4:0] \add_5s_5ns_5_2_1_U5.top_add_5s_5ns_5_2_1_Adder_4_U.a ;
wire [4:0] \add_5s_5ns_5_2_1_U5.top_add_5s_5ns_5_2_1_Adder_4_U.ain_s0 ;
wire [4:0] \add_5s_5ns_5_2_1_U5.top_add_5s_5ns_5_2_1_Adder_4_U.b ;
wire [4:0] \add_5s_5ns_5_2_1_U5.top_add_5s_5ns_5_2_1_Adder_4_U.bin_s0 ;
wire \add_5s_5ns_5_2_1_U5.top_add_5s_5ns_5_2_1_Adder_4_U.ce ;
wire \add_5s_5ns_5_2_1_U5.top_add_5s_5ns_5_2_1_Adder_4_U.clk ;
wire \add_5s_5ns_5_2_1_U5.top_add_5s_5ns_5_2_1_Adder_4_U.facout_s1 ;
wire \add_5s_5ns_5_2_1_U5.top_add_5s_5ns_5_2_1_Adder_4_U.facout_s2 ;
wire [1:0] \add_5s_5ns_5_2_1_U5.top_add_5s_5ns_5_2_1_Adder_4_U.fas_s1 ;
wire [2:0] \add_5s_5ns_5_2_1_U5.top_add_5s_5ns_5_2_1_Adder_4_U.fas_s2 ;
wire \add_5s_5ns_5_2_1_U5.top_add_5s_5ns_5_2_1_Adder_4_U.reset ;
wire [4:0] \add_5s_5ns_5_2_1_U5.top_add_5s_5ns_5_2_1_Adder_4_U.s ;
wire [1:0] \add_5s_5ns_5_2_1_U5.top_add_5s_5ns_5_2_1_Adder_4_U.u1.a ;
wire [1:0] \add_5s_5ns_5_2_1_U5.top_add_5s_5ns_5_2_1_Adder_4_U.u1.b ;
wire \add_5s_5ns_5_2_1_U5.top_add_5s_5ns_5_2_1_Adder_4_U.u1.cin ;
wire \add_5s_5ns_5_2_1_U5.top_add_5s_5ns_5_2_1_Adder_4_U.u1.cout ;
wire [1:0] \add_5s_5ns_5_2_1_U5.top_add_5s_5ns_5_2_1_Adder_4_U.u1.s ;
wire [2:0] \add_5s_5ns_5_2_1_U5.top_add_5s_5ns_5_2_1_Adder_4_U.u2.a ;
wire [2:0] \add_5s_5ns_5_2_1_U5.top_add_5s_5ns_5_2_1_Adder_4_U.u2.b ;
wire \add_5s_5ns_5_2_1_U5.top_add_5s_5ns_5_2_1_Adder_4_U.u2.cin ;
wire \add_5s_5ns_5_2_1_U5.top_add_5s_5ns_5_2_1_Adder_4_U.u2.cout ;
wire [2:0] \add_5s_5ns_5_2_1_U5.top_add_5s_5ns_5_2_1_Adder_4_U.u2.s ;
wire \add_5s_5s_5_2_1_U4.ce ;
wire \add_5s_5s_5_2_1_U4.clk ;
wire [4:0] \add_5s_5s_5_2_1_U4.din0 ;
wire [4:0] \add_5s_5s_5_2_1_U4.din1 ;
wire [4:0] \add_5s_5s_5_2_1_U4.dout ;
wire \add_5s_5s_5_2_1_U4.reset ;
wire [4:0] \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_3_U.a ;
wire [4:0] \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_3_U.ain_s0 ;
wire [4:0] \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_3_U.b ;
wire [4:0] \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_3_U.bin_s0 ;
wire \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_3_U.ce ;
wire \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_3_U.clk ;
wire \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_3_U.facout_s1 ;
wire \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_3_U.facout_s2 ;
wire [1:0] \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_3_U.fas_s1 ;
wire [2:0] \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_3_U.fas_s2 ;
wire \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_3_U.reset ;
wire [4:0] \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_3_U.s ;
wire [1:0] \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_3_U.u1.a ;
wire [1:0] \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_3_U.u1.b ;
wire \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_3_U.u1.cin ;
wire \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_3_U.u1.cout ;
wire [1:0] \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_3_U.u1.s ;
wire [2:0] \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_3_U.u2.a ;
wire [2:0] \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_3_U.u2.b ;
wire \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_3_U.u2.cin ;
wire \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_3_U.u2.cout ;
wire [2:0] \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_3_U.u2.s ;
wire ap_CS_fsm_state1;
wire ap_CS_fsm_state10;
wire ap_CS_fsm_state11;
wire ap_CS_fsm_state12;
wire ap_CS_fsm_state13;
wire ap_CS_fsm_state14;
wire ap_CS_fsm_state15;
wire ap_CS_fsm_state16;
wire ap_CS_fsm_state17;
wire ap_CS_fsm_state18;
wire ap_CS_fsm_state19;
wire ap_CS_fsm_state2;
wire ap_CS_fsm_state20;
wire ap_CS_fsm_state21;
wire ap_CS_fsm_state22;
wire ap_CS_fsm_state23;
wire ap_CS_fsm_state24;
wire ap_CS_fsm_state25;
wire ap_CS_fsm_state26;
wire ap_CS_fsm_state27;
wire ap_CS_fsm_state28;
wire ap_CS_fsm_state29;
wire ap_CS_fsm_state3;
wire ap_CS_fsm_state30;
wire ap_CS_fsm_state4;
wire ap_CS_fsm_state5;
wire ap_CS_fsm_state6;
wire ap_CS_fsm_state7;
wire ap_CS_fsm_state8;
wire ap_CS_fsm_state9;
wire [29:0] ap_NS_fsm;
wire ap_clk;
wire ap_done;
wire ap_idle;
wire ap_ready;
wire ap_rst;
wire ap_start;
wire [31:0] conv_i270_fu_408_p1;
wire [4:0] grp_fu_199_p0;
wire [4:0] grp_fu_199_p1;
wire [4:0] grp_fu_199_p2;
wire [2:0] grp_fu_228_p0;
wire [2:0] grp_fu_228_p2;
wire [2:0] grp_fu_253_p2;
wire [4:0] grp_fu_273_p0;
wire [4:0] grp_fu_273_p1;
wire [4:0] grp_fu_273_p2;
wire [4:0] grp_fu_292_p0;
wire [4:0] grp_fu_292_p2;
wire [2:0] grp_fu_324_p1;
wire [2:0] grp_fu_324_p2;
wire [4:0] grp_fu_386_p1;
wire [4:0] grp_fu_386_p2;
wire [31:0] grp_fu_411_p1;
wire [31:0] grp_fu_411_p2;
wire [31:0] grp_fu_420_p1;
wire [31:0] grp_fu_420_p2;
wire [33:0] grp_fu_447_p0;
wire [33:0] grp_fu_447_p1;
wire [33:0] grp_fu_447_p2;
wire [31:0] grp_fu_463_p2;
wire [31:0] grp_fu_503_p1;
wire [31:0] grp_fu_503_p2;
wire [34:0] grp_fu_532_p0;
wire [34:0] grp_fu_532_p1;
wire [34:0] grp_fu_532_p2;
wire [1:0] grp_fu_551_p1;
wire [1:0] grp_fu_551_p2;
wire [31:0] grp_fu_566_p2;
wire [31:0] grp_fu_604_p1;
wire [31:0] grp_fu_604_p2;
wire [31:0] grp_fu_612_p0;
wire [31:0] grp_fu_612_p2;
wire icmp_ln1495_fu_426_p2;
wire [1:0] icmp_ln1498_1_fu_337_p1;
wire icmp_ln1498_1_fu_337_p2;
wire icmp_ln1498_fu_377_p2;
wire icmp_ln851_1_fu_542_p2;
wire icmp_ln851_fu_209_p2;
wire \lshr_32ns_32s_32_7_1_U9.ce ;
wire \lshr_32ns_32s_32_7_1_U9.clk ;
wire [31:0] \lshr_32ns_32s_32_7_1_U9.din0 ;
wire [31:0] \lshr_32ns_32s_32_7_1_U9.din1 ;
wire [31:0] \lshr_32ns_32s_32_7_1_U9.din1_cast ;
wire [31:0] \lshr_32ns_32s_32_7_1_U9.din1_mask ;
wire [31:0] \lshr_32ns_32s_32_7_1_U9.dout ;
wire \lshr_32ns_32s_32_7_1_U9.reset ;
wire [3:0] op_0;
wire [7:0] op_1;
wire [1:0] op_10;
wire [7:0] op_14;
wire [3:0] op_15;
wire [7:0] op_16;
wire [1:0] op_17_V_fu_511_p3;
wire [1:0] op_2;
wire [31:0] op_29;
wire op_29_ap_vld;
wire op_3;
wire [31:0] op_4;
wire op_6_V_fu_306_p2;
wire [1:0] op_7;
wire op_8;
wire p_Result_1_fu_343_p3;
wire p_Result_2_fu_468_p3;
wire p_Result_3_fu_578_p3;
wire p_Result_s_fu_234_p3;
wire [1:0] ret_V_11_fu_571_p1;
wire [1:0] ret_V_11_fu_571_p3;
wire [2:0] ret_V_13_fu_246_p3;
wire [4:0] ret_V_15_fu_359_p3;
wire [31:0] ret_V_17_fu_484_p3;
wire [31:0] ret_V_19_fu_590_p3;
wire [33:0] rhs_5_fu_521_p3;
wire [3:0] rhs_fu_187_p3;
wire [1:0] select_ln1498_fu_330_p3;
wire [4:0] select_ln850_1_fu_353_p3;
wire [31:0] select_ln850_2_fu_478_p3;
wire [31:0] select_ln850_3_fu_585_p3;
wire [2:0] select_ln850_fu_241_p3;
wire [1:0] sext_ln1192_1_fu_258_p0;
wire [3:0] sext_ln1192_fu_183_p0;
wire [1:0] sext_ln1497_fu_312_p0;
wire [7:0] sext_ln1498_fu_373_p1;
wire [1:0] sext_ln545_fu_405_p0;
wire [3:0] sext_ln69_1_fu_597_p1;
wire [7:0] sext_ln703_1_fu_517_p0;
wire [7:0] sext_ln703_fu_432_p0;
wire [1:0] sext_ln727_fu_391_p0;
wire [2:0] sext_ln727_fu_391_p1;
wire [2:0] sext_ln835_fu_225_p1;
wire [4:0] sext_ln850_fu_289_p1;
wire \shl_32ns_32s_32_7_1_U8.ce ;
wire \shl_32ns_32s_32_7_1_U8.clk ;
wire [31:0] \shl_32ns_32s_32_7_1_U8.din0 ;
wire [31:0] \shl_32ns_32s_32_7_1_U8.din1 ;
wire [31:0] \shl_32ns_32s_32_7_1_U8.din1_cast ;
wire [31:0] \shl_32ns_32s_32_7_1_U8.din1_mask ;
wire [31:0] \shl_32ns_32s_32_7_1_U8.dout ;
wire \shl_32ns_32s_32_7_1_U8.reset ;
wire [1:0] shl_ln728_1_fu_298_p1;
wire [31:0] shl_ln728_1_fu_298_p3;
wire [1:0] shl_ln728_3_fu_394_p3;
wire [1:0] shl_ln_fu_366_p1;
wire [5:0] shl_ln_fu_366_p3;
wire \sub_3ns_3s_3_2_1_U6.ce ;
wire \sub_3ns_3s_3_2_1_U6.clk ;
wire [2:0] \sub_3ns_3s_3_2_1_U6.din0 ;
wire [2:0] \sub_3ns_3s_3_2_1_U6.din1 ;
wire [2:0] \sub_3ns_3s_3_2_1_U6.dout ;
wire \sub_3ns_3s_3_2_1_U6.reset ;
wire [2:0] \sub_3ns_3s_3_2_1_U6.top_sub_3ns_3s_3_2_1_Adder_5_U.a ;
wire [2:0] \sub_3ns_3s_3_2_1_U6.top_sub_3ns_3s_3_2_1_Adder_5_U.ain_s0 ;
wire [2:0] \sub_3ns_3s_3_2_1_U6.top_sub_3ns_3s_3_2_1_Adder_5_U.b ;
wire [2:0] \sub_3ns_3s_3_2_1_U6.top_sub_3ns_3s_3_2_1_Adder_5_U.bin_s0 ;
wire \sub_3ns_3s_3_2_1_U6.top_sub_3ns_3s_3_2_1_Adder_5_U.ce ;
wire \sub_3ns_3s_3_2_1_U6.top_sub_3ns_3s_3_2_1_Adder_5_U.clk ;
wire \sub_3ns_3s_3_2_1_U6.top_sub_3ns_3s_3_2_1_Adder_5_U.facout_s1 ;
wire \sub_3ns_3s_3_2_1_U6.top_sub_3ns_3s_3_2_1_Adder_5_U.facout_s2 ;
wire \sub_3ns_3s_3_2_1_U6.top_sub_3ns_3s_3_2_1_Adder_5_U.fas_s1 ;
wire [1:0] \sub_3ns_3s_3_2_1_U6.top_sub_3ns_3s_3_2_1_Adder_5_U.fas_s2 ;
wire \sub_3ns_3s_3_2_1_U6.top_sub_3ns_3s_3_2_1_Adder_5_U.reset ;
wire [2:0] \sub_3ns_3s_3_2_1_U6.top_sub_3ns_3s_3_2_1_Adder_5_U.s ;
wire \sub_3ns_3s_3_2_1_U6.top_sub_3ns_3s_3_2_1_Adder_5_U.u1.a ;
wire \sub_3ns_3s_3_2_1_U6.top_sub_3ns_3s_3_2_1_Adder_5_U.u1.b ;
wire \sub_3ns_3s_3_2_1_U6.top_sub_3ns_3s_3_2_1_Adder_5_U.u1.cin ;
wire \sub_3ns_3s_3_2_1_U6.top_sub_3ns_3s_3_2_1_Adder_5_U.u1.cout ;
wire \sub_3ns_3s_3_2_1_U6.top_sub_3ns_3s_3_2_1_Adder_5_U.u1.s ;
wire [1:0] \sub_3ns_3s_3_2_1_U6.top_sub_3ns_3s_3_2_1_Adder_5_U.u2.a ;
wire [1:0] \sub_3ns_3s_3_2_1_U6.top_sub_3ns_3s_3_2_1_Adder_5_U.u2.b ;
wire \sub_3ns_3s_3_2_1_U6.top_sub_3ns_3s_3_2_1_Adder_5_U.u2.cin ;
wire \sub_3ns_3s_3_2_1_U6.top_sub_3ns_3s_3_2_1_Adder_5_U.u2.cout ;
wire [1:0] \sub_3ns_3s_3_2_1_U6.top_sub_3ns_3s_3_2_1_Adder_5_U.u2.s ;
wire [3:0] tmp_1_fu_262_p3;
wire [5:0] tmp_4_fu_436_p3;
wire [1:0] tmp_fu_316_p1;
wire trunc_ln1497_1_fu_495_p1;
wire [1:0] trunc_ln1497_fu_491_p1;
wire [1:0] trunc_ln851_1_fu_350_p0;
wire trunc_ln851_1_fu_350_p1;
wire [7:0] trunc_ln851_2_fu_475_p0;
wire trunc_ln851_2_fu_475_p1;
wire [7:0] trunc_ln851_3_fu_538_p0;
wire [1:0] trunc_ln851_3_fu_538_p1;
wire [3:0] trunc_ln851_fu_205_p0;
wire [2:0] trunc_ln851_fu_205_p1;
wire [1:0] zext_ln1497_fu_508_p1;
wire [2:0] zext_ln835_fu_401_p1;


assign _037_ = icmp_ln851_1_reg_853 & ap_CS_fsm[24];
assign _038_ = _043_ & ap_CS_fsm[3];
assign _039_ = ap_CS_fsm[19] & tmp_reg_724;
assign _040_ = ap_CS_fsm[19] & _044_;
assign _041_ = _045_ & ap_CS_fsm[0];
assign _042_ = ap_start & ap_CS_fsm[0];
assign _043_ = ~ icmp_ln851_reg_628;
assign _044_ = ~ tmp_reg_724;
assign _045_ = ~ ap_start;
assign _046_ = select_ln1498_fu_330_p3 == op_7;
assign _047_ = { op_2[1], op_2[1], op_2, 4'h0 } == op_1;
assign _048_ = ! op_0[2:0];
always @(posedge \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_11_U.clk )
\add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_11_U.bin_s1  <= _050_;
always @(posedge \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_11_U.clk )
\add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_11_U.ain_s1  <= _049_;
always @(posedge \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_11_U.clk )
\add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_11_U.sum_s1  <= _052_;
always @(posedge \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_11_U.clk )
\add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_11_U.carry_s1  <= _051_;
assign _050_ = \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_11_U.ce  ? \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_11_U.b [1] : \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_11_U.bin_s1 ;
assign _049_ = \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_11_U.ce  ? \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_11_U.a [1] : \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_11_U.ain_s1 ;
assign _051_ = \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_11_U.ce  ? \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_11_U.facout_s1  : \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_11_U.carry_s1 ;
assign _052_ = \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_11_U.ce  ? \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_11_U.fas_s1  : \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_11_U.sum_s1 ;
assign _053_ = \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_11_U.u1.a  + \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_11_U.u1.b ;
assign { \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_11_U.u1.cout , \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_11_U.u1.s  } = _053_ + \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_11_U.u1.cin ;
assign _054_ = \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_11_U.u2.a  + \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_11_U.u2.b ;
assign { \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_11_U.u2.cout , \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_11_U.u2.s  } = _054_ + \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_11_U.u2.cin ;
always @(posedge \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.clk )
\add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.bin_s1  <= _056_;
always @(posedge \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.clk )
\add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.ain_s1  <= _055_;
always @(posedge \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.clk )
\add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.sum_s1  <= _058_;
always @(posedge \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.clk )
\add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.carry_s1  <= _057_;
assign _056_ = \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.ce  ? \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.b [31:16] : \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.bin_s1 ;
assign _055_ = \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.ce  ? \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.a [31:16] : \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.ain_s1 ;
assign _057_ = \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.ce  ? \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.facout_s1  : \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.carry_s1 ;
assign _058_ = \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.ce  ? \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.fas_s1  : \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.sum_s1 ;
assign _059_ = \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.u1.a  + \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.u1.b ;
assign { \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.u1.cout , \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.u1.s  } = _059_ + \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.u1.cin ;
assign _060_ = \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.u2.a  + \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.u2.b ;
assign { \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.u2.cout , \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.u2.s  } = _060_ + \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.u2.cin ;
always @(posedge \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_8_U.clk )
\add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_8_U.bin_s1  <= _062_;
always @(posedge \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_8_U.clk )
\add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_8_U.ain_s1  <= _061_;
always @(posedge \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_8_U.clk )
\add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_8_U.sum_s1  <= _064_;
always @(posedge \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_8_U.clk )
\add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_8_U.carry_s1  <= _063_;
assign _062_ = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_8_U.ce  ? \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_8_U.b [31:16] : \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_8_U.bin_s1 ;
assign _061_ = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_8_U.ce  ? \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_8_U.a [31:16] : \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_8_U.ain_s1 ;
assign _063_ = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_8_U.ce  ? \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_8_U.facout_s1  : \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_8_U.carry_s1 ;
assign _064_ = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_8_U.ce  ? \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_8_U.fas_s1  : \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_8_U.sum_s1 ;
assign _065_ = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_8_U.u1.a  + \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_8_U.u1.b ;
assign { \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_8_U.u1.cout , \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_8_U.u1.s  } = _065_ + \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_8_U.u1.cin ;
assign _066_ = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_8_U.u2.a  + \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_8_U.u2.b ;
assign { \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_8_U.u2.cout , \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_8_U.u2.s  } = _066_ + \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_8_U.u2.cin ;
always @(posedge \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_8_U.clk )
\add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_8_U.bin_s1  <= _068_;
always @(posedge \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_8_U.clk )
\add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_8_U.ain_s1  <= _067_;
always @(posedge \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_8_U.clk )
\add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_8_U.sum_s1  <= _070_;
always @(posedge \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_8_U.clk )
\add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_8_U.carry_s1  <= _069_;
assign _068_ = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_8_U.ce  ? \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_8_U.b [31:16] : \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_8_U.bin_s1 ;
assign _067_ = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_8_U.ce  ? \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_8_U.a [31:16] : \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_8_U.ain_s1 ;
assign _069_ = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_8_U.ce  ? \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_8_U.facout_s1  : \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_8_U.carry_s1 ;
assign _070_ = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_8_U.ce  ? \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_8_U.fas_s1  : \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_8_U.sum_s1 ;
assign _071_ = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_8_U.u1.a  + \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_8_U.u1.b ;
assign { \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_8_U.u1.cout , \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_8_U.u1.s  } = _071_ + \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_8_U.u1.cin ;
assign _072_ = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_8_U.u2.a  + \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_8_U.u2.b ;
assign { \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_8_U.u2.cout , \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_8_U.u2.s  } = _072_ + \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_8_U.u2.cin ;
always @(posedge \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.clk )
\add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.bin_s1  <= _074_;
always @(posedge \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.clk )
\add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.ain_s1  <= _073_;
always @(posedge \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.clk )
\add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.sum_s1  <= _076_;
always @(posedge \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.clk )
\add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.carry_s1  <= _075_;
assign _074_ = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.ce  ? \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.b [31:16] : \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.bin_s1 ;
assign _073_ = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.ce  ? \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.a [31:16] : \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.ain_s1 ;
assign _075_ = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.ce  ? \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.facout_s1  : \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.carry_s1 ;
assign _076_ = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.ce  ? \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.fas_s1  : \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.sum_s1 ;
assign _077_ = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.u1.a  + \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.u1.b ;
assign { \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.u1.cout , \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.u1.s  } = _077_ + \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.u1.cin ;
assign _078_ = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.u2.a  + \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.u2.b ;
assign { \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.u2.cout , \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.u2.s  } = _078_ + \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.u2.cin ;
always @(posedge \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_9_U.clk )
\add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_9_U.bin_s1  <= _080_;
always @(posedge \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_9_U.clk )
\add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_9_U.ain_s1  <= _079_;
always @(posedge \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_9_U.clk )
\add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_9_U.sum_s1  <= _082_;
always @(posedge \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_9_U.clk )
\add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_9_U.carry_s1  <= _081_;
assign _080_ = \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_9_U.ce  ? \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_9_U.b [31:16] : \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_9_U.bin_s1 ;
assign _079_ = \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_9_U.ce  ? \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_9_U.a [31:16] : \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_9_U.ain_s1 ;
assign _081_ = \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_9_U.ce  ? \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_9_U.facout_s1  : \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_9_U.carry_s1 ;
assign _082_ = \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_9_U.ce  ? \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_9_U.fas_s1  : \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_9_U.sum_s1 ;
assign _083_ = \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_9_U.u1.a  + \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_9_U.u1.b ;
assign { \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_9_U.u1.cout , \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_9_U.u1.s  } = _083_ + \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_9_U.u1.cin ;
assign _084_ = \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_9_U.u2.a  + \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_9_U.u2.b ;
assign { \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_9_U.u2.cout , \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_9_U.u2.s  } = _084_ + \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_9_U.u2.cin ;
always @(posedge \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_7_U.clk )
\add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_7_U.bin_s1  <= _086_;
always @(posedge \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_7_U.clk )
\add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_7_U.ain_s1  <= _085_;
always @(posedge \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_7_U.clk )
\add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_7_U.sum_s1  <= _088_;
always @(posedge \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_7_U.clk )
\add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_7_U.carry_s1  <= _087_;
assign _086_ = \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_7_U.ce  ? \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_7_U.b [33:17] : \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_7_U.bin_s1 ;
assign _085_ = \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_7_U.ce  ? \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_7_U.a [33:17] : \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_7_U.ain_s1 ;
assign _087_ = \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_7_U.ce  ? \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_7_U.facout_s1  : \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_7_U.carry_s1 ;
assign _088_ = \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_7_U.ce  ? \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_7_U.fas_s1  : \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_7_U.sum_s1 ;
assign _089_ = \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_7_U.u1.a  + \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_7_U.u1.b ;
assign { \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_7_U.u1.cout , \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_7_U.u1.s  } = _089_ + \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_7_U.u1.cin ;
assign _090_ = \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_7_U.u2.a  + \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_7_U.u2.b ;
assign { \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_7_U.u2.cout , \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_7_U.u2.s  } = _090_ + \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_7_U.u2.cin ;
always @(posedge \add_35s_35s_35_2_1_U13.top_add_35s_35s_35_2_1_Adder_10_U.clk )
\add_35s_35s_35_2_1_U13.top_add_35s_35s_35_2_1_Adder_10_U.bin_s1  <= _092_;
always @(posedge \add_35s_35s_35_2_1_U13.top_add_35s_35s_35_2_1_Adder_10_U.clk )
\add_35s_35s_35_2_1_U13.top_add_35s_35s_35_2_1_Adder_10_U.ain_s1  <= _091_;
always @(posedge \add_35s_35s_35_2_1_U13.top_add_35s_35s_35_2_1_Adder_10_U.clk )
\add_35s_35s_35_2_1_U13.top_add_35s_35s_35_2_1_Adder_10_U.sum_s1  <= _094_;
always @(posedge \add_35s_35s_35_2_1_U13.top_add_35s_35s_35_2_1_Adder_10_U.clk )
\add_35s_35s_35_2_1_U13.top_add_35s_35s_35_2_1_Adder_10_U.carry_s1  <= _093_;
assign _092_ = \add_35s_35s_35_2_1_U13.top_add_35s_35s_35_2_1_Adder_10_U.ce  ? \add_35s_35s_35_2_1_U13.top_add_35s_35s_35_2_1_Adder_10_U.b [34:17] : \add_35s_35s_35_2_1_U13.top_add_35s_35s_35_2_1_Adder_10_U.bin_s1 ;
assign _091_ = \add_35s_35s_35_2_1_U13.top_add_35s_35s_35_2_1_Adder_10_U.ce  ? \add_35s_35s_35_2_1_U13.top_add_35s_35s_35_2_1_Adder_10_U.a [34:17] : \add_35s_35s_35_2_1_U13.top_add_35s_35s_35_2_1_Adder_10_U.ain_s1 ;
assign _093_ = \add_35s_35s_35_2_1_U13.top_add_35s_35s_35_2_1_Adder_10_U.ce  ? \add_35s_35s_35_2_1_U13.top_add_35s_35s_35_2_1_Adder_10_U.facout_s1  : \add_35s_35s_35_2_1_U13.top_add_35s_35s_35_2_1_Adder_10_U.carry_s1 ;
assign _094_ = \add_35s_35s_35_2_1_U13.top_add_35s_35s_35_2_1_Adder_10_U.ce  ? \add_35s_35s_35_2_1_U13.top_add_35s_35s_35_2_1_Adder_10_U.fas_s1  : \add_35s_35s_35_2_1_U13.top_add_35s_35s_35_2_1_Adder_10_U.sum_s1 ;
assign _095_ = \add_35s_35s_35_2_1_U13.top_add_35s_35s_35_2_1_Adder_10_U.u1.a  + \add_35s_35s_35_2_1_U13.top_add_35s_35s_35_2_1_Adder_10_U.u1.b ;
assign { \add_35s_35s_35_2_1_U13.top_add_35s_35s_35_2_1_Adder_10_U.u1.cout , \add_35s_35s_35_2_1_U13.top_add_35s_35s_35_2_1_Adder_10_U.u1.s  } = _095_ + \add_35s_35s_35_2_1_U13.top_add_35s_35s_35_2_1_Adder_10_U.u1.cin ;
assign _096_ = \add_35s_35s_35_2_1_U13.top_add_35s_35s_35_2_1_Adder_10_U.u2.a  + \add_35s_35s_35_2_1_U13.top_add_35s_35s_35_2_1_Adder_10_U.u2.b ;
assign { \add_35s_35s_35_2_1_U13.top_add_35s_35s_35_2_1_Adder_10_U.u2.cout , \add_35s_35s_35_2_1_U13.top_add_35s_35s_35_2_1_Adder_10_U.u2.s  } = _096_ + \add_35s_35s_35_2_1_U13.top_add_35s_35s_35_2_1_Adder_10_U.u2.cin ;
always @(posedge \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_2_U.clk )
\add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_2_U.bin_s1  <= _098_;
always @(posedge \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_2_U.clk )
\add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_2_U.ain_s1  <= _097_;
always @(posedge \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_2_U.clk )
\add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_2_U.sum_s1  <= _100_;
always @(posedge \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_2_U.clk )
\add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_2_U.carry_s1  <= _099_;
assign _098_ = \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_2_U.ce  ? \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_2_U.b [2:1] : \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_2_U.bin_s1 ;
assign _097_ = \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_2_U.ce  ? \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_2_U.a [2:1] : \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_2_U.ain_s1 ;
assign _099_ = \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_2_U.ce  ? \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_2_U.facout_s1  : \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_2_U.carry_s1 ;
assign _100_ = \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_2_U.ce  ? \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_2_U.fas_s1  : \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_2_U.sum_s1 ;
assign _101_ = \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_2_U.u1.a  + \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_2_U.u1.b ;
assign { \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_2_U.u1.cout , \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_2_U.u1.s  } = _101_ + \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_2_U.u1.cin ;
assign _102_ = \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_2_U.u2.a  + \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_2_U.u2.b ;
assign { \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_2_U.u2.cout , \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_2_U.u2.s  } = _102_ + \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_2_U.u2.cin ;
always @(posedge \add_3s_3ns_3_2_1_U2.top_add_3s_3ns_3_2_1_Adder_1_U.clk )
\add_3s_3ns_3_2_1_U2.top_add_3s_3ns_3_2_1_Adder_1_U.bin_s1  <= _104_;
always @(posedge \add_3s_3ns_3_2_1_U2.top_add_3s_3ns_3_2_1_Adder_1_U.clk )
\add_3s_3ns_3_2_1_U2.top_add_3s_3ns_3_2_1_Adder_1_U.ain_s1  <= _103_;
always @(posedge \add_3s_3ns_3_2_1_U2.top_add_3s_3ns_3_2_1_Adder_1_U.clk )
\add_3s_3ns_3_2_1_U2.top_add_3s_3ns_3_2_1_Adder_1_U.sum_s1  <= _106_;
always @(posedge \add_3s_3ns_3_2_1_U2.top_add_3s_3ns_3_2_1_Adder_1_U.clk )
\add_3s_3ns_3_2_1_U2.top_add_3s_3ns_3_2_1_Adder_1_U.carry_s1  <= _105_;
assign _104_ = \add_3s_3ns_3_2_1_U2.top_add_3s_3ns_3_2_1_Adder_1_U.ce  ? \add_3s_3ns_3_2_1_U2.top_add_3s_3ns_3_2_1_Adder_1_U.b [2:1] : \add_3s_3ns_3_2_1_U2.top_add_3s_3ns_3_2_1_Adder_1_U.bin_s1 ;
assign _103_ = \add_3s_3ns_3_2_1_U2.top_add_3s_3ns_3_2_1_Adder_1_U.ce  ? \add_3s_3ns_3_2_1_U2.top_add_3s_3ns_3_2_1_Adder_1_U.a [2:1] : \add_3s_3ns_3_2_1_U2.top_add_3s_3ns_3_2_1_Adder_1_U.ain_s1 ;
assign _105_ = \add_3s_3ns_3_2_1_U2.top_add_3s_3ns_3_2_1_Adder_1_U.ce  ? \add_3s_3ns_3_2_1_U2.top_add_3s_3ns_3_2_1_Adder_1_U.facout_s1  : \add_3s_3ns_3_2_1_U2.top_add_3s_3ns_3_2_1_Adder_1_U.carry_s1 ;
assign _106_ = \add_3s_3ns_3_2_1_U2.top_add_3s_3ns_3_2_1_Adder_1_U.ce  ? \add_3s_3ns_3_2_1_U2.top_add_3s_3ns_3_2_1_Adder_1_U.fas_s1  : \add_3s_3ns_3_2_1_U2.top_add_3s_3ns_3_2_1_Adder_1_U.sum_s1 ;
assign _107_ = \add_3s_3ns_3_2_1_U2.top_add_3s_3ns_3_2_1_Adder_1_U.u1.a  + \add_3s_3ns_3_2_1_U2.top_add_3s_3ns_3_2_1_Adder_1_U.u1.b ;
assign { \add_3s_3ns_3_2_1_U2.top_add_3s_3ns_3_2_1_Adder_1_U.u1.cout , \add_3s_3ns_3_2_1_U2.top_add_3s_3ns_3_2_1_Adder_1_U.u1.s  } = _107_ + \add_3s_3ns_3_2_1_U2.top_add_3s_3ns_3_2_1_Adder_1_U.u1.cin ;
assign _108_ = \add_3s_3ns_3_2_1_U2.top_add_3s_3ns_3_2_1_Adder_1_U.u2.a  + \add_3s_3ns_3_2_1_U2.top_add_3s_3ns_3_2_1_Adder_1_U.u2.b ;
assign { \add_3s_3ns_3_2_1_U2.top_add_3s_3ns_3_2_1_Adder_1_U.u2.cout , \add_3s_3ns_3_2_1_U2.top_add_3s_3ns_3_2_1_Adder_1_U.u2.s  } = _108_ + \add_3s_3ns_3_2_1_U2.top_add_3s_3ns_3_2_1_Adder_1_U.u2.cin ;
always @(posedge \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_6_U.clk )
\add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_6_U.bin_s1  <= _110_;
always @(posedge \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_6_U.clk )
\add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_6_U.ain_s1  <= _109_;
always @(posedge \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_6_U.clk )
\add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_6_U.sum_s1  <= _112_;
always @(posedge \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_6_U.clk )
\add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_6_U.carry_s1  <= _111_;
assign _110_ = \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_6_U.ce  ? \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_6_U.b [4:2] : \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_6_U.bin_s1 ;
assign _109_ = \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_6_U.ce  ? \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_6_U.a [4:2] : \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_6_U.ain_s1 ;
assign _111_ = \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_6_U.ce  ? \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_6_U.facout_s1  : \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_6_U.carry_s1 ;
assign _112_ = \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_6_U.ce  ? \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_6_U.fas_s1  : \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_6_U.sum_s1 ;
assign _113_ = \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_6_U.u1.a  + \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_6_U.u1.b ;
assign { \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_6_U.u1.cout , \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_6_U.u1.s  } = _113_ + \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_6_U.u1.cin ;
assign _114_ = \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_6_U.u2.a  + \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_6_U.u2.b ;
assign { \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_6_U.u2.cout , \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_6_U.u2.s  } = _114_ + \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_6_U.u2.cin ;
always @(posedge \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.clk )
\add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.bin_s1  <= _116_;
always @(posedge \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.clk )
\add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.ain_s1  <= _115_;
always @(posedge \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.clk )
\add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.sum_s1  <= _118_;
always @(posedge \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.clk )
\add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.carry_s1  <= _117_;
assign _116_ = \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.ce  ? \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.b [4:2] : \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.bin_s1 ;
assign _115_ = \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.ce  ? \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.a [4:2] : \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.ain_s1 ;
assign _117_ = \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.ce  ? \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.facout_s1  : \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.carry_s1 ;
assign _118_ = \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.ce  ? \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.fas_s1  : \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.sum_s1 ;
assign _119_ = \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.u1.a  + \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.u1.b ;
assign { \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.u1.cout , \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.u1.s  } = _119_ + \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.u1.cin ;
assign _120_ = \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.u2.a  + \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.u2.b ;
assign { \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.u2.cout , \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.u2.s  } = _120_ + \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.u2.cin ;
always @(posedge \add_5s_5ns_5_2_1_U5.top_add_5s_5ns_5_2_1_Adder_4_U.clk )
\add_5s_5ns_5_2_1_U5.top_add_5s_5ns_5_2_1_Adder_4_U.bin_s1  <= _122_;
always @(posedge \add_5s_5ns_5_2_1_U5.top_add_5s_5ns_5_2_1_Adder_4_U.clk )
\add_5s_5ns_5_2_1_U5.top_add_5s_5ns_5_2_1_Adder_4_U.ain_s1  <= _121_;
always @(posedge \add_5s_5ns_5_2_1_U5.top_add_5s_5ns_5_2_1_Adder_4_U.clk )
\add_5s_5ns_5_2_1_U5.top_add_5s_5ns_5_2_1_Adder_4_U.sum_s1  <= _124_;
always @(posedge \add_5s_5ns_5_2_1_U5.top_add_5s_5ns_5_2_1_Adder_4_U.clk )
\add_5s_5ns_5_2_1_U5.top_add_5s_5ns_5_2_1_Adder_4_U.carry_s1  <= _123_;
assign _122_ = \add_5s_5ns_5_2_1_U5.top_add_5s_5ns_5_2_1_Adder_4_U.ce  ? \add_5s_5ns_5_2_1_U5.top_add_5s_5ns_5_2_1_Adder_4_U.b [4:2] : \add_5s_5ns_5_2_1_U5.top_add_5s_5ns_5_2_1_Adder_4_U.bin_s1 ;
assign _121_ = \add_5s_5ns_5_2_1_U5.top_add_5s_5ns_5_2_1_Adder_4_U.ce  ? \add_5s_5ns_5_2_1_U5.top_add_5s_5ns_5_2_1_Adder_4_U.a [4:2] : \add_5s_5ns_5_2_1_U5.top_add_5s_5ns_5_2_1_Adder_4_U.ain_s1 ;
assign _123_ = \add_5s_5ns_5_2_1_U5.top_add_5s_5ns_5_2_1_Adder_4_U.ce  ? \add_5s_5ns_5_2_1_U5.top_add_5s_5ns_5_2_1_Adder_4_U.facout_s1  : \add_5s_5ns_5_2_1_U5.top_add_5s_5ns_5_2_1_Adder_4_U.carry_s1 ;
assign _124_ = \add_5s_5ns_5_2_1_U5.top_add_5s_5ns_5_2_1_Adder_4_U.ce  ? \add_5s_5ns_5_2_1_U5.top_add_5s_5ns_5_2_1_Adder_4_U.fas_s1  : \add_5s_5ns_5_2_1_U5.top_add_5s_5ns_5_2_1_Adder_4_U.sum_s1 ;
assign _125_ = \add_5s_5ns_5_2_1_U5.top_add_5s_5ns_5_2_1_Adder_4_U.u1.a  + \add_5s_5ns_5_2_1_U5.top_add_5s_5ns_5_2_1_Adder_4_U.u1.b ;
assign { \add_5s_5ns_5_2_1_U5.top_add_5s_5ns_5_2_1_Adder_4_U.u1.cout , \add_5s_5ns_5_2_1_U5.top_add_5s_5ns_5_2_1_Adder_4_U.u1.s  } = _125_ + \add_5s_5ns_5_2_1_U5.top_add_5s_5ns_5_2_1_Adder_4_U.u1.cin ;
assign _126_ = \add_5s_5ns_5_2_1_U5.top_add_5s_5ns_5_2_1_Adder_4_U.u2.a  + \add_5s_5ns_5_2_1_U5.top_add_5s_5ns_5_2_1_Adder_4_U.u2.b ;
assign { \add_5s_5ns_5_2_1_U5.top_add_5s_5ns_5_2_1_Adder_4_U.u2.cout , \add_5s_5ns_5_2_1_U5.top_add_5s_5ns_5_2_1_Adder_4_U.u2.s  } = _126_ + \add_5s_5ns_5_2_1_U5.top_add_5s_5ns_5_2_1_Adder_4_U.u2.cin ;
always @(posedge \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_3_U.clk )
\add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_3_U.bin_s1  <= _128_;
always @(posedge \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_3_U.clk )
\add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_3_U.ain_s1  <= _127_;
always @(posedge \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_3_U.clk )
\add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_3_U.sum_s1  <= _130_;
always @(posedge \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_3_U.clk )
\add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_3_U.carry_s1  <= _129_;
assign _128_ = \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_3_U.ce  ? \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_3_U.b [4:2] : \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_3_U.bin_s1 ;
assign _127_ = \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_3_U.ce  ? \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_3_U.a [4:2] : \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_3_U.ain_s1 ;
assign _129_ = \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_3_U.ce  ? \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_3_U.facout_s1  : \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_3_U.carry_s1 ;
assign _130_ = \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_3_U.ce  ? \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_3_U.fas_s1  : \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_3_U.sum_s1 ;
assign _131_ = \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_3_U.u1.a  + \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_3_U.u1.b ;
assign { \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_3_U.u1.cout , \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_3_U.u1.s  } = _131_ + \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_3_U.u1.cin ;
assign _132_ = \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_3_U.u2.a  + \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_3_U.u2.b ;
assign { \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_3_U.u2.cout , \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_3_U.u2.s  } = _132_ + \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_3_U.u2.cin ;
always @(posedge \lshr_32ns_32s_32_7_1_U9.clk )
\lshr_32ns_32s_32_7_1_U9.dout_array[5]  <= _144_;
always @(posedge \lshr_32ns_32s_32_7_1_U9.clk )
\lshr_32ns_32s_32_7_1_U9.din1_cast_array[5]  <= _138_;
always @(posedge \lshr_32ns_32s_32_7_1_U9.clk )
\lshr_32ns_32s_32_7_1_U9.dout_array[4]  <= _143_;
always @(posedge \lshr_32ns_32s_32_7_1_U9.clk )
\lshr_32ns_32s_32_7_1_U9.din1_cast_array[4]  <= _137_;
always @(posedge \lshr_32ns_32s_32_7_1_U9.clk )
\lshr_32ns_32s_32_7_1_U9.dout_array[3]  <= _142_;
always @(posedge \lshr_32ns_32s_32_7_1_U9.clk )
\lshr_32ns_32s_32_7_1_U9.din1_cast_array[3]  <= _136_;
always @(posedge \lshr_32ns_32s_32_7_1_U9.clk )
\lshr_32ns_32s_32_7_1_U9.dout_array[2]  <= _141_;
always @(posedge \lshr_32ns_32s_32_7_1_U9.clk )
\lshr_32ns_32s_32_7_1_U9.din1_cast_array[2]  <= _135_;
always @(posedge \lshr_32ns_32s_32_7_1_U9.clk )
\lshr_32ns_32s_32_7_1_U9.dout_array[1]  <= _140_;
always @(posedge \lshr_32ns_32s_32_7_1_U9.clk )
\lshr_32ns_32s_32_7_1_U9.din1_cast_array[1]  <= _134_;
always @(posedge \lshr_32ns_32s_32_7_1_U9.clk )
\lshr_32ns_32s_32_7_1_U9.dout_array[0]  <= _139_;
always @(posedge \lshr_32ns_32s_32_7_1_U9.clk )
\lshr_32ns_32s_32_7_1_U9.din1_cast_array[0]  <= _133_;
assign _145_ = \lshr_32ns_32s_32_7_1_U9.ce  ? \lshr_32ns_32s_32_7_1_U9.din1_cast_array[4]  : \lshr_32ns_32s_32_7_1_U9.din1_cast_array[5] ;
assign _138_ = \lshr_32ns_32s_32_7_1_U9.reset  ? 32'd0 : _145_;
assign _146_ = \lshr_32ns_32s_32_7_1_U9.ce  ? _162_ : \lshr_32ns_32s_32_7_1_U9.dout_array[5] ;
assign _144_ = \lshr_32ns_32s_32_7_1_U9.reset  ? 32'd0 : _146_;
assign _147_ = \lshr_32ns_32s_32_7_1_U9.ce  ? \lshr_32ns_32s_32_7_1_U9.din1_cast_array[3]  : \lshr_32ns_32s_32_7_1_U9.din1_cast_array[4] ;
assign _137_ = \lshr_32ns_32s_32_7_1_U9.reset  ? 32'd0 : _147_;
assign _148_ = \lshr_32ns_32s_32_7_1_U9.ce  ? _161_ : \lshr_32ns_32s_32_7_1_U9.dout_array[4] ;
assign _143_ = \lshr_32ns_32s_32_7_1_U9.reset  ? 32'd0 : _148_;
assign _149_ = \lshr_32ns_32s_32_7_1_U9.ce  ? \lshr_32ns_32s_32_7_1_U9.din1_cast_array[2]  : \lshr_32ns_32s_32_7_1_U9.din1_cast_array[3] ;
assign _136_ = \lshr_32ns_32s_32_7_1_U9.reset  ? 32'd0 : _149_;
assign _150_ = \lshr_32ns_32s_32_7_1_U9.ce  ? _160_ : \lshr_32ns_32s_32_7_1_U9.dout_array[3] ;
assign _142_ = \lshr_32ns_32s_32_7_1_U9.reset  ? 32'd0 : _150_;
assign _151_ = \lshr_32ns_32s_32_7_1_U9.ce  ? \lshr_32ns_32s_32_7_1_U9.din1_cast_array[1]  : \lshr_32ns_32s_32_7_1_U9.din1_cast_array[2] ;
assign _135_ = \lshr_32ns_32s_32_7_1_U9.reset  ? 32'd0 : _151_;
assign _152_ = \lshr_32ns_32s_32_7_1_U9.ce  ? _159_ : \lshr_32ns_32s_32_7_1_U9.dout_array[2] ;
assign _141_ = \lshr_32ns_32s_32_7_1_U9.reset  ? 32'd0 : _152_;
assign _153_ = \lshr_32ns_32s_32_7_1_U9.ce  ? \lshr_32ns_32s_32_7_1_U9.din1_cast_array[0]  : \lshr_32ns_32s_32_7_1_U9.din1_cast_array[1] ;
assign _134_ = \lshr_32ns_32s_32_7_1_U9.reset  ? 32'd0 : _153_;
assign _154_ = \lshr_32ns_32s_32_7_1_U9.ce  ? _158_ : \lshr_32ns_32s_32_7_1_U9.dout_array[1] ;
assign _140_ = \lshr_32ns_32s_32_7_1_U9.reset  ? 32'd0 : _154_;
assign _155_ = \lshr_32ns_32s_32_7_1_U9.ce  ? \lshr_32ns_32s_32_7_1_U9.din1  : \lshr_32ns_32s_32_7_1_U9.din1_cast_array[0] ;
assign _133_ = \lshr_32ns_32s_32_7_1_U9.reset  ? 32'd0 : _155_;
assign _156_ = \lshr_32ns_32s_32_7_1_U9.ce  ? _157_ : \lshr_32ns_32s_32_7_1_U9.dout_array[0] ;
assign _139_ = \lshr_32ns_32s_32_7_1_U9.reset  ? 32'd0 : _156_;
assign _157_ = \lshr_32ns_32s_32_7_1_U9.din0  >> { \lshr_32ns_32s_32_7_1_U9.din1 [31:30], 30'h00000000 };
assign _158_ = \lshr_32ns_32s_32_7_1_U9.dout_array[0]  >> { \lshr_32ns_32s_32_7_1_U9.din1_cast_array[0] [29:25], 25'h0000000 };
assign _159_ = \lshr_32ns_32s_32_7_1_U9.dout_array[1]  >> { \lshr_32ns_32s_32_7_1_U9.din1_cast_array[1] [24:20], 20'h00000 };
assign _160_ = \lshr_32ns_32s_32_7_1_U9.dout_array[2]  >> { \lshr_32ns_32s_32_7_1_U9.din1_cast_array[2] [19:15], 15'h0000 };
assign _161_ = \lshr_32ns_32s_32_7_1_U9.dout_array[3]  >> { \lshr_32ns_32s_32_7_1_U9.din1_cast_array[3] [14:10], 10'h000 };
assign _162_ = \lshr_32ns_32s_32_7_1_U9.dout_array[4]  >> { \lshr_32ns_32s_32_7_1_U9.din1_cast_array[4] [9:5], 5'h00 };
assign \lshr_32ns_32s_32_7_1_U9.dout  = \lshr_32ns_32s_32_7_1_U9.dout_array[5]  >> \lshr_32ns_32s_32_7_1_U9.din1_cast_array[5] [4:0];
always @(posedge \shl_32ns_32s_32_7_1_U8.clk )
\shl_32ns_32s_32_7_1_U8.dout_array[5]  <= _174_;
always @(posedge \shl_32ns_32s_32_7_1_U8.clk )
\shl_32ns_32s_32_7_1_U8.din1_cast_array[5]  <= _168_;
always @(posedge \shl_32ns_32s_32_7_1_U8.clk )
\shl_32ns_32s_32_7_1_U8.dout_array[4]  <= _173_;
always @(posedge \shl_32ns_32s_32_7_1_U8.clk )
\shl_32ns_32s_32_7_1_U8.din1_cast_array[4]  <= _167_;
always @(posedge \shl_32ns_32s_32_7_1_U8.clk )
\shl_32ns_32s_32_7_1_U8.dout_array[3]  <= _172_;
always @(posedge \shl_32ns_32s_32_7_1_U8.clk )
\shl_32ns_32s_32_7_1_U8.din1_cast_array[3]  <= _166_;
always @(posedge \shl_32ns_32s_32_7_1_U8.clk )
\shl_32ns_32s_32_7_1_U8.dout_array[2]  <= _171_;
always @(posedge \shl_32ns_32s_32_7_1_U8.clk )
\shl_32ns_32s_32_7_1_U8.din1_cast_array[2]  <= _165_;
always @(posedge \shl_32ns_32s_32_7_1_U8.clk )
\shl_32ns_32s_32_7_1_U8.dout_array[1]  <= _170_;
always @(posedge \shl_32ns_32s_32_7_1_U8.clk )
\shl_32ns_32s_32_7_1_U8.din1_cast_array[1]  <= _164_;
always @(posedge \shl_32ns_32s_32_7_1_U8.clk )
\shl_32ns_32s_32_7_1_U8.dout_array[0]  <= _169_;
always @(posedge \shl_32ns_32s_32_7_1_U8.clk )
\shl_32ns_32s_32_7_1_U8.din1_cast_array[0]  <= _163_;
assign _175_ = \shl_32ns_32s_32_7_1_U8.ce  ? \shl_32ns_32s_32_7_1_U8.din1_cast_array[4]  : \shl_32ns_32s_32_7_1_U8.din1_cast_array[5] ;
assign _168_ = \shl_32ns_32s_32_7_1_U8.reset  ? 32'd0 : _175_;
assign _176_ = \shl_32ns_32s_32_7_1_U8.ce  ? _192_ : \shl_32ns_32s_32_7_1_U8.dout_array[5] ;
assign _174_ = \shl_32ns_32s_32_7_1_U8.reset  ? 32'd0 : _176_;
assign _177_ = \shl_32ns_32s_32_7_1_U8.ce  ? \shl_32ns_32s_32_7_1_U8.din1_cast_array[3]  : \shl_32ns_32s_32_7_1_U8.din1_cast_array[4] ;
assign _167_ = \shl_32ns_32s_32_7_1_U8.reset  ? 32'd0 : _177_;
assign _178_ = \shl_32ns_32s_32_7_1_U8.ce  ? _191_ : \shl_32ns_32s_32_7_1_U8.dout_array[4] ;
assign _173_ = \shl_32ns_32s_32_7_1_U8.reset  ? 32'd0 : _178_;
assign _179_ = \shl_32ns_32s_32_7_1_U8.ce  ? \shl_32ns_32s_32_7_1_U8.din1_cast_array[2]  : \shl_32ns_32s_32_7_1_U8.din1_cast_array[3] ;
assign _166_ = \shl_32ns_32s_32_7_1_U8.reset  ? 32'd0 : _179_;
assign _180_ = \shl_32ns_32s_32_7_1_U8.ce  ? _190_ : \shl_32ns_32s_32_7_1_U8.dout_array[3] ;
assign _172_ = \shl_32ns_32s_32_7_1_U8.reset  ? 32'd0 : _180_;
assign _181_ = \shl_32ns_32s_32_7_1_U8.ce  ? \shl_32ns_32s_32_7_1_U8.din1_cast_array[1]  : \shl_32ns_32s_32_7_1_U8.din1_cast_array[2] ;
assign _165_ = \shl_32ns_32s_32_7_1_U8.reset  ? 32'd0 : _181_;
assign _182_ = \shl_32ns_32s_32_7_1_U8.ce  ? _189_ : \shl_32ns_32s_32_7_1_U8.dout_array[2] ;
assign _171_ = \shl_32ns_32s_32_7_1_U8.reset  ? 32'd0 : _182_;
assign _183_ = \shl_32ns_32s_32_7_1_U8.ce  ? \shl_32ns_32s_32_7_1_U8.din1_cast_array[0]  : \shl_32ns_32s_32_7_1_U8.din1_cast_array[1] ;
assign _164_ = \shl_32ns_32s_32_7_1_U8.reset  ? 32'd0 : _183_;
assign _184_ = \shl_32ns_32s_32_7_1_U8.ce  ? _188_ : \shl_32ns_32s_32_7_1_U8.dout_array[1] ;
assign _170_ = \shl_32ns_32s_32_7_1_U8.reset  ? 32'd0 : _184_;
assign _185_ = \shl_32ns_32s_32_7_1_U8.ce  ? \shl_32ns_32s_32_7_1_U8.din1  : \shl_32ns_32s_32_7_1_U8.din1_cast_array[0] ;
assign _163_ = \shl_32ns_32s_32_7_1_U8.reset  ? 32'd0 : _185_;
assign _186_ = \shl_32ns_32s_32_7_1_U8.ce  ? _187_ : \shl_32ns_32s_32_7_1_U8.dout_array[0] ;
assign _169_ = \shl_32ns_32s_32_7_1_U8.reset  ? 32'd0 : _186_;
assign _187_ = \shl_32ns_32s_32_7_1_U8.din0  << { \shl_32ns_32s_32_7_1_U8.din1 [31:30], 30'h00000000 };
assign _188_ = \shl_32ns_32s_32_7_1_U8.dout_array[0]  << { \shl_32ns_32s_32_7_1_U8.din1_cast_array[0] [29:25], 25'h0000000 };
assign _189_ = \shl_32ns_32s_32_7_1_U8.dout_array[1]  << { \shl_32ns_32s_32_7_1_U8.din1_cast_array[1] [24:20], 20'h00000 };
assign _190_ = \shl_32ns_32s_32_7_1_U8.dout_array[2]  << { \shl_32ns_32s_32_7_1_U8.din1_cast_array[2] [19:15], 15'h0000 };
assign _191_ = \shl_32ns_32s_32_7_1_U8.dout_array[3]  << { \shl_32ns_32s_32_7_1_U8.din1_cast_array[3] [14:10], 10'h000 };
assign _192_ = \shl_32ns_32s_32_7_1_U8.dout_array[4]  << { \shl_32ns_32s_32_7_1_U8.din1_cast_array[4] [9:5], 5'h00 };
assign \shl_32ns_32s_32_7_1_U8.dout  = \shl_32ns_32s_32_7_1_U8.dout_array[5]  << \shl_32ns_32s_32_7_1_U8.din1_cast_array[5] [4:0];
assign \sub_3ns_3s_3_2_1_U6.top_sub_3ns_3s_3_2_1_Adder_5_U.bin_s0  = ~ \sub_3ns_3s_3_2_1_U6.top_sub_3ns_3s_3_2_1_Adder_5_U.b ;
always @(posedge \sub_3ns_3s_3_2_1_U6.top_sub_3ns_3s_3_2_1_Adder_5_U.clk )
\sub_3ns_3s_3_2_1_U6.top_sub_3ns_3s_3_2_1_Adder_5_U.bin_s1  <= _194_;
always @(posedge \sub_3ns_3s_3_2_1_U6.top_sub_3ns_3s_3_2_1_Adder_5_U.clk )
\sub_3ns_3s_3_2_1_U6.top_sub_3ns_3s_3_2_1_Adder_5_U.ain_s1  <= _193_;
always @(posedge \sub_3ns_3s_3_2_1_U6.top_sub_3ns_3s_3_2_1_Adder_5_U.clk )
\sub_3ns_3s_3_2_1_U6.top_sub_3ns_3s_3_2_1_Adder_5_U.sum_s1  <= _196_;
always @(posedge \sub_3ns_3s_3_2_1_U6.top_sub_3ns_3s_3_2_1_Adder_5_U.clk )
\sub_3ns_3s_3_2_1_U6.top_sub_3ns_3s_3_2_1_Adder_5_U.carry_s1  <= _195_;
assign _194_ = \sub_3ns_3s_3_2_1_U6.top_sub_3ns_3s_3_2_1_Adder_5_U.ce  ? \sub_3ns_3s_3_2_1_U6.top_sub_3ns_3s_3_2_1_Adder_5_U.bin_s0 [2:1] : \sub_3ns_3s_3_2_1_U6.top_sub_3ns_3s_3_2_1_Adder_5_U.bin_s1 ;
assign _193_ = \sub_3ns_3s_3_2_1_U6.top_sub_3ns_3s_3_2_1_Adder_5_U.ce  ? \sub_3ns_3s_3_2_1_U6.top_sub_3ns_3s_3_2_1_Adder_5_U.a [2:1] : \sub_3ns_3s_3_2_1_U6.top_sub_3ns_3s_3_2_1_Adder_5_U.ain_s1 ;
assign _195_ = \sub_3ns_3s_3_2_1_U6.top_sub_3ns_3s_3_2_1_Adder_5_U.ce  ? \sub_3ns_3s_3_2_1_U6.top_sub_3ns_3s_3_2_1_Adder_5_U.facout_s1  : \sub_3ns_3s_3_2_1_U6.top_sub_3ns_3s_3_2_1_Adder_5_U.carry_s1 ;
assign _196_ = \sub_3ns_3s_3_2_1_U6.top_sub_3ns_3s_3_2_1_Adder_5_U.ce  ? \sub_3ns_3s_3_2_1_U6.top_sub_3ns_3s_3_2_1_Adder_5_U.fas_s1  : \sub_3ns_3s_3_2_1_U6.top_sub_3ns_3s_3_2_1_Adder_5_U.sum_s1 ;
assign _197_ = \sub_3ns_3s_3_2_1_U6.top_sub_3ns_3s_3_2_1_Adder_5_U.u1.a  + \sub_3ns_3s_3_2_1_U6.top_sub_3ns_3s_3_2_1_Adder_5_U.u1.b ;
assign { \sub_3ns_3s_3_2_1_U6.top_sub_3ns_3s_3_2_1_Adder_5_U.u1.cout , \sub_3ns_3s_3_2_1_U6.top_sub_3ns_3s_3_2_1_Adder_5_U.u1.s  } = _197_ + \sub_3ns_3s_3_2_1_U6.top_sub_3ns_3s_3_2_1_Adder_5_U.u1.cin ;
assign _198_ = \sub_3ns_3s_3_2_1_U6.top_sub_3ns_3s_3_2_1_Adder_5_U.u2.a  + \sub_3ns_3s_3_2_1_U6.top_sub_3ns_3s_3_2_1_Adder_5_U.u2.b ;
assign { \sub_3ns_3s_3_2_1_U6.top_sub_3ns_3s_3_2_1_Adder_5_U.u2.cout , \sub_3ns_3s_3_2_1_U6.top_sub_3ns_3s_3_2_1_Adder_5_U.u2.s  } = _198_ + \sub_3ns_3s_3_2_1_U6.top_sub_3ns_3s_3_2_1_Adder_5_U.u2.cin ;
assign _199_ = $signed({ op_2, 30'h00000000 }) > $signed(op_4);
assign _200_ = $signed(op_2) < $signed({ 1'h0, icmp_ln1498_reg_739, 1'h0 });
assign _201_ = | op_16[1:0];
always @(posedge ap_clk)
trunc_ln1497_reg_818 <= _035_;
always @(posedge ap_clk)
trunc_ln1497_1_reg_823 <= _034_;
always @(posedge ap_clk)
sext_ln850_reg_690 <= _030_;
always @(posedge ap_clk)
sext_ln835_reg_643 <= _029_;
always @(posedge ap_clk)
ret_V_3_reg_650 <= _026_;
always @(posedge ap_clk)
ret_V_17_reg_813 <= _023_;
always @(posedge ap_clk)
ret_V_16_reg_796 <= _022_;
always @(posedge ap_clk)
ret_V_7_cast_reg_801 <= _027_;
always @(posedge ap_clk)
ret_V_14_reg_680 <= _019_;
always @(posedge ap_clk)
tmp_2_reg_685 <= _032_;
always @(posedge ap_clk)
ret_V_13_reg_655 <= _018_;
always @(posedge ap_clk)
ret_V_12_reg_633 <= _017_;
always @(posedge ap_clk)
ret_V_reg_638 <= _028_;
always @(posedge ap_clk)
ret_V_11_reg_885 <= _016_;
always @(posedge ap_clk)
ret_V_19_reg_890 <= _025_;
always @(posedge ap_clk)
op_21_V_reg_660 <= _012_;
always @(posedge ap_clk)
op_17_V_reg_833 <= _011_;
always @(posedge ap_clk)
op_25_V_reg_838 <= _014_;
always @(posedge ap_clk)
icmp_ln851_reg_628 <= _010_;
always @(posedge ap_clk)
icmp_ln851_1_reg_853 <= _009_;
always @(posedge ap_clk)
icmp_ln1498_reg_739 <= _008_;
always @(posedge ap_clk)
sub_ln1497_reg_745 <= _031_;
always @(posedge ap_clk)
tmp_reg_724 <= _033_;
always @(posedge ap_clk)
icmp_ln1498_1_reg_729 <= _007_;
always @(posedge ap_clk)
ret_V_15_reg_734 <= _021_;
always @(posedge ap_clk)
icmp_ln1495_reg_771 <= _006_;
always @(posedge ap_clk)
op_23_V_reg_776 <= _013_;
always @(posedge ap_clk)
add_ln69_reg_900 <= _004_;
always @(posedge ap_clk)
ret_V_18_reg_863 <= _024_;
always @(posedge ap_clk)
ret_V_15_cast_reg_868 <= _020_;
always @(posedge ap_clk)
add_ln69_1_reg_875 <= _003_;
always @(posedge ap_clk)
op_6_V_reg_703 <= _015_;
always @(posedge ap_clk)
add_ln691_reg_708 <= _002_;
always @(posedge ap_clk)
add_ln691_2_reg_880 <= _001_;
always @(posedge ap_clk)
add_ln691_1_reg_808 <= _000_;
always @(posedge ap_clk)
ap_CS_fsm <= _005_;
assign _036_ = _042_ ? 2'h2 : 2'h1;
assign _202_ = ap_CS_fsm == 1'h1;
function [29:0] _552_;
input [29:0] a;
input [899:0] b;
input [29:0] s;
case (s)
30'b000000000000000000000000000001:
_552_ = b[29:0];
30'b000000000000000000000000000010:
_552_ = b[59:30];
30'b000000000000000000000000000100:
_552_ = b[89:60];
30'b000000000000000000000000001000:
_552_ = b[119:90];
30'b000000000000000000000000010000:
_552_ = b[149:120];
30'b000000000000000000000000100000:
_552_ = b[179:150];
30'b000000000000000000000001000000:
_552_ = b[209:180];
30'b000000000000000000000010000000:
_552_ = b[239:210];
30'b000000000000000000000100000000:
_552_ = b[269:240];
30'b000000000000000000001000000000:
_552_ = b[299:270];
30'b000000000000000000010000000000:
_552_ = b[329:300];
30'b000000000000000000100000000000:
_552_ = b[359:330];
30'b000000000000000001000000000000:
_552_ = b[389:360];
30'b000000000000000010000000000000:
_552_ = b[419:390];
30'b000000000000000100000000000000:
_552_ = b[449:420];
30'b000000000000001000000000000000:
_552_ = b[479:450];
30'b000000000000010000000000000000:
_552_ = b[509:480];
30'b000000000000100000000000000000:
_552_ = b[539:510];
30'b000000000001000000000000000000:
_552_ = b[569:540];
30'b000000000010000000000000000000:
_552_ = b[599:570];
30'b000000000100000000000000000000:
_552_ = b[629:600];
30'b000000001000000000000000000000:
_552_ = b[659:630];
30'b000000010000000000000000000000:
_552_ = b[689:660];
30'b000000100000000000000000000000:
_552_ = b[719:690];
30'b000001000000000000000000000000:
_552_ = b[749:720];
30'b000010000000000000000000000000:
_552_ = b[779:750];
30'b000100000000000000000000000000:
_552_ = b[809:780];
30'b001000000000000000000000000000:
_552_ = b[839:810];
30'b010000000000000000000000000000:
_552_ = b[869:840];
30'b100000000000000000000000000000:
_552_ = b[899:870];
30'b000000000000000000000000000000:
_552_ = a;
default:
_552_ = 30'bx;
endcase
endfunction
assign ap_NS_fsm = _552_(30'hxxxxxxxx, { 28'h0000000, _036_, 870'h00000004000000200000010000000800000040000002000000100000008000000400000020000001000000080000004000000200000010000000800000040000002000000100000008000000400000020000001000000080000004000000200000010000000800000000000001 }, { _202_, _231_, _230_, _229_, _228_, _227_, _226_, _225_, _224_, _223_, _222_, _221_, _220_, _219_, _218_, _217_, _216_, _215_, _214_, _213_, _212_, _211_, _210_, _209_, _208_, _207_, _206_, _205_, _204_, _203_ });
assign _203_ = ap_CS_fsm == 30'h20000000;
assign _204_ = ap_CS_fsm == 29'h10000000;
assign _205_ = ap_CS_fsm == 28'h8000000;
assign _206_ = ap_CS_fsm == 27'h4000000;
assign _207_ = ap_CS_fsm == 26'h2000000;
assign _208_ = ap_CS_fsm == 25'h1000000;
assign _209_ = ap_CS_fsm == 24'h800000;
assign _210_ = ap_CS_fsm == 23'h400000;
assign _211_ = ap_CS_fsm == 22'h200000;
assign _212_ = ap_CS_fsm == 21'h100000;
assign _213_ = ap_CS_fsm == 20'h80000;
assign _214_ = ap_CS_fsm == 19'h40000;
assign _215_ = ap_CS_fsm == 18'h20000;
assign _216_ = ap_CS_fsm == 17'h10000;
assign _217_ = ap_CS_fsm == 16'h8000;
assign _218_ = ap_CS_fsm == 15'h4000;
assign _219_ = ap_CS_fsm == 14'h2000;
assign _220_ = ap_CS_fsm == 13'h1000;
assign _221_ = ap_CS_fsm == 12'h800;
assign _222_ = ap_CS_fsm == 11'h400;
assign _223_ = ap_CS_fsm == 10'h200;
assign _224_ = ap_CS_fsm == 9'h100;
assign _225_ = ap_CS_fsm == 8'h80;
assign _226_ = ap_CS_fsm == 7'h40;
assign _227_ = ap_CS_fsm == 6'h20;
assign _228_ = ap_CS_fsm == 5'h10;
assign _229_ = ap_CS_fsm == 4'h8;
assign _230_ = ap_CS_fsm == 3'h4;
assign _231_ = ap_CS_fsm == 2'h2;
assign op_29_ap_vld = ap_CS_fsm[29] ? 1'h1 : 1'h0;
assign ap_idle = _041_ ? 1'h1 : 1'h0;
assign _035_ = _040_ ? grp_fu_411_p2[1:0] : trunc_ln1497_reg_818;
assign _034_ = _039_ ? grp_fu_420_p2[0] : trunc_ln1497_1_reg_823;
assign _030_ = ap_CS_fsm[9] ? { tmp_2_reg_685[3], tmp_2_reg_685 } : sext_ln850_reg_690;
assign _029_ = ap_CS_fsm[2] ? { ret_V_reg_638[1], ret_V_reg_638 } : sext_ln835_reg_643;
assign _026_ = _038_ ? grp_fu_228_p2 : ret_V_3_reg_650;
assign _023_ = ap_CS_fsm[18] ? ret_V_17_fu_484_p3 : ret_V_17_reg_813;
assign _027_ = ap_CS_fsm[15] ? grp_fu_447_p2[32:1] : ret_V_7_cast_reg_801;
assign _022_ = ap_CS_fsm[15] ? grp_fu_447_p2 : ret_V_16_reg_796;
assign _032_ = ap_CS_fsm[8] ? grp_fu_273_p2[4:1] : tmp_2_reg_685;
assign _019_ = ap_CS_fsm[8] ? grp_fu_273_p2 : ret_V_14_reg_680;
assign _018_ = ap_CS_fsm[4] ? ret_V_13_fu_246_p3 : ret_V_13_reg_655;
assign _028_ = ap_CS_fsm[1] ? grp_fu_199_p2[4:3] : ret_V_reg_638;
assign _017_ = ap_CS_fsm[1] ? grp_fu_199_p2 : ret_V_12_reg_633;
assign _025_ = ap_CS_fsm[25] ? ret_V_19_fu_590_p3 : ret_V_19_reg_890;
assign _016_ = ap_CS_fsm[25] ? ret_V_11_fu_571_p3 : ret_V_11_reg_885;
assign _012_ = ap_CS_fsm[6] ? grp_fu_253_p2 : op_21_V_reg_660;
assign _014_ = ap_CS_fsm[20] ? grp_fu_503_p2 : op_25_V_reg_838;
assign _011_ = ap_CS_fsm[20] ? op_17_V_fu_511_p3 : op_17_V_reg_833;
assign _010_ = ap_CS_fsm[0] ? icmp_ln851_fu_209_p2 : icmp_ln851_reg_628;
assign _009_ = ap_CS_fsm[21] ? icmp_ln851_1_fu_542_p2 : icmp_ln851_1_reg_853;
assign _031_ = ap_CS_fsm[12] ? grp_fu_324_p2 : sub_ln1497_reg_745;
assign _008_ = ap_CS_fsm[12] ? icmp_ln1498_fu_377_p2 : icmp_ln1498_reg_739;
assign _021_ = ap_CS_fsm[11] ? ret_V_15_fu_359_p3 : ret_V_15_reg_734;
assign _007_ = ap_CS_fsm[11] ? icmp_ln1498_1_fu_337_p2 : icmp_ln1498_1_reg_729;
assign _033_ = ap_CS_fsm[11] ? op_7[1] : tmp_reg_724;
assign _013_ = ap_CS_fsm[13] ? grp_fu_386_p2 : op_23_V_reg_776;
assign _006_ = ap_CS_fsm[13] ? icmp_ln1495_fu_426_p2 : icmp_ln1495_reg_771;
assign _004_ = ap_CS_fsm[27] ? grp_fu_604_p2 : add_ln69_reg_900;
assign _003_ = ap_CS_fsm[22] ? grp_fu_551_p2 : add_ln69_1_reg_875;
assign _020_ = ap_CS_fsm[22] ? grp_fu_532_p2[33:2] : ret_V_15_cast_reg_868;
assign _024_ = ap_CS_fsm[22] ? grp_fu_532_p2 : ret_V_18_reg_863;
assign _002_ = ap_CS_fsm[10] ? grp_fu_292_p2 : add_ln691_reg_708;
assign _015_ = ap_CS_fsm[10] ? op_6_V_fu_306_p2 : op_6_V_reg_703;
assign _001_ = _037_ ? grp_fu_566_p2 : add_ln691_2_reg_880;
assign _000_ = ap_CS_fsm[17] ? grp_fu_463_p2 : add_ln691_1_reg_808;
assign _005_ = ap_rst ? 30'h00000001 : ap_NS_fsm;
assign icmp_ln1495_fu_426_p2 = _200_ ? 1'h1 : 1'h0;
assign icmp_ln1498_1_fu_337_p2 = _046_ ? 1'h1 : 1'h0;
assign icmp_ln1498_fu_377_p2 = _047_ ? 1'h1 : 1'h0;
assign icmp_ln851_1_fu_542_p2 = _201_ ? 1'h1 : 1'h0;
assign icmp_ln851_fu_209_p2 = _048_ ? 1'h1 : 1'h0;
assign op_17_V_fu_511_p3 = tmp_reg_724 ? { 1'h0, trunc_ln1497_1_reg_823 } : trunc_ln1497_reg_818;
assign op_6_V_fu_306_p2 = _199_ ? 1'h1 : 1'h0;
assign ret_V_11_fu_571_p3 = op_3 ? op_7 : 2'h0;
assign ret_V_13_fu_246_p3 = ret_V_12_reg_633[4] ? select_ln850_fu_241_p3 : sext_ln835_reg_643;
assign ret_V_15_fu_359_p3 = ret_V_14_reg_680[4] ? select_ln850_1_fu_353_p3 : sext_ln850_reg_690;
assign ret_V_17_fu_484_p3 = ret_V_16_reg_796[33] ? select_ln850_2_fu_478_p3 : ret_V_7_cast_reg_801;
assign ret_V_19_fu_590_p3 = ret_V_18_reg_863[34] ? select_ln850_3_fu_585_p3 : ret_V_15_cast_reg_868;
assign select_ln1498_fu_330_p3 = op_6_V_reg_703 ? 2'h3 : 2'h0;
assign select_ln850_1_fu_353_p3 = op_10[0] ? add_ln691_reg_708 : sext_ln850_reg_690;
assign select_ln850_2_fu_478_p3 = op_14[0] ? add_ln691_1_reg_808 : ret_V_7_cast_reg_801;
assign select_ln850_3_fu_585_p3 = icmp_ln851_1_reg_853 ? add_ln691_2_reg_880 : ret_V_15_cast_reg_868;
assign select_ln850_fu_241_p3 = icmp_ln851_reg_628 ? sext_ln835_reg_643 : ret_V_3_reg_650;
assign ap_CS_fsm_state1 = ap_CS_fsm[0];
assign ap_CS_fsm_state10 = ap_CS_fsm[9];
assign ap_CS_fsm_state11 = ap_CS_fsm[10];
assign ap_CS_fsm_state12 = ap_CS_fsm[11];
assign ap_CS_fsm_state13 = ap_CS_fsm[12];
assign ap_CS_fsm_state14 = ap_CS_fsm[13];
assign ap_CS_fsm_state15 = ap_CS_fsm[14];
assign ap_CS_fsm_state16 = ap_CS_fsm[15];
assign ap_CS_fsm_state17 = ap_CS_fsm[16];
assign ap_CS_fsm_state18 = ap_CS_fsm[17];
assign ap_CS_fsm_state19 = ap_CS_fsm[18];
assign ap_CS_fsm_state2 = ap_CS_fsm[1];
assign ap_CS_fsm_state20 = ap_CS_fsm[19];
assign ap_CS_fsm_state21 = ap_CS_fsm[20];
assign ap_CS_fsm_state22 = ap_CS_fsm[21];
assign ap_CS_fsm_state23 = ap_CS_fsm[22];
assign ap_CS_fsm_state24 = ap_CS_fsm[23];
assign ap_CS_fsm_state25 = ap_CS_fsm[24];
assign ap_CS_fsm_state26 = ap_CS_fsm[25];
assign ap_CS_fsm_state27 = ap_CS_fsm[26];
assign ap_CS_fsm_state28 = ap_CS_fsm[27];
assign ap_CS_fsm_state29 = ap_CS_fsm[28];
assign ap_CS_fsm_state3 = ap_CS_fsm[2];
assign ap_CS_fsm_state30 = ap_CS_fsm[29];
assign ap_CS_fsm_state4 = ap_CS_fsm[3];
assign ap_CS_fsm_state5 = ap_CS_fsm[4];
assign ap_CS_fsm_state6 = ap_CS_fsm[5];
assign ap_CS_fsm_state7 = ap_CS_fsm[6];
assign ap_CS_fsm_state8 = ap_CS_fsm[7];
assign ap_CS_fsm_state9 = ap_CS_fsm[8];
assign ap_done = op_29_ap_vld;
assign ap_ready = op_29_ap_vld;
assign conv_i270_fu_408_p1 = { 31'h00000000, icmp_ln1498_reg_739 };
assign grp_fu_199_p0 = { 1'h0, op_8, 3'h0 };
assign grp_fu_199_p1 = { op_0[3], op_0 };
assign grp_fu_228_p0 = { ret_V_reg_638[1], ret_V_reg_638 };
assign grp_fu_273_p0 = { op_21_V_reg_660[2], op_21_V_reg_660, 1'h0 };
assign grp_fu_273_p1 = { op_10[1], op_10[1], op_10[1], op_10 };
assign grp_fu_292_p0 = { tmp_2_reg_685[3], tmp_2_reg_685 };
assign grp_fu_324_p1 = { op_7[1], op_7 };
assign grp_fu_386_p1 = { 4'h0, icmp_ln1498_1_reg_729 };
assign grp_fu_411_p1 = { op_7[1], op_7[1], op_7[1], op_7[1], op_7[1], op_7[1], op_7[1], op_7[1], op_7[1], op_7[1], op_7[1], op_7[1], op_7[1], op_7[1], op_7[1], op_7[1], op_7[1], op_7[1], op_7[1], op_7[1], op_7[1], op_7[1], op_7[1], op_7[1], op_7[1], op_7[1], op_7[1], op_7[1], op_7[1], op_7[1], op_7 };
assign grp_fu_420_p1 = { sub_ln1497_reg_745[2], sub_ln1497_reg_745[2], sub_ln1497_reg_745[2], sub_ln1497_reg_745[2], sub_ln1497_reg_745[2], sub_ln1497_reg_745[2], sub_ln1497_reg_745[2], sub_ln1497_reg_745[2], sub_ln1497_reg_745[2], sub_ln1497_reg_745[2], sub_ln1497_reg_745[2], sub_ln1497_reg_745[2], sub_ln1497_reg_745[2], sub_ln1497_reg_745[2], sub_ln1497_reg_745[2], sub_ln1497_reg_745[2], sub_ln1497_reg_745[2], sub_ln1497_reg_745[2], sub_ln1497_reg_745[2], sub_ln1497_reg_745[2], sub_ln1497_reg_745[2], sub_ln1497_reg_745[2], sub_ln1497_reg_745[2], sub_ln1497_reg_745[2], sub_ln1497_reg_745[2], sub_ln1497_reg_745[2], sub_ln1497_reg_745[2], sub_ln1497_reg_745[2], sub_ln1497_reg_745[2], sub_ln1497_reg_745 };
assign grp_fu_447_p0 = { op_23_V_reg_776[4], op_23_V_reg_776[4], op_23_V_reg_776[4], op_23_V_reg_776[4], op_23_V_reg_776[4], op_23_V_reg_776[4], op_23_V_reg_776[4], op_23_V_reg_776[4], op_23_V_reg_776[4], op_23_V_reg_776[4], op_23_V_reg_776[4], op_23_V_reg_776[4], op_23_V_reg_776[4], op_23_V_reg_776[4], op_23_V_reg_776[4], op_23_V_reg_776[4], op_23_V_reg_776[4], op_23_V_reg_776[4], op_23_V_reg_776[4], op_23_V_reg_776[4], op_23_V_reg_776[4], op_23_V_reg_776[4], op_23_V_reg_776[4], op_23_V_reg_776[4], op_23_V_reg_776[4], op_23_V_reg_776[4], op_23_V_reg_776[4], op_23_V_reg_776[4], op_23_V_reg_776, 1'h0 };
assign grp_fu_447_p1 = { op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14 };
assign grp_fu_503_p1 = { op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15 };
assign grp_fu_532_p0 = { op_25_V_reg_838[31], op_25_V_reg_838, 2'h0 };
assign grp_fu_532_p1 = { op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16 };
assign grp_fu_551_p1 = { 1'h0, icmp_ln1495_reg_771 };
assign grp_fu_604_p1 = { 28'h0000000, ret_V_11_reg_885[1], ret_V_11_reg_885[1], ret_V_11_reg_885 };
assign grp_fu_612_p0 = { 30'h00000000, add_ln69_1_reg_875 };
assign icmp_ln1498_1_fu_337_p1 = op_7;
assign op_29 = grp_fu_612_p2;
assign p_Result_1_fu_343_p3 = ret_V_14_reg_680[4];
assign p_Result_2_fu_468_p3 = ret_V_16_reg_796[33];
assign p_Result_3_fu_578_p3 = ret_V_18_reg_863[34];
assign p_Result_s_fu_234_p3 = ret_V_12_reg_633[4];
assign ret_V_11_fu_571_p1 = op_7;
assign rhs_5_fu_521_p3 = { op_25_V_reg_838, 2'h0 };
assign rhs_fu_187_p3 = { op_8, 3'h0 };
assign sext_ln1192_1_fu_258_p0 = op_10;
assign sext_ln1192_fu_183_p0 = op_0;
assign sext_ln1497_fu_312_p0 = op_7;
assign sext_ln1498_fu_373_p1 = { op_2[1], op_2[1], op_2, 4'h0 };
assign sext_ln545_fu_405_p0 = op_7;
assign sext_ln69_1_fu_597_p1 = { ret_V_11_reg_885[1], ret_V_11_reg_885[1], ret_V_11_reg_885 };
assign sext_ln703_1_fu_517_p0 = op_16;
assign sext_ln703_fu_432_p0 = op_14;
assign sext_ln727_fu_391_p0 = op_2;
assign sext_ln727_fu_391_p1 = { op_2[1], op_2 };
assign sext_ln835_fu_225_p1 = { ret_V_reg_638[1], ret_V_reg_638 };
assign sext_ln850_fu_289_p1 = { tmp_2_reg_685[3], tmp_2_reg_685 };
assign shl_ln728_1_fu_298_p1 = op_2;
assign shl_ln728_1_fu_298_p3 = { op_2, 30'h00000000 };
assign shl_ln728_3_fu_394_p3 = { icmp_ln1498_reg_739, 1'h0 };
assign shl_ln_fu_366_p1 = op_2;
assign shl_ln_fu_366_p3 = { op_2, 4'h0 };
assign tmp_1_fu_262_p3 = { op_21_V_reg_660, 1'h0 };
assign tmp_4_fu_436_p3 = { op_23_V_reg_776, 1'h0 };
assign tmp_fu_316_p1 = op_7;
assign trunc_ln1497_1_fu_495_p1 = grp_fu_420_p2[0];
assign trunc_ln1497_fu_491_p1 = grp_fu_411_p2[1:0];
assign trunc_ln851_1_fu_350_p0 = op_10;
assign trunc_ln851_1_fu_350_p1 = op_10[0];
assign trunc_ln851_2_fu_475_p0 = op_14;
assign trunc_ln851_2_fu_475_p1 = op_14[0];
assign trunc_ln851_3_fu_538_p0 = op_16;
assign trunc_ln851_3_fu_538_p1 = op_16[1:0];
assign trunc_ln851_fu_205_p0 = op_0;
assign trunc_ln851_fu_205_p1 = op_0[2:0];
assign zext_ln1497_fu_508_p1 = { 1'h0, trunc_ln1497_1_reg_823 };
assign zext_ln835_fu_401_p1 = { 1'h0, icmp_ln1498_reg_739, 1'h0 };
assign \sub_3ns_3s_3_2_1_U6.top_sub_3ns_3s_3_2_1_Adder_5_U.ain_s0  = \sub_3ns_3s_3_2_1_U6.top_sub_3ns_3s_3_2_1_Adder_5_U.a ;
assign \sub_3ns_3s_3_2_1_U6.top_sub_3ns_3s_3_2_1_Adder_5_U.s  = { \sub_3ns_3s_3_2_1_U6.top_sub_3ns_3s_3_2_1_Adder_5_U.fas_s2 , \sub_3ns_3s_3_2_1_U6.top_sub_3ns_3s_3_2_1_Adder_5_U.sum_s1  };
assign \sub_3ns_3s_3_2_1_U6.top_sub_3ns_3s_3_2_1_Adder_5_U.u2.a  = \sub_3ns_3s_3_2_1_U6.top_sub_3ns_3s_3_2_1_Adder_5_U.ain_s1 ;
assign \sub_3ns_3s_3_2_1_U6.top_sub_3ns_3s_3_2_1_Adder_5_U.u2.b  = \sub_3ns_3s_3_2_1_U6.top_sub_3ns_3s_3_2_1_Adder_5_U.bin_s1 ;
assign \sub_3ns_3s_3_2_1_U6.top_sub_3ns_3s_3_2_1_Adder_5_U.u2.cin  = \sub_3ns_3s_3_2_1_U6.top_sub_3ns_3s_3_2_1_Adder_5_U.carry_s1 ;
assign \sub_3ns_3s_3_2_1_U6.top_sub_3ns_3s_3_2_1_Adder_5_U.facout_s2  = \sub_3ns_3s_3_2_1_U6.top_sub_3ns_3s_3_2_1_Adder_5_U.u2.cout ;
assign \sub_3ns_3s_3_2_1_U6.top_sub_3ns_3s_3_2_1_Adder_5_U.fas_s2  = \sub_3ns_3s_3_2_1_U6.top_sub_3ns_3s_3_2_1_Adder_5_U.u2.s ;
assign \sub_3ns_3s_3_2_1_U6.top_sub_3ns_3s_3_2_1_Adder_5_U.u1.a  = \sub_3ns_3s_3_2_1_U6.top_sub_3ns_3s_3_2_1_Adder_5_U.a [0];
assign \sub_3ns_3s_3_2_1_U6.top_sub_3ns_3s_3_2_1_Adder_5_U.u1.b  = \sub_3ns_3s_3_2_1_U6.top_sub_3ns_3s_3_2_1_Adder_5_U.bin_s0 [0];
assign \sub_3ns_3s_3_2_1_U6.top_sub_3ns_3s_3_2_1_Adder_5_U.u1.cin  = 1'h1;
assign \sub_3ns_3s_3_2_1_U6.top_sub_3ns_3s_3_2_1_Adder_5_U.facout_s1  = \sub_3ns_3s_3_2_1_U6.top_sub_3ns_3s_3_2_1_Adder_5_U.u1.cout ;
assign \sub_3ns_3s_3_2_1_U6.top_sub_3ns_3s_3_2_1_Adder_5_U.fas_s1  = \sub_3ns_3s_3_2_1_U6.top_sub_3ns_3s_3_2_1_Adder_5_U.u1.s ;
assign \sub_3ns_3s_3_2_1_U6.top_sub_3ns_3s_3_2_1_Adder_5_U.a  = \sub_3ns_3s_3_2_1_U6.din0 ;
assign \sub_3ns_3s_3_2_1_U6.top_sub_3ns_3s_3_2_1_Adder_5_U.b  = \sub_3ns_3s_3_2_1_U6.din1 ;
assign \sub_3ns_3s_3_2_1_U6.top_sub_3ns_3s_3_2_1_Adder_5_U.ce  = \sub_3ns_3s_3_2_1_U6.ce ;
assign \sub_3ns_3s_3_2_1_U6.top_sub_3ns_3s_3_2_1_Adder_5_U.clk  = \sub_3ns_3s_3_2_1_U6.clk ;
assign \sub_3ns_3s_3_2_1_U6.top_sub_3ns_3s_3_2_1_Adder_5_U.reset  = \sub_3ns_3s_3_2_1_U6.reset ;
assign \sub_3ns_3s_3_2_1_U6.dout  = \sub_3ns_3s_3_2_1_U6.top_sub_3ns_3s_3_2_1_Adder_5_U.s ;
assign \sub_3ns_3s_3_2_1_U6.ce  = 1'h1;
assign \sub_3ns_3s_3_2_1_U6.clk  = ap_clk;
assign \sub_3ns_3s_3_2_1_U6.din0  = 3'h0;
assign \sub_3ns_3s_3_2_1_U6.din1  = { op_7[1], op_7 };
assign grp_fu_324_p2 = \sub_3ns_3s_3_2_1_U6.dout ;
assign \sub_3ns_3s_3_2_1_U6.reset  = ap_rst;
assign \shl_32ns_32s_32_7_1_U8.din1_cast  = \shl_32ns_32s_32_7_1_U8.din1 ;
assign \shl_32ns_32s_32_7_1_U8.din1_mask  = 32'd31;
assign \shl_32ns_32s_32_7_1_U8.ce  = 1'h1;
assign \shl_32ns_32s_32_7_1_U8.clk  = ap_clk;
assign \shl_32ns_32s_32_7_1_U8.din0  = { 31'h00000000, icmp_ln1498_reg_739 };
assign \shl_32ns_32s_32_7_1_U8.din1  = { op_7[1], op_7[1], op_7[1], op_7[1], op_7[1], op_7[1], op_7[1], op_7[1], op_7[1], op_7[1], op_7[1], op_7[1], op_7[1], op_7[1], op_7[1], op_7[1], op_7[1], op_7[1], op_7[1], op_7[1], op_7[1], op_7[1], op_7[1], op_7[1], op_7[1], op_7[1], op_7[1], op_7[1], op_7[1], op_7[1], op_7 };
assign grp_fu_411_p2 = \shl_32ns_32s_32_7_1_U8.dout ;
assign \shl_32ns_32s_32_7_1_U8.reset  = ap_rst;
assign \lshr_32ns_32s_32_7_1_U9.din1_cast  = \lshr_32ns_32s_32_7_1_U9.din1 ;
assign \lshr_32ns_32s_32_7_1_U9.din1_mask  = 32'd31;
assign \lshr_32ns_32s_32_7_1_U9.ce  = 1'h1;
assign \lshr_32ns_32s_32_7_1_U9.clk  = ap_clk;
assign \lshr_32ns_32s_32_7_1_U9.din0  = { 31'h00000000, icmp_ln1498_reg_739 };
assign \lshr_32ns_32s_32_7_1_U9.din1  = { sub_ln1497_reg_745[2], sub_ln1497_reg_745[2], sub_ln1497_reg_745[2], sub_ln1497_reg_745[2], sub_ln1497_reg_745[2], sub_ln1497_reg_745[2], sub_ln1497_reg_745[2], sub_ln1497_reg_745[2], sub_ln1497_reg_745[2], sub_ln1497_reg_745[2], sub_ln1497_reg_745[2], sub_ln1497_reg_745[2], sub_ln1497_reg_745[2], sub_ln1497_reg_745[2], sub_ln1497_reg_745[2], sub_ln1497_reg_745[2], sub_ln1497_reg_745[2], sub_ln1497_reg_745[2], sub_ln1497_reg_745[2], sub_ln1497_reg_745[2], sub_ln1497_reg_745[2], sub_ln1497_reg_745[2], sub_ln1497_reg_745[2], sub_ln1497_reg_745[2], sub_ln1497_reg_745[2], sub_ln1497_reg_745[2], sub_ln1497_reg_745[2], sub_ln1497_reg_745[2], sub_ln1497_reg_745[2], sub_ln1497_reg_745 };
assign grp_fu_420_p2 = \lshr_32ns_32s_32_7_1_U9.dout ;
assign \lshr_32ns_32s_32_7_1_U9.reset  = ap_rst;
assign \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_3_U.ain_s0  = \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_3_U.a ;
assign \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_3_U.bin_s0  = \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_3_U.b ;
assign \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_3_U.s  = { \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_3_U.fas_s2 , \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_3_U.sum_s1  };
assign \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_3_U.u2.a  = \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_3_U.ain_s1 ;
assign \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_3_U.u2.b  = \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_3_U.bin_s1 ;
assign \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_3_U.u2.cin  = \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_3_U.carry_s1 ;
assign \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_3_U.facout_s2  = \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_3_U.u2.cout ;
assign \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_3_U.fas_s2  = \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_3_U.u2.s ;
assign \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_3_U.u1.a  = \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_3_U.a [1:0];
assign \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_3_U.u1.b  = \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_3_U.b [1:0];
assign \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_3_U.u1.cin  = 1'h0;
assign \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_3_U.facout_s1  = \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_3_U.u1.cout ;
assign \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_3_U.fas_s1  = \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_3_U.u1.s ;
assign \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_3_U.a  = \add_5s_5s_5_2_1_U4.din0 ;
assign \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_3_U.b  = \add_5s_5s_5_2_1_U4.din1 ;
assign \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_3_U.ce  = \add_5s_5s_5_2_1_U4.ce ;
assign \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_3_U.clk  = \add_5s_5s_5_2_1_U4.clk ;
assign \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_3_U.reset  = \add_5s_5s_5_2_1_U4.reset ;
assign \add_5s_5s_5_2_1_U4.dout  = \add_5s_5s_5_2_1_U4.top_add_5s_5s_5_2_1_Adder_3_U.s ;
assign \add_5s_5s_5_2_1_U4.ce  = 1'h1;
assign \add_5s_5s_5_2_1_U4.clk  = ap_clk;
assign \add_5s_5s_5_2_1_U4.din0  = { op_21_V_reg_660[2], op_21_V_reg_660, 1'h0 };
assign \add_5s_5s_5_2_1_U4.din1  = { op_10[1], op_10[1], op_10[1], op_10 };
assign grp_fu_273_p2 = \add_5s_5s_5_2_1_U4.dout ;
assign \add_5s_5s_5_2_1_U4.reset  = ap_rst;
assign \add_5s_5ns_5_2_1_U5.top_add_5s_5ns_5_2_1_Adder_4_U.ain_s0  = \add_5s_5ns_5_2_1_U5.top_add_5s_5ns_5_2_1_Adder_4_U.a ;
assign \add_5s_5ns_5_2_1_U5.top_add_5s_5ns_5_2_1_Adder_4_U.bin_s0  = \add_5s_5ns_5_2_1_U5.top_add_5s_5ns_5_2_1_Adder_4_U.b ;
assign \add_5s_5ns_5_2_1_U5.top_add_5s_5ns_5_2_1_Adder_4_U.s  = { \add_5s_5ns_5_2_1_U5.top_add_5s_5ns_5_2_1_Adder_4_U.fas_s2 , \add_5s_5ns_5_2_1_U5.top_add_5s_5ns_5_2_1_Adder_4_U.sum_s1  };
assign \add_5s_5ns_5_2_1_U5.top_add_5s_5ns_5_2_1_Adder_4_U.u2.a  = \add_5s_5ns_5_2_1_U5.top_add_5s_5ns_5_2_1_Adder_4_U.ain_s1 ;
assign \add_5s_5ns_5_2_1_U5.top_add_5s_5ns_5_2_1_Adder_4_U.u2.b  = \add_5s_5ns_5_2_1_U5.top_add_5s_5ns_5_2_1_Adder_4_U.bin_s1 ;
assign \add_5s_5ns_5_2_1_U5.top_add_5s_5ns_5_2_1_Adder_4_U.u2.cin  = \add_5s_5ns_5_2_1_U5.top_add_5s_5ns_5_2_1_Adder_4_U.carry_s1 ;
assign \add_5s_5ns_5_2_1_U5.top_add_5s_5ns_5_2_1_Adder_4_U.facout_s2  = \add_5s_5ns_5_2_1_U5.top_add_5s_5ns_5_2_1_Adder_4_U.u2.cout ;
assign \add_5s_5ns_5_2_1_U5.top_add_5s_5ns_5_2_1_Adder_4_U.fas_s2  = \add_5s_5ns_5_2_1_U5.top_add_5s_5ns_5_2_1_Adder_4_U.u2.s ;
assign \add_5s_5ns_5_2_1_U5.top_add_5s_5ns_5_2_1_Adder_4_U.u1.a  = \add_5s_5ns_5_2_1_U5.top_add_5s_5ns_5_2_1_Adder_4_U.a [1:0];
assign \add_5s_5ns_5_2_1_U5.top_add_5s_5ns_5_2_1_Adder_4_U.u1.b  = \add_5s_5ns_5_2_1_U5.top_add_5s_5ns_5_2_1_Adder_4_U.b [1:0];
assign \add_5s_5ns_5_2_1_U5.top_add_5s_5ns_5_2_1_Adder_4_U.u1.cin  = 1'h0;
assign \add_5s_5ns_5_2_1_U5.top_add_5s_5ns_5_2_1_Adder_4_U.facout_s1  = \add_5s_5ns_5_2_1_U5.top_add_5s_5ns_5_2_1_Adder_4_U.u1.cout ;
assign \add_5s_5ns_5_2_1_U5.top_add_5s_5ns_5_2_1_Adder_4_U.fas_s1  = \add_5s_5ns_5_2_1_U5.top_add_5s_5ns_5_2_1_Adder_4_U.u1.s ;
assign \add_5s_5ns_5_2_1_U5.top_add_5s_5ns_5_2_1_Adder_4_U.a  = \add_5s_5ns_5_2_1_U5.din0 ;
assign \add_5s_5ns_5_2_1_U5.top_add_5s_5ns_5_2_1_Adder_4_U.b  = \add_5s_5ns_5_2_1_U5.din1 ;
assign \add_5s_5ns_5_2_1_U5.top_add_5s_5ns_5_2_1_Adder_4_U.ce  = \add_5s_5ns_5_2_1_U5.ce ;
assign \add_5s_5ns_5_2_1_U5.top_add_5s_5ns_5_2_1_Adder_4_U.clk  = \add_5s_5ns_5_2_1_U5.clk ;
assign \add_5s_5ns_5_2_1_U5.top_add_5s_5ns_5_2_1_Adder_4_U.reset  = \add_5s_5ns_5_2_1_U5.reset ;
assign \add_5s_5ns_5_2_1_U5.dout  = \add_5s_5ns_5_2_1_U5.top_add_5s_5ns_5_2_1_Adder_4_U.s ;
assign \add_5s_5ns_5_2_1_U5.ce  = 1'h1;
assign \add_5s_5ns_5_2_1_U5.clk  = ap_clk;
assign \add_5s_5ns_5_2_1_U5.din0  = { tmp_2_reg_685[3], tmp_2_reg_685 };
assign \add_5s_5ns_5_2_1_U5.din1  = 5'h01;
assign grp_fu_292_p2 = \add_5s_5ns_5_2_1_U5.dout ;
assign \add_5s_5ns_5_2_1_U5.reset  = ap_rst;
assign \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.ain_s0  = \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.a ;
assign \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.bin_s0  = \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.b ;
assign \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.s  = { \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.fas_s2 , \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.sum_s1  };
assign \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.u2.a  = \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.ain_s1 ;
assign \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.u2.b  = \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.bin_s1 ;
assign \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.u2.cin  = \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.carry_s1 ;
assign \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.facout_s2  = \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.u2.cout ;
assign \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.fas_s2  = \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.u2.s ;
assign \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.u1.a  = \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.a [1:0];
assign \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.u1.b  = \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.b [1:0];
assign \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.u1.cin  = 1'h0;
assign \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.facout_s1  = \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.u1.cout ;
assign \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.fas_s1  = \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.u1.s ;
assign \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.a  = \add_5ns_5s_5_2_1_U1.din0 ;
assign \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.b  = \add_5ns_5s_5_2_1_U1.din1 ;
assign \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.ce  = \add_5ns_5s_5_2_1_U1.ce ;
assign \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.clk  = \add_5ns_5s_5_2_1_U1.clk ;
assign \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.reset  = \add_5ns_5s_5_2_1_U1.reset ;
assign \add_5ns_5s_5_2_1_U1.dout  = \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.s ;
assign \add_5ns_5s_5_2_1_U1.ce  = 1'h1;
assign \add_5ns_5s_5_2_1_U1.clk  = ap_clk;
assign \add_5ns_5s_5_2_1_U1.din0  = { 1'h0, op_8, 3'h0 };
assign \add_5ns_5s_5_2_1_U1.din1  = { op_0[3], op_0 };
assign grp_fu_199_p2 = \add_5ns_5s_5_2_1_U1.dout ;
assign \add_5ns_5s_5_2_1_U1.reset  = ap_rst;
assign \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_6_U.ain_s0  = \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_6_U.a ;
assign \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_6_U.bin_s0  = \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_6_U.b ;
assign \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_6_U.s  = { \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_6_U.fas_s2 , \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_6_U.sum_s1  };
assign \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_6_U.u2.a  = \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_6_U.ain_s1 ;
assign \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_6_U.u2.b  = \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_6_U.bin_s1 ;
assign \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_6_U.u2.cin  = \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_6_U.carry_s1 ;
assign \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_6_U.facout_s2  = \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_6_U.u2.cout ;
assign \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_6_U.fas_s2  = \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_6_U.u2.s ;
assign \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_6_U.u1.a  = \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_6_U.a [1:0];
assign \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_6_U.u1.b  = \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_6_U.b [1:0];
assign \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_6_U.u1.cin  = 1'h0;
assign \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_6_U.facout_s1  = \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_6_U.u1.cout ;
assign \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_6_U.fas_s1  = \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_6_U.u1.s ;
assign \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_6_U.a  = \add_5ns_5ns_5_2_1_U7.din0 ;
assign \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_6_U.b  = \add_5ns_5ns_5_2_1_U7.din1 ;
assign \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_6_U.ce  = \add_5ns_5ns_5_2_1_U7.ce ;
assign \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_6_U.clk  = \add_5ns_5ns_5_2_1_U7.clk ;
assign \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_6_U.reset  = \add_5ns_5ns_5_2_1_U7.reset ;
assign \add_5ns_5ns_5_2_1_U7.dout  = \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_6_U.s ;
assign \add_5ns_5ns_5_2_1_U7.ce  = 1'h1;
assign \add_5ns_5ns_5_2_1_U7.clk  = ap_clk;
assign \add_5ns_5ns_5_2_1_U7.din0  = ret_V_15_reg_734;
assign \add_5ns_5ns_5_2_1_U7.din1  = { 4'h0, icmp_ln1498_1_reg_729 };
assign grp_fu_386_p2 = \add_5ns_5ns_5_2_1_U7.dout ;
assign \add_5ns_5ns_5_2_1_U7.reset  = ap_rst;
assign \add_3s_3ns_3_2_1_U2.top_add_3s_3ns_3_2_1_Adder_1_U.ain_s0  = \add_3s_3ns_3_2_1_U2.top_add_3s_3ns_3_2_1_Adder_1_U.a ;
assign \add_3s_3ns_3_2_1_U2.top_add_3s_3ns_3_2_1_Adder_1_U.bin_s0  = \add_3s_3ns_3_2_1_U2.top_add_3s_3ns_3_2_1_Adder_1_U.b ;
assign \add_3s_3ns_3_2_1_U2.top_add_3s_3ns_3_2_1_Adder_1_U.s  = { \add_3s_3ns_3_2_1_U2.top_add_3s_3ns_3_2_1_Adder_1_U.fas_s2 , \add_3s_3ns_3_2_1_U2.top_add_3s_3ns_3_2_1_Adder_1_U.sum_s1  };
assign \add_3s_3ns_3_2_1_U2.top_add_3s_3ns_3_2_1_Adder_1_U.u2.a  = \add_3s_3ns_3_2_1_U2.top_add_3s_3ns_3_2_1_Adder_1_U.ain_s1 ;
assign \add_3s_3ns_3_2_1_U2.top_add_3s_3ns_3_2_1_Adder_1_U.u2.b  = \add_3s_3ns_3_2_1_U2.top_add_3s_3ns_3_2_1_Adder_1_U.bin_s1 ;
assign \add_3s_3ns_3_2_1_U2.top_add_3s_3ns_3_2_1_Adder_1_U.u2.cin  = \add_3s_3ns_3_2_1_U2.top_add_3s_3ns_3_2_1_Adder_1_U.carry_s1 ;
assign \add_3s_3ns_3_2_1_U2.top_add_3s_3ns_3_2_1_Adder_1_U.facout_s2  = \add_3s_3ns_3_2_1_U2.top_add_3s_3ns_3_2_1_Adder_1_U.u2.cout ;
assign \add_3s_3ns_3_2_1_U2.top_add_3s_3ns_3_2_1_Adder_1_U.fas_s2  = \add_3s_3ns_3_2_1_U2.top_add_3s_3ns_3_2_1_Adder_1_U.u2.s ;
assign \add_3s_3ns_3_2_1_U2.top_add_3s_3ns_3_2_1_Adder_1_U.u1.a  = \add_3s_3ns_3_2_1_U2.top_add_3s_3ns_3_2_1_Adder_1_U.a [0];
assign \add_3s_3ns_3_2_1_U2.top_add_3s_3ns_3_2_1_Adder_1_U.u1.b  = \add_3s_3ns_3_2_1_U2.top_add_3s_3ns_3_2_1_Adder_1_U.b [0];
assign \add_3s_3ns_3_2_1_U2.top_add_3s_3ns_3_2_1_Adder_1_U.u1.cin  = 1'h0;
assign \add_3s_3ns_3_2_1_U2.top_add_3s_3ns_3_2_1_Adder_1_U.facout_s1  = \add_3s_3ns_3_2_1_U2.top_add_3s_3ns_3_2_1_Adder_1_U.u1.cout ;
assign \add_3s_3ns_3_2_1_U2.top_add_3s_3ns_3_2_1_Adder_1_U.fas_s1  = \add_3s_3ns_3_2_1_U2.top_add_3s_3ns_3_2_1_Adder_1_U.u1.s ;
assign \add_3s_3ns_3_2_1_U2.top_add_3s_3ns_3_2_1_Adder_1_U.a  = \add_3s_3ns_3_2_1_U2.din0 ;
assign \add_3s_3ns_3_2_1_U2.top_add_3s_3ns_3_2_1_Adder_1_U.b  = \add_3s_3ns_3_2_1_U2.din1 ;
assign \add_3s_3ns_3_2_1_U2.top_add_3s_3ns_3_2_1_Adder_1_U.ce  = \add_3s_3ns_3_2_1_U2.ce ;
assign \add_3s_3ns_3_2_1_U2.top_add_3s_3ns_3_2_1_Adder_1_U.clk  = \add_3s_3ns_3_2_1_U2.clk ;
assign \add_3s_3ns_3_2_1_U2.top_add_3s_3ns_3_2_1_Adder_1_U.reset  = \add_3s_3ns_3_2_1_U2.reset ;
assign \add_3s_3ns_3_2_1_U2.dout  = \add_3s_3ns_3_2_1_U2.top_add_3s_3ns_3_2_1_Adder_1_U.s ;
assign \add_3s_3ns_3_2_1_U2.ce  = 1'h1;
assign \add_3s_3ns_3_2_1_U2.clk  = ap_clk;
assign \add_3s_3ns_3_2_1_U2.din0  = { ret_V_reg_638[1], ret_V_reg_638 };
assign \add_3s_3ns_3_2_1_U2.din1  = 3'h1;
assign grp_fu_228_p2 = \add_3s_3ns_3_2_1_U2.dout ;
assign \add_3s_3ns_3_2_1_U2.reset  = ap_rst;
assign \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_2_U.ain_s0  = \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_2_U.a ;
assign \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_2_U.bin_s0  = \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_2_U.b ;
assign \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_2_U.s  = { \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_2_U.fas_s2 , \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_2_U.sum_s1  };
assign \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_2_U.u2.a  = \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_2_U.ain_s1 ;
assign \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_2_U.u2.b  = \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_2_U.bin_s1 ;
assign \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_2_U.u2.cin  = \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_2_U.carry_s1 ;
assign \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_2_U.facout_s2  = \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_2_U.u2.cout ;
assign \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_2_U.fas_s2  = \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_2_U.u2.s ;
assign \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_2_U.u1.a  = \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_2_U.a [0];
assign \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_2_U.u1.b  = \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_2_U.b [0];
assign \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_2_U.u1.cin  = 1'h0;
assign \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_2_U.facout_s1  = \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_2_U.u1.cout ;
assign \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_2_U.fas_s1  = \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_2_U.u1.s ;
assign \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_2_U.a  = \add_3ns_3ns_3_2_1_U3.din0 ;
assign \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_2_U.b  = \add_3ns_3ns_3_2_1_U3.din1 ;
assign \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_2_U.ce  = \add_3ns_3ns_3_2_1_U3.ce ;
assign \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_2_U.clk  = \add_3ns_3ns_3_2_1_U3.clk ;
assign \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_2_U.reset  = \add_3ns_3ns_3_2_1_U3.reset ;
assign \add_3ns_3ns_3_2_1_U3.dout  = \add_3ns_3ns_3_2_1_U3.top_add_3ns_3ns_3_2_1_Adder_2_U.s ;
assign \add_3ns_3ns_3_2_1_U3.ce  = 1'h1;
assign \add_3ns_3ns_3_2_1_U3.clk  = ap_clk;
assign \add_3ns_3ns_3_2_1_U3.din0  = ret_V_13_reg_655;
assign \add_3ns_3ns_3_2_1_U3.din1  = 3'h1;
assign grp_fu_253_p2 = \add_3ns_3ns_3_2_1_U3.dout ;
assign \add_3ns_3ns_3_2_1_U3.reset  = ap_rst;
assign \add_35s_35s_35_2_1_U13.top_add_35s_35s_35_2_1_Adder_10_U.ain_s0  = \add_35s_35s_35_2_1_U13.top_add_35s_35s_35_2_1_Adder_10_U.a ;
assign \add_35s_35s_35_2_1_U13.top_add_35s_35s_35_2_1_Adder_10_U.bin_s0  = \add_35s_35s_35_2_1_U13.top_add_35s_35s_35_2_1_Adder_10_U.b ;
assign \add_35s_35s_35_2_1_U13.top_add_35s_35s_35_2_1_Adder_10_U.s  = { \add_35s_35s_35_2_1_U13.top_add_35s_35s_35_2_1_Adder_10_U.fas_s2 , \add_35s_35s_35_2_1_U13.top_add_35s_35s_35_2_1_Adder_10_U.sum_s1  };
assign \add_35s_35s_35_2_1_U13.top_add_35s_35s_35_2_1_Adder_10_U.u2.a  = \add_35s_35s_35_2_1_U13.top_add_35s_35s_35_2_1_Adder_10_U.ain_s1 ;
assign \add_35s_35s_35_2_1_U13.top_add_35s_35s_35_2_1_Adder_10_U.u2.b  = \add_35s_35s_35_2_1_U13.top_add_35s_35s_35_2_1_Adder_10_U.bin_s1 ;
assign \add_35s_35s_35_2_1_U13.top_add_35s_35s_35_2_1_Adder_10_U.u2.cin  = \add_35s_35s_35_2_1_U13.top_add_35s_35s_35_2_1_Adder_10_U.carry_s1 ;
assign \add_35s_35s_35_2_1_U13.top_add_35s_35s_35_2_1_Adder_10_U.facout_s2  = \add_35s_35s_35_2_1_U13.top_add_35s_35s_35_2_1_Adder_10_U.u2.cout ;
assign \add_35s_35s_35_2_1_U13.top_add_35s_35s_35_2_1_Adder_10_U.fas_s2  = \add_35s_35s_35_2_1_U13.top_add_35s_35s_35_2_1_Adder_10_U.u2.s ;
assign \add_35s_35s_35_2_1_U13.top_add_35s_35s_35_2_1_Adder_10_U.u1.a  = \add_35s_35s_35_2_1_U13.top_add_35s_35s_35_2_1_Adder_10_U.a [16:0];
assign \add_35s_35s_35_2_1_U13.top_add_35s_35s_35_2_1_Adder_10_U.u1.b  = \add_35s_35s_35_2_1_U13.top_add_35s_35s_35_2_1_Adder_10_U.b [16:0];
assign \add_35s_35s_35_2_1_U13.top_add_35s_35s_35_2_1_Adder_10_U.u1.cin  = 1'h0;
assign \add_35s_35s_35_2_1_U13.top_add_35s_35s_35_2_1_Adder_10_U.facout_s1  = \add_35s_35s_35_2_1_U13.top_add_35s_35s_35_2_1_Adder_10_U.u1.cout ;
assign \add_35s_35s_35_2_1_U13.top_add_35s_35s_35_2_1_Adder_10_U.fas_s1  = \add_35s_35s_35_2_1_U13.top_add_35s_35s_35_2_1_Adder_10_U.u1.s ;
assign \add_35s_35s_35_2_1_U13.top_add_35s_35s_35_2_1_Adder_10_U.a  = \add_35s_35s_35_2_1_U13.din0 ;
assign \add_35s_35s_35_2_1_U13.top_add_35s_35s_35_2_1_Adder_10_U.b  = \add_35s_35s_35_2_1_U13.din1 ;
assign \add_35s_35s_35_2_1_U13.top_add_35s_35s_35_2_1_Adder_10_U.ce  = \add_35s_35s_35_2_1_U13.ce ;
assign \add_35s_35s_35_2_1_U13.top_add_35s_35s_35_2_1_Adder_10_U.clk  = \add_35s_35s_35_2_1_U13.clk ;
assign \add_35s_35s_35_2_1_U13.top_add_35s_35s_35_2_1_Adder_10_U.reset  = \add_35s_35s_35_2_1_U13.reset ;
assign \add_35s_35s_35_2_1_U13.dout  = \add_35s_35s_35_2_1_U13.top_add_35s_35s_35_2_1_Adder_10_U.s ;
assign \add_35s_35s_35_2_1_U13.ce  = 1'h1;
assign \add_35s_35s_35_2_1_U13.clk  = ap_clk;
assign \add_35s_35s_35_2_1_U13.din0  = { op_25_V_reg_838[31], op_25_V_reg_838, 2'h0 };
assign \add_35s_35s_35_2_1_U13.din1  = { op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16 };
assign grp_fu_532_p2 = \add_35s_35s_35_2_1_U13.dout ;
assign \add_35s_35s_35_2_1_U13.reset  = ap_rst;
assign \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_7_U.ain_s0  = \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_7_U.a ;
assign \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_7_U.bin_s0  = \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_7_U.b ;
assign \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_7_U.s  = { \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_7_U.fas_s2 , \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_7_U.sum_s1  };
assign \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_7_U.u2.a  = \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_7_U.ain_s1 ;
assign \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_7_U.u2.b  = \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_7_U.bin_s1 ;
assign \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_7_U.u2.cin  = \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_7_U.carry_s1 ;
assign \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_7_U.facout_s2  = \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_7_U.u2.cout ;
assign \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_7_U.fas_s2  = \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_7_U.u2.s ;
assign \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_7_U.u1.a  = \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_7_U.a [16:0];
assign \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_7_U.u1.b  = \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_7_U.b [16:0];
assign \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_7_U.u1.cin  = 1'h0;
assign \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_7_U.facout_s1  = \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_7_U.u1.cout ;
assign \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_7_U.fas_s1  = \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_7_U.u1.s ;
assign \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_7_U.a  = \add_34s_34s_34_2_1_U10.din0 ;
assign \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_7_U.b  = \add_34s_34s_34_2_1_U10.din1 ;
assign \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_7_U.ce  = \add_34s_34s_34_2_1_U10.ce ;
assign \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_7_U.clk  = \add_34s_34s_34_2_1_U10.clk ;
assign \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_7_U.reset  = \add_34s_34s_34_2_1_U10.reset ;
assign \add_34s_34s_34_2_1_U10.dout  = \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_7_U.s ;
assign \add_34s_34s_34_2_1_U10.ce  = 1'h1;
assign \add_34s_34s_34_2_1_U10.clk  = ap_clk;
assign \add_34s_34s_34_2_1_U10.din0  = { op_23_V_reg_776[4], op_23_V_reg_776[4], op_23_V_reg_776[4], op_23_V_reg_776[4], op_23_V_reg_776[4], op_23_V_reg_776[4], op_23_V_reg_776[4], op_23_V_reg_776[4], op_23_V_reg_776[4], op_23_V_reg_776[4], op_23_V_reg_776[4], op_23_V_reg_776[4], op_23_V_reg_776[4], op_23_V_reg_776[4], op_23_V_reg_776[4], op_23_V_reg_776[4], op_23_V_reg_776[4], op_23_V_reg_776[4], op_23_V_reg_776[4], op_23_V_reg_776[4], op_23_V_reg_776[4], op_23_V_reg_776[4], op_23_V_reg_776[4], op_23_V_reg_776[4], op_23_V_reg_776[4], op_23_V_reg_776[4], op_23_V_reg_776[4], op_23_V_reg_776[4], op_23_V_reg_776, 1'h0 };
assign \add_34s_34s_34_2_1_U10.din1  = { op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14 };
assign grp_fu_447_p2 = \add_34s_34s_34_2_1_U10.dout ;
assign \add_34s_34s_34_2_1_U10.reset  = ap_rst;
assign \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_9_U.ain_s0  = \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_9_U.a ;
assign \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_9_U.bin_s0  = \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_9_U.b ;
assign \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_9_U.s  = { \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_9_U.fas_s2 , \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_9_U.sum_s1  };
assign \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_9_U.u2.a  = \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_9_U.ain_s1 ;
assign \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_9_U.u2.b  = \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_9_U.bin_s1 ;
assign \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_9_U.u2.cin  = \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_9_U.carry_s1 ;
assign \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_9_U.facout_s2  = \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_9_U.u2.cout ;
assign \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_9_U.fas_s2  = \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_9_U.u2.s ;
assign \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_9_U.u1.a  = \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_9_U.a [15:0];
assign \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_9_U.u1.b  = \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_9_U.b [15:0];
assign \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_9_U.u1.cin  = 1'h0;
assign \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_9_U.facout_s1  = \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_9_U.u1.cout ;
assign \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_9_U.fas_s1  = \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_9_U.u1.s ;
assign \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_9_U.a  = \add_32ns_32s_32_2_1_U12.din0 ;
assign \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_9_U.b  = \add_32ns_32s_32_2_1_U12.din1 ;
assign \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_9_U.ce  = \add_32ns_32s_32_2_1_U12.ce ;
assign \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_9_U.clk  = \add_32ns_32s_32_2_1_U12.clk ;
assign \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_9_U.reset  = \add_32ns_32s_32_2_1_U12.reset ;
assign \add_32ns_32s_32_2_1_U12.dout  = \add_32ns_32s_32_2_1_U12.top_add_32ns_32s_32_2_1_Adder_9_U.s ;
assign \add_32ns_32s_32_2_1_U12.ce  = 1'h1;
assign \add_32ns_32s_32_2_1_U12.clk  = ap_clk;
assign \add_32ns_32s_32_2_1_U12.din0  = ret_V_17_reg_813;
assign \add_32ns_32s_32_2_1_U12.din1  = { op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15 };
assign grp_fu_503_p2 = \add_32ns_32s_32_2_1_U12.dout ;
assign \add_32ns_32s_32_2_1_U12.reset  = ap_rst;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.ain_s0  = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.a ;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.bin_s0  = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.b ;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.s  = { \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.fas_s2 , \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.sum_s1  };
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.u2.a  = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.ain_s1 ;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.u2.b  = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.bin_s1 ;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.u2.cin  = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.carry_s1 ;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.facout_s2  = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.u2.cout ;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.fas_s2  = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.u2.s ;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.u1.a  = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.a [15:0];
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.u1.b  = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.b [15:0];
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.u1.cin  = 1'h0;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.facout_s1  = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.u1.cout ;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.fas_s1  = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.u1.s ;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.a  = \add_32ns_32ns_32_2_1_U17.din0 ;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.b  = \add_32ns_32ns_32_2_1_U17.din1 ;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.ce  = \add_32ns_32ns_32_2_1_U17.ce ;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.clk  = \add_32ns_32ns_32_2_1_U17.clk ;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.reset  = \add_32ns_32ns_32_2_1_U17.reset ;
assign \add_32ns_32ns_32_2_1_U17.dout  = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.s ;
assign \add_32ns_32ns_32_2_1_U17.ce  = 1'h1;
assign \add_32ns_32ns_32_2_1_U17.clk  = ap_clk;
assign \add_32ns_32ns_32_2_1_U17.din0  = { 30'h00000000, add_ln69_1_reg_875 };
assign \add_32ns_32ns_32_2_1_U17.din1  = add_ln69_reg_900;
assign grp_fu_612_p2 = \add_32ns_32ns_32_2_1_U17.dout ;
assign \add_32ns_32ns_32_2_1_U17.reset  = ap_rst;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_8_U.ain_s0  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_8_U.a ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_8_U.bin_s0  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_8_U.b ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_8_U.s  = { \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_8_U.fas_s2 , \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_8_U.sum_s1  };
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_8_U.u2.a  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_8_U.ain_s1 ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_8_U.u2.b  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_8_U.bin_s1 ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_8_U.u2.cin  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_8_U.carry_s1 ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_8_U.facout_s2  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_8_U.u2.cout ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_8_U.fas_s2  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_8_U.u2.s ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_8_U.u1.a  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_8_U.a [15:0];
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_8_U.u1.b  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_8_U.b [15:0];
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_8_U.u1.cin  = 1'h0;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_8_U.facout_s1  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_8_U.u1.cout ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_8_U.fas_s1  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_8_U.u1.s ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_8_U.a  = \add_32ns_32ns_32_2_1_U16.din0 ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_8_U.b  = \add_32ns_32ns_32_2_1_U16.din1 ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_8_U.ce  = \add_32ns_32ns_32_2_1_U16.ce ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_8_U.clk  = \add_32ns_32ns_32_2_1_U16.clk ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_8_U.reset  = \add_32ns_32ns_32_2_1_U16.reset ;
assign \add_32ns_32ns_32_2_1_U16.dout  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_8_U.s ;
assign \add_32ns_32ns_32_2_1_U16.ce  = 1'h1;
assign \add_32ns_32ns_32_2_1_U16.clk  = ap_clk;
assign \add_32ns_32ns_32_2_1_U16.din0  = ret_V_19_reg_890;
assign \add_32ns_32ns_32_2_1_U16.din1  = { 28'h0000000, ret_V_11_reg_885[1], ret_V_11_reg_885[1], ret_V_11_reg_885 };
assign grp_fu_604_p2 = \add_32ns_32ns_32_2_1_U16.dout ;
assign \add_32ns_32ns_32_2_1_U16.reset  = ap_rst;
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_8_U.ain_s0  = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_8_U.a ;
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_8_U.bin_s0  = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_8_U.b ;
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_8_U.s  = { \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_8_U.fas_s2 , \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_8_U.sum_s1  };
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_8_U.u2.a  = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_8_U.ain_s1 ;
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_8_U.u2.b  = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_8_U.bin_s1 ;
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_8_U.u2.cin  = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_8_U.carry_s1 ;
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_8_U.facout_s2  = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_8_U.u2.cout ;
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_8_U.fas_s2  = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_8_U.u2.s ;
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_8_U.u1.a  = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_8_U.a [15:0];
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_8_U.u1.b  = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_8_U.b [15:0];
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_8_U.u1.cin  = 1'h0;
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_8_U.facout_s1  = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_8_U.u1.cout ;
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_8_U.fas_s1  = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_8_U.u1.s ;
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_8_U.a  = \add_32ns_32ns_32_2_1_U15.din0 ;
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_8_U.b  = \add_32ns_32ns_32_2_1_U15.din1 ;
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_8_U.ce  = \add_32ns_32ns_32_2_1_U15.ce ;
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_8_U.clk  = \add_32ns_32ns_32_2_1_U15.clk ;
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_8_U.reset  = \add_32ns_32ns_32_2_1_U15.reset ;
assign \add_32ns_32ns_32_2_1_U15.dout  = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_8_U.s ;
assign \add_32ns_32ns_32_2_1_U15.ce  = 1'h1;
assign \add_32ns_32ns_32_2_1_U15.clk  = ap_clk;
assign \add_32ns_32ns_32_2_1_U15.din0  = ret_V_15_cast_reg_868;
assign \add_32ns_32ns_32_2_1_U15.din1  = 32'd1;
assign grp_fu_566_p2 = \add_32ns_32ns_32_2_1_U15.dout ;
assign \add_32ns_32ns_32_2_1_U15.reset  = ap_rst;
assign \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.ain_s0  = \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.a ;
assign \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.bin_s0  = \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.b ;
assign \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.s  = { \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.fas_s2 , \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.sum_s1  };
assign \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.u2.a  = \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.ain_s1 ;
assign \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.u2.b  = \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.bin_s1 ;
assign \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.u2.cin  = \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.carry_s1 ;
assign \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.facout_s2  = \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.u2.cout ;
assign \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.fas_s2  = \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.u2.s ;
assign \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.u1.a  = \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.a [15:0];
assign \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.u1.b  = \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.b [15:0];
assign \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.u1.cin  = 1'h0;
assign \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.facout_s1  = \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.u1.cout ;
assign \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.fas_s1  = \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.u1.s ;
assign \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.a  = \add_32ns_32ns_32_2_1_U11.din0 ;
assign \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.b  = \add_32ns_32ns_32_2_1_U11.din1 ;
assign \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.ce  = \add_32ns_32ns_32_2_1_U11.ce ;
assign \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.clk  = \add_32ns_32ns_32_2_1_U11.clk ;
assign \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.reset  = \add_32ns_32ns_32_2_1_U11.reset ;
assign \add_32ns_32ns_32_2_1_U11.dout  = \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.s ;
assign \add_32ns_32ns_32_2_1_U11.ce  = 1'h1;
assign \add_32ns_32ns_32_2_1_U11.clk  = ap_clk;
assign \add_32ns_32ns_32_2_1_U11.din0  = ret_V_7_cast_reg_801;
assign \add_32ns_32ns_32_2_1_U11.din1  = 32'd1;
assign grp_fu_463_p2 = \add_32ns_32ns_32_2_1_U11.dout ;
assign \add_32ns_32ns_32_2_1_U11.reset  = ap_rst;
assign \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_11_U.ain_s0  = \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_11_U.a ;
assign \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_11_U.bin_s0  = \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_11_U.b ;
assign \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_11_U.s  = { \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_11_U.fas_s2 , \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_11_U.sum_s1  };
assign \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_11_U.u2.a  = \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_11_U.ain_s1 ;
assign \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_11_U.u2.b  = \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_11_U.bin_s1 ;
assign \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_11_U.u2.cin  = \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_11_U.carry_s1 ;
assign \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_11_U.facout_s2  = \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_11_U.u2.cout ;
assign \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_11_U.fas_s2  = \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_11_U.u2.s ;
assign \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_11_U.u1.a  = \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_11_U.a [0];
assign \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_11_U.u1.b  = \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_11_U.b [0];
assign \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_11_U.u1.cin  = 1'h0;
assign \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_11_U.facout_s1  = \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_11_U.u1.cout ;
assign \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_11_U.fas_s1  = \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_11_U.u1.s ;
assign \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_11_U.a  = \add_2ns_2ns_2_2_1_U14.din0 ;
assign \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_11_U.b  = \add_2ns_2ns_2_2_1_U14.din1 ;
assign \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_11_U.ce  = \add_2ns_2ns_2_2_1_U14.ce ;
assign \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_11_U.clk  = \add_2ns_2ns_2_2_1_U14.clk ;
assign \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_11_U.reset  = \add_2ns_2ns_2_2_1_U14.reset ;
assign \add_2ns_2ns_2_2_1_U14.dout  = \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_11_U.s ;
assign \add_2ns_2ns_2_2_1_U14.ce  = 1'h1;
assign \add_2ns_2ns_2_2_1_U14.clk  = ap_clk;
assign \add_2ns_2ns_2_2_1_U14.din0  = op_17_V_reg_833;
assign \add_2ns_2ns_2_2_1_U14.din1  = { 1'h0, icmp_ln1495_reg_771 };
assign grp_fu_551_p2 = \add_2ns_2ns_2_2_1_U14.dout ;
assign \add_2ns_2ns_2_2_1_U14.reset  = ap_rst;
endmodule


// Machine B:
// Processed by function `add_clk_enable_signal` in `verilog_tricks.py`.
// Processed by function `remove_reset_signal` in `verilog_tricks.py`.
module top_B (
  ap_clk,
  ap_start,
  ap_done,
  ap_idle,
  ap_ready,
  op_0,
  op_1,
  op_2,
  op_3,
  op_4,
  op_7,
  op_8,
  op_10,
  op_14,
  op_15,
  op_16,
  op_29,
  op_29_ap_vld,
clk_enable
);
input clk_enable;


input ap_clk;
wire ap_rst;
assign ap_rst = op_29_ap_vld;
input ap_start;
input [3:0] op_0;
input [7:0] op_1;
input [1:0] op_10;
input [7:0] op_14;
input [3:0] op_15;
input [7:0] op_16;
input [1:0] op_2;
input op_3;
input [31:0] op_4;
input [1:0] op_7;
input op_8;
output ap_done;
output ap_idle;
output ap_ready;
output [31:0] op_29;
output op_29_ap_vld;


reg [31:0] add_ln691_1_reg_709;
reg [1:0] add_ln69_1_reg_761;
reg [8:0] ap_CS_fsm = 9'h001;
reg icmp_ln1495_reg_729;
reg icmp_ln1498_reg_719;
reg icmp_ln851_1_reg_746;
reg icmp_ln851_reg_643;
reg [4:0] op_23_V_reg_687;
reg [31:0] op_25_V_reg_714;
reg op_6_V_reg_664;
reg [1:0] ret_V_11_reg_751;
reg [4:0] ret_V_12_reg_632;
reg [4:0] ret_V_14_reg_669;
reg [31:0] ret_V_15_cast_reg_739;
reg [33:0] ret_V_16_reg_697;
reg [34:0] ret_V_18_reg_734;
reg [31:0] ret_V_19_reg_756;
reg [2:0] ret_V_3_reg_648;
reg [31:0] ret_V_7_cast_reg_702;
reg [2:0] sext_ln835_reg_637;
reg [2:0] sub_ln1497_reg_724;
reg [3:0] tmp_2_reg_674;
wire [31:0] _000_;
wire [1:0] _001_;
wire [8:0] _002_;
wire _003_;
wire _004_;
wire _005_;
wire _006_;
wire [4:0] _007_;
wire [31:0] _008_;
wire _009_;
wire [1:0] _010_;
wire [4:0] _011_;
wire [4:0] _012_;
wire [31:0] _013_;
wire [33:0] _014_;
wire [34:0] _015_;
wire [31:0] _016_;
wire [2:0] _017_;
wire [31:0] _018_;
wire [2:0] _019_;
wire [2:0] _020_;
wire [3:0] _021_;
wire [1:0] _022_;
wire _023_;
wire _024_;
wire _025_;
wire _026_;
wire _027_;
wire _028_;
wire _029_;
wire _030_;
wire _031_;
wire _032_;
wire _033_;
wire _034_;
wire _035_;
wire _036_;
wire _037_;
wire _038_;
wire _039_;
wire _040_;
wire [31:0] add_ln691_1_fu_395_p2;
wire [31:0] add_ln691_2_fu_583_p2;
wire [4:0] add_ln691_fu_332_p2;
wire [1:0] add_ln69_1_fu_604_p2;
wire [31:0] add_ln69_fu_617_p2;
wire ap_CS_fsm_state1;
wire ap_CS_fsm_state2;
wire ap_CS_fsm_state3;
wire ap_CS_fsm_state4;
wire ap_CS_fsm_state5;
wire ap_CS_fsm_state6;
wire ap_CS_fsm_state7;
wire ap_CS_fsm_state8;
wire ap_CS_fsm_state9;
wire [8:0] ap_NS_fsm;
wire ap_clk;
wire ap_done;
wire ap_idle;
wire ap_ready;
wire ap_rst;
wire ap_start;
wire [31:0] conv_i270_fu_538_p1;
wire icmp_ln1495_fu_474_p2;
wire [1:0] icmp_ln1498_1_fu_313_p1;
wire icmp_ln1498_1_fu_313_p2;
wire icmp_ln1498_fu_444_p2;
wire icmp_ln851_1_fu_515_p2;
wire icmp_ln851_fu_223_p2;
wire [31:0] lshr_ln1497_fu_554_p2;
wire [3:0] op_0;
wire [7:0] op_1;
wire [1:0] op_10;
wire [7:0] op_14;
wire [3:0] op_15;
wire [7:0] op_16;
wire [1:0] op_17_V_fu_568_p3;
wire [1:0] op_2;
wire [2:0] op_21_V_fu_268_p2;
wire [4:0] op_23_V_fu_358_p2;
wire [31:0] op_25_V_fu_427_p2;
wire [31:0] op_29;
wire op_29_ap_vld;
wire op_3;
wire [31:0] op_4;
wire op_6_V_fu_243_p2;
wire [1:0] op_7;
wire op_8;
wire p_Result_1_fu_322_p3;
wire p_Result_2_fu_400_p3;
wire p_Result_3_fu_576_p3;
wire p_Result_s_fu_249_p3;
wire [1:0] ret_V_11_fu_521_p1;
wire [1:0] ret_V_11_fu_521_p3;
wire [4:0] ret_V_12_fu_199_p2;
wire [2:0] ret_V_13_fu_261_p3;
wire [4:0] ret_V_14_fu_290_p2;
wire [4:0] ret_V_15_fu_346_p3;
wire [33:0] ret_V_16_fu_379_p2;
wire [31:0] ret_V_17_fu_416_p3;
wire [34:0] ret_V_18_fu_495_p2;
wire [31:0] ret_V_19_fu_594_p3;
wire [2:0] ret_V_3_fu_229_p2;
wire [1:0] ret_V_fu_205_p4;
wire [4:0] rhs_2_fu_286_p1;
wire [33:0] rhs_5_fu_484_p3;
wire [3:0] rhs_fu_187_p3;
wire [1:0] select_ln1498_fu_306_p3;
wire [4:0] select_ln850_1_fu_338_p3;
wire [31:0] select_ln850_2_fu_410_p3;
wire [31:0] select_ln850_3_fu_588_p3;
wire [2:0] select_ln850_fu_256_p3;
wire [1:0] sext_ln1192_1_fu_274_p0;
wire [4:0] sext_ln1192_1_fu_274_p1;
wire [33:0] sext_ln1192_2_fu_375_p1;
wire [34:0] sext_ln1192_3_fu_491_p1;
wire [3:0] sext_ln1192_fu_183_p0;
wire [4:0] sext_ln1192_fu_183_p1;
wire [31:0] sext_ln1497_1_fu_551_p1;
wire [1:0] sext_ln1497_fu_465_p0;
wire [2:0] sext_ln1497_fu_465_p1;
wire [7:0] sext_ln1498_fu_440_p1;
wire [1:0] sext_ln545_fu_528_p0;
wire [31:0] sext_ln545_fu_528_p1;
wire [3:0] sext_ln69_1_fu_610_p1;
wire [31:0] sext_ln69_fu_423_p1;
wire [7:0] sext_ln703_1_fu_480_p0;
wire [34:0] sext_ln703_1_fu_480_p1;
wire [7:0] sext_ln703_fu_364_p0;
wire [33:0] sext_ln703_fu_364_p1;
wire [1:0] sext_ln727_fu_450_p0;
wire [2:0] sext_ln727_fu_450_p1;
wire [2:0] sext_ln835_fu_215_p1;
wire [4:0] sext_ln850_fu_319_p1;
wire [31:0] shl_ln1497_fu_541_p2;
wire [1:0] shl_ln728_1_fu_235_p1;
wire [31:0] shl_ln728_1_fu_235_p3;
wire [1:0] shl_ln728_3_fu_453_p3;
wire [1:0] shl_ln_fu_433_p1;
wire [5:0] shl_ln_fu_433_p3;
wire [2:0] sub_ln1497_fu_468_p2;
wire [3:0] tmp_1_fu_278_p3;
wire [5:0] tmp_4_fu_368_p3;
wire [1:0] tmp_fu_531_p1;
wire tmp_fu_531_p3;
wire trunc_ln1497_1_fu_560_p1;
wire [1:0] trunc_ln1497_fu_547_p1;
wire [1:0] trunc_ln851_1_fu_329_p0;
wire trunc_ln851_1_fu_329_p1;
wire [7:0] trunc_ln851_2_fu_407_p0;
wire trunc_ln851_2_fu_407_p1;
wire [7:0] trunc_ln851_3_fu_511_p0;
wire [1:0] trunc_ln851_3_fu_511_p1;
wire [3:0] trunc_ln851_fu_219_p0;
wire [2:0] trunc_ln851_fu_219_p1;
wire [4:0] zext_ln1192_fu_195_p1;
wire [1:0] zext_ln1497_fu_564_p1;
wire [31:0] zext_ln69_1_fu_613_p1;
wire [1:0] zext_ln69_2_fu_601_p1;
wire [31:0] zext_ln69_3_fu_622_p1;
wire [4:0] zext_ln69_fu_354_p1;
wire [2:0] zext_ln835_fu_461_p1;


assign add_ln691_1_fu_395_p2 = ret_V_7_cast_reg_702 + 1'h1;
assign add_ln691_2_fu_583_p2 = ret_V_15_cast_reg_739 + 1'h1;
assign add_ln691_fu_332_p2 = $signed(tmp_2_reg_674) + $signed(2'h1);
assign add_ln69_1_fu_604_p2 = op_17_V_fu_568_p3 + icmp_ln1495_reg_729;
assign add_ln69_fu_617_p2 = ret_V_19_reg_756 + { ret_V_11_reg_751[1], ret_V_11_reg_751[1], ret_V_11_reg_751 };
assign op_21_V_fu_268_p2 = ret_V_13_fu_261_p3 + 1'h1;
assign op_23_V_fu_358_p2 = ret_V_15_fu_346_p3 + icmp_ln1498_1_fu_313_p2;
assign op_25_V_fu_427_p2 = $signed(ret_V_17_fu_416_p3) + $signed(op_15);
assign op_29 = add_ln69_1_reg_761 + add_ln69_fu_617_p2;
assign ret_V_12_fu_199_p2 = $signed({ 1'h0, op_8, 3'h0 }) + $signed(op_0);
assign ret_V_14_fu_290_p2 = $signed({ op_21_V_fu_268_p2, 1'h0 }) + $signed(op_10);
assign { ret_V_16_fu_379_p2[33], ret_V_16_fu_379_p2[7:0] } = $signed({ op_23_V_reg_687, 1'h0 }) + $signed(op_14);
assign ret_V_18_fu_495_p2 = $signed({ op_25_V_reg_714, 2'h0 }) + $signed(op_16);
assign ret_V_3_fu_229_p2 = $signed(ret_V_12_fu_199_p2[4:3]) + $signed(2'h1);
assign _023_ = ap_CS_fsm[0] & _025_;
assign _024_ = ap_CS_fsm[0] & ap_start;
assign _025_ = ~ ap_start;
assign _026_ = select_ln1498_fu_306_p3 == op_7;
assign _027_ = { op_2[1], op_2[1], op_2, 4'h0 } == op_1;
assign _028_ = ! op_0[2:0];
assign _029_ = $signed({ op_2, 30'h00000000 }) > $signed(op_4);
assign _030_ = $signed(op_2) < $signed({ 1'h0, icmp_ln1498_fu_444_p2, 1'h0 });
assign _031_ = | op_16[1:0];
always @(posedge ap_clk)
ret_V_16_reg_697 <= _014_;
always @(posedge ap_clk)
ret_V_7_cast_reg_702 <= _018_;
always @(posedge ap_clk)
op_6_V_reg_664 <= _009_;
always @(posedge ap_clk)
ret_V_14_reg_669 <= _012_;
always @(posedge ap_clk)
tmp_2_reg_674 <= _021_;
always @(posedge ap_clk)
op_25_V_reg_714 <= _008_;
always @(posedge ap_clk)
op_23_V_reg_687 <= _007_;
always @(posedge ap_clk)
ret_V_12_reg_632 <= _011_;
always @(posedge ap_clk)
sext_ln835_reg_637 <= _019_;
always @(posedge ap_clk)
icmp_ln851_reg_643 <= _006_;
always @(posedge ap_clk)
ret_V_3_reg_648 <= _017_;
always @(posedge ap_clk)
icmp_ln1498_reg_719 <= _004_;
always @(posedge ap_clk)
sub_ln1497_reg_724 <= _020_;
always @(posedge ap_clk)
icmp_ln1495_reg_729 <= _003_;
always @(posedge ap_clk)
ret_V_18_reg_734 <= _015_;
always @(posedge ap_clk)
ret_V_15_cast_reg_739 <= _013_;
always @(posedge ap_clk)
icmp_ln851_1_reg_746 <= _005_;
always @(posedge ap_clk)
ret_V_11_reg_751 <= _010_;
always @(posedge ap_clk)
ret_V_19_reg_756 <= _016_;
always @(posedge ap_clk)
add_ln69_1_reg_761 <= _001_;
always @(posedge ap_clk)
add_ln691_1_reg_709 <= _000_;
always @(posedge ap_clk)
ap_CS_fsm <= _002_;
function [8:0] _086_;
input [8:0] a;
input [80:0] b;
input [8:0] s;
case (s)
9'b000000001:
_086_ = b[8:0];
9'b000000010:
_086_ = b[17:9];
9'b000000100:
_086_ = b[26:18];
9'b000001000:
_086_ = b[35:27];
9'b000010000:
_086_ = b[44:36];
9'b000100000:
_086_ = b[53:45];
9'b001000000:
_086_ = b[62:54];
9'b010000000:
_086_ = b[71:63];
9'b100000000:
_086_ = b[80:72];
9'b000000000:
_086_ = a;
default:
_086_ = 9'bx;
endcase
endfunction
assign ap_NS_fsm = _086_(9'hxxx, { 7'h00, _022_, 72'h020202020202020001 }, { _040_, _039_, _038_, _037_, _036_, _035_, _034_, _033_, _032_ });
assign _032_ = ap_CS_fsm == 9'h100;
assign _033_ = ap_CS_fsm == 8'h80;
assign _034_ = ap_CS_fsm == 7'h40;
assign _035_ = ap_CS_fsm == 6'h20;
assign _036_ = ap_CS_fsm == 5'h10;
assign _037_ = ap_CS_fsm == 4'h8;
assign _038_ = ap_CS_fsm == 3'h4;
assign _039_ = ap_CS_fsm == 2'h2;
assign _040_ = ap_CS_fsm == 1'h1;
assign op_29_ap_vld = ap_CS_fsm[8] ? 1'h1 : 1'h0;
assign ap_idle = _023_ ? 1'h1 : 1'h0;
assign _018_ = ap_CS_fsm[3] ? { ret_V_16_fu_379_p2[33], ret_V_16_fu_379_p2[33], ret_V_16_fu_379_p2[33], ret_V_16_fu_379_p2[33], ret_V_16_fu_379_p2[33], ret_V_16_fu_379_p2[33], ret_V_16_fu_379_p2[33], ret_V_16_fu_379_p2[33], ret_V_16_fu_379_p2[33], ret_V_16_fu_379_p2[33], ret_V_16_fu_379_p2[33], ret_V_16_fu_379_p2[33], ret_V_16_fu_379_p2[33], ret_V_16_fu_379_p2[33], ret_V_16_fu_379_p2[33], ret_V_16_fu_379_p2[33], ret_V_16_fu_379_p2[33], ret_V_16_fu_379_p2[33], ret_V_16_fu_379_p2[33], ret_V_16_fu_379_p2[33], ret_V_16_fu_379_p2[33], ret_V_16_fu_379_p2[33], ret_V_16_fu_379_p2[33], ret_V_16_fu_379_p2[33], ret_V_16_fu_379_p2[33], ret_V_16_fu_379_p2[7:1] } : ret_V_7_cast_reg_702;
assign _014_ = ap_CS_fsm[3] ? { ret_V_16_fu_379_p2[33], ret_V_16_fu_379_p2[33], ret_V_16_fu_379_p2[33], ret_V_16_fu_379_p2[33], ret_V_16_fu_379_p2[33], ret_V_16_fu_379_p2[33], ret_V_16_fu_379_p2[33], ret_V_16_fu_379_p2[33], ret_V_16_fu_379_p2[33], ret_V_16_fu_379_p2[33], ret_V_16_fu_379_p2[33], ret_V_16_fu_379_p2[33], ret_V_16_fu_379_p2[33], ret_V_16_fu_379_p2[33], ret_V_16_fu_379_p2[33], ret_V_16_fu_379_p2[33], ret_V_16_fu_379_p2[33], ret_V_16_fu_379_p2[33], ret_V_16_fu_379_p2[33], ret_V_16_fu_379_p2[33], ret_V_16_fu_379_p2[33], ret_V_16_fu_379_p2[33], ret_V_16_fu_379_p2[33], ret_V_16_fu_379_p2[33], ret_V_16_fu_379_p2[33], ret_V_16_fu_379_p2[33], ret_V_16_fu_379_p2[7:0] } : ret_V_16_reg_697;
assign _021_ = ap_CS_fsm[1] ? ret_V_14_fu_290_p2[4:1] : tmp_2_reg_674;
assign _012_ = ap_CS_fsm[1] ? ret_V_14_fu_290_p2 : ret_V_14_reg_669;
assign _009_ = ap_CS_fsm[1] ? op_6_V_fu_243_p2 : op_6_V_reg_664;
assign _008_ = ap_CS_fsm[5] ? op_25_V_fu_427_p2 : op_25_V_reg_714;
assign _007_ = ap_CS_fsm[2] ? op_23_V_fu_358_p2 : op_23_V_reg_687;
assign _017_ = ap_CS_fsm[0] ? ret_V_3_fu_229_p2 : ret_V_3_reg_648;
assign _006_ = ap_CS_fsm[0] ? icmp_ln851_fu_223_p2 : icmp_ln851_reg_643;
assign _019_ = ap_CS_fsm[0] ? { ret_V_12_fu_199_p2[4], ret_V_12_fu_199_p2[4:3] } : sext_ln835_reg_637;
assign _011_ = ap_CS_fsm[0] ? ret_V_12_fu_199_p2 : ret_V_12_reg_632;
assign _005_ = ap_CS_fsm[6] ? icmp_ln851_1_fu_515_p2 : icmp_ln851_1_reg_746;
assign _013_ = ap_CS_fsm[6] ? ret_V_18_fu_495_p2[33:2] : ret_V_15_cast_reg_739;
assign _015_ = ap_CS_fsm[6] ? ret_V_18_fu_495_p2 : ret_V_18_reg_734;
assign _003_ = ap_CS_fsm[6] ? icmp_ln1495_fu_474_p2 : icmp_ln1495_reg_729;
assign _020_ = ap_CS_fsm[6] ? sub_ln1497_fu_468_p2 : sub_ln1497_reg_724;
assign _004_ = ap_CS_fsm[6] ? icmp_ln1498_fu_444_p2 : icmp_ln1498_reg_719;
assign _001_ = ap_CS_fsm[7] ? add_ln69_1_fu_604_p2 : add_ln69_1_reg_761;
assign _016_ = ap_CS_fsm[7] ? ret_V_19_fu_594_p3 : ret_V_19_reg_756;
assign _010_ = ap_CS_fsm[7] ? ret_V_11_fu_521_p3 : ret_V_11_reg_751;
assign _000_ = ap_CS_fsm[4] ? add_ln691_1_fu_395_p2 : add_ln691_1_reg_709;
assign _002_ = ap_rst ? 9'h001 : ap_NS_fsm;
assign _022_ = _024_ ? 2'h2 : 2'h1;
assign trunc_ln1497_fu_547_p1 = icmp_ln1498_reg_719 << { op_7[1], op_7[1], op_7[1], op_7[1], op_7[1], op_7[1], op_7[1], op_7[1], op_7[1], op_7[1], op_7[1], op_7[1], op_7[1], op_7[1], op_7[1], op_7[1], op_7[1], op_7[1], op_7[1], op_7[1], op_7[1], op_7[1], op_7[1], op_7[1], op_7[1], op_7[1], op_7[1], op_7[1], op_7[1], op_7[1], op_7 };
assign trunc_ln1497_1_fu_560_p1 = icmp_ln1498_reg_719 >> { sub_ln1497_reg_724[2], sub_ln1497_reg_724[2], sub_ln1497_reg_724[2], sub_ln1497_reg_724[2], sub_ln1497_reg_724[2], sub_ln1497_reg_724[2], sub_ln1497_reg_724[2], sub_ln1497_reg_724[2], sub_ln1497_reg_724[2], sub_ln1497_reg_724[2], sub_ln1497_reg_724[2], sub_ln1497_reg_724[2], sub_ln1497_reg_724[2], sub_ln1497_reg_724[2], sub_ln1497_reg_724[2], sub_ln1497_reg_724[2], sub_ln1497_reg_724[2], sub_ln1497_reg_724[2], sub_ln1497_reg_724[2], sub_ln1497_reg_724[2], sub_ln1497_reg_724[2], sub_ln1497_reg_724[2], sub_ln1497_reg_724[2], sub_ln1497_reg_724[2], sub_ln1497_reg_724[2], sub_ln1497_reg_724[2], sub_ln1497_reg_724[2], sub_ln1497_reg_724[2], sub_ln1497_reg_724[2], sub_ln1497_reg_724 };
assign sub_ln1497_fu_468_p2 = $signed(1'h0) - $signed(op_7);
assign icmp_ln1495_fu_474_p2 = _030_ ? 1'h1 : 1'h0;
assign icmp_ln1498_1_fu_313_p2 = _026_ ? 1'h1 : 1'h0;
assign icmp_ln1498_fu_444_p2 = _027_ ? 1'h1 : 1'h0;
assign icmp_ln851_1_fu_515_p2 = _031_ ? 1'h1 : 1'h0;
assign icmp_ln851_fu_223_p2 = _028_ ? 1'h1 : 1'h0;
assign op_17_V_fu_568_p3 = op_7[1] ? { 1'h0, trunc_ln1497_1_fu_560_p1 } : trunc_ln1497_fu_547_p1;
assign op_6_V_fu_243_p2 = _029_ ? 1'h1 : 1'h0;
assign ret_V_11_fu_521_p3 = op_3 ? op_7 : 2'h0;
assign ret_V_13_fu_261_p3 = ret_V_12_reg_632[4] ? select_ln850_fu_256_p3 : sext_ln835_reg_637;
assign ret_V_15_fu_346_p3 = ret_V_14_reg_669[4] ? select_ln850_1_fu_338_p3 : { tmp_2_reg_674[3], tmp_2_reg_674 };
assign ret_V_17_fu_416_p3 = ret_V_16_reg_697[33] ? select_ln850_2_fu_410_p3 : ret_V_7_cast_reg_702;
assign ret_V_19_fu_594_p3 = ret_V_18_reg_734[34] ? select_ln850_3_fu_588_p3 : ret_V_15_cast_reg_739;
assign select_ln1498_fu_306_p3 = op_6_V_reg_664 ? 2'h3 : 2'h0;
assign select_ln850_1_fu_338_p3 = op_10[0] ? add_ln691_fu_332_p2 : { tmp_2_reg_674[3], tmp_2_reg_674 };
assign select_ln850_2_fu_410_p3 = op_14[0] ? add_ln691_1_reg_709 : ret_V_7_cast_reg_702;
assign select_ln850_3_fu_588_p3 = icmp_ln851_1_reg_746 ? add_ln691_2_fu_583_p2 : ret_V_15_cast_reg_739;
assign select_ln850_fu_256_p3 = icmp_ln851_reg_643 ? sext_ln835_reg_637 : ret_V_3_reg_648;
assign ap_CS_fsm_state1 = ap_CS_fsm[0];
assign ap_CS_fsm_state2 = ap_CS_fsm[1];
assign ap_CS_fsm_state3 = ap_CS_fsm[2];
assign ap_CS_fsm_state4 = ap_CS_fsm[3];
assign ap_CS_fsm_state5 = ap_CS_fsm[4];
assign ap_CS_fsm_state6 = ap_CS_fsm[5];
assign ap_CS_fsm_state7 = ap_CS_fsm[6];
assign ap_CS_fsm_state8 = ap_CS_fsm[7];
assign ap_CS_fsm_state9 = ap_CS_fsm[8];
assign ap_done = op_29_ap_vld;
assign ap_ready = op_29_ap_vld;
assign conv_i270_fu_538_p1 = { 31'h00000000, icmp_ln1498_reg_719 };
assign icmp_ln1498_1_fu_313_p1 = op_7;
assign lshr_ln1497_fu_554_p2[0] = trunc_ln1497_1_fu_560_p1;
assign p_Result_1_fu_322_p3 = ret_V_14_reg_669[4];
assign p_Result_2_fu_400_p3 = ret_V_16_reg_697[33];
assign p_Result_3_fu_576_p3 = ret_V_18_reg_734[34];
assign p_Result_s_fu_249_p3 = ret_V_12_reg_632[4];
assign ret_V_11_fu_521_p1 = op_7;
assign ret_V_16_fu_379_p2[32:8] = { ret_V_16_fu_379_p2[33], ret_V_16_fu_379_p2[33], ret_V_16_fu_379_p2[33], ret_V_16_fu_379_p2[33], ret_V_16_fu_379_p2[33], ret_V_16_fu_379_p2[33], ret_V_16_fu_379_p2[33], ret_V_16_fu_379_p2[33], ret_V_16_fu_379_p2[33], ret_V_16_fu_379_p2[33], ret_V_16_fu_379_p2[33], ret_V_16_fu_379_p2[33], ret_V_16_fu_379_p2[33], ret_V_16_fu_379_p2[33], ret_V_16_fu_379_p2[33], ret_V_16_fu_379_p2[33], ret_V_16_fu_379_p2[33], ret_V_16_fu_379_p2[33], ret_V_16_fu_379_p2[33], ret_V_16_fu_379_p2[33], ret_V_16_fu_379_p2[33], ret_V_16_fu_379_p2[33], ret_V_16_fu_379_p2[33], ret_V_16_fu_379_p2[33], ret_V_16_fu_379_p2[33] };
assign ret_V_fu_205_p4 = ret_V_12_fu_199_p2[4:3];
assign rhs_2_fu_286_p1 = { op_21_V_fu_268_p2[2], op_21_V_fu_268_p2, 1'h0 };
assign rhs_5_fu_484_p3 = { op_25_V_reg_714, 2'h0 };
assign rhs_fu_187_p3 = { op_8, 3'h0 };
assign sext_ln1192_1_fu_274_p0 = op_10;
assign sext_ln1192_1_fu_274_p1 = { op_10[1], op_10[1], op_10[1], op_10 };
assign sext_ln1192_2_fu_375_p1 = { op_23_V_reg_687[4], op_23_V_reg_687[4], op_23_V_reg_687[4], op_23_V_reg_687[4], op_23_V_reg_687[4], op_23_V_reg_687[4], op_23_V_reg_687[4], op_23_V_reg_687[4], op_23_V_reg_687[4], op_23_V_reg_687[4], op_23_V_reg_687[4], op_23_V_reg_687[4], op_23_V_reg_687[4], op_23_V_reg_687[4], op_23_V_reg_687[4], op_23_V_reg_687[4], op_23_V_reg_687[4], op_23_V_reg_687[4], op_23_V_reg_687[4], op_23_V_reg_687[4], op_23_V_reg_687[4], op_23_V_reg_687[4], op_23_V_reg_687[4], op_23_V_reg_687[4], op_23_V_reg_687[4], op_23_V_reg_687[4], op_23_V_reg_687[4], op_23_V_reg_687[4], op_23_V_reg_687, 1'h0 };
assign sext_ln1192_3_fu_491_p1 = { op_25_V_reg_714[31], op_25_V_reg_714, 2'h0 };
assign sext_ln1192_fu_183_p0 = op_0;
assign sext_ln1192_fu_183_p1 = { op_0[3], op_0 };
assign sext_ln1497_1_fu_551_p1 = { sub_ln1497_reg_724[2], sub_ln1497_reg_724[2], sub_ln1497_reg_724[2], sub_ln1497_reg_724[2], sub_ln1497_reg_724[2], sub_ln1497_reg_724[2], sub_ln1497_reg_724[2], sub_ln1497_reg_724[2], sub_ln1497_reg_724[2], sub_ln1497_reg_724[2], sub_ln1497_reg_724[2], sub_ln1497_reg_724[2], sub_ln1497_reg_724[2], sub_ln1497_reg_724[2], sub_ln1497_reg_724[2], sub_ln1497_reg_724[2], sub_ln1497_reg_724[2], sub_ln1497_reg_724[2], sub_ln1497_reg_724[2], sub_ln1497_reg_724[2], sub_ln1497_reg_724[2], sub_ln1497_reg_724[2], sub_ln1497_reg_724[2], sub_ln1497_reg_724[2], sub_ln1497_reg_724[2], sub_ln1497_reg_724[2], sub_ln1497_reg_724[2], sub_ln1497_reg_724[2], sub_ln1497_reg_724[2], sub_ln1497_reg_724 };
assign sext_ln1497_fu_465_p0 = op_7;
assign sext_ln1497_fu_465_p1 = { op_7[1], op_7 };
assign sext_ln1498_fu_440_p1 = { op_2[1], op_2[1], op_2, 4'h0 };
assign sext_ln545_fu_528_p0 = op_7;
assign sext_ln545_fu_528_p1 = { op_7[1], op_7[1], op_7[1], op_7[1], op_7[1], op_7[1], op_7[1], op_7[1], op_7[1], op_7[1], op_7[1], op_7[1], op_7[1], op_7[1], op_7[1], op_7[1], op_7[1], op_7[1], op_7[1], op_7[1], op_7[1], op_7[1], op_7[1], op_7[1], op_7[1], op_7[1], op_7[1], op_7[1], op_7[1], op_7[1], op_7 };
assign sext_ln69_1_fu_610_p1 = { ret_V_11_reg_751[1], ret_V_11_reg_751[1], ret_V_11_reg_751 };
assign sext_ln69_fu_423_p1 = { op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15 };
assign sext_ln703_1_fu_480_p0 = op_16;
assign sext_ln703_1_fu_480_p1 = { op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16 };
assign sext_ln703_fu_364_p0 = op_14;
assign sext_ln703_fu_364_p1 = { op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14 };
assign sext_ln727_fu_450_p0 = op_2;
assign sext_ln727_fu_450_p1 = { op_2[1], op_2 };
assign sext_ln835_fu_215_p1 = { ret_V_12_fu_199_p2[4], ret_V_12_fu_199_p2[4:3] };
assign sext_ln850_fu_319_p1 = { tmp_2_reg_674[3], tmp_2_reg_674 };
assign shl_ln1497_fu_541_p2[1:0] = trunc_ln1497_fu_547_p1;
assign shl_ln728_1_fu_235_p1 = op_2;
assign shl_ln728_1_fu_235_p3 = { op_2, 30'h00000000 };
assign shl_ln728_3_fu_453_p3 = { icmp_ln1498_fu_444_p2, 1'h0 };
assign shl_ln_fu_433_p1 = op_2;
assign shl_ln_fu_433_p3 = { op_2, 4'h0 };
assign tmp_1_fu_278_p3 = { op_21_V_fu_268_p2, 1'h0 };
assign tmp_4_fu_368_p3 = { op_23_V_reg_687, 1'h0 };
assign tmp_fu_531_p1 = op_7;
assign tmp_fu_531_p3 = op_7[1];
assign trunc_ln851_1_fu_329_p0 = op_10;
assign trunc_ln851_1_fu_329_p1 = op_10[0];
assign trunc_ln851_2_fu_407_p0 = op_14;
assign trunc_ln851_2_fu_407_p1 = op_14[0];
assign trunc_ln851_3_fu_511_p0 = op_16;
assign trunc_ln851_3_fu_511_p1 = op_16[1:0];
assign trunc_ln851_fu_219_p0 = op_0;
assign trunc_ln851_fu_219_p1 = op_0[2:0];
assign zext_ln1192_fu_195_p1 = { 1'h0, op_8, 3'h0 };
assign zext_ln1497_fu_564_p1 = { 1'h0, trunc_ln1497_1_fu_560_p1 };
assign zext_ln69_1_fu_613_p1 = { 28'h0000000, ret_V_11_reg_751[1], ret_V_11_reg_751[1], ret_V_11_reg_751 };
assign zext_ln69_2_fu_601_p1 = { 1'h0, icmp_ln1495_reg_729 };
assign zext_ln69_3_fu_622_p1 = { 30'h00000000, add_ln69_1_reg_761 };
assign zext_ln69_fu_354_p1 = { 4'h0, icmp_ln1498_1_fu_313_p2 };
assign zext_ln835_fu_461_p1 = { 1'h0, icmp_ln1498_fu_444_p2, 1'h0 };
endmodule


// Product machine:
module top_A_times_top_B (ap_start, op_0, op_1, op_10, op_14, op_15, op_16, op_2, op_3, op_4, op_7, op_8, ap_clk, unsafe_signal);
input ap_start;
input [3:0] op_0;
input [7:0] op_1;
input [1:0] op_10;
input [7:0] op_14;
input [3:0] op_15;
input [7:0] op_16;
input [1:0] op_2;
input op_3;
input [31:0] op_4;
input [1:0] op_7;
input op_8;
input ap_clk;
output unsafe_signal;
reg _setup;
initial _setup = 1'b0;
always @ (posedge ap_clk) _setup <= 1'b1;
reg ap_start_internal;
always @ (posedge ap_clk) if (!_setup) ap_start_internal <= ap_start;
reg [3:0] op_0_internal;
always @ (posedge ap_clk) if (!_setup) op_0_internal <= op_0;
reg [7:0] op_1_internal;
always @ (posedge ap_clk) if (!_setup) op_1_internal <= op_1;
reg [1:0] op_10_internal;
always @ (posedge ap_clk) if (!_setup) op_10_internal <= op_10;
reg [7:0] op_14_internal;
always @ (posedge ap_clk) if (!_setup) op_14_internal <= op_14;
reg [3:0] op_15_internal;
always @ (posedge ap_clk) if (!_setup) op_15_internal <= op_15;
reg [7:0] op_16_internal;
always @ (posedge ap_clk) if (!_setup) op_16_internal <= op_16;
reg [1:0] op_2_internal;
always @ (posedge ap_clk) if (!_setup) op_2_internal <= op_2;
reg op_3_internal;
always @ (posedge ap_clk) if (!_setup) op_3_internal <= op_3;
reg [31:0] op_4_internal;
always @ (posedge ap_clk) if (!_setup) op_4_internal <= op_4;
reg [1:0] op_7_internal;
always @ (posedge ap_clk) if (!_setup) op_7_internal <= op_7;
reg op_8_internal;
always @ (posedge ap_clk) if (!_setup) op_8_internal <= op_8;
wire ap_done_A;
wire ap_done_B;
wire ap_done_eq;
assign ap_done_eq = ap_done_A == ap_done_B;
wire ap_idle_A;
wire ap_idle_B;
wire ap_idle_eq;
assign ap_idle_eq = ap_idle_A == ap_idle_B;
wire ap_ready_A;
wire ap_ready_B;
wire ap_ready_eq;
assign ap_ready_eq = ap_ready_A == ap_ready_B;
wire [31:0] op_29_A;
wire [31:0] op_29_B;
wire op_29_eq;
assign op_29_eq = op_29_A == op_29_B;
wire op_29_ap_vld_A;
wire op_29_ap_vld_B;
wire clk_enable_A;
wire clk_enable_B;
assign clk_enable_A = _setup & (~op_29_ap_vld_A | op_29_ap_vld_B);
assign clk_enable_B = _setup;
wire divergent;
assign divergent = ~(ap_done_eq & ap_idle_eq & ap_ready_eq & op_29_eq);
assign unsafe_signal = op_29_ap_vld_A & op_29_ap_vld_B & divergent;
top_A instance_A (
    .ap_clk(ap_clk),
    .clk_enable(clk_enable_A),
    .ap_start(ap_start_internal),
    .op_0(op_0_internal),
    .op_1(op_1_internal),
    .op_10(op_10_internal),
    .op_14(op_14_internal),
    .op_15(op_15_internal),
    .op_16(op_16_internal),
    .op_2(op_2_internal),
    .op_3(op_3_internal),
    .op_4(op_4_internal),
    .op_7(op_7_internal),
    .op_8(op_8_internal),
    .ap_done(ap_done_A),
    .ap_idle(ap_idle_A),
    .ap_ready(ap_ready_A),
    .op_29(op_29_A),
    .op_29_ap_vld(op_29_ap_vld_A)
);
top_B instance_B (
    .ap_clk(ap_clk),
    .clk_enable(clk_enable_B),
    .ap_start(ap_start_internal),
    .op_0(op_0_internal),
    .op_1(op_1_internal),
    .op_10(op_10_internal),
    .op_14(op_14_internal),
    .op_15(op_15_internal),
    .op_16(op_16_internal),
    .op_2(op_2_internal),
    .op_3(op_3_internal),
    .op_4(op_4_internal),
    .op_7(op_7_internal),
    .op_8(op_8_internal),
    .ap_done(ap_done_B),
    .ap_idle(ap_idle_B),
    .ap_ready(ap_ready_B),
    .op_29(op_29_B),
    .op_29_ap_vld(op_29_ap_vld_B)
);
endmodule
