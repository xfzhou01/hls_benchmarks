// Processed by function `construct_kairos` in `verilog_tricks.py`.
// Machine A:
// Processed by function `add_clk_enable_signal` in `verilog_tricks.py`.
// Processed by function `remove_reset_signal` in `verilog_tricks.py`.
module top_A (
  ap_clk,
  ap_start,
  ap_done,
  ap_idle,
  ap_ready,
  op_0,
  op_1,
  op_2,
  op_4,
  op_5,
  op_13,
  op_14,
  op_15,
  op_16,
  op_17,
  op_18,
  op_29,
  op_29_ap_vld,
clk_enable
);
input clk_enable;


input ap_clk;
wire ap_rst;
assign ap_rst = op_29_ap_vld;
input ap_start;
input [7:0] op_0;
input [7:0] op_1;
input [15:0] op_13;
input [7:0] op_14;
input [3:0] op_15;
input [1:0] op_16;
input [1:0] op_17;
input [3:0] op_18;
input [3:0] op_2;
input [31:0] op_4;
input op_5;
output ap_done;
output ap_idle;
output ap_ready;
output [31:0] op_29;
output op_29_ap_vld;


reg Range1_all_ones_reg_1119;
reg [8:0] \add_17s_17ns_17_2_1_U18.top_add_17s_17ns_17_2_1_Adder_12_U.ain_s1 ;
reg [8:0] \add_17s_17ns_17_2_1_U18.top_add_17s_17ns_17_2_1_Adder_12_U.bin_s1 ;
reg \add_17s_17ns_17_2_1_U18.top_add_17s_17ns_17_2_1_Adder_12_U.carry_s1 ;
reg [7:0] \add_17s_17ns_17_2_1_U18.top_add_17s_17ns_17_2_1_Adder_12_U.sum_s1 ;
reg [8:0] \add_17s_17s_17_2_1_U15.top_add_17s_17s_17_2_1_Adder_11_U.ain_s1 ;
reg [8:0] \add_17s_17s_17_2_1_U15.top_add_17s_17s_17_2_1_Adder_11_U.bin_s1 ;
reg \add_17s_17s_17_2_1_U15.top_add_17s_17s_17_2_1_Adder_11_U.carry_s1 ;
reg [7:0] \add_17s_17s_17_2_1_U15.top_add_17s_17s_17_2_1_Adder_11_U.sum_s1 ;
reg [14:0] \add_29s_29ns_29_2_1_U12.top_add_29s_29ns_29_2_1_Adder_9_U.ain_s1 ;
reg [14:0] \add_29s_29ns_29_2_1_U12.top_add_29s_29ns_29_2_1_Adder_9_U.bin_s1 ;
reg \add_29s_29ns_29_2_1_U12.top_add_29s_29ns_29_2_1_Adder_9_U.carry_s1 ;
reg [13:0] \add_29s_29ns_29_2_1_U12.top_add_29s_29ns_29_2_1_Adder_9_U.sum_s1 ;
reg \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.ain_s1 ;
reg \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.bin_s1 ;
reg \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.carry_s1 ;
reg \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.sum_s1 ;
reg \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_0_U.ain_s1 ;
reg \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_0_U.bin_s1 ;
reg \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_0_U.carry_s1 ;
reg \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_0_U.sum_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_14_U.ain_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_14_U.bin_s1 ;
reg \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_14_U.carry_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_14_U.sum_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_14_U.ain_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_14_U.bin_s1 ;
reg \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_14_U.carry_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_14_U.sum_s1 ;
reg [15:0] \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_16_U.ain_s1 ;
reg [15:0] \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_16_U.bin_s1 ;
reg \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_16_U.carry_s1 ;
reg [15:0] \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_16_U.sum_s1 ;
reg [16:0] \add_34s_34s_34_2_1_U19.top_add_34s_34s_34_2_1_Adder_13_U.ain_s1 ;
reg [16:0] \add_34s_34s_34_2_1_U19.top_add_34s_34s_34_2_1_Adder_13_U.bin_s1 ;
reg \add_34s_34s_34_2_1_U19.top_add_34s_34s_34_2_1_Adder_13_U.carry_s1 ;
reg [16:0] \add_34s_34s_34_2_1_U19.top_add_34s_34s_34_2_1_Adder_13_U.sum_s1 ;
reg [1:0] \add_3ns_3ns_3_2_1_U8.top_add_3ns_3ns_3_2_1_Adder_6_U.ain_s1 ;
reg [1:0] \add_3ns_3ns_3_2_1_U8.top_add_3ns_3ns_3_2_1_Adder_6_U.bin_s1 ;
reg \add_3ns_3ns_3_2_1_U8.top_add_3ns_3ns_3_2_1_Adder_6_U.carry_s1 ;
reg \add_3ns_3ns_3_2_1_U8.top_add_3ns_3ns_3_2_1_Adder_6_U.sum_s1 ;
reg [2:0] \add_5ns_5ns_5_2_1_U9.top_add_5ns_5ns_5_2_1_Adder_7_U.ain_s1 ;
reg [2:0] \add_5ns_5ns_5_2_1_U9.top_add_5ns_5ns_5_2_1_Adder_7_U.bin_s1 ;
reg \add_5ns_5ns_5_2_1_U9.top_add_5ns_5ns_5_2_1_Adder_7_U.carry_s1 ;
reg [1:0] \add_5ns_5ns_5_2_1_U9.top_add_5ns_5ns_5_2_1_Adder_7_U.sum_s1 ;
reg [2:0] \add_5s_5ns_5_2_1_U10.top_add_5s_5ns_5_2_1_Adder_8_U.ain_s1 ;
reg [2:0] \add_5s_5ns_5_2_1_U10.top_add_5s_5ns_5_2_1_Adder_8_U.bin_s1 ;
reg \add_5s_5ns_5_2_1_U10.top_add_5s_5ns_5_2_1_Adder_8_U.carry_s1 ;
reg [1:0] \add_5s_5ns_5_2_1_U10.top_add_5s_5ns_5_2_1_Adder_8_U.sum_s1 ;
reg [2:0] \add_5s_5s_5_2_1_U22.top_add_5s_5s_5_2_1_Adder_15_U.ain_s1 ;
reg [2:0] \add_5s_5s_5_2_1_U22.top_add_5s_5s_5_2_1_Adder_15_U.bin_s1 ;
reg \add_5s_5s_5_2_1_U22.top_add_5s_5s_5_2_1_Adder_15_U.carry_s1 ;
reg [1:0] \add_5s_5s_5_2_1_U22.top_add_5s_5s_5_2_1_Adder_15_U.sum_s1 ;
reg [3:0] \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_5_U.ain_s1 ;
reg [3:0] \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_5_U.bin_s1 ;
reg \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_5_U.carry_s1 ;
reg [3:0] \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_5_U.sum_s1 ;
reg [4:0] \add_9s_9s_9_2_1_U13.top_add_9s_9s_9_2_1_Adder_4_U.ain_s1 ;
reg [4:0] \add_9s_9s_9_2_1_U13.top_add_9s_9s_9_2_1_Adder_4_U.bin_s1 ;
reg \add_9s_9s_9_2_1_U13.top_add_9s_9s_9_2_1_Adder_4_U.carry_s1 ;
reg [3:0] \add_9s_9s_9_2_1_U13.top_add_9s_9s_9_2_1_Adder_4_U.sum_s1 ;
reg [4:0] \add_9s_9s_9_2_1_U6.top_add_9s_9s_9_2_1_Adder_4_U.ain_s1 ;
reg [4:0] \add_9s_9s_9_2_1_U6.top_add_9s_9s_9_2_1_Adder_4_U.bin_s1 ;
reg \add_9s_9s_9_2_1_U6.top_add_9s_9s_9_2_1_Adder_4_U.carry_s1 ;
reg [3:0] \add_9s_9s_9_2_1_U6.top_add_9s_9s_9_2_1_Adder_4_U.sum_s1 ;
reg [31:0] add_ln691_reg_1506;
reg [4:0] add_ln69_1_reg_1357;
reg [8:0] add_ln69_2_reg_1413;
reg [31:0] add_ln69_4_reg_1536;
reg [4:0] add_ln69_5_reg_1541;
reg [16:0] add_ln69_reg_1454;
reg [1:0] add_ln731_reg_1053;
reg [27:0] ap_CS_fsm = 28'h0000001;
reg [31:0] \ashr_32s_32s_32_7_1_U16.din1_cast_array[0] ;
reg [31:0] \ashr_32s_32s_32_7_1_U16.din1_cast_array[1] ;
reg [31:0] \ashr_32s_32s_32_7_1_U16.din1_cast_array[2] ;
reg [31:0] \ashr_32s_32s_32_7_1_U16.din1_cast_array[3] ;
reg [31:0] \ashr_32s_32s_32_7_1_U16.din1_cast_array[4] ;
reg [31:0] \ashr_32s_32s_32_7_1_U16.din1_cast_array[5] ;
reg [31:0] \ashr_32s_32s_32_7_1_U16.dout_array[0] ;
reg [31:0] \ashr_32s_32s_32_7_1_U16.dout_array[1] ;
reg [31:0] \ashr_32s_32s_32_7_1_U16.dout_array[2] ;
reg [31:0] \ashr_32s_32s_32_7_1_U16.dout_array[3] ;
reg [31:0] \ashr_32s_32s_32_7_1_U16.dout_array[4] ;
reg [31:0] \ashr_32s_32s_32_7_1_U16.dout_array[5] ;
reg icmp_ln785_reg_1124;
reg icmp_ln790_reg_1194;
reg icmp_ln850_reg_1209;
reg icmp_ln851_1_reg_1362;
reg icmp_ln851_2_reg_1249;
reg icmp_ln851_3_reg_1315;
reg icmp_ln851_reg_1288;
reg [31:0] \mul_32s_4s_36_7_1_U4.top_mul_32s_4s_36_7_1_Mul_DSP_0_U.a_reg0 ;
reg [3:0] \mul_32s_4s_36_7_1_U4.top_mul_32s_4s_36_7_1_Mul_DSP_0_U.b_reg0 ;
reg [35:0] \mul_32s_4s_36_7_1_U4.top_mul_32s_4s_36_7_1_Mul_DSP_0_U.buff0 ;
reg [35:0] \mul_32s_4s_36_7_1_U4.top_mul_32s_4s_36_7_1_Mul_DSP_0_U.buff1 ;
reg [35:0] \mul_32s_4s_36_7_1_U4.top_mul_32s_4s_36_7_1_Mul_DSP_0_U.buff2 ;
reg [35:0] \mul_32s_4s_36_7_1_U4.top_mul_32s_4s_36_7_1_Mul_DSP_0_U.buff3 ;
reg [35:0] \mul_32s_4s_36_7_1_U4.top_mul_32s_4s_36_7_1_Mul_DSP_0_U.buff4 ;
reg [3:0] op_21_V_reg_1408;
reg [16:0] op_25_V_reg_1464;
reg [7:0] op_3_V_reg_1058;
reg [3:0] op_6_V_reg_1113;
reg [7:0] op_8_V_reg_1214;
reg [25:0] or_ln1195_reg_1168;
reg or_ln384_reg_1183;
reg overflow_1_reg_1188;
reg overflow_reg_1134;
reg p_Result_11_reg_1085;
reg p_Result_12_reg_1091;
reg p_Result_13_reg_1145;
reg p_Result_14_reg_1151;
reg [7:0] p_Result_s_20_reg_1097;
reg [35:0] r_V_reg_1330;
reg [1:0] r_reg_1511;
reg [1:0] ret_V_10_reg_1398;
reg [2:0] ret_V_13_reg_1303;
reg [4:0] ret_V_14_reg_1347;
reg [4:0] ret_V_15_reg_1367;
reg [15:0] ret_V_21_reg_1079;
reg [8:0] ret_V_22_reg_1140;
reg [32:0] ret_V_23_reg_1259;
reg [1:0] ret_V_24_cast_reg_1335;
reg [1:0] ret_V_24_reg_1418;
reg [8:0] ret_V_25_reg_1276;
reg [33:0] ret_V_26_reg_1484;
reg [31:0] ret_V_27_reg_1516;
reg [31:0] ret_V_34_cast_reg_1489;
reg [2:0] ret_V_6_reg_1281;
reg [7:0] ret_V_7_reg_1298;
reg [7:0] ret_V_8_reg_1325;
reg [4:0] ret_V_9_reg_1308;
reg [7:0] ret_V_reg_1264;
reg [8:0] select_ln1193_reg_1103;
reg [1:0] select_ln384_3_reg_1219;
reg [4:0] select_ln69_reg_1254;
reg [2:0] select_ln850_7_reg_1352;
reg [31:0] \shl_32s_32s_32_7_1_U17.din1_cast_array[0] ;
reg [31:0] \shl_32s_32s_32_7_1_U17.din1_cast_array[1] ;
reg [31:0] \shl_32s_32s_32_7_1_U17.din1_cast_array[2] ;
reg [31:0] \shl_32s_32s_32_7_1_U17.din1_cast_array[3] ;
reg [31:0] \shl_32s_32s_32_7_1_U17.din1_cast_array[4] ;
reg [31:0] \shl_32s_32s_32_7_1_U17.din1_cast_array[5] ;
reg [31:0] \shl_32s_32s_32_7_1_U17.dout_array[0] ;
reg [31:0] \shl_32s_32s_32_7_1_U17.dout_array[1] ;
reg [31:0] \shl_32s_32s_32_7_1_U17.dout_array[2] ;
reg [31:0] \shl_32s_32s_32_7_1_U17.dout_array[3] ;
reg [31:0] \shl_32s_32s_32_7_1_U17.dout_array[4] ;
reg [31:0] \shl_32s_32s_32_7_1_U17.dout_array[5] ;
reg signbit_reg_1178;
reg [7:0] \sub_16ns_16s_16_2_1_U2.top_sub_16ns_16s_16_2_1_Adder_1_U.ain_s1 ;
reg [7:0] \sub_16ns_16s_16_2_1_U2.top_sub_16ns_16s_16_2_1_Adder_1_U.bin_s1 ;
reg \sub_16ns_16s_16_2_1_U2.top_sub_16ns_16s_16_2_1_Adder_1_U.carry_s1 ;
reg [7:0] \sub_16ns_16s_16_2_1_U2.top_sub_16ns_16s_16_2_1_Adder_1_U.sum_s1 ;
reg [16:0] \sub_33s_33s_33_2_1_U5.top_sub_33s_33s_33_2_1_Adder_3_U.ain_s1 ;
reg [16:0] \sub_33s_33s_33_2_1_U5.top_sub_33s_33s_33_2_1_Adder_3_U.bin_s1 ;
reg \sub_33s_33s_33_2_1_U5.top_sub_33s_33s_33_2_1_Adder_3_U.carry_s1 ;
reg [15:0] \sub_33s_33s_33_2_1_U5.top_sub_33s_33s_33_2_1_Adder_3_U.sum_s1 ;
reg [2:0] \sub_6ns_6s_6_2_1_U14.top_sub_6ns_6s_6_2_1_Adder_10_U.ain_s1 ;
reg [2:0] \sub_6ns_6s_6_2_1_U14.top_sub_6ns_6s_6_2_1_Adder_10_U.bin_s1 ;
reg \sub_6ns_6s_6_2_1_U14.top_sub_6ns_6s_6_2_1_Adder_10_U.carry_s1 ;
reg [2:0] \sub_6ns_6s_6_2_1_U14.top_sub_6ns_6s_6_2_1_Adder_10_U.sum_s1 ;
reg [4:0] \sub_9s_9ns_9_2_1_U3.top_sub_9s_9ns_9_2_1_Adder_2_U.ain_s1 ;
reg [4:0] \sub_9s_9ns_9_2_1_U3.top_sub_9s_9ns_9_2_1_Adder_2_U.bin_s1 ;
reg \sub_9s_9ns_9_2_1_U3.top_sub_9s_9ns_9_2_1_Adder_2_U.carry_s1 ;
reg [3:0] \sub_9s_9ns_9_2_1_U3.top_sub_9s_9ns_9_2_1_Adder_2_U.sum_s1 ;
reg [5:0] sub_ln1497_reg_1423;
reg tmp_13_reg_1373;
reg [1:0] trunc_ln1497_1_reg_1501;
reg [1:0] trunc_ln1497_reg_1496;
reg trunc_ln728_reg_1108;
reg [6:0] trunc_ln790_reg_1157;
reg [24:0] trunc_ln851_1_reg_1271;
reg [24:0] trunc_ln851_2_reg_1342;
reg [5:0] trunc_ln851_3_reg_1224;
reg [24:0] trunc_ln851_reg_1173;
wire _000_;
wire [31:0] _001_;
wire [4:0] _002_;
wire [8:0] _003_;
wire [31:0] _004_;
wire [4:0] _005_;
wire [16:0] _006_;
wire [1:0] _007_;
wire [27:0] _008_;
wire _009_;
wire _010_;
wire _011_;
wire _012_;
wire _013_;
wire _014_;
wire _015_;
wire [3:0] _016_;
wire [16:0] _017_;
wire [1:0] _018_;
wire [3:0] _019_;
wire [7:0] _020_;
wire [25:0] _021_;
wire _022_;
wire _023_;
wire _024_;
wire _025_;
wire _026_;
wire _027_;
wire _028_;
wire [7:0] _029_;
wire [35:0] _030_;
wire [1:0] _031_;
wire [1:0] _032_;
wire [2:0] _033_;
wire [4:0] _034_;
wire [4:0] _035_;
wire [15:0] _036_;
wire [8:0] _037_;
wire [32:0] _038_;
wire [1:0] _039_;
wire [1:0] _040_;
wire [8:0] _041_;
wire [33:0] _042_;
wire [31:0] _043_;
wire [31:0] _044_;
wire [2:0] _045_;
wire [7:0] _046_;
wire [7:0] _047_;
wire [4:0] _048_;
wire [7:0] _049_;
wire [2:0] _050_;
wire [1:0] _051_;
wire [4:0] _052_;
wire [2:0] _053_;
wire _054_;
wire [5:0] _055_;
wire _056_;
wire [1:0] _057_;
wire [1:0] _058_;
wire _059_;
wire [6:0] _060_;
wire [24:0] _061_;
wire [24:0] _062_;
wire [5:0] _063_;
wire [24:0] _064_;
wire [1:0] _065_;
wire _066_;
wire _067_;
wire _068_;
wire _069_;
wire _070_;
wire _071_;
wire _072_;
wire _073_;
wire _074_;
wire _075_;
wire _076_;
wire _077_;
wire _078_;
wire _079_;
wire _080_;
wire _081_;
wire [8:0] _082_;
wire [8:0] _083_;
wire _084_;
wire [7:0] _085_;
wire [8:0] _086_;
wire [9:0] _087_;
wire [8:0] _088_;
wire [8:0] _089_;
wire _090_;
wire [7:0] _091_;
wire [8:0] _092_;
wire [9:0] _093_;
wire [14:0] _094_;
wire [14:0] _095_;
wire _096_;
wire [13:0] _097_;
wire [14:0] _098_;
wire [15:0] _099_;
wire _100_;
wire _101_;
wire _102_;
wire _103_;
wire [1:0] _104_;
wire [1:0] _105_;
wire _106_;
wire _107_;
wire _108_;
wire _109_;
wire [1:0] _110_;
wire [1:0] _111_;
wire [15:0] _112_;
wire [15:0] _113_;
wire _114_;
wire [15:0] _115_;
wire [16:0] _116_;
wire [16:0] _117_;
wire [15:0] _118_;
wire [15:0] _119_;
wire _120_;
wire [15:0] _121_;
wire [16:0] _122_;
wire [16:0] _123_;
wire [15:0] _124_;
wire [15:0] _125_;
wire _126_;
wire [15:0] _127_;
wire [16:0] _128_;
wire [16:0] _129_;
wire [16:0] _130_;
wire [16:0] _131_;
wire _132_;
wire [16:0] _133_;
wire [17:0] _134_;
wire [17:0] _135_;
wire [1:0] _136_;
wire [1:0] _137_;
wire _138_;
wire _139_;
wire [1:0] _140_;
wire [2:0] _141_;
wire [2:0] _142_;
wire [2:0] _143_;
wire _144_;
wire [1:0] _145_;
wire [2:0] _146_;
wire [3:0] _147_;
wire [2:0] _148_;
wire [2:0] _149_;
wire _150_;
wire [1:0] _151_;
wire [2:0] _152_;
wire [3:0] _153_;
wire [2:0] _154_;
wire [2:0] _155_;
wire _156_;
wire [1:0] _157_;
wire [2:0] _158_;
wire [3:0] _159_;
wire [3:0] _160_;
wire [3:0] _161_;
wire _162_;
wire [3:0] _163_;
wire [4:0] _164_;
wire [4:0] _165_;
wire [4:0] _166_;
wire [4:0] _167_;
wire _168_;
wire [3:0] _169_;
wire [4:0] _170_;
wire [5:0] _171_;
wire [4:0] _172_;
wire [4:0] _173_;
wire _174_;
wire [3:0] _175_;
wire [4:0] _176_;
wire [5:0] _177_;
wire [31:0] _178_;
wire [31:0] _179_;
wire [31:0] _180_;
wire [31:0] _181_;
wire [31:0] _182_;
wire [31:0] _183_;
wire [31:0] _184_;
wire [31:0] _185_;
wire [31:0] _186_;
wire [31:0] _187_;
wire [31:0] _188_;
wire [31:0] _189_;
wire [31:0] _190_;
wire [31:0] _191_;
wire [31:0] _192_;
wire [31:0] _193_;
wire [31:0] _194_;
wire [31:0] _195_;
wire [31:0] _196_;
wire [31:0] _197_;
wire [31:0] _198_;
wire [31:0] _199_;
wire [31:0] _200_;
wire [31:0] _201_;
wire [31:0] _202_;
wire [31:0] _203_;
wire [31:0] _204_;
wire [31:0] _205_;
wire [31:0] _206_;
wire [31:0] _207_;
wire [31:0] _208_;
wire [3:0] _209_;
wire [35:0] _210_;
wire [35:0] _211_;
wire [35:0] _212_;
wire [35:0] _213_;
wire [35:0] _214_;
wire [31:0] _215_;
wire [31:0] _216_;
wire [31:0] _217_;
wire [31:0] _218_;
wire [31:0] _219_;
wire [31:0] _220_;
wire [31:0] _221_;
wire [31:0] _222_;
wire [31:0] _223_;
wire [31:0] _224_;
wire [31:0] _225_;
wire [31:0] _226_;
wire [31:0] _227_;
wire [31:0] _228_;
wire [31:0] _229_;
wire [31:0] _230_;
wire [31:0] _231_;
wire [31:0] _232_;
wire [31:0] _233_;
wire [31:0] _234_;
wire [31:0] _235_;
wire [31:0] _236_;
wire [31:0] _237_;
wire [31:0] _238_;
wire [31:0] _239_;
wire [31:0] _240_;
wire [31:0] _241_;
wire [31:0] _242_;
wire [31:0] _243_;
wire [31:0] _244_;
wire [7:0] _245_;
wire [7:0] _246_;
wire _247_;
wire [7:0] _248_;
wire [8:0] _249_;
wire [8:0] _250_;
wire [16:0] _251_;
wire [16:0] _252_;
wire _253_;
wire [15:0] _254_;
wire [16:0] _255_;
wire [17:0] _256_;
wire [2:0] _257_;
wire [2:0] _258_;
wire _259_;
wire [2:0] _260_;
wire [3:0] _261_;
wire [3:0] _262_;
wire [4:0] _263_;
wire [4:0] _264_;
wire _265_;
wire [3:0] _266_;
wire [4:0] _267_;
wire [5:0] _268_;
wire _269_;
wire _270_;
wire _271_;
wire _272_;
wire _273_;
wire _274_;
wire _275_;
wire _276_;
wire _277_;
wire _278_;
wire _279_;
wire _280_;
wire _281_;
wire _282_;
wire _283_;
wire _284_;
wire _285_;
wire _286_;
wire _287_;
wire _288_;
wire _289_;
wire _290_;
wire _291_;
wire _292_;
wire _293_;
wire _294_;
wire _295_;
wire _296_;
wire _297_;
wire _298_;
wire Range1_all_ones_fu_352_p2;
wire \add_17s_17ns_17_2_1_U18.ce ;
wire \add_17s_17ns_17_2_1_U18.clk ;
wire [16:0] \add_17s_17ns_17_2_1_U18.din0 ;
wire [16:0] \add_17s_17ns_17_2_1_U18.din1 ;
wire [16:0] \add_17s_17ns_17_2_1_U18.dout ;
wire \add_17s_17ns_17_2_1_U18.reset ;
wire [16:0] \add_17s_17ns_17_2_1_U18.top_add_17s_17ns_17_2_1_Adder_12_U.a ;
wire [16:0] \add_17s_17ns_17_2_1_U18.top_add_17s_17ns_17_2_1_Adder_12_U.ain_s0 ;
wire [16:0] \add_17s_17ns_17_2_1_U18.top_add_17s_17ns_17_2_1_Adder_12_U.b ;
wire [16:0] \add_17s_17ns_17_2_1_U18.top_add_17s_17ns_17_2_1_Adder_12_U.bin_s0 ;
wire \add_17s_17ns_17_2_1_U18.top_add_17s_17ns_17_2_1_Adder_12_U.ce ;
wire \add_17s_17ns_17_2_1_U18.top_add_17s_17ns_17_2_1_Adder_12_U.clk ;
wire \add_17s_17ns_17_2_1_U18.top_add_17s_17ns_17_2_1_Adder_12_U.facout_s1 ;
wire \add_17s_17ns_17_2_1_U18.top_add_17s_17ns_17_2_1_Adder_12_U.facout_s2 ;
wire [7:0] \add_17s_17ns_17_2_1_U18.top_add_17s_17ns_17_2_1_Adder_12_U.fas_s1 ;
wire [8:0] \add_17s_17ns_17_2_1_U18.top_add_17s_17ns_17_2_1_Adder_12_U.fas_s2 ;
wire \add_17s_17ns_17_2_1_U18.top_add_17s_17ns_17_2_1_Adder_12_U.reset ;
wire [16:0] \add_17s_17ns_17_2_1_U18.top_add_17s_17ns_17_2_1_Adder_12_U.s ;
wire [7:0] \add_17s_17ns_17_2_1_U18.top_add_17s_17ns_17_2_1_Adder_12_U.u1.a ;
wire [7:0] \add_17s_17ns_17_2_1_U18.top_add_17s_17ns_17_2_1_Adder_12_U.u1.b ;
wire \add_17s_17ns_17_2_1_U18.top_add_17s_17ns_17_2_1_Adder_12_U.u1.cin ;
wire \add_17s_17ns_17_2_1_U18.top_add_17s_17ns_17_2_1_Adder_12_U.u1.cout ;
wire [7:0] \add_17s_17ns_17_2_1_U18.top_add_17s_17ns_17_2_1_Adder_12_U.u1.s ;
wire [8:0] \add_17s_17ns_17_2_1_U18.top_add_17s_17ns_17_2_1_Adder_12_U.u2.a ;
wire [8:0] \add_17s_17ns_17_2_1_U18.top_add_17s_17ns_17_2_1_Adder_12_U.u2.b ;
wire \add_17s_17ns_17_2_1_U18.top_add_17s_17ns_17_2_1_Adder_12_U.u2.cin ;
wire \add_17s_17ns_17_2_1_U18.top_add_17s_17ns_17_2_1_Adder_12_U.u2.cout ;
wire [8:0] \add_17s_17ns_17_2_1_U18.top_add_17s_17ns_17_2_1_Adder_12_U.u2.s ;
wire \add_17s_17s_17_2_1_U15.ce ;
wire \add_17s_17s_17_2_1_U15.clk ;
wire [16:0] \add_17s_17s_17_2_1_U15.din0 ;
wire [16:0] \add_17s_17s_17_2_1_U15.din1 ;
wire [16:0] \add_17s_17s_17_2_1_U15.dout ;
wire \add_17s_17s_17_2_1_U15.reset ;
wire [16:0] \add_17s_17s_17_2_1_U15.top_add_17s_17s_17_2_1_Adder_11_U.a ;
wire [16:0] \add_17s_17s_17_2_1_U15.top_add_17s_17s_17_2_1_Adder_11_U.ain_s0 ;
wire [16:0] \add_17s_17s_17_2_1_U15.top_add_17s_17s_17_2_1_Adder_11_U.b ;
wire [16:0] \add_17s_17s_17_2_1_U15.top_add_17s_17s_17_2_1_Adder_11_U.bin_s0 ;
wire \add_17s_17s_17_2_1_U15.top_add_17s_17s_17_2_1_Adder_11_U.ce ;
wire \add_17s_17s_17_2_1_U15.top_add_17s_17s_17_2_1_Adder_11_U.clk ;
wire \add_17s_17s_17_2_1_U15.top_add_17s_17s_17_2_1_Adder_11_U.facout_s1 ;
wire \add_17s_17s_17_2_1_U15.top_add_17s_17s_17_2_1_Adder_11_U.facout_s2 ;
wire [7:0] \add_17s_17s_17_2_1_U15.top_add_17s_17s_17_2_1_Adder_11_U.fas_s1 ;
wire [8:0] \add_17s_17s_17_2_1_U15.top_add_17s_17s_17_2_1_Adder_11_U.fas_s2 ;
wire \add_17s_17s_17_2_1_U15.top_add_17s_17s_17_2_1_Adder_11_U.reset ;
wire [16:0] \add_17s_17s_17_2_1_U15.top_add_17s_17s_17_2_1_Adder_11_U.s ;
wire [7:0] \add_17s_17s_17_2_1_U15.top_add_17s_17s_17_2_1_Adder_11_U.u1.a ;
wire [7:0] \add_17s_17s_17_2_1_U15.top_add_17s_17s_17_2_1_Adder_11_U.u1.b ;
wire \add_17s_17s_17_2_1_U15.top_add_17s_17s_17_2_1_Adder_11_U.u1.cin ;
wire \add_17s_17s_17_2_1_U15.top_add_17s_17s_17_2_1_Adder_11_U.u1.cout ;
wire [7:0] \add_17s_17s_17_2_1_U15.top_add_17s_17s_17_2_1_Adder_11_U.u1.s ;
wire [8:0] \add_17s_17s_17_2_1_U15.top_add_17s_17s_17_2_1_Adder_11_U.u2.a ;
wire [8:0] \add_17s_17s_17_2_1_U15.top_add_17s_17s_17_2_1_Adder_11_U.u2.b ;
wire \add_17s_17s_17_2_1_U15.top_add_17s_17s_17_2_1_Adder_11_U.u2.cin ;
wire \add_17s_17s_17_2_1_U15.top_add_17s_17s_17_2_1_Adder_11_U.u2.cout ;
wire [8:0] \add_17s_17s_17_2_1_U15.top_add_17s_17s_17_2_1_Adder_11_U.u2.s ;
wire \add_29s_29ns_29_2_1_U12.ce ;
wire \add_29s_29ns_29_2_1_U12.clk ;
wire [28:0] \add_29s_29ns_29_2_1_U12.din0 ;
wire [28:0] \add_29s_29ns_29_2_1_U12.din1 ;
wire [28:0] \add_29s_29ns_29_2_1_U12.dout ;
wire \add_29s_29ns_29_2_1_U12.reset ;
wire [28:0] \add_29s_29ns_29_2_1_U12.top_add_29s_29ns_29_2_1_Adder_9_U.a ;
wire [28:0] \add_29s_29ns_29_2_1_U12.top_add_29s_29ns_29_2_1_Adder_9_U.ain_s0 ;
wire [28:0] \add_29s_29ns_29_2_1_U12.top_add_29s_29ns_29_2_1_Adder_9_U.b ;
wire [28:0] \add_29s_29ns_29_2_1_U12.top_add_29s_29ns_29_2_1_Adder_9_U.bin_s0 ;
wire \add_29s_29ns_29_2_1_U12.top_add_29s_29ns_29_2_1_Adder_9_U.ce ;
wire \add_29s_29ns_29_2_1_U12.top_add_29s_29ns_29_2_1_Adder_9_U.clk ;
wire \add_29s_29ns_29_2_1_U12.top_add_29s_29ns_29_2_1_Adder_9_U.facout_s1 ;
wire \add_29s_29ns_29_2_1_U12.top_add_29s_29ns_29_2_1_Adder_9_U.facout_s2 ;
wire [13:0] \add_29s_29ns_29_2_1_U12.top_add_29s_29ns_29_2_1_Adder_9_U.fas_s1 ;
wire [14:0] \add_29s_29ns_29_2_1_U12.top_add_29s_29ns_29_2_1_Adder_9_U.fas_s2 ;
wire \add_29s_29ns_29_2_1_U12.top_add_29s_29ns_29_2_1_Adder_9_U.reset ;
wire [28:0] \add_29s_29ns_29_2_1_U12.top_add_29s_29ns_29_2_1_Adder_9_U.s ;
wire [13:0] \add_29s_29ns_29_2_1_U12.top_add_29s_29ns_29_2_1_Adder_9_U.u1.a ;
wire [13:0] \add_29s_29ns_29_2_1_U12.top_add_29s_29ns_29_2_1_Adder_9_U.u1.b ;
wire \add_29s_29ns_29_2_1_U12.top_add_29s_29ns_29_2_1_Adder_9_U.u1.cin ;
wire \add_29s_29ns_29_2_1_U12.top_add_29s_29ns_29_2_1_Adder_9_U.u1.cout ;
wire [13:0] \add_29s_29ns_29_2_1_U12.top_add_29s_29ns_29_2_1_Adder_9_U.u1.s ;
wire [14:0] \add_29s_29ns_29_2_1_U12.top_add_29s_29ns_29_2_1_Adder_9_U.u2.a ;
wire [14:0] \add_29s_29ns_29_2_1_U12.top_add_29s_29ns_29_2_1_Adder_9_U.u2.b ;
wire \add_29s_29ns_29_2_1_U12.top_add_29s_29ns_29_2_1_Adder_9_U.u2.cin ;
wire \add_29s_29ns_29_2_1_U12.top_add_29s_29ns_29_2_1_Adder_9_U.u2.cout ;
wire [14:0] \add_29s_29ns_29_2_1_U12.top_add_29s_29ns_29_2_1_Adder_9_U.u2.s ;
wire \add_2ns_2ns_2_2_1_U1.ce ;
wire \add_2ns_2ns_2_2_1_U1.clk ;
wire [1:0] \add_2ns_2ns_2_2_1_U1.din0 ;
wire [1:0] \add_2ns_2ns_2_2_1_U1.din1 ;
wire [1:0] \add_2ns_2ns_2_2_1_U1.dout ;
wire \add_2ns_2ns_2_2_1_U1.reset ;
wire [1:0] \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.a ;
wire [1:0] \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.ain_s0 ;
wire [1:0] \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.b ;
wire [1:0] \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.bin_s0 ;
wire \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.ce ;
wire \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.clk ;
wire \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.facout_s1 ;
wire \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.facout_s2 ;
wire \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.fas_s1 ;
wire \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.fas_s2 ;
wire \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.reset ;
wire [1:0] \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.s ;
wire \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.u1.a ;
wire \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.u1.b ;
wire \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.u1.cin ;
wire \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.u1.cout ;
wire \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.u1.s ;
wire \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.u2.a ;
wire \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.u2.b ;
wire \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.u2.cin ;
wire \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.u2.cout ;
wire \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.u2.s ;
wire \add_2ns_2ns_2_2_1_U11.ce ;
wire \add_2ns_2ns_2_2_1_U11.clk ;
wire [1:0] \add_2ns_2ns_2_2_1_U11.din0 ;
wire [1:0] \add_2ns_2ns_2_2_1_U11.din1 ;
wire [1:0] \add_2ns_2ns_2_2_1_U11.dout ;
wire \add_2ns_2ns_2_2_1_U11.reset ;
wire [1:0] \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_0_U.a ;
wire [1:0] \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_0_U.ain_s0 ;
wire [1:0] \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_0_U.b ;
wire [1:0] \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_0_U.bin_s0 ;
wire \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_0_U.ce ;
wire \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_0_U.clk ;
wire \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_0_U.facout_s1 ;
wire \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_0_U.facout_s2 ;
wire \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_0_U.fas_s1 ;
wire \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_0_U.fas_s2 ;
wire \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_0_U.reset ;
wire [1:0] \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_0_U.s ;
wire \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_0_U.u1.a ;
wire \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_0_U.u1.b ;
wire \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_0_U.u1.cin ;
wire \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_0_U.u1.cout ;
wire \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_0_U.u1.s ;
wire \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_0_U.u2.a ;
wire \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_0_U.u2.b ;
wire \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_0_U.u2.cin ;
wire \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_0_U.u2.cout ;
wire \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_0_U.u2.s ;
wire \add_32ns_32ns_32_2_1_U20.ce ;
wire \add_32ns_32ns_32_2_1_U20.clk ;
wire [31:0] \add_32ns_32ns_32_2_1_U20.din0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U20.din1 ;
wire [31:0] \add_32ns_32ns_32_2_1_U20.dout ;
wire \add_32ns_32ns_32_2_1_U20.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_14_U.a ;
wire [31:0] \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_14_U.ain_s0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_14_U.b ;
wire [31:0] \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_14_U.bin_s0 ;
wire \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_14_U.ce ;
wire \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_14_U.clk ;
wire \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_14_U.facout_s1 ;
wire \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_14_U.facout_s2 ;
wire [15:0] \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_14_U.fas_s1 ;
wire [15:0] \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_14_U.fas_s2 ;
wire \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_14_U.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_14_U.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_14_U.u1.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_14_U.u1.b ;
wire \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_14_U.u1.cin ;
wire \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_14_U.u1.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_14_U.u1.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_14_U.u2.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_14_U.u2.b ;
wire \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_14_U.u2.cin ;
wire \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_14_U.u2.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_14_U.u2.s ;
wire \add_32ns_32ns_32_2_1_U21.ce ;
wire \add_32ns_32ns_32_2_1_U21.clk ;
wire [31:0] \add_32ns_32ns_32_2_1_U21.din0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U21.din1 ;
wire [31:0] \add_32ns_32ns_32_2_1_U21.dout ;
wire \add_32ns_32ns_32_2_1_U21.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_14_U.a ;
wire [31:0] \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_14_U.ain_s0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_14_U.b ;
wire [31:0] \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_14_U.bin_s0 ;
wire \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_14_U.ce ;
wire \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_14_U.clk ;
wire \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_14_U.facout_s1 ;
wire \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_14_U.facout_s2 ;
wire [15:0] \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_14_U.fas_s1 ;
wire [15:0] \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_14_U.fas_s2 ;
wire \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_14_U.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_14_U.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_14_U.u1.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_14_U.u1.b ;
wire \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_14_U.u1.cin ;
wire \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_14_U.u1.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_14_U.u1.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_14_U.u2.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_14_U.u2.b ;
wire \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_14_U.u2.cin ;
wire \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_14_U.u2.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_14_U.u2.s ;
wire \add_32s_32ns_32_2_1_U23.ce ;
wire \add_32s_32ns_32_2_1_U23.clk ;
wire [31:0] \add_32s_32ns_32_2_1_U23.din0 ;
wire [31:0] \add_32s_32ns_32_2_1_U23.din1 ;
wire [31:0] \add_32s_32ns_32_2_1_U23.dout ;
wire \add_32s_32ns_32_2_1_U23.reset ;
wire [31:0] \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_16_U.a ;
wire [31:0] \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_16_U.ain_s0 ;
wire [31:0] \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_16_U.b ;
wire [31:0] \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_16_U.bin_s0 ;
wire \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_16_U.ce ;
wire \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_16_U.clk ;
wire \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_16_U.facout_s1 ;
wire \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_16_U.facout_s2 ;
wire [15:0] \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_16_U.fas_s1 ;
wire [15:0] \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_16_U.fas_s2 ;
wire \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_16_U.reset ;
wire [31:0] \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_16_U.s ;
wire [15:0] \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_16_U.u1.a ;
wire [15:0] \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_16_U.u1.b ;
wire \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_16_U.u1.cin ;
wire \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_16_U.u1.cout ;
wire [15:0] \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_16_U.u1.s ;
wire [15:0] \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_16_U.u2.a ;
wire [15:0] \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_16_U.u2.b ;
wire \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_16_U.u2.cin ;
wire \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_16_U.u2.cout ;
wire [15:0] \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_16_U.u2.s ;
wire \add_34s_34s_34_2_1_U19.ce ;
wire \add_34s_34s_34_2_1_U19.clk ;
wire [33:0] \add_34s_34s_34_2_1_U19.din0 ;
wire [33:0] \add_34s_34s_34_2_1_U19.din1 ;
wire [33:0] \add_34s_34s_34_2_1_U19.dout ;
wire \add_34s_34s_34_2_1_U19.reset ;
wire [33:0] \add_34s_34s_34_2_1_U19.top_add_34s_34s_34_2_1_Adder_13_U.a ;
wire [33:0] \add_34s_34s_34_2_1_U19.top_add_34s_34s_34_2_1_Adder_13_U.ain_s0 ;
wire [33:0] \add_34s_34s_34_2_1_U19.top_add_34s_34s_34_2_1_Adder_13_U.b ;
wire [33:0] \add_34s_34s_34_2_1_U19.top_add_34s_34s_34_2_1_Adder_13_U.bin_s0 ;
wire \add_34s_34s_34_2_1_U19.top_add_34s_34s_34_2_1_Adder_13_U.ce ;
wire \add_34s_34s_34_2_1_U19.top_add_34s_34s_34_2_1_Adder_13_U.clk ;
wire \add_34s_34s_34_2_1_U19.top_add_34s_34s_34_2_1_Adder_13_U.facout_s1 ;
wire \add_34s_34s_34_2_1_U19.top_add_34s_34s_34_2_1_Adder_13_U.facout_s2 ;
wire [16:0] \add_34s_34s_34_2_1_U19.top_add_34s_34s_34_2_1_Adder_13_U.fas_s1 ;
wire [16:0] \add_34s_34s_34_2_1_U19.top_add_34s_34s_34_2_1_Adder_13_U.fas_s2 ;
wire \add_34s_34s_34_2_1_U19.top_add_34s_34s_34_2_1_Adder_13_U.reset ;
wire [33:0] \add_34s_34s_34_2_1_U19.top_add_34s_34s_34_2_1_Adder_13_U.s ;
wire [16:0] \add_34s_34s_34_2_1_U19.top_add_34s_34s_34_2_1_Adder_13_U.u1.a ;
wire [16:0] \add_34s_34s_34_2_1_U19.top_add_34s_34s_34_2_1_Adder_13_U.u1.b ;
wire \add_34s_34s_34_2_1_U19.top_add_34s_34s_34_2_1_Adder_13_U.u1.cin ;
wire \add_34s_34s_34_2_1_U19.top_add_34s_34s_34_2_1_Adder_13_U.u1.cout ;
wire [16:0] \add_34s_34s_34_2_1_U19.top_add_34s_34s_34_2_1_Adder_13_U.u1.s ;
wire [16:0] \add_34s_34s_34_2_1_U19.top_add_34s_34s_34_2_1_Adder_13_U.u2.a ;
wire [16:0] \add_34s_34s_34_2_1_U19.top_add_34s_34s_34_2_1_Adder_13_U.u2.b ;
wire \add_34s_34s_34_2_1_U19.top_add_34s_34s_34_2_1_Adder_13_U.u2.cin ;
wire \add_34s_34s_34_2_1_U19.top_add_34s_34s_34_2_1_Adder_13_U.u2.cout ;
wire [16:0] \add_34s_34s_34_2_1_U19.top_add_34s_34s_34_2_1_Adder_13_U.u2.s ;
wire \add_3ns_3ns_3_2_1_U8.ce ;
wire \add_3ns_3ns_3_2_1_U8.clk ;
wire [2:0] \add_3ns_3ns_3_2_1_U8.din0 ;
wire [2:0] \add_3ns_3ns_3_2_1_U8.din1 ;
wire [2:0] \add_3ns_3ns_3_2_1_U8.dout ;
wire \add_3ns_3ns_3_2_1_U8.reset ;
wire [2:0] \add_3ns_3ns_3_2_1_U8.top_add_3ns_3ns_3_2_1_Adder_6_U.a ;
wire [2:0] \add_3ns_3ns_3_2_1_U8.top_add_3ns_3ns_3_2_1_Adder_6_U.ain_s0 ;
wire [2:0] \add_3ns_3ns_3_2_1_U8.top_add_3ns_3ns_3_2_1_Adder_6_U.b ;
wire [2:0] \add_3ns_3ns_3_2_1_U8.top_add_3ns_3ns_3_2_1_Adder_6_U.bin_s0 ;
wire \add_3ns_3ns_3_2_1_U8.top_add_3ns_3ns_3_2_1_Adder_6_U.ce ;
wire \add_3ns_3ns_3_2_1_U8.top_add_3ns_3ns_3_2_1_Adder_6_U.clk ;
wire \add_3ns_3ns_3_2_1_U8.top_add_3ns_3ns_3_2_1_Adder_6_U.facout_s1 ;
wire \add_3ns_3ns_3_2_1_U8.top_add_3ns_3ns_3_2_1_Adder_6_U.facout_s2 ;
wire \add_3ns_3ns_3_2_1_U8.top_add_3ns_3ns_3_2_1_Adder_6_U.fas_s1 ;
wire [1:0] \add_3ns_3ns_3_2_1_U8.top_add_3ns_3ns_3_2_1_Adder_6_U.fas_s2 ;
wire \add_3ns_3ns_3_2_1_U8.top_add_3ns_3ns_3_2_1_Adder_6_U.reset ;
wire [2:0] \add_3ns_3ns_3_2_1_U8.top_add_3ns_3ns_3_2_1_Adder_6_U.s ;
wire \add_3ns_3ns_3_2_1_U8.top_add_3ns_3ns_3_2_1_Adder_6_U.u1.a ;
wire \add_3ns_3ns_3_2_1_U8.top_add_3ns_3ns_3_2_1_Adder_6_U.u1.b ;
wire \add_3ns_3ns_3_2_1_U8.top_add_3ns_3ns_3_2_1_Adder_6_U.u1.cin ;
wire \add_3ns_3ns_3_2_1_U8.top_add_3ns_3ns_3_2_1_Adder_6_U.u1.cout ;
wire \add_3ns_3ns_3_2_1_U8.top_add_3ns_3ns_3_2_1_Adder_6_U.u1.s ;
wire [1:0] \add_3ns_3ns_3_2_1_U8.top_add_3ns_3ns_3_2_1_Adder_6_U.u2.a ;
wire [1:0] \add_3ns_3ns_3_2_1_U8.top_add_3ns_3ns_3_2_1_Adder_6_U.u2.b ;
wire \add_3ns_3ns_3_2_1_U8.top_add_3ns_3ns_3_2_1_Adder_6_U.u2.cin ;
wire \add_3ns_3ns_3_2_1_U8.top_add_3ns_3ns_3_2_1_Adder_6_U.u2.cout ;
wire [1:0] \add_3ns_3ns_3_2_1_U8.top_add_3ns_3ns_3_2_1_Adder_6_U.u2.s ;
wire \add_5ns_5ns_5_2_1_U9.ce ;
wire \add_5ns_5ns_5_2_1_U9.clk ;
wire [4:0] \add_5ns_5ns_5_2_1_U9.din0 ;
wire [4:0] \add_5ns_5ns_5_2_1_U9.din1 ;
wire [4:0] \add_5ns_5ns_5_2_1_U9.dout ;
wire \add_5ns_5ns_5_2_1_U9.reset ;
wire [4:0] \add_5ns_5ns_5_2_1_U9.top_add_5ns_5ns_5_2_1_Adder_7_U.a ;
wire [4:0] \add_5ns_5ns_5_2_1_U9.top_add_5ns_5ns_5_2_1_Adder_7_U.ain_s0 ;
wire [4:0] \add_5ns_5ns_5_2_1_U9.top_add_5ns_5ns_5_2_1_Adder_7_U.b ;
wire [4:0] \add_5ns_5ns_5_2_1_U9.top_add_5ns_5ns_5_2_1_Adder_7_U.bin_s0 ;
wire \add_5ns_5ns_5_2_1_U9.top_add_5ns_5ns_5_2_1_Adder_7_U.ce ;
wire \add_5ns_5ns_5_2_1_U9.top_add_5ns_5ns_5_2_1_Adder_7_U.clk ;
wire \add_5ns_5ns_5_2_1_U9.top_add_5ns_5ns_5_2_1_Adder_7_U.facout_s1 ;
wire \add_5ns_5ns_5_2_1_U9.top_add_5ns_5ns_5_2_1_Adder_7_U.facout_s2 ;
wire [1:0] \add_5ns_5ns_5_2_1_U9.top_add_5ns_5ns_5_2_1_Adder_7_U.fas_s1 ;
wire [2:0] \add_5ns_5ns_5_2_1_U9.top_add_5ns_5ns_5_2_1_Adder_7_U.fas_s2 ;
wire \add_5ns_5ns_5_2_1_U9.top_add_5ns_5ns_5_2_1_Adder_7_U.reset ;
wire [4:0] \add_5ns_5ns_5_2_1_U9.top_add_5ns_5ns_5_2_1_Adder_7_U.s ;
wire [1:0] \add_5ns_5ns_5_2_1_U9.top_add_5ns_5ns_5_2_1_Adder_7_U.u1.a ;
wire [1:0] \add_5ns_5ns_5_2_1_U9.top_add_5ns_5ns_5_2_1_Adder_7_U.u1.b ;
wire \add_5ns_5ns_5_2_1_U9.top_add_5ns_5ns_5_2_1_Adder_7_U.u1.cin ;
wire \add_5ns_5ns_5_2_1_U9.top_add_5ns_5ns_5_2_1_Adder_7_U.u1.cout ;
wire [1:0] \add_5ns_5ns_5_2_1_U9.top_add_5ns_5ns_5_2_1_Adder_7_U.u1.s ;
wire [2:0] \add_5ns_5ns_5_2_1_U9.top_add_5ns_5ns_5_2_1_Adder_7_U.u2.a ;
wire [2:0] \add_5ns_5ns_5_2_1_U9.top_add_5ns_5ns_5_2_1_Adder_7_U.u2.b ;
wire \add_5ns_5ns_5_2_1_U9.top_add_5ns_5ns_5_2_1_Adder_7_U.u2.cin ;
wire \add_5ns_5ns_5_2_1_U9.top_add_5ns_5ns_5_2_1_Adder_7_U.u2.cout ;
wire [2:0] \add_5ns_5ns_5_2_1_U9.top_add_5ns_5ns_5_2_1_Adder_7_U.u2.s ;
wire \add_5s_5ns_5_2_1_U10.ce ;
wire \add_5s_5ns_5_2_1_U10.clk ;
wire [4:0] \add_5s_5ns_5_2_1_U10.din0 ;
wire [4:0] \add_5s_5ns_5_2_1_U10.din1 ;
wire [4:0] \add_5s_5ns_5_2_1_U10.dout ;
wire \add_5s_5ns_5_2_1_U10.reset ;
wire [4:0] \add_5s_5ns_5_2_1_U10.top_add_5s_5ns_5_2_1_Adder_8_U.a ;
wire [4:0] \add_5s_5ns_5_2_1_U10.top_add_5s_5ns_5_2_1_Adder_8_U.ain_s0 ;
wire [4:0] \add_5s_5ns_5_2_1_U10.top_add_5s_5ns_5_2_1_Adder_8_U.b ;
wire [4:0] \add_5s_5ns_5_2_1_U10.top_add_5s_5ns_5_2_1_Adder_8_U.bin_s0 ;
wire \add_5s_5ns_5_2_1_U10.top_add_5s_5ns_5_2_1_Adder_8_U.ce ;
wire \add_5s_5ns_5_2_1_U10.top_add_5s_5ns_5_2_1_Adder_8_U.clk ;
wire \add_5s_5ns_5_2_1_U10.top_add_5s_5ns_5_2_1_Adder_8_U.facout_s1 ;
wire \add_5s_5ns_5_2_1_U10.top_add_5s_5ns_5_2_1_Adder_8_U.facout_s2 ;
wire [1:0] \add_5s_5ns_5_2_1_U10.top_add_5s_5ns_5_2_1_Adder_8_U.fas_s1 ;
wire [2:0] \add_5s_5ns_5_2_1_U10.top_add_5s_5ns_5_2_1_Adder_8_U.fas_s2 ;
wire \add_5s_5ns_5_2_1_U10.top_add_5s_5ns_5_2_1_Adder_8_U.reset ;
wire [4:0] \add_5s_5ns_5_2_1_U10.top_add_5s_5ns_5_2_1_Adder_8_U.s ;
wire [1:0] \add_5s_5ns_5_2_1_U10.top_add_5s_5ns_5_2_1_Adder_8_U.u1.a ;
wire [1:0] \add_5s_5ns_5_2_1_U10.top_add_5s_5ns_5_2_1_Adder_8_U.u1.b ;
wire \add_5s_5ns_5_2_1_U10.top_add_5s_5ns_5_2_1_Adder_8_U.u1.cin ;
wire \add_5s_5ns_5_2_1_U10.top_add_5s_5ns_5_2_1_Adder_8_U.u1.cout ;
wire [1:0] \add_5s_5ns_5_2_1_U10.top_add_5s_5ns_5_2_1_Adder_8_U.u1.s ;
wire [2:0] \add_5s_5ns_5_2_1_U10.top_add_5s_5ns_5_2_1_Adder_8_U.u2.a ;
wire [2:0] \add_5s_5ns_5_2_1_U10.top_add_5s_5ns_5_2_1_Adder_8_U.u2.b ;
wire \add_5s_5ns_5_2_1_U10.top_add_5s_5ns_5_2_1_Adder_8_U.u2.cin ;
wire \add_5s_5ns_5_2_1_U10.top_add_5s_5ns_5_2_1_Adder_8_U.u2.cout ;
wire [2:0] \add_5s_5ns_5_2_1_U10.top_add_5s_5ns_5_2_1_Adder_8_U.u2.s ;
wire \add_5s_5s_5_2_1_U22.ce ;
wire \add_5s_5s_5_2_1_U22.clk ;
wire [4:0] \add_5s_5s_5_2_1_U22.din0 ;
wire [4:0] \add_5s_5s_5_2_1_U22.din1 ;
wire [4:0] \add_5s_5s_5_2_1_U22.dout ;
wire \add_5s_5s_5_2_1_U22.reset ;
wire [4:0] \add_5s_5s_5_2_1_U22.top_add_5s_5s_5_2_1_Adder_15_U.a ;
wire [4:0] \add_5s_5s_5_2_1_U22.top_add_5s_5s_5_2_1_Adder_15_U.ain_s0 ;
wire [4:0] \add_5s_5s_5_2_1_U22.top_add_5s_5s_5_2_1_Adder_15_U.b ;
wire [4:0] \add_5s_5s_5_2_1_U22.top_add_5s_5s_5_2_1_Adder_15_U.bin_s0 ;
wire \add_5s_5s_5_2_1_U22.top_add_5s_5s_5_2_1_Adder_15_U.ce ;
wire \add_5s_5s_5_2_1_U22.top_add_5s_5s_5_2_1_Adder_15_U.clk ;
wire \add_5s_5s_5_2_1_U22.top_add_5s_5s_5_2_1_Adder_15_U.facout_s1 ;
wire \add_5s_5s_5_2_1_U22.top_add_5s_5s_5_2_1_Adder_15_U.facout_s2 ;
wire [1:0] \add_5s_5s_5_2_1_U22.top_add_5s_5s_5_2_1_Adder_15_U.fas_s1 ;
wire [2:0] \add_5s_5s_5_2_1_U22.top_add_5s_5s_5_2_1_Adder_15_U.fas_s2 ;
wire \add_5s_5s_5_2_1_U22.top_add_5s_5s_5_2_1_Adder_15_U.reset ;
wire [4:0] \add_5s_5s_5_2_1_U22.top_add_5s_5s_5_2_1_Adder_15_U.s ;
wire [1:0] \add_5s_5s_5_2_1_U22.top_add_5s_5s_5_2_1_Adder_15_U.u1.a ;
wire [1:0] \add_5s_5s_5_2_1_U22.top_add_5s_5s_5_2_1_Adder_15_U.u1.b ;
wire \add_5s_5s_5_2_1_U22.top_add_5s_5s_5_2_1_Adder_15_U.u1.cin ;
wire \add_5s_5s_5_2_1_U22.top_add_5s_5s_5_2_1_Adder_15_U.u1.cout ;
wire [1:0] \add_5s_5s_5_2_1_U22.top_add_5s_5s_5_2_1_Adder_15_U.u1.s ;
wire [2:0] \add_5s_5s_5_2_1_U22.top_add_5s_5s_5_2_1_Adder_15_U.u2.a ;
wire [2:0] \add_5s_5s_5_2_1_U22.top_add_5s_5s_5_2_1_Adder_15_U.u2.b ;
wire \add_5s_5s_5_2_1_U22.top_add_5s_5s_5_2_1_Adder_15_U.u2.cin ;
wire \add_5s_5s_5_2_1_U22.top_add_5s_5s_5_2_1_Adder_15_U.u2.cout ;
wire [2:0] \add_5s_5s_5_2_1_U22.top_add_5s_5s_5_2_1_Adder_15_U.u2.s ;
wire \add_8ns_8ns_8_2_1_U7.ce ;
wire \add_8ns_8ns_8_2_1_U7.clk ;
wire [7:0] \add_8ns_8ns_8_2_1_U7.din0 ;
wire [7:0] \add_8ns_8ns_8_2_1_U7.din1 ;
wire [7:0] \add_8ns_8ns_8_2_1_U7.dout ;
wire \add_8ns_8ns_8_2_1_U7.reset ;
wire [7:0] \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_5_U.a ;
wire [7:0] \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_5_U.ain_s0 ;
wire [7:0] \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_5_U.b ;
wire [7:0] \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_5_U.bin_s0 ;
wire \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_5_U.ce ;
wire \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_5_U.clk ;
wire \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_5_U.facout_s1 ;
wire \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_5_U.facout_s2 ;
wire [3:0] \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_5_U.fas_s1 ;
wire [3:0] \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_5_U.fas_s2 ;
wire \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_5_U.reset ;
wire [7:0] \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_5_U.s ;
wire [3:0] \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_5_U.u1.a ;
wire [3:0] \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_5_U.u1.b ;
wire \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_5_U.u1.cin ;
wire \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_5_U.u1.cout ;
wire [3:0] \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_5_U.u1.s ;
wire [3:0] \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_5_U.u2.a ;
wire [3:0] \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_5_U.u2.b ;
wire \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_5_U.u2.cin ;
wire \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_5_U.u2.cout ;
wire [3:0] \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_5_U.u2.s ;
wire \add_9s_9s_9_2_1_U13.ce ;
wire \add_9s_9s_9_2_1_U13.clk ;
wire [8:0] \add_9s_9s_9_2_1_U13.din0 ;
wire [8:0] \add_9s_9s_9_2_1_U13.din1 ;
wire [8:0] \add_9s_9s_9_2_1_U13.dout ;
wire \add_9s_9s_9_2_1_U13.reset ;
wire [8:0] \add_9s_9s_9_2_1_U13.top_add_9s_9s_9_2_1_Adder_4_U.a ;
wire [8:0] \add_9s_9s_9_2_1_U13.top_add_9s_9s_9_2_1_Adder_4_U.ain_s0 ;
wire [8:0] \add_9s_9s_9_2_1_U13.top_add_9s_9s_9_2_1_Adder_4_U.b ;
wire [8:0] \add_9s_9s_9_2_1_U13.top_add_9s_9s_9_2_1_Adder_4_U.bin_s0 ;
wire \add_9s_9s_9_2_1_U13.top_add_9s_9s_9_2_1_Adder_4_U.ce ;
wire \add_9s_9s_9_2_1_U13.top_add_9s_9s_9_2_1_Adder_4_U.clk ;
wire \add_9s_9s_9_2_1_U13.top_add_9s_9s_9_2_1_Adder_4_U.facout_s1 ;
wire \add_9s_9s_9_2_1_U13.top_add_9s_9s_9_2_1_Adder_4_U.facout_s2 ;
wire [3:0] \add_9s_9s_9_2_1_U13.top_add_9s_9s_9_2_1_Adder_4_U.fas_s1 ;
wire [4:0] \add_9s_9s_9_2_1_U13.top_add_9s_9s_9_2_1_Adder_4_U.fas_s2 ;
wire \add_9s_9s_9_2_1_U13.top_add_9s_9s_9_2_1_Adder_4_U.reset ;
wire [8:0] \add_9s_9s_9_2_1_U13.top_add_9s_9s_9_2_1_Adder_4_U.s ;
wire [3:0] \add_9s_9s_9_2_1_U13.top_add_9s_9s_9_2_1_Adder_4_U.u1.a ;
wire [3:0] \add_9s_9s_9_2_1_U13.top_add_9s_9s_9_2_1_Adder_4_U.u1.b ;
wire \add_9s_9s_9_2_1_U13.top_add_9s_9s_9_2_1_Adder_4_U.u1.cin ;
wire \add_9s_9s_9_2_1_U13.top_add_9s_9s_9_2_1_Adder_4_U.u1.cout ;
wire [3:0] \add_9s_9s_9_2_1_U13.top_add_9s_9s_9_2_1_Adder_4_U.u1.s ;
wire [4:0] \add_9s_9s_9_2_1_U13.top_add_9s_9s_9_2_1_Adder_4_U.u2.a ;
wire [4:0] \add_9s_9s_9_2_1_U13.top_add_9s_9s_9_2_1_Adder_4_U.u2.b ;
wire \add_9s_9s_9_2_1_U13.top_add_9s_9s_9_2_1_Adder_4_U.u2.cin ;
wire \add_9s_9s_9_2_1_U13.top_add_9s_9s_9_2_1_Adder_4_U.u2.cout ;
wire [4:0] \add_9s_9s_9_2_1_U13.top_add_9s_9s_9_2_1_Adder_4_U.u2.s ;
wire \add_9s_9s_9_2_1_U6.ce ;
wire \add_9s_9s_9_2_1_U6.clk ;
wire [8:0] \add_9s_9s_9_2_1_U6.din0 ;
wire [8:0] \add_9s_9s_9_2_1_U6.din1 ;
wire [8:0] \add_9s_9s_9_2_1_U6.dout ;
wire \add_9s_9s_9_2_1_U6.reset ;
wire [8:0] \add_9s_9s_9_2_1_U6.top_add_9s_9s_9_2_1_Adder_4_U.a ;
wire [8:0] \add_9s_9s_9_2_1_U6.top_add_9s_9s_9_2_1_Adder_4_U.ain_s0 ;
wire [8:0] \add_9s_9s_9_2_1_U6.top_add_9s_9s_9_2_1_Adder_4_U.b ;
wire [8:0] \add_9s_9s_9_2_1_U6.top_add_9s_9s_9_2_1_Adder_4_U.bin_s0 ;
wire \add_9s_9s_9_2_1_U6.top_add_9s_9s_9_2_1_Adder_4_U.ce ;
wire \add_9s_9s_9_2_1_U6.top_add_9s_9s_9_2_1_Adder_4_U.clk ;
wire \add_9s_9s_9_2_1_U6.top_add_9s_9s_9_2_1_Adder_4_U.facout_s1 ;
wire \add_9s_9s_9_2_1_U6.top_add_9s_9s_9_2_1_Adder_4_U.facout_s2 ;
wire [3:0] \add_9s_9s_9_2_1_U6.top_add_9s_9s_9_2_1_Adder_4_U.fas_s1 ;
wire [4:0] \add_9s_9s_9_2_1_U6.top_add_9s_9s_9_2_1_Adder_4_U.fas_s2 ;
wire \add_9s_9s_9_2_1_U6.top_add_9s_9s_9_2_1_Adder_4_U.reset ;
wire [8:0] \add_9s_9s_9_2_1_U6.top_add_9s_9s_9_2_1_Adder_4_U.s ;
wire [3:0] \add_9s_9s_9_2_1_U6.top_add_9s_9s_9_2_1_Adder_4_U.u1.a ;
wire [3:0] \add_9s_9s_9_2_1_U6.top_add_9s_9s_9_2_1_Adder_4_U.u1.b ;
wire \add_9s_9s_9_2_1_U6.top_add_9s_9s_9_2_1_Adder_4_U.u1.cin ;
wire \add_9s_9s_9_2_1_U6.top_add_9s_9s_9_2_1_Adder_4_U.u1.cout ;
wire [3:0] \add_9s_9s_9_2_1_U6.top_add_9s_9s_9_2_1_Adder_4_U.u1.s ;
wire [4:0] \add_9s_9s_9_2_1_U6.top_add_9s_9s_9_2_1_Adder_4_U.u2.a ;
wire [4:0] \add_9s_9s_9_2_1_U6.top_add_9s_9s_9_2_1_Adder_4_U.u2.b ;
wire \add_9s_9s_9_2_1_U6.top_add_9s_9s_9_2_1_Adder_4_U.u2.cin ;
wire \add_9s_9s_9_2_1_U6.top_add_9s_9s_9_2_1_Adder_4_U.u2.cout ;
wire [4:0] \add_9s_9s_9_2_1_U6.top_add_9s_9s_9_2_1_Adder_4_U.u2.s ;
wire and_ln353_fu_584_p2;
wire and_ln788_1_fu_451_p2;
wire and_ln788_fu_446_p2;
wire ap_CS_fsm_state1;
wire ap_CS_fsm_state10;
wire ap_CS_fsm_state11;
wire ap_CS_fsm_state12;
wire ap_CS_fsm_state13;
wire ap_CS_fsm_state14;
wire ap_CS_fsm_state15;
wire ap_CS_fsm_state16;
wire ap_CS_fsm_state17;
wire ap_CS_fsm_state18;
wire ap_CS_fsm_state19;
wire ap_CS_fsm_state2;
wire ap_CS_fsm_state20;
wire ap_CS_fsm_state21;
wire ap_CS_fsm_state22;
wire ap_CS_fsm_state23;
wire ap_CS_fsm_state24;
wire ap_CS_fsm_state25;
wire ap_CS_fsm_state26;
wire ap_CS_fsm_state27;
wire ap_CS_fsm_state28;
wire ap_CS_fsm_state3;
wire ap_CS_fsm_state4;
wire ap_CS_fsm_state5;
wire ap_CS_fsm_state6;
wire ap_CS_fsm_state7;
wire ap_CS_fsm_state8;
wire ap_CS_fsm_state9;
wire [27:0] ap_NS_fsm;
wire ap_clk;
wire ap_done;
wire ap_idle;
wire ap_ready;
wire ap_rst;
wire ap_start;
wire \ashr_32s_32s_32_7_1_U16.ce ;
wire \ashr_32s_32s_32_7_1_U16.clk ;
wire [31:0] \ashr_32s_32s_32_7_1_U16.din0 ;
wire [31:0] \ashr_32s_32s_32_7_1_U16.din1 ;
wire [31:0] \ashr_32s_32s_32_7_1_U16.din1_cast ;
wire [31:0] \ashr_32s_32s_32_7_1_U16.din1_mask ;
wire [31:0] \ashr_32s_32s_32_7_1_U16.dout ;
wire \ashr_32s_32s_32_7_1_U16.reset ;
wire [31:0] conv_i188_fu_905_p1;
wire [31:0] grp_fu_1018_p1;
wire [31:0] grp_fu_1018_p2;
wire [4:0] grp_fu_1023_p0;
wire [4:0] grp_fu_1023_p1;
wire [4:0] grp_fu_1023_p2;
wire [31:0] grp_fu_1032_p0;
wire [31:0] grp_fu_1032_p2;
wire [1:0] grp_fu_253_p0;
wire [1:0] grp_fu_253_p1;
wire [1:0] grp_fu_253_p2;
wire [15:0] grp_fu_281_p0;
wire [15:0] grp_fu_281_p1;
wire [15:0] grp_fu_281_p2;
wire [8:0] grp_fu_365_p0;
wire [8:0] grp_fu_365_p2;
wire [35:0] grp_fu_494_p2;
wire [32:0] grp_fu_609_p0;
wire [32:0] grp_fu_609_p1;
wire [32:0] grp_fu_609_p2;
wire [8:0] grp_fu_629_p0;
wire [8:0] grp_fu_629_p1;
wire [8:0] grp_fu_629_p2;
wire [7:0] grp_fu_677_p2;
wire [2:0] grp_fu_682_p2;
wire [4:0] grp_fu_707_p0;
wire [4:0] grp_fu_707_p2;
wire [4:0] grp_fu_717_p0;
wire [4:0] grp_fu_717_p2;
wire [1:0] grp_fu_786_p2;
wire [28:0] grp_fu_833_p0;
wire [28:0] grp_fu_833_p1;
wire [28:0] grp_fu_833_p2;
wire [8:0] grp_fu_845_p0;
wire [8:0] grp_fu_845_p1;
wire [8:0] grp_fu_845_p2;
wire [5:0] grp_fu_854_p1;
wire [5:0] grp_fu_854_p2;
wire [16:0] grp_fu_896_p0;
wire [16:0] grp_fu_896_p1;
wire [16:0] grp_fu_896_p2;
wire [31:0] grp_fu_908_p1;
wire [31:0] grp_fu_908_p2;
wire [31:0] grp_fu_917_p1;
wire [31:0] grp_fu_917_p2;
wire [16:0] grp_fu_926_p0;
wire [16:0] grp_fu_926_p2;
wire [33:0] grp_fu_946_p0;
wire [33:0] grp_fu_946_p1;
wire [33:0] grp_fu_946_p2;
wire [31:0] grp_fu_962_p2;
wire icmp_ln785_fu_357_p2;
wire icmp_ln790_fu_482_p2;
wire icmp_ln850_fu_500_p2;
wire icmp_ln851_1_fu_781_p2;
wire icmp_ln851_2_fu_635_p2;
wire icmp_ln851_3_fu_701_p2;
wire icmp_ln851_fu_672_p2;
wire [7:0] lhs_V_2_fu_615_p3;
wire [13:0] lhs_V_fu_266_p3;
wire [25:0] lhs_cast_fu_405_p3;
wire [9:0] lhs_fu_325_p3;
wire \mul_32s_4s_36_7_1_U4.ce ;
wire \mul_32s_4s_36_7_1_U4.clk ;
wire [31:0] \mul_32s_4s_36_7_1_U4.din0 ;
wire [3:0] \mul_32s_4s_36_7_1_U4.din1 ;
wire [35:0] \mul_32s_4s_36_7_1_U4.dout ;
wire \mul_32s_4s_36_7_1_U4.reset ;
wire [31:0] \mul_32s_4s_36_7_1_U4.top_mul_32s_4s_36_7_1_Mul_DSP_0_U.a ;
wire [3:0] \mul_32s_4s_36_7_1_U4.top_mul_32s_4s_36_7_1_Mul_DSP_0_U.b ;
wire \mul_32s_4s_36_7_1_U4.top_mul_32s_4s_36_7_1_Mul_DSP_0_U.ce ;
wire \mul_32s_4s_36_7_1_U4.top_mul_32s_4s_36_7_1_Mul_DSP_0_U.clk ;
wire [35:0] \mul_32s_4s_36_7_1_U4.top_mul_32s_4s_36_7_1_Mul_DSP_0_U.p ;
wire [35:0] \mul_32s_4s_36_7_1_U4.top_mul_32s_4s_36_7_1_Mul_DSP_0_U.tmp_product ;
wire [7:0] op_0;
wire [7:0] op_1;
wire [15:0] op_13;
wire [7:0] op_14;
wire [3:0] op_15;
wire [1:0] op_16;
wire [1:0] op_17;
wire [3:0] op_18;
wire [3:0] op_2;
wire [31:0] op_29;
wire op_29_ap_vld;
wire [7:0] op_3_V_fu_259_p3;
wire [31:0] op_4;
wire op_5;
wire [7:0] op_8_V_fu_544_p3;
wire [25:0] op_9_V_fu_774_p3;
wire [25:0] or_ln1195_fu_416_p2;
wire or_ln384_1_fu_539_p2;
wire or_ln384_fu_467_p2;
wire or_ln785_fu_370_p2;
wire or_ln788_fu_522_p2;
wire overflow_1_fu_477_p2;
wire overflow_fu_379_p2;
wire p_Result_10_fu_980_p3;
wire p_Result_6_fu_722_p3;
wire p_Result_7_fu_870_p3;
wire p_Result_8_fu_755_p3;
wire p_Result_9_fu_791_p3;
wire [31:0] p_Result_s_fu_577_p1;
wire p_Result_s_fu_577_p3;
wire [1:0] p_Val2_2_fu_505_p4;
wire [7:0] p_Val2_4_fu_514_p1;
wire [1:0] r_fu_975_p3;
wire [4:0] ret_V_15_fu_803_p3;
wire ret_V_19_fu_589_p2;
wire [9:0] ret_V_20_fu_336_p2;
wire [1:0] ret_V_24_fu_882_p3;
wire [31:0] ret_V_27_fu_996_p3;
wire [7:0] ret_V_8_fu_734_p3;
wire [28:0] rhs_1_fu_598_p3;
wire [27:0] rhs_3_fu_822_p3;
wire select_ln1193_fu_313_p0;
wire [8:0] select_ln1193_fu_313_p3;
wire select_ln1498_fu_426_p0;
wire [31:0] select_ln1498_fu_426_p3;
wire [1:0] select_ln384_2_fu_552_p3;
wire [1:0] select_ln384_3_fu_559_p3;
wire [7:0] select_ln384_fu_532_p3;
wire [4:0] select_ln69_fu_640_p3;
wire [1:0] select_ln850_2_fu_877_p3;
wire [4:0] select_ln850_3_fu_798_p3;
wire [31:0] select_ln850_5_fu_990_p3;
wire [2:0] select_ln850_6_fu_762_p3;
wire [2:0] select_ln850_7_fu_767_p3;
wire [7:0] select_ln850_fu_729_p3;
wire [9:0] sext_ln1196_fu_333_p1;
wire [15:0] sext_ln69_7_fu_1011_p1;
wire [31:0] sext_ln703_2_fu_595_p0;
wire [1:0] sext_ln703_4_fu_931_p0;
wire \shl_32s_32s_32_7_1_U17.ce ;
wire \shl_32s_32s_32_7_1_U17.clk ;
wire [31:0] \shl_32s_32s_32_7_1_U17.din0 ;
wire [31:0] \shl_32s_32s_32_7_1_U17.din1 ;
wire [31:0] \shl_32s_32s_32_7_1_U17.din1_cast ;
wire [31:0] \shl_32s_32s_32_7_1_U17.din1_mask ;
wire [31:0] \shl_32s_32s_32_7_1_U17.dout ;
wire \shl_32s_32s_32_7_1_U17.reset ;
wire [31:0] signbit_fu_433_p1;
wire signbit_fu_433_p2;
wire \sub_16ns_16s_16_2_1_U2.ce ;
wire \sub_16ns_16s_16_2_1_U2.clk ;
wire [15:0] \sub_16ns_16s_16_2_1_U2.din0 ;
wire [15:0] \sub_16ns_16s_16_2_1_U2.din1 ;
wire [15:0] \sub_16ns_16s_16_2_1_U2.dout ;
wire \sub_16ns_16s_16_2_1_U2.reset ;
wire [15:0] \sub_16ns_16s_16_2_1_U2.top_sub_16ns_16s_16_2_1_Adder_1_U.a ;
wire [15:0] \sub_16ns_16s_16_2_1_U2.top_sub_16ns_16s_16_2_1_Adder_1_U.ain_s0 ;
wire [15:0] \sub_16ns_16s_16_2_1_U2.top_sub_16ns_16s_16_2_1_Adder_1_U.b ;
wire [15:0] \sub_16ns_16s_16_2_1_U2.top_sub_16ns_16s_16_2_1_Adder_1_U.bin_s0 ;
wire \sub_16ns_16s_16_2_1_U2.top_sub_16ns_16s_16_2_1_Adder_1_U.ce ;
wire \sub_16ns_16s_16_2_1_U2.top_sub_16ns_16s_16_2_1_Adder_1_U.clk ;
wire \sub_16ns_16s_16_2_1_U2.top_sub_16ns_16s_16_2_1_Adder_1_U.facout_s1 ;
wire \sub_16ns_16s_16_2_1_U2.top_sub_16ns_16s_16_2_1_Adder_1_U.facout_s2 ;
wire [7:0] \sub_16ns_16s_16_2_1_U2.top_sub_16ns_16s_16_2_1_Adder_1_U.fas_s1 ;
wire [7:0] \sub_16ns_16s_16_2_1_U2.top_sub_16ns_16s_16_2_1_Adder_1_U.fas_s2 ;
wire \sub_16ns_16s_16_2_1_U2.top_sub_16ns_16s_16_2_1_Adder_1_U.reset ;
wire [15:0] \sub_16ns_16s_16_2_1_U2.top_sub_16ns_16s_16_2_1_Adder_1_U.s ;
wire [7:0] \sub_16ns_16s_16_2_1_U2.top_sub_16ns_16s_16_2_1_Adder_1_U.u1.a ;
wire [7:0] \sub_16ns_16s_16_2_1_U2.top_sub_16ns_16s_16_2_1_Adder_1_U.u1.b ;
wire \sub_16ns_16s_16_2_1_U2.top_sub_16ns_16s_16_2_1_Adder_1_U.u1.cin ;
wire \sub_16ns_16s_16_2_1_U2.top_sub_16ns_16s_16_2_1_Adder_1_U.u1.cout ;
wire [7:0] \sub_16ns_16s_16_2_1_U2.top_sub_16ns_16s_16_2_1_Adder_1_U.u1.s ;
wire [7:0] \sub_16ns_16s_16_2_1_U2.top_sub_16ns_16s_16_2_1_Adder_1_U.u2.a ;
wire [7:0] \sub_16ns_16s_16_2_1_U2.top_sub_16ns_16s_16_2_1_Adder_1_U.u2.b ;
wire \sub_16ns_16s_16_2_1_U2.top_sub_16ns_16s_16_2_1_Adder_1_U.u2.cin ;
wire \sub_16ns_16s_16_2_1_U2.top_sub_16ns_16s_16_2_1_Adder_1_U.u2.cout ;
wire [7:0] \sub_16ns_16s_16_2_1_U2.top_sub_16ns_16s_16_2_1_Adder_1_U.u2.s ;
wire \sub_33s_33s_33_2_1_U5.ce ;
wire \sub_33s_33s_33_2_1_U5.clk ;
wire [32:0] \sub_33s_33s_33_2_1_U5.din0 ;
wire [32:0] \sub_33s_33s_33_2_1_U5.din1 ;
wire [32:0] \sub_33s_33s_33_2_1_U5.dout ;
wire \sub_33s_33s_33_2_1_U5.reset ;
wire [32:0] \sub_33s_33s_33_2_1_U5.top_sub_33s_33s_33_2_1_Adder_3_U.a ;
wire [32:0] \sub_33s_33s_33_2_1_U5.top_sub_33s_33s_33_2_1_Adder_3_U.ain_s0 ;
wire [32:0] \sub_33s_33s_33_2_1_U5.top_sub_33s_33s_33_2_1_Adder_3_U.b ;
wire [32:0] \sub_33s_33s_33_2_1_U5.top_sub_33s_33s_33_2_1_Adder_3_U.bin_s0 ;
wire \sub_33s_33s_33_2_1_U5.top_sub_33s_33s_33_2_1_Adder_3_U.ce ;
wire \sub_33s_33s_33_2_1_U5.top_sub_33s_33s_33_2_1_Adder_3_U.clk ;
wire \sub_33s_33s_33_2_1_U5.top_sub_33s_33s_33_2_1_Adder_3_U.facout_s1 ;
wire \sub_33s_33s_33_2_1_U5.top_sub_33s_33s_33_2_1_Adder_3_U.facout_s2 ;
wire [15:0] \sub_33s_33s_33_2_1_U5.top_sub_33s_33s_33_2_1_Adder_3_U.fas_s1 ;
wire [16:0] \sub_33s_33s_33_2_1_U5.top_sub_33s_33s_33_2_1_Adder_3_U.fas_s2 ;
wire \sub_33s_33s_33_2_1_U5.top_sub_33s_33s_33_2_1_Adder_3_U.reset ;
wire [32:0] \sub_33s_33s_33_2_1_U5.top_sub_33s_33s_33_2_1_Adder_3_U.s ;
wire [15:0] \sub_33s_33s_33_2_1_U5.top_sub_33s_33s_33_2_1_Adder_3_U.u1.a ;
wire [15:0] \sub_33s_33s_33_2_1_U5.top_sub_33s_33s_33_2_1_Adder_3_U.u1.b ;
wire \sub_33s_33s_33_2_1_U5.top_sub_33s_33s_33_2_1_Adder_3_U.u1.cin ;
wire \sub_33s_33s_33_2_1_U5.top_sub_33s_33s_33_2_1_Adder_3_U.u1.cout ;
wire [15:0] \sub_33s_33s_33_2_1_U5.top_sub_33s_33s_33_2_1_Adder_3_U.u1.s ;
wire [16:0] \sub_33s_33s_33_2_1_U5.top_sub_33s_33s_33_2_1_Adder_3_U.u2.a ;
wire [16:0] \sub_33s_33s_33_2_1_U5.top_sub_33s_33s_33_2_1_Adder_3_U.u2.b ;
wire \sub_33s_33s_33_2_1_U5.top_sub_33s_33s_33_2_1_Adder_3_U.u2.cin ;
wire \sub_33s_33s_33_2_1_U5.top_sub_33s_33s_33_2_1_Adder_3_U.u2.cout ;
wire [16:0] \sub_33s_33s_33_2_1_U5.top_sub_33s_33s_33_2_1_Adder_3_U.u2.s ;
wire \sub_6ns_6s_6_2_1_U14.ce ;
wire \sub_6ns_6s_6_2_1_U14.clk ;
wire [5:0] \sub_6ns_6s_6_2_1_U14.din0 ;
wire [5:0] \sub_6ns_6s_6_2_1_U14.din1 ;
wire [5:0] \sub_6ns_6s_6_2_1_U14.dout ;
wire \sub_6ns_6s_6_2_1_U14.reset ;
wire [5:0] \sub_6ns_6s_6_2_1_U14.top_sub_6ns_6s_6_2_1_Adder_10_U.a ;
wire [5:0] \sub_6ns_6s_6_2_1_U14.top_sub_6ns_6s_6_2_1_Adder_10_U.ain_s0 ;
wire [5:0] \sub_6ns_6s_6_2_1_U14.top_sub_6ns_6s_6_2_1_Adder_10_U.b ;
wire [5:0] \sub_6ns_6s_6_2_1_U14.top_sub_6ns_6s_6_2_1_Adder_10_U.bin_s0 ;
wire \sub_6ns_6s_6_2_1_U14.top_sub_6ns_6s_6_2_1_Adder_10_U.ce ;
wire \sub_6ns_6s_6_2_1_U14.top_sub_6ns_6s_6_2_1_Adder_10_U.clk ;
wire \sub_6ns_6s_6_2_1_U14.top_sub_6ns_6s_6_2_1_Adder_10_U.facout_s1 ;
wire \sub_6ns_6s_6_2_1_U14.top_sub_6ns_6s_6_2_1_Adder_10_U.facout_s2 ;
wire [2:0] \sub_6ns_6s_6_2_1_U14.top_sub_6ns_6s_6_2_1_Adder_10_U.fas_s1 ;
wire [2:0] \sub_6ns_6s_6_2_1_U14.top_sub_6ns_6s_6_2_1_Adder_10_U.fas_s2 ;
wire \sub_6ns_6s_6_2_1_U14.top_sub_6ns_6s_6_2_1_Adder_10_U.reset ;
wire [5:0] \sub_6ns_6s_6_2_1_U14.top_sub_6ns_6s_6_2_1_Adder_10_U.s ;
wire [2:0] \sub_6ns_6s_6_2_1_U14.top_sub_6ns_6s_6_2_1_Adder_10_U.u1.a ;
wire [2:0] \sub_6ns_6s_6_2_1_U14.top_sub_6ns_6s_6_2_1_Adder_10_U.u1.b ;
wire \sub_6ns_6s_6_2_1_U14.top_sub_6ns_6s_6_2_1_Adder_10_U.u1.cin ;
wire \sub_6ns_6s_6_2_1_U14.top_sub_6ns_6s_6_2_1_Adder_10_U.u1.cout ;
wire [2:0] \sub_6ns_6s_6_2_1_U14.top_sub_6ns_6s_6_2_1_Adder_10_U.u1.s ;
wire [2:0] \sub_6ns_6s_6_2_1_U14.top_sub_6ns_6s_6_2_1_Adder_10_U.u2.a ;
wire [2:0] \sub_6ns_6s_6_2_1_U14.top_sub_6ns_6s_6_2_1_Adder_10_U.u2.b ;
wire \sub_6ns_6s_6_2_1_U14.top_sub_6ns_6s_6_2_1_Adder_10_U.u2.cin ;
wire \sub_6ns_6s_6_2_1_U14.top_sub_6ns_6s_6_2_1_Adder_10_U.u2.cout ;
wire [2:0] \sub_6ns_6s_6_2_1_U14.top_sub_6ns_6s_6_2_1_Adder_10_U.u2.s ;
wire \sub_9s_9ns_9_2_1_U3.ce ;
wire \sub_9s_9ns_9_2_1_U3.clk ;
wire [8:0] \sub_9s_9ns_9_2_1_U3.din0 ;
wire [8:0] \sub_9s_9ns_9_2_1_U3.din1 ;
wire [8:0] \sub_9s_9ns_9_2_1_U3.dout ;
wire \sub_9s_9ns_9_2_1_U3.reset ;
wire [8:0] \sub_9s_9ns_9_2_1_U3.top_sub_9s_9ns_9_2_1_Adder_2_U.a ;
wire [8:0] \sub_9s_9ns_9_2_1_U3.top_sub_9s_9ns_9_2_1_Adder_2_U.ain_s0 ;
wire [8:0] \sub_9s_9ns_9_2_1_U3.top_sub_9s_9ns_9_2_1_Adder_2_U.b ;
wire [8:0] \sub_9s_9ns_9_2_1_U3.top_sub_9s_9ns_9_2_1_Adder_2_U.bin_s0 ;
wire \sub_9s_9ns_9_2_1_U3.top_sub_9s_9ns_9_2_1_Adder_2_U.ce ;
wire \sub_9s_9ns_9_2_1_U3.top_sub_9s_9ns_9_2_1_Adder_2_U.clk ;
wire \sub_9s_9ns_9_2_1_U3.top_sub_9s_9ns_9_2_1_Adder_2_U.facout_s1 ;
wire \sub_9s_9ns_9_2_1_U3.top_sub_9s_9ns_9_2_1_Adder_2_U.facout_s2 ;
wire [3:0] \sub_9s_9ns_9_2_1_U3.top_sub_9s_9ns_9_2_1_Adder_2_U.fas_s1 ;
wire [4:0] \sub_9s_9ns_9_2_1_U3.top_sub_9s_9ns_9_2_1_Adder_2_U.fas_s2 ;
wire \sub_9s_9ns_9_2_1_U3.top_sub_9s_9ns_9_2_1_Adder_2_U.reset ;
wire [8:0] \sub_9s_9ns_9_2_1_U3.top_sub_9s_9ns_9_2_1_Adder_2_U.s ;
wire [3:0] \sub_9s_9ns_9_2_1_U3.top_sub_9s_9ns_9_2_1_Adder_2_U.u1.a ;
wire [3:0] \sub_9s_9ns_9_2_1_U3.top_sub_9s_9ns_9_2_1_Adder_2_U.u1.b ;
wire \sub_9s_9ns_9_2_1_U3.top_sub_9s_9ns_9_2_1_Adder_2_U.u1.cin ;
wire \sub_9s_9ns_9_2_1_U3.top_sub_9s_9ns_9_2_1_Adder_2_U.u1.cout ;
wire [3:0] \sub_9s_9ns_9_2_1_U3.top_sub_9s_9ns_9_2_1_Adder_2_U.u1.s ;
wire [4:0] \sub_9s_9ns_9_2_1_U3.top_sub_9s_9ns_9_2_1_Adder_2_U.u2.a ;
wire [4:0] \sub_9s_9ns_9_2_1_U3.top_sub_9s_9ns_9_2_1_Adder_2_U.u2.b ;
wire \sub_9s_9ns_9_2_1_U3.top_sub_9s_9ns_9_2_1_Adder_2_U.u2.cin ;
wire \sub_9s_9ns_9_2_1_U3.top_sub_9s_9ns_9_2_1_Adder_2_U.u2.cout ;
wire [4:0] \sub_9s_9ns_9_2_1_U3.top_sub_9s_9ns_9_2_1_Adder_2_U.u2.s ;
wire tmp_1_fu_570_p3;
wire tmp_6_fu_439_p3;
wire [17:0] tmp_fu_935_p3;
wire [31:0] trunc_ln1195_fu_412_p0;
wire [25:0] trunc_ln1195_fu_412_p1;
wire [1:0] trunc_ln1497_1_fu_971_p1;
wire [1:0] trunc_ln1497_fu_967_p1;
wire trunc_ln728_fu_321_p1;
wire [6:0] trunc_ln790_fu_401_p1;
wire [24:0] trunc_ln851_1_fu_658_p1;
wire [24:0] trunc_ln851_2_fu_751_p1;
wire [5:0] trunc_ln851_3_fu_566_p1;
wire [2:0] trunc_ln851_4_fu_697_p1;
wire [1:0] trunc_ln851_5_fu_987_p0;
wire trunc_ln851_5_fu_987_p1;
wire [24:0] trunc_ln851_fu_422_p1;
wire underflow_1_fu_527_p2;
wire underflow_fu_462_p2;
wire xor_ln785_1_fu_472_p2;
wire xor_ln785_fu_374_p2;
wire xor_ln786_fu_517_p2;
wire xor_ln788_fu_456_p2;


assign _066_ = ap_CS_fsm[11] & _072_;
assign _067_ = tmp_13_reg_1373 & ap_CS_fsm[15];
assign _068_ = _073_ & ap_CS_fsm[22];
assign _069_ = tmp_13_reg_1373 & ap_CS_fsm[22];
assign _070_ = _074_ & ap_CS_fsm[0];
assign _071_ = ap_start & ap_CS_fsm[0];
assign and_ln353_fu_584_p2 = op_4[31] & icmp_ln850_reg_1209;
assign and_ln788_1_fu_451_p2 = p_Result_12_reg_1091 & and_ln788_fu_446_p2;
assign and_ln788_fu_446_p2 = ret_V_21_reg_1079[6] & Range1_all_ones_reg_1119;
assign overflow_1_fu_477_p2 = xor_ln785_1_fu_472_p2 & p_Result_14_reg_1151;
assign overflow_fu_379_p2 = xor_ln785_fu_374_p2 & or_ln785_fu_370_p2;
assign underflow_1_fu_527_p2 = p_Result_13_reg_1145 & or_ln788_fu_522_p2;
assign underflow_fu_462_p2 = xor_ln788_fu_456_p2 & p_Result_11_reg_1085;
assign xor_ln786_fu_517_p2 = ~ p_Result_14_reg_1151;
assign xor_ln788_fu_456_p2 = ~ and_ln788_1_fu_451_p2;
assign xor_ln785_1_fu_472_p2 = ~ p_Result_13_reg_1145;
assign xor_ln785_fu_374_p2 = ~ p_Result_11_reg_1085;
assign _072_ = ~ icmp_ln851_2_reg_1249;
assign _073_ = ~ tmp_13_reg_1373;
assign _074_ = ~ ap_start;
assign _075_ = p_Result_s_20_reg_1097 == 8'hff;
assign _076_ = ! trunc_ln790_reg_1157;
assign _077_ = ! trunc_ln851_2_reg_1342;
assign _078_ = ! trunc_ln851_3_reg_1224;
assign _079_ = ! op_14[2:0];
assign _080_ = ! trunc_ln851_1_reg_1271;
assign _081_ = select_ln1498_fu_426_p3 == op_4;
always @(posedge \add_17s_17ns_17_2_1_U18.top_add_17s_17ns_17_2_1_Adder_12_U.clk )
\add_17s_17ns_17_2_1_U18.top_add_17s_17ns_17_2_1_Adder_12_U.bin_s1  <= _083_;
always @(posedge \add_17s_17ns_17_2_1_U18.top_add_17s_17ns_17_2_1_Adder_12_U.clk )
\add_17s_17ns_17_2_1_U18.top_add_17s_17ns_17_2_1_Adder_12_U.ain_s1  <= _082_;
always @(posedge \add_17s_17ns_17_2_1_U18.top_add_17s_17ns_17_2_1_Adder_12_U.clk )
\add_17s_17ns_17_2_1_U18.top_add_17s_17ns_17_2_1_Adder_12_U.sum_s1  <= _085_;
always @(posedge \add_17s_17ns_17_2_1_U18.top_add_17s_17ns_17_2_1_Adder_12_U.clk )
\add_17s_17ns_17_2_1_U18.top_add_17s_17ns_17_2_1_Adder_12_U.carry_s1  <= _084_;
assign _083_ = \add_17s_17ns_17_2_1_U18.top_add_17s_17ns_17_2_1_Adder_12_U.ce  ? \add_17s_17ns_17_2_1_U18.top_add_17s_17ns_17_2_1_Adder_12_U.b [16:8] : \add_17s_17ns_17_2_1_U18.top_add_17s_17ns_17_2_1_Adder_12_U.bin_s1 ;
assign _082_ = \add_17s_17ns_17_2_1_U18.top_add_17s_17ns_17_2_1_Adder_12_U.ce  ? \add_17s_17ns_17_2_1_U18.top_add_17s_17ns_17_2_1_Adder_12_U.a [16:8] : \add_17s_17ns_17_2_1_U18.top_add_17s_17ns_17_2_1_Adder_12_U.ain_s1 ;
assign _084_ = \add_17s_17ns_17_2_1_U18.top_add_17s_17ns_17_2_1_Adder_12_U.ce  ? \add_17s_17ns_17_2_1_U18.top_add_17s_17ns_17_2_1_Adder_12_U.facout_s1  : \add_17s_17ns_17_2_1_U18.top_add_17s_17ns_17_2_1_Adder_12_U.carry_s1 ;
assign _085_ = \add_17s_17ns_17_2_1_U18.top_add_17s_17ns_17_2_1_Adder_12_U.ce  ? \add_17s_17ns_17_2_1_U18.top_add_17s_17ns_17_2_1_Adder_12_U.fas_s1  : \add_17s_17ns_17_2_1_U18.top_add_17s_17ns_17_2_1_Adder_12_U.sum_s1 ;
assign _086_ = \add_17s_17ns_17_2_1_U18.top_add_17s_17ns_17_2_1_Adder_12_U.u1.a  + \add_17s_17ns_17_2_1_U18.top_add_17s_17ns_17_2_1_Adder_12_U.u1.b ;
assign { \add_17s_17ns_17_2_1_U18.top_add_17s_17ns_17_2_1_Adder_12_U.u1.cout , \add_17s_17ns_17_2_1_U18.top_add_17s_17ns_17_2_1_Adder_12_U.u1.s  } = _086_ + \add_17s_17ns_17_2_1_U18.top_add_17s_17ns_17_2_1_Adder_12_U.u1.cin ;
assign _087_ = \add_17s_17ns_17_2_1_U18.top_add_17s_17ns_17_2_1_Adder_12_U.u2.a  + \add_17s_17ns_17_2_1_U18.top_add_17s_17ns_17_2_1_Adder_12_U.u2.b ;
assign { \add_17s_17ns_17_2_1_U18.top_add_17s_17ns_17_2_1_Adder_12_U.u2.cout , \add_17s_17ns_17_2_1_U18.top_add_17s_17ns_17_2_1_Adder_12_U.u2.s  } = _087_ + \add_17s_17ns_17_2_1_U18.top_add_17s_17ns_17_2_1_Adder_12_U.u2.cin ;
always @(posedge \add_17s_17s_17_2_1_U15.top_add_17s_17s_17_2_1_Adder_11_U.clk )
\add_17s_17s_17_2_1_U15.top_add_17s_17s_17_2_1_Adder_11_U.bin_s1  <= _089_;
always @(posedge \add_17s_17s_17_2_1_U15.top_add_17s_17s_17_2_1_Adder_11_U.clk )
\add_17s_17s_17_2_1_U15.top_add_17s_17s_17_2_1_Adder_11_U.ain_s1  <= _088_;
always @(posedge \add_17s_17s_17_2_1_U15.top_add_17s_17s_17_2_1_Adder_11_U.clk )
\add_17s_17s_17_2_1_U15.top_add_17s_17s_17_2_1_Adder_11_U.sum_s1  <= _091_;
always @(posedge \add_17s_17s_17_2_1_U15.top_add_17s_17s_17_2_1_Adder_11_U.clk )
\add_17s_17s_17_2_1_U15.top_add_17s_17s_17_2_1_Adder_11_U.carry_s1  <= _090_;
assign _089_ = \add_17s_17s_17_2_1_U15.top_add_17s_17s_17_2_1_Adder_11_U.ce  ? \add_17s_17s_17_2_1_U15.top_add_17s_17s_17_2_1_Adder_11_U.b [16:8] : \add_17s_17s_17_2_1_U15.top_add_17s_17s_17_2_1_Adder_11_U.bin_s1 ;
assign _088_ = \add_17s_17s_17_2_1_U15.top_add_17s_17s_17_2_1_Adder_11_U.ce  ? \add_17s_17s_17_2_1_U15.top_add_17s_17s_17_2_1_Adder_11_U.a [16:8] : \add_17s_17s_17_2_1_U15.top_add_17s_17s_17_2_1_Adder_11_U.ain_s1 ;
assign _090_ = \add_17s_17s_17_2_1_U15.top_add_17s_17s_17_2_1_Adder_11_U.ce  ? \add_17s_17s_17_2_1_U15.top_add_17s_17s_17_2_1_Adder_11_U.facout_s1  : \add_17s_17s_17_2_1_U15.top_add_17s_17s_17_2_1_Adder_11_U.carry_s1 ;
assign _091_ = \add_17s_17s_17_2_1_U15.top_add_17s_17s_17_2_1_Adder_11_U.ce  ? \add_17s_17s_17_2_1_U15.top_add_17s_17s_17_2_1_Adder_11_U.fas_s1  : \add_17s_17s_17_2_1_U15.top_add_17s_17s_17_2_1_Adder_11_U.sum_s1 ;
assign _092_ = \add_17s_17s_17_2_1_U15.top_add_17s_17s_17_2_1_Adder_11_U.u1.a  + \add_17s_17s_17_2_1_U15.top_add_17s_17s_17_2_1_Adder_11_U.u1.b ;
assign { \add_17s_17s_17_2_1_U15.top_add_17s_17s_17_2_1_Adder_11_U.u1.cout , \add_17s_17s_17_2_1_U15.top_add_17s_17s_17_2_1_Adder_11_U.u1.s  } = _092_ + \add_17s_17s_17_2_1_U15.top_add_17s_17s_17_2_1_Adder_11_U.u1.cin ;
assign _093_ = \add_17s_17s_17_2_1_U15.top_add_17s_17s_17_2_1_Adder_11_U.u2.a  + \add_17s_17s_17_2_1_U15.top_add_17s_17s_17_2_1_Adder_11_U.u2.b ;
assign { \add_17s_17s_17_2_1_U15.top_add_17s_17s_17_2_1_Adder_11_U.u2.cout , \add_17s_17s_17_2_1_U15.top_add_17s_17s_17_2_1_Adder_11_U.u2.s  } = _093_ + \add_17s_17s_17_2_1_U15.top_add_17s_17s_17_2_1_Adder_11_U.u2.cin ;
always @(posedge \add_29s_29ns_29_2_1_U12.top_add_29s_29ns_29_2_1_Adder_9_U.clk )
\add_29s_29ns_29_2_1_U12.top_add_29s_29ns_29_2_1_Adder_9_U.bin_s1  <= _095_;
always @(posedge \add_29s_29ns_29_2_1_U12.top_add_29s_29ns_29_2_1_Adder_9_U.clk )
\add_29s_29ns_29_2_1_U12.top_add_29s_29ns_29_2_1_Adder_9_U.ain_s1  <= _094_;
always @(posedge \add_29s_29ns_29_2_1_U12.top_add_29s_29ns_29_2_1_Adder_9_U.clk )
\add_29s_29ns_29_2_1_U12.top_add_29s_29ns_29_2_1_Adder_9_U.sum_s1  <= _097_;
always @(posedge \add_29s_29ns_29_2_1_U12.top_add_29s_29ns_29_2_1_Adder_9_U.clk )
\add_29s_29ns_29_2_1_U12.top_add_29s_29ns_29_2_1_Adder_9_U.carry_s1  <= _096_;
assign _095_ = \add_29s_29ns_29_2_1_U12.top_add_29s_29ns_29_2_1_Adder_9_U.ce  ? \add_29s_29ns_29_2_1_U12.top_add_29s_29ns_29_2_1_Adder_9_U.b [28:14] : \add_29s_29ns_29_2_1_U12.top_add_29s_29ns_29_2_1_Adder_9_U.bin_s1 ;
assign _094_ = \add_29s_29ns_29_2_1_U12.top_add_29s_29ns_29_2_1_Adder_9_U.ce  ? \add_29s_29ns_29_2_1_U12.top_add_29s_29ns_29_2_1_Adder_9_U.a [28:14] : \add_29s_29ns_29_2_1_U12.top_add_29s_29ns_29_2_1_Adder_9_U.ain_s1 ;
assign _096_ = \add_29s_29ns_29_2_1_U12.top_add_29s_29ns_29_2_1_Adder_9_U.ce  ? \add_29s_29ns_29_2_1_U12.top_add_29s_29ns_29_2_1_Adder_9_U.facout_s1  : \add_29s_29ns_29_2_1_U12.top_add_29s_29ns_29_2_1_Adder_9_U.carry_s1 ;
assign _097_ = \add_29s_29ns_29_2_1_U12.top_add_29s_29ns_29_2_1_Adder_9_U.ce  ? \add_29s_29ns_29_2_1_U12.top_add_29s_29ns_29_2_1_Adder_9_U.fas_s1  : \add_29s_29ns_29_2_1_U12.top_add_29s_29ns_29_2_1_Adder_9_U.sum_s1 ;
assign _098_ = \add_29s_29ns_29_2_1_U12.top_add_29s_29ns_29_2_1_Adder_9_U.u1.a  + \add_29s_29ns_29_2_1_U12.top_add_29s_29ns_29_2_1_Adder_9_U.u1.b ;
assign { \add_29s_29ns_29_2_1_U12.top_add_29s_29ns_29_2_1_Adder_9_U.u1.cout , \add_29s_29ns_29_2_1_U12.top_add_29s_29ns_29_2_1_Adder_9_U.u1.s  } = _098_ + \add_29s_29ns_29_2_1_U12.top_add_29s_29ns_29_2_1_Adder_9_U.u1.cin ;
assign _099_ = \add_29s_29ns_29_2_1_U12.top_add_29s_29ns_29_2_1_Adder_9_U.u2.a  + \add_29s_29ns_29_2_1_U12.top_add_29s_29ns_29_2_1_Adder_9_U.u2.b ;
assign { \add_29s_29ns_29_2_1_U12.top_add_29s_29ns_29_2_1_Adder_9_U.u2.cout , \add_29s_29ns_29_2_1_U12.top_add_29s_29ns_29_2_1_Adder_9_U.u2.s  } = _099_ + \add_29s_29ns_29_2_1_U12.top_add_29s_29ns_29_2_1_Adder_9_U.u2.cin ;
always @(posedge \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.clk )
\add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.bin_s1  <= _101_;
always @(posedge \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.clk )
\add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.ain_s1  <= _100_;
always @(posedge \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.clk )
\add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.sum_s1  <= _103_;
always @(posedge \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.clk )
\add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.carry_s1  <= _102_;
assign _101_ = \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.ce  ? \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.b [1] : \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.bin_s1 ;
assign _100_ = \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.ce  ? \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.a [1] : \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.ain_s1 ;
assign _102_ = \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.ce  ? \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.facout_s1  : \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.carry_s1 ;
assign _103_ = \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.ce  ? \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.fas_s1  : \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.sum_s1 ;
assign _104_ = \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.u1.a  + \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.u1.b ;
assign { \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.u1.cout , \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.u1.s  } = _104_ + \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.u1.cin ;
assign _105_ = \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.u2.a  + \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.u2.b ;
assign { \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.u2.cout , \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.u2.s  } = _105_ + \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.u2.cin ;
always @(posedge \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_0_U.clk )
\add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_0_U.bin_s1  <= _107_;
always @(posedge \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_0_U.clk )
\add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_0_U.ain_s1  <= _106_;
always @(posedge \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_0_U.clk )
\add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_0_U.sum_s1  <= _109_;
always @(posedge \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_0_U.clk )
\add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_0_U.carry_s1  <= _108_;
assign _107_ = \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_0_U.ce  ? \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_0_U.b [1] : \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_0_U.bin_s1 ;
assign _106_ = \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_0_U.ce  ? \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_0_U.a [1] : \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_0_U.ain_s1 ;
assign _108_ = \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_0_U.ce  ? \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_0_U.facout_s1  : \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_0_U.carry_s1 ;
assign _109_ = \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_0_U.ce  ? \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_0_U.fas_s1  : \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_0_U.sum_s1 ;
assign _110_ = \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_0_U.u1.a  + \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_0_U.u1.b ;
assign { \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_0_U.u1.cout , \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_0_U.u1.s  } = _110_ + \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_0_U.u1.cin ;
assign _111_ = \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_0_U.u2.a  + \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_0_U.u2.b ;
assign { \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_0_U.u2.cout , \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_0_U.u2.s  } = _111_ + \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_0_U.u2.cin ;
always @(posedge \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_14_U.clk )
\add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_14_U.bin_s1  <= _113_;
always @(posedge \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_14_U.clk )
\add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_14_U.ain_s1  <= _112_;
always @(posedge \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_14_U.clk )
\add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_14_U.sum_s1  <= _115_;
always @(posedge \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_14_U.clk )
\add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_14_U.carry_s1  <= _114_;
assign _113_ = \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_14_U.ce  ? \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_14_U.b [31:16] : \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_14_U.bin_s1 ;
assign _112_ = \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_14_U.ce  ? \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_14_U.a [31:16] : \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_14_U.ain_s1 ;
assign _114_ = \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_14_U.ce  ? \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_14_U.facout_s1  : \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_14_U.carry_s1 ;
assign _115_ = \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_14_U.ce  ? \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_14_U.fas_s1  : \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_14_U.sum_s1 ;
assign _116_ = \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_14_U.u1.a  + \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_14_U.u1.b ;
assign { \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_14_U.u1.cout , \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_14_U.u1.s  } = _116_ + \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_14_U.u1.cin ;
assign _117_ = \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_14_U.u2.a  + \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_14_U.u2.b ;
assign { \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_14_U.u2.cout , \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_14_U.u2.s  } = _117_ + \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_14_U.u2.cin ;
always @(posedge \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_14_U.clk )
\add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_14_U.bin_s1  <= _119_;
always @(posedge \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_14_U.clk )
\add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_14_U.ain_s1  <= _118_;
always @(posedge \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_14_U.clk )
\add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_14_U.sum_s1  <= _121_;
always @(posedge \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_14_U.clk )
\add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_14_U.carry_s1  <= _120_;
assign _119_ = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_14_U.ce  ? \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_14_U.b [31:16] : \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_14_U.bin_s1 ;
assign _118_ = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_14_U.ce  ? \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_14_U.a [31:16] : \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_14_U.ain_s1 ;
assign _120_ = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_14_U.ce  ? \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_14_U.facout_s1  : \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_14_U.carry_s1 ;
assign _121_ = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_14_U.ce  ? \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_14_U.fas_s1  : \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_14_U.sum_s1 ;
assign _122_ = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_14_U.u1.a  + \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_14_U.u1.b ;
assign { \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_14_U.u1.cout , \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_14_U.u1.s  } = _122_ + \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_14_U.u1.cin ;
assign _123_ = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_14_U.u2.a  + \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_14_U.u2.b ;
assign { \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_14_U.u2.cout , \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_14_U.u2.s  } = _123_ + \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_14_U.u2.cin ;
always @(posedge \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_16_U.clk )
\add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_16_U.bin_s1  <= _125_;
always @(posedge \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_16_U.clk )
\add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_16_U.ain_s1  <= _124_;
always @(posedge \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_16_U.clk )
\add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_16_U.sum_s1  <= _127_;
always @(posedge \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_16_U.clk )
\add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_16_U.carry_s1  <= _126_;
assign _125_ = \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_16_U.ce  ? \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_16_U.b [31:16] : \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_16_U.bin_s1 ;
assign _124_ = \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_16_U.ce  ? \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_16_U.a [31:16] : \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_16_U.ain_s1 ;
assign _126_ = \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_16_U.ce  ? \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_16_U.facout_s1  : \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_16_U.carry_s1 ;
assign _127_ = \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_16_U.ce  ? \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_16_U.fas_s1  : \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_16_U.sum_s1 ;
assign _128_ = \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_16_U.u1.a  + \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_16_U.u1.b ;
assign { \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_16_U.u1.cout , \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_16_U.u1.s  } = _128_ + \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_16_U.u1.cin ;
assign _129_ = \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_16_U.u2.a  + \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_16_U.u2.b ;
assign { \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_16_U.u2.cout , \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_16_U.u2.s  } = _129_ + \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_16_U.u2.cin ;
always @(posedge \add_34s_34s_34_2_1_U19.top_add_34s_34s_34_2_1_Adder_13_U.clk )
\add_34s_34s_34_2_1_U19.top_add_34s_34s_34_2_1_Adder_13_U.bin_s1  <= _131_;
always @(posedge \add_34s_34s_34_2_1_U19.top_add_34s_34s_34_2_1_Adder_13_U.clk )
\add_34s_34s_34_2_1_U19.top_add_34s_34s_34_2_1_Adder_13_U.ain_s1  <= _130_;
always @(posedge \add_34s_34s_34_2_1_U19.top_add_34s_34s_34_2_1_Adder_13_U.clk )
\add_34s_34s_34_2_1_U19.top_add_34s_34s_34_2_1_Adder_13_U.sum_s1  <= _133_;
always @(posedge \add_34s_34s_34_2_1_U19.top_add_34s_34s_34_2_1_Adder_13_U.clk )
\add_34s_34s_34_2_1_U19.top_add_34s_34s_34_2_1_Adder_13_U.carry_s1  <= _132_;
assign _131_ = \add_34s_34s_34_2_1_U19.top_add_34s_34s_34_2_1_Adder_13_U.ce  ? \add_34s_34s_34_2_1_U19.top_add_34s_34s_34_2_1_Adder_13_U.b [33:17] : \add_34s_34s_34_2_1_U19.top_add_34s_34s_34_2_1_Adder_13_U.bin_s1 ;
assign _130_ = \add_34s_34s_34_2_1_U19.top_add_34s_34s_34_2_1_Adder_13_U.ce  ? \add_34s_34s_34_2_1_U19.top_add_34s_34s_34_2_1_Adder_13_U.a [33:17] : \add_34s_34s_34_2_1_U19.top_add_34s_34s_34_2_1_Adder_13_U.ain_s1 ;
assign _132_ = \add_34s_34s_34_2_1_U19.top_add_34s_34s_34_2_1_Adder_13_U.ce  ? \add_34s_34s_34_2_1_U19.top_add_34s_34s_34_2_1_Adder_13_U.facout_s1  : \add_34s_34s_34_2_1_U19.top_add_34s_34s_34_2_1_Adder_13_U.carry_s1 ;
assign _133_ = \add_34s_34s_34_2_1_U19.top_add_34s_34s_34_2_1_Adder_13_U.ce  ? \add_34s_34s_34_2_1_U19.top_add_34s_34s_34_2_1_Adder_13_U.fas_s1  : \add_34s_34s_34_2_1_U19.top_add_34s_34s_34_2_1_Adder_13_U.sum_s1 ;
assign _134_ = \add_34s_34s_34_2_1_U19.top_add_34s_34s_34_2_1_Adder_13_U.u1.a  + \add_34s_34s_34_2_1_U19.top_add_34s_34s_34_2_1_Adder_13_U.u1.b ;
assign { \add_34s_34s_34_2_1_U19.top_add_34s_34s_34_2_1_Adder_13_U.u1.cout , \add_34s_34s_34_2_1_U19.top_add_34s_34s_34_2_1_Adder_13_U.u1.s  } = _134_ + \add_34s_34s_34_2_1_U19.top_add_34s_34s_34_2_1_Adder_13_U.u1.cin ;
assign _135_ = \add_34s_34s_34_2_1_U19.top_add_34s_34s_34_2_1_Adder_13_U.u2.a  + \add_34s_34s_34_2_1_U19.top_add_34s_34s_34_2_1_Adder_13_U.u2.b ;
assign { \add_34s_34s_34_2_1_U19.top_add_34s_34s_34_2_1_Adder_13_U.u2.cout , \add_34s_34s_34_2_1_U19.top_add_34s_34s_34_2_1_Adder_13_U.u2.s  } = _135_ + \add_34s_34s_34_2_1_U19.top_add_34s_34s_34_2_1_Adder_13_U.u2.cin ;
always @(posedge \add_3ns_3ns_3_2_1_U8.top_add_3ns_3ns_3_2_1_Adder_6_U.clk )
\add_3ns_3ns_3_2_1_U8.top_add_3ns_3ns_3_2_1_Adder_6_U.bin_s1  <= _137_;
always @(posedge \add_3ns_3ns_3_2_1_U8.top_add_3ns_3ns_3_2_1_Adder_6_U.clk )
\add_3ns_3ns_3_2_1_U8.top_add_3ns_3ns_3_2_1_Adder_6_U.ain_s1  <= _136_;
always @(posedge \add_3ns_3ns_3_2_1_U8.top_add_3ns_3ns_3_2_1_Adder_6_U.clk )
\add_3ns_3ns_3_2_1_U8.top_add_3ns_3ns_3_2_1_Adder_6_U.sum_s1  <= _139_;
always @(posedge \add_3ns_3ns_3_2_1_U8.top_add_3ns_3ns_3_2_1_Adder_6_U.clk )
\add_3ns_3ns_3_2_1_U8.top_add_3ns_3ns_3_2_1_Adder_6_U.carry_s1  <= _138_;
assign _137_ = \add_3ns_3ns_3_2_1_U8.top_add_3ns_3ns_3_2_1_Adder_6_U.ce  ? \add_3ns_3ns_3_2_1_U8.top_add_3ns_3ns_3_2_1_Adder_6_U.b [2:1] : \add_3ns_3ns_3_2_1_U8.top_add_3ns_3ns_3_2_1_Adder_6_U.bin_s1 ;
assign _136_ = \add_3ns_3ns_3_2_1_U8.top_add_3ns_3ns_3_2_1_Adder_6_U.ce  ? \add_3ns_3ns_3_2_1_U8.top_add_3ns_3ns_3_2_1_Adder_6_U.a [2:1] : \add_3ns_3ns_3_2_1_U8.top_add_3ns_3ns_3_2_1_Adder_6_U.ain_s1 ;
assign _138_ = \add_3ns_3ns_3_2_1_U8.top_add_3ns_3ns_3_2_1_Adder_6_U.ce  ? \add_3ns_3ns_3_2_1_U8.top_add_3ns_3ns_3_2_1_Adder_6_U.facout_s1  : \add_3ns_3ns_3_2_1_U8.top_add_3ns_3ns_3_2_1_Adder_6_U.carry_s1 ;
assign _139_ = \add_3ns_3ns_3_2_1_U8.top_add_3ns_3ns_3_2_1_Adder_6_U.ce  ? \add_3ns_3ns_3_2_1_U8.top_add_3ns_3ns_3_2_1_Adder_6_U.fas_s1  : \add_3ns_3ns_3_2_1_U8.top_add_3ns_3ns_3_2_1_Adder_6_U.sum_s1 ;
assign _140_ = \add_3ns_3ns_3_2_1_U8.top_add_3ns_3ns_3_2_1_Adder_6_U.u1.a  + \add_3ns_3ns_3_2_1_U8.top_add_3ns_3ns_3_2_1_Adder_6_U.u1.b ;
assign { \add_3ns_3ns_3_2_1_U8.top_add_3ns_3ns_3_2_1_Adder_6_U.u1.cout , \add_3ns_3ns_3_2_1_U8.top_add_3ns_3ns_3_2_1_Adder_6_U.u1.s  } = _140_ + \add_3ns_3ns_3_2_1_U8.top_add_3ns_3ns_3_2_1_Adder_6_U.u1.cin ;
assign _141_ = \add_3ns_3ns_3_2_1_U8.top_add_3ns_3ns_3_2_1_Adder_6_U.u2.a  + \add_3ns_3ns_3_2_1_U8.top_add_3ns_3ns_3_2_1_Adder_6_U.u2.b ;
assign { \add_3ns_3ns_3_2_1_U8.top_add_3ns_3ns_3_2_1_Adder_6_U.u2.cout , \add_3ns_3ns_3_2_1_U8.top_add_3ns_3ns_3_2_1_Adder_6_U.u2.s  } = _141_ + \add_3ns_3ns_3_2_1_U8.top_add_3ns_3ns_3_2_1_Adder_6_U.u2.cin ;
always @(posedge \add_5ns_5ns_5_2_1_U9.top_add_5ns_5ns_5_2_1_Adder_7_U.clk )
\add_5ns_5ns_5_2_1_U9.top_add_5ns_5ns_5_2_1_Adder_7_U.bin_s1  <= _143_;
always @(posedge \add_5ns_5ns_5_2_1_U9.top_add_5ns_5ns_5_2_1_Adder_7_U.clk )
\add_5ns_5ns_5_2_1_U9.top_add_5ns_5ns_5_2_1_Adder_7_U.ain_s1  <= _142_;
always @(posedge \add_5ns_5ns_5_2_1_U9.top_add_5ns_5ns_5_2_1_Adder_7_U.clk )
\add_5ns_5ns_5_2_1_U9.top_add_5ns_5ns_5_2_1_Adder_7_U.sum_s1  <= _145_;
always @(posedge \add_5ns_5ns_5_2_1_U9.top_add_5ns_5ns_5_2_1_Adder_7_U.clk )
\add_5ns_5ns_5_2_1_U9.top_add_5ns_5ns_5_2_1_Adder_7_U.carry_s1  <= _144_;
assign _143_ = \add_5ns_5ns_5_2_1_U9.top_add_5ns_5ns_5_2_1_Adder_7_U.ce  ? \add_5ns_5ns_5_2_1_U9.top_add_5ns_5ns_5_2_1_Adder_7_U.b [4:2] : \add_5ns_5ns_5_2_1_U9.top_add_5ns_5ns_5_2_1_Adder_7_U.bin_s1 ;
assign _142_ = \add_5ns_5ns_5_2_1_U9.top_add_5ns_5ns_5_2_1_Adder_7_U.ce  ? \add_5ns_5ns_5_2_1_U9.top_add_5ns_5ns_5_2_1_Adder_7_U.a [4:2] : \add_5ns_5ns_5_2_1_U9.top_add_5ns_5ns_5_2_1_Adder_7_U.ain_s1 ;
assign _144_ = \add_5ns_5ns_5_2_1_U9.top_add_5ns_5ns_5_2_1_Adder_7_U.ce  ? \add_5ns_5ns_5_2_1_U9.top_add_5ns_5ns_5_2_1_Adder_7_U.facout_s1  : \add_5ns_5ns_5_2_1_U9.top_add_5ns_5ns_5_2_1_Adder_7_U.carry_s1 ;
assign _145_ = \add_5ns_5ns_5_2_1_U9.top_add_5ns_5ns_5_2_1_Adder_7_U.ce  ? \add_5ns_5ns_5_2_1_U9.top_add_5ns_5ns_5_2_1_Adder_7_U.fas_s1  : \add_5ns_5ns_5_2_1_U9.top_add_5ns_5ns_5_2_1_Adder_7_U.sum_s1 ;
assign _146_ = \add_5ns_5ns_5_2_1_U9.top_add_5ns_5ns_5_2_1_Adder_7_U.u1.a  + \add_5ns_5ns_5_2_1_U9.top_add_5ns_5ns_5_2_1_Adder_7_U.u1.b ;
assign { \add_5ns_5ns_5_2_1_U9.top_add_5ns_5ns_5_2_1_Adder_7_U.u1.cout , \add_5ns_5ns_5_2_1_U9.top_add_5ns_5ns_5_2_1_Adder_7_U.u1.s  } = _146_ + \add_5ns_5ns_5_2_1_U9.top_add_5ns_5ns_5_2_1_Adder_7_U.u1.cin ;
assign _147_ = \add_5ns_5ns_5_2_1_U9.top_add_5ns_5ns_5_2_1_Adder_7_U.u2.a  + \add_5ns_5ns_5_2_1_U9.top_add_5ns_5ns_5_2_1_Adder_7_U.u2.b ;
assign { \add_5ns_5ns_5_2_1_U9.top_add_5ns_5ns_5_2_1_Adder_7_U.u2.cout , \add_5ns_5ns_5_2_1_U9.top_add_5ns_5ns_5_2_1_Adder_7_U.u2.s  } = _147_ + \add_5ns_5ns_5_2_1_U9.top_add_5ns_5ns_5_2_1_Adder_7_U.u2.cin ;
always @(posedge \add_5s_5ns_5_2_1_U10.top_add_5s_5ns_5_2_1_Adder_8_U.clk )
\add_5s_5ns_5_2_1_U10.top_add_5s_5ns_5_2_1_Adder_8_U.bin_s1  <= _149_;
always @(posedge \add_5s_5ns_5_2_1_U10.top_add_5s_5ns_5_2_1_Adder_8_U.clk )
\add_5s_5ns_5_2_1_U10.top_add_5s_5ns_5_2_1_Adder_8_U.ain_s1  <= _148_;
always @(posedge \add_5s_5ns_5_2_1_U10.top_add_5s_5ns_5_2_1_Adder_8_U.clk )
\add_5s_5ns_5_2_1_U10.top_add_5s_5ns_5_2_1_Adder_8_U.sum_s1  <= _151_;
always @(posedge \add_5s_5ns_5_2_1_U10.top_add_5s_5ns_5_2_1_Adder_8_U.clk )
\add_5s_5ns_5_2_1_U10.top_add_5s_5ns_5_2_1_Adder_8_U.carry_s1  <= _150_;
assign _149_ = \add_5s_5ns_5_2_1_U10.top_add_5s_5ns_5_2_1_Adder_8_U.ce  ? \add_5s_5ns_5_2_1_U10.top_add_5s_5ns_5_2_1_Adder_8_U.b [4:2] : \add_5s_5ns_5_2_1_U10.top_add_5s_5ns_5_2_1_Adder_8_U.bin_s1 ;
assign _148_ = \add_5s_5ns_5_2_1_U10.top_add_5s_5ns_5_2_1_Adder_8_U.ce  ? \add_5s_5ns_5_2_1_U10.top_add_5s_5ns_5_2_1_Adder_8_U.a [4:2] : \add_5s_5ns_5_2_1_U10.top_add_5s_5ns_5_2_1_Adder_8_U.ain_s1 ;
assign _150_ = \add_5s_5ns_5_2_1_U10.top_add_5s_5ns_5_2_1_Adder_8_U.ce  ? \add_5s_5ns_5_2_1_U10.top_add_5s_5ns_5_2_1_Adder_8_U.facout_s1  : \add_5s_5ns_5_2_1_U10.top_add_5s_5ns_5_2_1_Adder_8_U.carry_s1 ;
assign _151_ = \add_5s_5ns_5_2_1_U10.top_add_5s_5ns_5_2_1_Adder_8_U.ce  ? \add_5s_5ns_5_2_1_U10.top_add_5s_5ns_5_2_1_Adder_8_U.fas_s1  : \add_5s_5ns_5_2_1_U10.top_add_5s_5ns_5_2_1_Adder_8_U.sum_s1 ;
assign _152_ = \add_5s_5ns_5_2_1_U10.top_add_5s_5ns_5_2_1_Adder_8_U.u1.a  + \add_5s_5ns_5_2_1_U10.top_add_5s_5ns_5_2_1_Adder_8_U.u1.b ;
assign { \add_5s_5ns_5_2_1_U10.top_add_5s_5ns_5_2_1_Adder_8_U.u1.cout , \add_5s_5ns_5_2_1_U10.top_add_5s_5ns_5_2_1_Adder_8_U.u1.s  } = _152_ + \add_5s_5ns_5_2_1_U10.top_add_5s_5ns_5_2_1_Adder_8_U.u1.cin ;
assign _153_ = \add_5s_5ns_5_2_1_U10.top_add_5s_5ns_5_2_1_Adder_8_U.u2.a  + \add_5s_5ns_5_2_1_U10.top_add_5s_5ns_5_2_1_Adder_8_U.u2.b ;
assign { \add_5s_5ns_5_2_1_U10.top_add_5s_5ns_5_2_1_Adder_8_U.u2.cout , \add_5s_5ns_5_2_1_U10.top_add_5s_5ns_5_2_1_Adder_8_U.u2.s  } = _153_ + \add_5s_5ns_5_2_1_U10.top_add_5s_5ns_5_2_1_Adder_8_U.u2.cin ;
always @(posedge \add_5s_5s_5_2_1_U22.top_add_5s_5s_5_2_1_Adder_15_U.clk )
\add_5s_5s_5_2_1_U22.top_add_5s_5s_5_2_1_Adder_15_U.bin_s1  <= _155_;
always @(posedge \add_5s_5s_5_2_1_U22.top_add_5s_5s_5_2_1_Adder_15_U.clk )
\add_5s_5s_5_2_1_U22.top_add_5s_5s_5_2_1_Adder_15_U.ain_s1  <= _154_;
always @(posedge \add_5s_5s_5_2_1_U22.top_add_5s_5s_5_2_1_Adder_15_U.clk )
\add_5s_5s_5_2_1_U22.top_add_5s_5s_5_2_1_Adder_15_U.sum_s1  <= _157_;
always @(posedge \add_5s_5s_5_2_1_U22.top_add_5s_5s_5_2_1_Adder_15_U.clk )
\add_5s_5s_5_2_1_U22.top_add_5s_5s_5_2_1_Adder_15_U.carry_s1  <= _156_;
assign _155_ = \add_5s_5s_5_2_1_U22.top_add_5s_5s_5_2_1_Adder_15_U.ce  ? \add_5s_5s_5_2_1_U22.top_add_5s_5s_5_2_1_Adder_15_U.b [4:2] : \add_5s_5s_5_2_1_U22.top_add_5s_5s_5_2_1_Adder_15_U.bin_s1 ;
assign _154_ = \add_5s_5s_5_2_1_U22.top_add_5s_5s_5_2_1_Adder_15_U.ce  ? \add_5s_5s_5_2_1_U22.top_add_5s_5s_5_2_1_Adder_15_U.a [4:2] : \add_5s_5s_5_2_1_U22.top_add_5s_5s_5_2_1_Adder_15_U.ain_s1 ;
assign _156_ = \add_5s_5s_5_2_1_U22.top_add_5s_5s_5_2_1_Adder_15_U.ce  ? \add_5s_5s_5_2_1_U22.top_add_5s_5s_5_2_1_Adder_15_U.facout_s1  : \add_5s_5s_5_2_1_U22.top_add_5s_5s_5_2_1_Adder_15_U.carry_s1 ;
assign _157_ = \add_5s_5s_5_2_1_U22.top_add_5s_5s_5_2_1_Adder_15_U.ce  ? \add_5s_5s_5_2_1_U22.top_add_5s_5s_5_2_1_Adder_15_U.fas_s1  : \add_5s_5s_5_2_1_U22.top_add_5s_5s_5_2_1_Adder_15_U.sum_s1 ;
assign _158_ = \add_5s_5s_5_2_1_U22.top_add_5s_5s_5_2_1_Adder_15_U.u1.a  + \add_5s_5s_5_2_1_U22.top_add_5s_5s_5_2_1_Adder_15_U.u1.b ;
assign { \add_5s_5s_5_2_1_U22.top_add_5s_5s_5_2_1_Adder_15_U.u1.cout , \add_5s_5s_5_2_1_U22.top_add_5s_5s_5_2_1_Adder_15_U.u1.s  } = _158_ + \add_5s_5s_5_2_1_U22.top_add_5s_5s_5_2_1_Adder_15_U.u1.cin ;
assign _159_ = \add_5s_5s_5_2_1_U22.top_add_5s_5s_5_2_1_Adder_15_U.u2.a  + \add_5s_5s_5_2_1_U22.top_add_5s_5s_5_2_1_Adder_15_U.u2.b ;
assign { \add_5s_5s_5_2_1_U22.top_add_5s_5s_5_2_1_Adder_15_U.u2.cout , \add_5s_5s_5_2_1_U22.top_add_5s_5s_5_2_1_Adder_15_U.u2.s  } = _159_ + \add_5s_5s_5_2_1_U22.top_add_5s_5s_5_2_1_Adder_15_U.u2.cin ;
always @(posedge \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_5_U.clk )
\add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_5_U.bin_s1  <= _161_;
always @(posedge \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_5_U.clk )
\add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_5_U.ain_s1  <= _160_;
always @(posedge \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_5_U.clk )
\add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_5_U.sum_s1  <= _163_;
always @(posedge \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_5_U.clk )
\add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_5_U.carry_s1  <= _162_;
assign _161_ = \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_5_U.ce  ? \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_5_U.b [7:4] : \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_5_U.bin_s1 ;
assign _160_ = \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_5_U.ce  ? \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_5_U.a [7:4] : \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_5_U.ain_s1 ;
assign _162_ = \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_5_U.ce  ? \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_5_U.facout_s1  : \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_5_U.carry_s1 ;
assign _163_ = \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_5_U.ce  ? \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_5_U.fas_s1  : \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_5_U.sum_s1 ;
assign _164_ = \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_5_U.u1.a  + \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_5_U.u1.b ;
assign { \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_5_U.u1.cout , \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_5_U.u1.s  } = _164_ + \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_5_U.u1.cin ;
assign _165_ = \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_5_U.u2.a  + \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_5_U.u2.b ;
assign { \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_5_U.u2.cout , \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_5_U.u2.s  } = _165_ + \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_5_U.u2.cin ;
always @(posedge \add_9s_9s_9_2_1_U13.top_add_9s_9s_9_2_1_Adder_4_U.clk )
\add_9s_9s_9_2_1_U13.top_add_9s_9s_9_2_1_Adder_4_U.bin_s1  <= _167_;
always @(posedge \add_9s_9s_9_2_1_U13.top_add_9s_9s_9_2_1_Adder_4_U.clk )
\add_9s_9s_9_2_1_U13.top_add_9s_9s_9_2_1_Adder_4_U.ain_s1  <= _166_;
always @(posedge \add_9s_9s_9_2_1_U13.top_add_9s_9s_9_2_1_Adder_4_U.clk )
\add_9s_9s_9_2_1_U13.top_add_9s_9s_9_2_1_Adder_4_U.sum_s1  <= _169_;
always @(posedge \add_9s_9s_9_2_1_U13.top_add_9s_9s_9_2_1_Adder_4_U.clk )
\add_9s_9s_9_2_1_U13.top_add_9s_9s_9_2_1_Adder_4_U.carry_s1  <= _168_;
assign _167_ = \add_9s_9s_9_2_1_U13.top_add_9s_9s_9_2_1_Adder_4_U.ce  ? \add_9s_9s_9_2_1_U13.top_add_9s_9s_9_2_1_Adder_4_U.b [8:4] : \add_9s_9s_9_2_1_U13.top_add_9s_9s_9_2_1_Adder_4_U.bin_s1 ;
assign _166_ = \add_9s_9s_9_2_1_U13.top_add_9s_9s_9_2_1_Adder_4_U.ce  ? \add_9s_9s_9_2_1_U13.top_add_9s_9s_9_2_1_Adder_4_U.a [8:4] : \add_9s_9s_9_2_1_U13.top_add_9s_9s_9_2_1_Adder_4_U.ain_s1 ;
assign _168_ = \add_9s_9s_9_2_1_U13.top_add_9s_9s_9_2_1_Adder_4_U.ce  ? \add_9s_9s_9_2_1_U13.top_add_9s_9s_9_2_1_Adder_4_U.facout_s1  : \add_9s_9s_9_2_1_U13.top_add_9s_9s_9_2_1_Adder_4_U.carry_s1 ;
assign _169_ = \add_9s_9s_9_2_1_U13.top_add_9s_9s_9_2_1_Adder_4_U.ce  ? \add_9s_9s_9_2_1_U13.top_add_9s_9s_9_2_1_Adder_4_U.fas_s1  : \add_9s_9s_9_2_1_U13.top_add_9s_9s_9_2_1_Adder_4_U.sum_s1 ;
assign _170_ = \add_9s_9s_9_2_1_U13.top_add_9s_9s_9_2_1_Adder_4_U.u1.a  + \add_9s_9s_9_2_1_U13.top_add_9s_9s_9_2_1_Adder_4_U.u1.b ;
assign { \add_9s_9s_9_2_1_U13.top_add_9s_9s_9_2_1_Adder_4_U.u1.cout , \add_9s_9s_9_2_1_U13.top_add_9s_9s_9_2_1_Adder_4_U.u1.s  } = _170_ + \add_9s_9s_9_2_1_U13.top_add_9s_9s_9_2_1_Adder_4_U.u1.cin ;
assign _171_ = \add_9s_9s_9_2_1_U13.top_add_9s_9s_9_2_1_Adder_4_U.u2.a  + \add_9s_9s_9_2_1_U13.top_add_9s_9s_9_2_1_Adder_4_U.u2.b ;
assign { \add_9s_9s_9_2_1_U13.top_add_9s_9s_9_2_1_Adder_4_U.u2.cout , \add_9s_9s_9_2_1_U13.top_add_9s_9s_9_2_1_Adder_4_U.u2.s  } = _171_ + \add_9s_9s_9_2_1_U13.top_add_9s_9s_9_2_1_Adder_4_U.u2.cin ;
always @(posedge \add_9s_9s_9_2_1_U6.top_add_9s_9s_9_2_1_Adder_4_U.clk )
\add_9s_9s_9_2_1_U6.top_add_9s_9s_9_2_1_Adder_4_U.bin_s1  <= _173_;
always @(posedge \add_9s_9s_9_2_1_U6.top_add_9s_9s_9_2_1_Adder_4_U.clk )
\add_9s_9s_9_2_1_U6.top_add_9s_9s_9_2_1_Adder_4_U.ain_s1  <= _172_;
always @(posedge \add_9s_9s_9_2_1_U6.top_add_9s_9s_9_2_1_Adder_4_U.clk )
\add_9s_9s_9_2_1_U6.top_add_9s_9s_9_2_1_Adder_4_U.sum_s1  <= _175_;
always @(posedge \add_9s_9s_9_2_1_U6.top_add_9s_9s_9_2_1_Adder_4_U.clk )
\add_9s_9s_9_2_1_U6.top_add_9s_9s_9_2_1_Adder_4_U.carry_s1  <= _174_;
assign _173_ = \add_9s_9s_9_2_1_U6.top_add_9s_9s_9_2_1_Adder_4_U.ce  ? \add_9s_9s_9_2_1_U6.top_add_9s_9s_9_2_1_Adder_4_U.b [8:4] : \add_9s_9s_9_2_1_U6.top_add_9s_9s_9_2_1_Adder_4_U.bin_s1 ;
assign _172_ = \add_9s_9s_9_2_1_U6.top_add_9s_9s_9_2_1_Adder_4_U.ce  ? \add_9s_9s_9_2_1_U6.top_add_9s_9s_9_2_1_Adder_4_U.a [8:4] : \add_9s_9s_9_2_1_U6.top_add_9s_9s_9_2_1_Adder_4_U.ain_s1 ;
assign _174_ = \add_9s_9s_9_2_1_U6.top_add_9s_9s_9_2_1_Adder_4_U.ce  ? \add_9s_9s_9_2_1_U6.top_add_9s_9s_9_2_1_Adder_4_U.facout_s1  : \add_9s_9s_9_2_1_U6.top_add_9s_9s_9_2_1_Adder_4_U.carry_s1 ;
assign _175_ = \add_9s_9s_9_2_1_U6.top_add_9s_9s_9_2_1_Adder_4_U.ce  ? \add_9s_9s_9_2_1_U6.top_add_9s_9s_9_2_1_Adder_4_U.fas_s1  : \add_9s_9s_9_2_1_U6.top_add_9s_9s_9_2_1_Adder_4_U.sum_s1 ;
assign _176_ = \add_9s_9s_9_2_1_U6.top_add_9s_9s_9_2_1_Adder_4_U.u1.a  + \add_9s_9s_9_2_1_U6.top_add_9s_9s_9_2_1_Adder_4_U.u1.b ;
assign { \add_9s_9s_9_2_1_U6.top_add_9s_9s_9_2_1_Adder_4_U.u1.cout , \add_9s_9s_9_2_1_U6.top_add_9s_9s_9_2_1_Adder_4_U.u1.s  } = _176_ + \add_9s_9s_9_2_1_U6.top_add_9s_9s_9_2_1_Adder_4_U.u1.cin ;
assign _177_ = \add_9s_9s_9_2_1_U6.top_add_9s_9s_9_2_1_Adder_4_U.u2.a  + \add_9s_9s_9_2_1_U6.top_add_9s_9s_9_2_1_Adder_4_U.u2.b ;
assign { \add_9s_9s_9_2_1_U6.top_add_9s_9s_9_2_1_Adder_4_U.u2.cout , \add_9s_9s_9_2_1_U6.top_add_9s_9s_9_2_1_Adder_4_U.u2.s  } = _177_ + \add_9s_9s_9_2_1_U6.top_add_9s_9s_9_2_1_Adder_4_U.u2.cin ;
always @(posedge \ashr_32s_32s_32_7_1_U16.clk )
\ashr_32s_32s_32_7_1_U16.dout_array[5]  <= _189_;
always @(posedge \ashr_32s_32s_32_7_1_U16.clk )
\ashr_32s_32s_32_7_1_U16.din1_cast_array[5]  <= _183_;
always @(posedge \ashr_32s_32s_32_7_1_U16.clk )
\ashr_32s_32s_32_7_1_U16.dout_array[4]  <= _188_;
always @(posedge \ashr_32s_32s_32_7_1_U16.clk )
\ashr_32s_32s_32_7_1_U16.din1_cast_array[4]  <= _182_;
always @(posedge \ashr_32s_32s_32_7_1_U16.clk )
\ashr_32s_32s_32_7_1_U16.dout_array[3]  <= _187_;
always @(posedge \ashr_32s_32s_32_7_1_U16.clk )
\ashr_32s_32s_32_7_1_U16.din1_cast_array[3]  <= _181_;
always @(posedge \ashr_32s_32s_32_7_1_U16.clk )
\ashr_32s_32s_32_7_1_U16.dout_array[2]  <= _186_;
always @(posedge \ashr_32s_32s_32_7_1_U16.clk )
\ashr_32s_32s_32_7_1_U16.din1_cast_array[2]  <= _180_;
always @(posedge \ashr_32s_32s_32_7_1_U16.clk )
\ashr_32s_32s_32_7_1_U16.dout_array[1]  <= _185_;
always @(posedge \ashr_32s_32s_32_7_1_U16.clk )
\ashr_32s_32s_32_7_1_U16.din1_cast_array[1]  <= _179_;
always @(posedge \ashr_32s_32s_32_7_1_U16.clk )
\ashr_32s_32s_32_7_1_U16.dout_array[0]  <= _184_;
always @(posedge \ashr_32s_32s_32_7_1_U16.clk )
\ashr_32s_32s_32_7_1_U16.din1_cast_array[0]  <= _178_;
assign _190_ = \ashr_32s_32s_32_7_1_U16.ce  ? \ashr_32s_32s_32_7_1_U16.din1_cast_array[4]  : \ashr_32s_32s_32_7_1_U16.din1_cast_array[5] ;
assign _183_ = \ashr_32s_32s_32_7_1_U16.reset  ? 32'd0 : _190_;
assign _191_ = \ashr_32s_32s_32_7_1_U16.ce  ? _207_ : \ashr_32s_32s_32_7_1_U16.dout_array[5] ;
assign _189_ = \ashr_32s_32s_32_7_1_U16.reset  ? 32'd0 : _191_;
assign _192_ = \ashr_32s_32s_32_7_1_U16.ce  ? \ashr_32s_32s_32_7_1_U16.din1_cast_array[3]  : \ashr_32s_32s_32_7_1_U16.din1_cast_array[4] ;
assign _182_ = \ashr_32s_32s_32_7_1_U16.reset  ? 32'd0 : _192_;
assign _193_ = \ashr_32s_32s_32_7_1_U16.ce  ? _206_ : \ashr_32s_32s_32_7_1_U16.dout_array[4] ;
assign _188_ = \ashr_32s_32s_32_7_1_U16.reset  ? 32'd0 : _193_;
assign _194_ = \ashr_32s_32s_32_7_1_U16.ce  ? \ashr_32s_32s_32_7_1_U16.din1_cast_array[2]  : \ashr_32s_32s_32_7_1_U16.din1_cast_array[3] ;
assign _181_ = \ashr_32s_32s_32_7_1_U16.reset  ? 32'd0 : _194_;
assign _195_ = \ashr_32s_32s_32_7_1_U16.ce  ? _205_ : \ashr_32s_32s_32_7_1_U16.dout_array[3] ;
assign _187_ = \ashr_32s_32s_32_7_1_U16.reset  ? 32'd0 : _195_;
assign _196_ = \ashr_32s_32s_32_7_1_U16.ce  ? \ashr_32s_32s_32_7_1_U16.din1_cast_array[1]  : \ashr_32s_32s_32_7_1_U16.din1_cast_array[2] ;
assign _180_ = \ashr_32s_32s_32_7_1_U16.reset  ? 32'd0 : _196_;
assign _197_ = \ashr_32s_32s_32_7_1_U16.ce  ? _204_ : \ashr_32s_32s_32_7_1_U16.dout_array[2] ;
assign _186_ = \ashr_32s_32s_32_7_1_U16.reset  ? 32'd0 : _197_;
assign _198_ = \ashr_32s_32s_32_7_1_U16.ce  ? \ashr_32s_32s_32_7_1_U16.din1_cast_array[0]  : \ashr_32s_32s_32_7_1_U16.din1_cast_array[1] ;
assign _179_ = \ashr_32s_32s_32_7_1_U16.reset  ? 32'd0 : _198_;
assign _199_ = \ashr_32s_32s_32_7_1_U16.ce  ? _203_ : \ashr_32s_32s_32_7_1_U16.dout_array[1] ;
assign _185_ = \ashr_32s_32s_32_7_1_U16.reset  ? 32'd0 : _199_;
assign _200_ = \ashr_32s_32s_32_7_1_U16.ce  ? \ashr_32s_32s_32_7_1_U16.din1  : \ashr_32s_32s_32_7_1_U16.din1_cast_array[0] ;
assign _178_ = \ashr_32s_32s_32_7_1_U16.reset  ? 32'd0 : _200_;
assign _201_ = \ashr_32s_32s_32_7_1_U16.ce  ? _202_ : \ashr_32s_32s_32_7_1_U16.dout_array[0] ;
assign _184_ = \ashr_32s_32s_32_7_1_U16.reset  ? 32'd0 : _201_;
assign _202_ = $signed(\ashr_32s_32s_32_7_1_U16.din0 ) >>> { \ashr_32s_32s_32_7_1_U16.din1 [31:30], 30'h00000000 };
assign _203_ = $signed(\ashr_32s_32s_32_7_1_U16.dout_array[0] ) >>> { \ashr_32s_32s_32_7_1_U16.din1_cast_array[0] [29:25], 25'h0000000 };
assign _204_ = $signed(\ashr_32s_32s_32_7_1_U16.dout_array[1] ) >>> { \ashr_32s_32s_32_7_1_U16.din1_cast_array[1] [24:20], 20'h00000 };
assign _205_ = $signed(\ashr_32s_32s_32_7_1_U16.dout_array[2] ) >>> { \ashr_32s_32s_32_7_1_U16.din1_cast_array[2] [19:15], 15'h0000 };
assign _206_ = $signed(\ashr_32s_32s_32_7_1_U16.dout_array[3] ) >>> { \ashr_32s_32s_32_7_1_U16.din1_cast_array[3] [14:10], 10'h000 };
assign _207_ = $signed(\ashr_32s_32s_32_7_1_U16.dout_array[4] ) >>> { \ashr_32s_32s_32_7_1_U16.din1_cast_array[4] [9:5], 5'h00 };
assign \ashr_32s_32s_32_7_1_U16.dout  = $signed(\ashr_32s_32s_32_7_1_U16.dout_array[5] ) >>> \ashr_32s_32s_32_7_1_U16.din1_cast_array[5] [4:0];
assign \mul_32s_4s_36_7_1_U4.top_mul_32s_4s_36_7_1_Mul_DSP_0_U.tmp_product  = $signed(\mul_32s_4s_36_7_1_U4.top_mul_32s_4s_36_7_1_Mul_DSP_0_U.a_reg0 ) * $signed(\mul_32s_4s_36_7_1_U4.top_mul_32s_4s_36_7_1_Mul_DSP_0_U.b_reg0 );
always @(posedge \mul_32s_4s_36_7_1_U4.top_mul_32s_4s_36_7_1_Mul_DSP_0_U.clk )
\mul_32s_4s_36_7_1_U4.top_mul_32s_4s_36_7_1_Mul_DSP_0_U.a_reg0  <= _208_;
always @(posedge \mul_32s_4s_36_7_1_U4.top_mul_32s_4s_36_7_1_Mul_DSP_0_U.clk )
\mul_32s_4s_36_7_1_U4.top_mul_32s_4s_36_7_1_Mul_DSP_0_U.b_reg0  <= _209_;
always @(posedge \mul_32s_4s_36_7_1_U4.top_mul_32s_4s_36_7_1_Mul_DSP_0_U.clk )
\mul_32s_4s_36_7_1_U4.top_mul_32s_4s_36_7_1_Mul_DSP_0_U.buff0  <= _210_;
always @(posedge \mul_32s_4s_36_7_1_U4.top_mul_32s_4s_36_7_1_Mul_DSP_0_U.clk )
\mul_32s_4s_36_7_1_U4.top_mul_32s_4s_36_7_1_Mul_DSP_0_U.buff1  <= _211_;
always @(posedge \mul_32s_4s_36_7_1_U4.top_mul_32s_4s_36_7_1_Mul_DSP_0_U.clk )
\mul_32s_4s_36_7_1_U4.top_mul_32s_4s_36_7_1_Mul_DSP_0_U.buff2  <= _212_;
always @(posedge \mul_32s_4s_36_7_1_U4.top_mul_32s_4s_36_7_1_Mul_DSP_0_U.clk )
\mul_32s_4s_36_7_1_U4.top_mul_32s_4s_36_7_1_Mul_DSP_0_U.buff3  <= _213_;
always @(posedge \mul_32s_4s_36_7_1_U4.top_mul_32s_4s_36_7_1_Mul_DSP_0_U.clk )
\mul_32s_4s_36_7_1_U4.top_mul_32s_4s_36_7_1_Mul_DSP_0_U.buff4  <= _214_;
assign _214_ = \mul_32s_4s_36_7_1_U4.top_mul_32s_4s_36_7_1_Mul_DSP_0_U.ce  ? \mul_32s_4s_36_7_1_U4.top_mul_32s_4s_36_7_1_Mul_DSP_0_U.buff3  : \mul_32s_4s_36_7_1_U4.top_mul_32s_4s_36_7_1_Mul_DSP_0_U.buff4 ;
assign _213_ = \mul_32s_4s_36_7_1_U4.top_mul_32s_4s_36_7_1_Mul_DSP_0_U.ce  ? \mul_32s_4s_36_7_1_U4.top_mul_32s_4s_36_7_1_Mul_DSP_0_U.buff2  : \mul_32s_4s_36_7_1_U4.top_mul_32s_4s_36_7_1_Mul_DSP_0_U.buff3 ;
assign _212_ = \mul_32s_4s_36_7_1_U4.top_mul_32s_4s_36_7_1_Mul_DSP_0_U.ce  ? \mul_32s_4s_36_7_1_U4.top_mul_32s_4s_36_7_1_Mul_DSP_0_U.buff1  : \mul_32s_4s_36_7_1_U4.top_mul_32s_4s_36_7_1_Mul_DSP_0_U.buff2 ;
assign _211_ = \mul_32s_4s_36_7_1_U4.top_mul_32s_4s_36_7_1_Mul_DSP_0_U.ce  ? \mul_32s_4s_36_7_1_U4.top_mul_32s_4s_36_7_1_Mul_DSP_0_U.buff0  : \mul_32s_4s_36_7_1_U4.top_mul_32s_4s_36_7_1_Mul_DSP_0_U.buff1 ;
assign _210_ = \mul_32s_4s_36_7_1_U4.top_mul_32s_4s_36_7_1_Mul_DSP_0_U.ce  ? \mul_32s_4s_36_7_1_U4.top_mul_32s_4s_36_7_1_Mul_DSP_0_U.tmp_product  : \mul_32s_4s_36_7_1_U4.top_mul_32s_4s_36_7_1_Mul_DSP_0_U.buff0 ;
assign _209_ = \mul_32s_4s_36_7_1_U4.top_mul_32s_4s_36_7_1_Mul_DSP_0_U.ce  ? \mul_32s_4s_36_7_1_U4.top_mul_32s_4s_36_7_1_Mul_DSP_0_U.b  : \mul_32s_4s_36_7_1_U4.top_mul_32s_4s_36_7_1_Mul_DSP_0_U.b_reg0 ;
assign _208_ = \mul_32s_4s_36_7_1_U4.top_mul_32s_4s_36_7_1_Mul_DSP_0_U.ce  ? \mul_32s_4s_36_7_1_U4.top_mul_32s_4s_36_7_1_Mul_DSP_0_U.a  : \mul_32s_4s_36_7_1_U4.top_mul_32s_4s_36_7_1_Mul_DSP_0_U.a_reg0 ;
always @(posedge \shl_32s_32s_32_7_1_U17.clk )
\shl_32s_32s_32_7_1_U17.dout_array[5]  <= _226_;
always @(posedge \shl_32s_32s_32_7_1_U17.clk )
\shl_32s_32s_32_7_1_U17.din1_cast_array[5]  <= _220_;
always @(posedge \shl_32s_32s_32_7_1_U17.clk )
\shl_32s_32s_32_7_1_U17.dout_array[4]  <= _225_;
always @(posedge \shl_32s_32s_32_7_1_U17.clk )
\shl_32s_32s_32_7_1_U17.din1_cast_array[4]  <= _219_;
always @(posedge \shl_32s_32s_32_7_1_U17.clk )
\shl_32s_32s_32_7_1_U17.dout_array[3]  <= _224_;
always @(posedge \shl_32s_32s_32_7_1_U17.clk )
\shl_32s_32s_32_7_1_U17.din1_cast_array[3]  <= _218_;
always @(posedge \shl_32s_32s_32_7_1_U17.clk )
\shl_32s_32s_32_7_1_U17.dout_array[2]  <= _223_;
always @(posedge \shl_32s_32s_32_7_1_U17.clk )
\shl_32s_32s_32_7_1_U17.din1_cast_array[2]  <= _217_;
always @(posedge \shl_32s_32s_32_7_1_U17.clk )
\shl_32s_32s_32_7_1_U17.dout_array[1]  <= _222_;
always @(posedge \shl_32s_32s_32_7_1_U17.clk )
\shl_32s_32s_32_7_1_U17.din1_cast_array[1]  <= _216_;
always @(posedge \shl_32s_32s_32_7_1_U17.clk )
\shl_32s_32s_32_7_1_U17.dout_array[0]  <= _221_;
always @(posedge \shl_32s_32s_32_7_1_U17.clk )
\shl_32s_32s_32_7_1_U17.din1_cast_array[0]  <= _215_;
assign _227_ = \shl_32s_32s_32_7_1_U17.ce  ? \shl_32s_32s_32_7_1_U17.din1_cast_array[4]  : \shl_32s_32s_32_7_1_U17.din1_cast_array[5] ;
assign _220_ = \shl_32s_32s_32_7_1_U17.reset  ? 32'd0 : _227_;
assign _228_ = \shl_32s_32s_32_7_1_U17.ce  ? _244_ : \shl_32s_32s_32_7_1_U17.dout_array[5] ;
assign _226_ = \shl_32s_32s_32_7_1_U17.reset  ? 32'd0 : _228_;
assign _229_ = \shl_32s_32s_32_7_1_U17.ce  ? \shl_32s_32s_32_7_1_U17.din1_cast_array[3]  : \shl_32s_32s_32_7_1_U17.din1_cast_array[4] ;
assign _219_ = \shl_32s_32s_32_7_1_U17.reset  ? 32'd0 : _229_;
assign _230_ = \shl_32s_32s_32_7_1_U17.ce  ? _243_ : \shl_32s_32s_32_7_1_U17.dout_array[4] ;
assign _225_ = \shl_32s_32s_32_7_1_U17.reset  ? 32'd0 : _230_;
assign _231_ = \shl_32s_32s_32_7_1_U17.ce  ? \shl_32s_32s_32_7_1_U17.din1_cast_array[2]  : \shl_32s_32s_32_7_1_U17.din1_cast_array[3] ;
assign _218_ = \shl_32s_32s_32_7_1_U17.reset  ? 32'd0 : _231_;
assign _232_ = \shl_32s_32s_32_7_1_U17.ce  ? _242_ : \shl_32s_32s_32_7_1_U17.dout_array[3] ;
assign _224_ = \shl_32s_32s_32_7_1_U17.reset  ? 32'd0 : _232_;
assign _233_ = \shl_32s_32s_32_7_1_U17.ce  ? \shl_32s_32s_32_7_1_U17.din1_cast_array[1]  : \shl_32s_32s_32_7_1_U17.din1_cast_array[2] ;
assign _217_ = \shl_32s_32s_32_7_1_U17.reset  ? 32'd0 : _233_;
assign _234_ = \shl_32s_32s_32_7_1_U17.ce  ? _241_ : \shl_32s_32s_32_7_1_U17.dout_array[2] ;
assign _223_ = \shl_32s_32s_32_7_1_U17.reset  ? 32'd0 : _234_;
assign _235_ = \shl_32s_32s_32_7_1_U17.ce  ? \shl_32s_32s_32_7_1_U17.din1_cast_array[0]  : \shl_32s_32s_32_7_1_U17.din1_cast_array[1] ;
assign _216_ = \shl_32s_32s_32_7_1_U17.reset  ? 32'd0 : _235_;
assign _236_ = \shl_32s_32s_32_7_1_U17.ce  ? _240_ : \shl_32s_32s_32_7_1_U17.dout_array[1] ;
assign _222_ = \shl_32s_32s_32_7_1_U17.reset  ? 32'd0 : _236_;
assign _237_ = \shl_32s_32s_32_7_1_U17.ce  ? \shl_32s_32s_32_7_1_U17.din1  : \shl_32s_32s_32_7_1_U17.din1_cast_array[0] ;
assign _215_ = \shl_32s_32s_32_7_1_U17.reset  ? 32'd0 : _237_;
assign _238_ = \shl_32s_32s_32_7_1_U17.ce  ? _239_ : \shl_32s_32s_32_7_1_U17.dout_array[0] ;
assign _221_ = \shl_32s_32s_32_7_1_U17.reset  ? 32'd0 : _238_;
assign _239_ = \shl_32s_32s_32_7_1_U17.din0  << { \shl_32s_32s_32_7_1_U17.din1 [31:30], 30'h00000000 };
assign _240_ = \shl_32s_32s_32_7_1_U17.dout_array[0]  << { \shl_32s_32s_32_7_1_U17.din1_cast_array[0] [29:25], 25'h0000000 };
assign _241_ = \shl_32s_32s_32_7_1_U17.dout_array[1]  << { \shl_32s_32s_32_7_1_U17.din1_cast_array[1] [24:20], 20'h00000 };
assign _242_ = \shl_32s_32s_32_7_1_U17.dout_array[2]  << { \shl_32s_32s_32_7_1_U17.din1_cast_array[2] [19:15], 15'h0000 };
assign _243_ = \shl_32s_32s_32_7_1_U17.dout_array[3]  << { \shl_32s_32s_32_7_1_U17.din1_cast_array[3] [14:10], 10'h000 };
assign _244_ = \shl_32s_32s_32_7_1_U17.dout_array[4]  << { \shl_32s_32s_32_7_1_U17.din1_cast_array[4] [9:5], 5'h00 };
assign \shl_32s_32s_32_7_1_U17.dout  = \shl_32s_32s_32_7_1_U17.dout_array[5]  << \shl_32s_32s_32_7_1_U17.din1_cast_array[5] [4:0];
assign \sub_16ns_16s_16_2_1_U2.top_sub_16ns_16s_16_2_1_Adder_1_U.bin_s0  = ~ \sub_16ns_16s_16_2_1_U2.top_sub_16ns_16s_16_2_1_Adder_1_U.b ;
always @(posedge \sub_16ns_16s_16_2_1_U2.top_sub_16ns_16s_16_2_1_Adder_1_U.clk )
\sub_16ns_16s_16_2_1_U2.top_sub_16ns_16s_16_2_1_Adder_1_U.bin_s1  <= _246_;
always @(posedge \sub_16ns_16s_16_2_1_U2.top_sub_16ns_16s_16_2_1_Adder_1_U.clk )
\sub_16ns_16s_16_2_1_U2.top_sub_16ns_16s_16_2_1_Adder_1_U.ain_s1  <= _245_;
always @(posedge \sub_16ns_16s_16_2_1_U2.top_sub_16ns_16s_16_2_1_Adder_1_U.clk )
\sub_16ns_16s_16_2_1_U2.top_sub_16ns_16s_16_2_1_Adder_1_U.sum_s1  <= _248_;
always @(posedge \sub_16ns_16s_16_2_1_U2.top_sub_16ns_16s_16_2_1_Adder_1_U.clk )
\sub_16ns_16s_16_2_1_U2.top_sub_16ns_16s_16_2_1_Adder_1_U.carry_s1  <= _247_;
assign _246_ = \sub_16ns_16s_16_2_1_U2.top_sub_16ns_16s_16_2_1_Adder_1_U.ce  ? \sub_16ns_16s_16_2_1_U2.top_sub_16ns_16s_16_2_1_Adder_1_U.bin_s0 [15:8] : \sub_16ns_16s_16_2_1_U2.top_sub_16ns_16s_16_2_1_Adder_1_U.bin_s1 ;
assign _245_ = \sub_16ns_16s_16_2_1_U2.top_sub_16ns_16s_16_2_1_Adder_1_U.ce  ? \sub_16ns_16s_16_2_1_U2.top_sub_16ns_16s_16_2_1_Adder_1_U.a [15:8] : \sub_16ns_16s_16_2_1_U2.top_sub_16ns_16s_16_2_1_Adder_1_U.ain_s1 ;
assign _247_ = \sub_16ns_16s_16_2_1_U2.top_sub_16ns_16s_16_2_1_Adder_1_U.ce  ? \sub_16ns_16s_16_2_1_U2.top_sub_16ns_16s_16_2_1_Adder_1_U.facout_s1  : \sub_16ns_16s_16_2_1_U2.top_sub_16ns_16s_16_2_1_Adder_1_U.carry_s1 ;
assign _248_ = \sub_16ns_16s_16_2_1_U2.top_sub_16ns_16s_16_2_1_Adder_1_U.ce  ? \sub_16ns_16s_16_2_1_U2.top_sub_16ns_16s_16_2_1_Adder_1_U.fas_s1  : \sub_16ns_16s_16_2_1_U2.top_sub_16ns_16s_16_2_1_Adder_1_U.sum_s1 ;
assign _249_ = \sub_16ns_16s_16_2_1_U2.top_sub_16ns_16s_16_2_1_Adder_1_U.u1.a  + \sub_16ns_16s_16_2_1_U2.top_sub_16ns_16s_16_2_1_Adder_1_U.u1.b ;
assign { \sub_16ns_16s_16_2_1_U2.top_sub_16ns_16s_16_2_1_Adder_1_U.u1.cout , \sub_16ns_16s_16_2_1_U2.top_sub_16ns_16s_16_2_1_Adder_1_U.u1.s  } = _249_ + \sub_16ns_16s_16_2_1_U2.top_sub_16ns_16s_16_2_1_Adder_1_U.u1.cin ;
assign _250_ = \sub_16ns_16s_16_2_1_U2.top_sub_16ns_16s_16_2_1_Adder_1_U.u2.a  + \sub_16ns_16s_16_2_1_U2.top_sub_16ns_16s_16_2_1_Adder_1_U.u2.b ;
assign { \sub_16ns_16s_16_2_1_U2.top_sub_16ns_16s_16_2_1_Adder_1_U.u2.cout , \sub_16ns_16s_16_2_1_U2.top_sub_16ns_16s_16_2_1_Adder_1_U.u2.s  } = _250_ + \sub_16ns_16s_16_2_1_U2.top_sub_16ns_16s_16_2_1_Adder_1_U.u2.cin ;
assign \sub_33s_33s_33_2_1_U5.top_sub_33s_33s_33_2_1_Adder_3_U.bin_s0  = ~ \sub_33s_33s_33_2_1_U5.top_sub_33s_33s_33_2_1_Adder_3_U.b ;
always @(posedge \sub_33s_33s_33_2_1_U5.top_sub_33s_33s_33_2_1_Adder_3_U.clk )
\sub_33s_33s_33_2_1_U5.top_sub_33s_33s_33_2_1_Adder_3_U.bin_s1  <= _252_;
always @(posedge \sub_33s_33s_33_2_1_U5.top_sub_33s_33s_33_2_1_Adder_3_U.clk )
\sub_33s_33s_33_2_1_U5.top_sub_33s_33s_33_2_1_Adder_3_U.ain_s1  <= _251_;
always @(posedge \sub_33s_33s_33_2_1_U5.top_sub_33s_33s_33_2_1_Adder_3_U.clk )
\sub_33s_33s_33_2_1_U5.top_sub_33s_33s_33_2_1_Adder_3_U.sum_s1  <= _254_;
always @(posedge \sub_33s_33s_33_2_1_U5.top_sub_33s_33s_33_2_1_Adder_3_U.clk )
\sub_33s_33s_33_2_1_U5.top_sub_33s_33s_33_2_1_Adder_3_U.carry_s1  <= _253_;
assign _252_ = \sub_33s_33s_33_2_1_U5.top_sub_33s_33s_33_2_1_Adder_3_U.ce  ? \sub_33s_33s_33_2_1_U5.top_sub_33s_33s_33_2_1_Adder_3_U.bin_s0 [32:16] : \sub_33s_33s_33_2_1_U5.top_sub_33s_33s_33_2_1_Adder_3_U.bin_s1 ;
assign _251_ = \sub_33s_33s_33_2_1_U5.top_sub_33s_33s_33_2_1_Adder_3_U.ce  ? \sub_33s_33s_33_2_1_U5.top_sub_33s_33s_33_2_1_Adder_3_U.a [32:16] : \sub_33s_33s_33_2_1_U5.top_sub_33s_33s_33_2_1_Adder_3_U.ain_s1 ;
assign _253_ = \sub_33s_33s_33_2_1_U5.top_sub_33s_33s_33_2_1_Adder_3_U.ce  ? \sub_33s_33s_33_2_1_U5.top_sub_33s_33s_33_2_1_Adder_3_U.facout_s1  : \sub_33s_33s_33_2_1_U5.top_sub_33s_33s_33_2_1_Adder_3_U.carry_s1 ;
assign _254_ = \sub_33s_33s_33_2_1_U5.top_sub_33s_33s_33_2_1_Adder_3_U.ce  ? \sub_33s_33s_33_2_1_U5.top_sub_33s_33s_33_2_1_Adder_3_U.fas_s1  : \sub_33s_33s_33_2_1_U5.top_sub_33s_33s_33_2_1_Adder_3_U.sum_s1 ;
assign _255_ = \sub_33s_33s_33_2_1_U5.top_sub_33s_33s_33_2_1_Adder_3_U.u1.a  + \sub_33s_33s_33_2_1_U5.top_sub_33s_33s_33_2_1_Adder_3_U.u1.b ;
assign { \sub_33s_33s_33_2_1_U5.top_sub_33s_33s_33_2_1_Adder_3_U.u1.cout , \sub_33s_33s_33_2_1_U5.top_sub_33s_33s_33_2_1_Adder_3_U.u1.s  } = _255_ + \sub_33s_33s_33_2_1_U5.top_sub_33s_33s_33_2_1_Adder_3_U.u1.cin ;
assign _256_ = \sub_33s_33s_33_2_1_U5.top_sub_33s_33s_33_2_1_Adder_3_U.u2.a  + \sub_33s_33s_33_2_1_U5.top_sub_33s_33s_33_2_1_Adder_3_U.u2.b ;
assign { \sub_33s_33s_33_2_1_U5.top_sub_33s_33s_33_2_1_Adder_3_U.u2.cout , \sub_33s_33s_33_2_1_U5.top_sub_33s_33s_33_2_1_Adder_3_U.u2.s  } = _256_ + \sub_33s_33s_33_2_1_U5.top_sub_33s_33s_33_2_1_Adder_3_U.u2.cin ;
assign \sub_6ns_6s_6_2_1_U14.top_sub_6ns_6s_6_2_1_Adder_10_U.bin_s0  = ~ \sub_6ns_6s_6_2_1_U14.top_sub_6ns_6s_6_2_1_Adder_10_U.b ;
always @(posedge \sub_6ns_6s_6_2_1_U14.top_sub_6ns_6s_6_2_1_Adder_10_U.clk )
\sub_6ns_6s_6_2_1_U14.top_sub_6ns_6s_6_2_1_Adder_10_U.bin_s1  <= _258_;
always @(posedge \sub_6ns_6s_6_2_1_U14.top_sub_6ns_6s_6_2_1_Adder_10_U.clk )
\sub_6ns_6s_6_2_1_U14.top_sub_6ns_6s_6_2_1_Adder_10_U.ain_s1  <= _257_;
always @(posedge \sub_6ns_6s_6_2_1_U14.top_sub_6ns_6s_6_2_1_Adder_10_U.clk )
\sub_6ns_6s_6_2_1_U14.top_sub_6ns_6s_6_2_1_Adder_10_U.sum_s1  <= _260_;
always @(posedge \sub_6ns_6s_6_2_1_U14.top_sub_6ns_6s_6_2_1_Adder_10_U.clk )
\sub_6ns_6s_6_2_1_U14.top_sub_6ns_6s_6_2_1_Adder_10_U.carry_s1  <= _259_;
assign _258_ = \sub_6ns_6s_6_2_1_U14.top_sub_6ns_6s_6_2_1_Adder_10_U.ce  ? \sub_6ns_6s_6_2_1_U14.top_sub_6ns_6s_6_2_1_Adder_10_U.bin_s0 [5:3] : \sub_6ns_6s_6_2_1_U14.top_sub_6ns_6s_6_2_1_Adder_10_U.bin_s1 ;
assign _257_ = \sub_6ns_6s_6_2_1_U14.top_sub_6ns_6s_6_2_1_Adder_10_U.ce  ? \sub_6ns_6s_6_2_1_U14.top_sub_6ns_6s_6_2_1_Adder_10_U.a [5:3] : \sub_6ns_6s_6_2_1_U14.top_sub_6ns_6s_6_2_1_Adder_10_U.ain_s1 ;
assign _259_ = \sub_6ns_6s_6_2_1_U14.top_sub_6ns_6s_6_2_1_Adder_10_U.ce  ? \sub_6ns_6s_6_2_1_U14.top_sub_6ns_6s_6_2_1_Adder_10_U.facout_s1  : \sub_6ns_6s_6_2_1_U14.top_sub_6ns_6s_6_2_1_Adder_10_U.carry_s1 ;
assign _260_ = \sub_6ns_6s_6_2_1_U14.top_sub_6ns_6s_6_2_1_Adder_10_U.ce  ? \sub_6ns_6s_6_2_1_U14.top_sub_6ns_6s_6_2_1_Adder_10_U.fas_s1  : \sub_6ns_6s_6_2_1_U14.top_sub_6ns_6s_6_2_1_Adder_10_U.sum_s1 ;
assign _261_ = \sub_6ns_6s_6_2_1_U14.top_sub_6ns_6s_6_2_1_Adder_10_U.u1.a  + \sub_6ns_6s_6_2_1_U14.top_sub_6ns_6s_6_2_1_Adder_10_U.u1.b ;
assign { \sub_6ns_6s_6_2_1_U14.top_sub_6ns_6s_6_2_1_Adder_10_U.u1.cout , \sub_6ns_6s_6_2_1_U14.top_sub_6ns_6s_6_2_1_Adder_10_U.u1.s  } = _261_ + \sub_6ns_6s_6_2_1_U14.top_sub_6ns_6s_6_2_1_Adder_10_U.u1.cin ;
assign _262_ = \sub_6ns_6s_6_2_1_U14.top_sub_6ns_6s_6_2_1_Adder_10_U.u2.a  + \sub_6ns_6s_6_2_1_U14.top_sub_6ns_6s_6_2_1_Adder_10_U.u2.b ;
assign { \sub_6ns_6s_6_2_1_U14.top_sub_6ns_6s_6_2_1_Adder_10_U.u2.cout , \sub_6ns_6s_6_2_1_U14.top_sub_6ns_6s_6_2_1_Adder_10_U.u2.s  } = _262_ + \sub_6ns_6s_6_2_1_U14.top_sub_6ns_6s_6_2_1_Adder_10_U.u2.cin ;
assign \sub_9s_9ns_9_2_1_U3.top_sub_9s_9ns_9_2_1_Adder_2_U.bin_s0  = ~ \sub_9s_9ns_9_2_1_U3.top_sub_9s_9ns_9_2_1_Adder_2_U.b ;
always @(posedge \sub_9s_9ns_9_2_1_U3.top_sub_9s_9ns_9_2_1_Adder_2_U.clk )
\sub_9s_9ns_9_2_1_U3.top_sub_9s_9ns_9_2_1_Adder_2_U.bin_s1  <= _264_;
always @(posedge \sub_9s_9ns_9_2_1_U3.top_sub_9s_9ns_9_2_1_Adder_2_U.clk )
\sub_9s_9ns_9_2_1_U3.top_sub_9s_9ns_9_2_1_Adder_2_U.ain_s1  <= _263_;
always @(posedge \sub_9s_9ns_9_2_1_U3.top_sub_9s_9ns_9_2_1_Adder_2_U.clk )
\sub_9s_9ns_9_2_1_U3.top_sub_9s_9ns_9_2_1_Adder_2_U.sum_s1  <= _266_;
always @(posedge \sub_9s_9ns_9_2_1_U3.top_sub_9s_9ns_9_2_1_Adder_2_U.clk )
\sub_9s_9ns_9_2_1_U3.top_sub_9s_9ns_9_2_1_Adder_2_U.carry_s1  <= _265_;
assign _264_ = \sub_9s_9ns_9_2_1_U3.top_sub_9s_9ns_9_2_1_Adder_2_U.ce  ? \sub_9s_9ns_9_2_1_U3.top_sub_9s_9ns_9_2_1_Adder_2_U.bin_s0 [8:4] : \sub_9s_9ns_9_2_1_U3.top_sub_9s_9ns_9_2_1_Adder_2_U.bin_s1 ;
assign _263_ = \sub_9s_9ns_9_2_1_U3.top_sub_9s_9ns_9_2_1_Adder_2_U.ce  ? \sub_9s_9ns_9_2_1_U3.top_sub_9s_9ns_9_2_1_Adder_2_U.a [8:4] : \sub_9s_9ns_9_2_1_U3.top_sub_9s_9ns_9_2_1_Adder_2_U.ain_s1 ;
assign _265_ = \sub_9s_9ns_9_2_1_U3.top_sub_9s_9ns_9_2_1_Adder_2_U.ce  ? \sub_9s_9ns_9_2_1_U3.top_sub_9s_9ns_9_2_1_Adder_2_U.facout_s1  : \sub_9s_9ns_9_2_1_U3.top_sub_9s_9ns_9_2_1_Adder_2_U.carry_s1 ;
assign _266_ = \sub_9s_9ns_9_2_1_U3.top_sub_9s_9ns_9_2_1_Adder_2_U.ce  ? \sub_9s_9ns_9_2_1_U3.top_sub_9s_9ns_9_2_1_Adder_2_U.fas_s1  : \sub_9s_9ns_9_2_1_U3.top_sub_9s_9ns_9_2_1_Adder_2_U.sum_s1 ;
assign _267_ = \sub_9s_9ns_9_2_1_U3.top_sub_9s_9ns_9_2_1_Adder_2_U.u1.a  + \sub_9s_9ns_9_2_1_U3.top_sub_9s_9ns_9_2_1_Adder_2_U.u1.b ;
assign { \sub_9s_9ns_9_2_1_U3.top_sub_9s_9ns_9_2_1_Adder_2_U.u1.cout , \sub_9s_9ns_9_2_1_U3.top_sub_9s_9ns_9_2_1_Adder_2_U.u1.s  } = _267_ + \sub_9s_9ns_9_2_1_U3.top_sub_9s_9ns_9_2_1_Adder_2_U.u1.cin ;
assign _268_ = \sub_9s_9ns_9_2_1_U3.top_sub_9s_9ns_9_2_1_Adder_2_U.u2.a  + \sub_9s_9ns_9_2_1_U3.top_sub_9s_9ns_9_2_1_Adder_2_U.u2.b ;
assign { \sub_9s_9ns_9_2_1_U3.top_sub_9s_9ns_9_2_1_Adder_2_U.u2.cout , \sub_9s_9ns_9_2_1_U3.top_sub_9s_9ns_9_2_1_Adder_2_U.u2.s  } = _268_ + \sub_9s_9ns_9_2_1_U3.top_sub_9s_9ns_9_2_1_Adder_2_U.u2.cin ;
assign _269_ = | p_Result_s_20_reg_1097;
assign _270_ = | trunc_ln851_reg_1173;
assign or_ln1195_fu_416_p2 = op_4[25:0] | { trunc_ln728_reg_1108, 25'h0000000 };
assign or_ln384_1_fu_539_p2 = underflow_1_fu_527_p2 | overflow_1_reg_1188;
assign or_ln384_fu_467_p2 = underflow_fu_462_p2 | overflow_reg_1134;
assign or_ln785_fu_370_p2 = p_Result_12_reg_1091 | icmp_ln785_reg_1124;
assign or_ln788_fu_522_p2 = xor_ln786_fu_517_p2 | icmp_ln790_reg_1194;
always @(posedge ap_clk)
op_3_V_reg_1058[5:0] <= 6'h00;
always @(posedge ap_clk)
select_ln1193_reg_1103[5:0] <= 6'h00;
always @(posedge ap_clk)
trunc_ln1497_reg_1496 <= _058_;
always @(posedge ap_clk)
trunc_ln1497_1_reg_1501 <= _057_;
always @(posedge ap_clk)
sub_ln1497_reg_1423 <= _055_;
always @(posedge ap_clk)
ret_V_26_reg_1484 <= _042_;
always @(posedge ap_clk)
ret_V_34_cast_reg_1489 <= _044_;
always @(posedge ap_clk)
ret_V_24_reg_1418 <= _040_;
always @(posedge ap_clk)
ret_V_23_reg_1259 <= _038_;
always @(posedge ap_clk)
ret_V_reg_1264 <= _049_;
always @(posedge ap_clk)
trunc_ln851_1_reg_1271 <= _061_;
always @(posedge ap_clk)
ret_V_25_reg_1276 <= _041_;
always @(posedge ap_clk)
ret_V_6_reg_1281 <= _045_;
always @(posedge ap_clk)
ret_V_13_reg_1303 <= _033_;
always @(posedge ap_clk)
r_reg_1511 <= _031_;
always @(posedge ap_clk)
ret_V_27_reg_1516 <= _043_;
always @(posedge ap_clk)
ret_V_21_reg_1079 <= _036_;
always @(posedge ap_clk)
p_Result_11_reg_1085 <= _025_;
always @(posedge ap_clk)
p_Result_12_reg_1091 <= _026_;
always @(posedge ap_clk)
p_Result_s_20_reg_1097 <= _029_;
always @(posedge ap_clk)
select_ln1193_reg_1103[8:6] <= _050_;
always @(posedge ap_clk)
overflow_reg_1134 <= _024_;
always @(posedge ap_clk)
ret_V_22_reg_1140 <= _037_;
always @(posedge ap_clk)
p_Result_13_reg_1145 <= _027_;
always @(posedge ap_clk)
p_Result_14_reg_1151 <= _028_;
always @(posedge ap_clk)
trunc_ln790_reg_1157 <= _060_;
always @(posedge ap_clk)
op_3_V_reg_1058[7:6] <= _018_;
always @(posedge ap_clk)
op_25_V_reg_1464 <= _017_;
always @(posedge ap_clk)
icmp_ln851_reg_1288 <= _015_;
always @(posedge ap_clk)
ret_V_7_reg_1298 <= _046_;
always @(posedge ap_clk)
ret_V_9_reg_1308 <= _048_;
always @(posedge ap_clk)
icmp_ln851_3_reg_1315 <= _014_;
always @(posedge ap_clk)
icmp_ln851_2_reg_1249 <= _013_;
always @(posedge ap_clk)
select_ln69_reg_1254 <= _052_;
always @(posedge ap_clk)
icmp_ln851_1_reg_1362 <= _012_;
always @(posedge ap_clk)
ret_V_15_reg_1367 <= _035_;
always @(posedge ap_clk)
tmp_13_reg_1373 <= _056_;
always @(posedge ap_clk)
icmp_ln850_reg_1209 <= _011_;
always @(posedge ap_clk)
op_8_V_reg_1214 <= _020_;
always @(posedge ap_clk)
select_ln384_3_reg_1219 <= _051_;
always @(posedge ap_clk)
trunc_ln851_3_reg_1224 <= _063_;
always @(posedge ap_clk)
or_ln1195_reg_1168 <= _021_;
always @(posedge ap_clk)
trunc_ln851_reg_1173 <= _064_;
always @(posedge ap_clk)
signbit_reg_1178 <= _054_;
always @(posedge ap_clk)
or_ln384_reg_1183 <= _022_;
always @(posedge ap_clk)
overflow_1_reg_1188 <= _023_;
always @(posedge ap_clk)
icmp_ln790_reg_1194 <= _010_;
always @(posedge ap_clk)
add_ln731_reg_1053 <= _007_;
always @(posedge ap_clk)
add_ln69_reg_1454 <= _006_;
always @(posedge ap_clk)
add_ln69_4_reg_1536 <= _004_;
always @(posedge ap_clk)
add_ln69_5_reg_1541 <= _005_;
always @(posedge ap_clk)
ret_V_10_reg_1398 <= _032_;
always @(posedge ap_clk)
op_21_V_reg_1408 <= _016_;
always @(posedge ap_clk)
add_ln69_2_reg_1413 <= _003_;
always @(posedge ap_clk)
ret_V_8_reg_1325 <= _047_;
always @(posedge ap_clk)
r_V_reg_1330 <= _030_;
always @(posedge ap_clk)
ret_V_24_cast_reg_1335 <= _039_;
always @(posedge ap_clk)
trunc_ln851_2_reg_1342 <= _062_;
always @(posedge ap_clk)
ret_V_14_reg_1347 <= _034_;
always @(posedge ap_clk)
select_ln850_7_reg_1352 <= _053_;
always @(posedge ap_clk)
add_ln69_1_reg_1357 <= _002_;
always @(posedge ap_clk)
add_ln691_reg_1506 <= _001_;
always @(posedge ap_clk)
trunc_ln728_reg_1108 <= _059_;
always @(posedge ap_clk)
op_6_V_reg_1113 <= _019_;
always @(posedge ap_clk)
Range1_all_ones_reg_1119 <= _000_;
always @(posedge ap_clk)
icmp_ln785_reg_1124 <= _009_;
always @(posedge ap_clk)
ap_CS_fsm <= _008_;
assign _065_ = _071_ ? 2'h2 : 2'h1;
assign _271_ = ap_CS_fsm == 1'h1;
function [27:0] _747_;
input [27:0] a;
input [783:0] b;
input [27:0] s;
case (s)
28'b0000000000000000000000000001:
_747_ = b[27:0];
28'b0000000000000000000000000010:
_747_ = b[55:28];
28'b0000000000000000000000000100:
_747_ = b[83:56];
28'b0000000000000000000000001000:
_747_ = b[111:84];
28'b0000000000000000000000010000:
_747_ = b[139:112];
28'b0000000000000000000000100000:
_747_ = b[167:140];
28'b0000000000000000000001000000:
_747_ = b[195:168];
28'b0000000000000000000010000000:
_747_ = b[223:196];
28'b0000000000000000000100000000:
_747_ = b[251:224];
28'b0000000000000000001000000000:
_747_ = b[279:252];
28'b0000000000000000010000000000:
_747_ = b[307:280];
28'b0000000000000000100000000000:
_747_ = b[335:308];
28'b0000000000000001000000000000:
_747_ = b[363:336];
28'b0000000000000010000000000000:
_747_ = b[391:364];
28'b0000000000000100000000000000:
_747_ = b[419:392];
28'b0000000000001000000000000000:
_747_ = b[447:420];
28'b0000000000010000000000000000:
_747_ = b[475:448];
28'b0000000000100000000000000000:
_747_ = b[503:476];
28'b0000000001000000000000000000:
_747_ = b[531:504];
28'b0000000010000000000000000000:
_747_ = b[559:532];
28'b0000000100000000000000000000:
_747_ = b[587:560];
28'b0000001000000000000000000000:
_747_ = b[615:588];
28'b0000010000000000000000000000:
_747_ = b[643:616];
28'b0000100000000000000000000000:
_747_ = b[671:644];
28'b0001000000000000000000000000:
_747_ = b[699:672];
28'b0010000000000000000000000000:
_747_ = b[727:700];
28'b0100000000000000000000000000:
_747_ = b[755:728];
28'b1000000000000000000000000000:
_747_ = b[783:756];
28'b0000000000000000000000000000:
_747_ = a;
default:
_747_ = 28'bx;
endcase
endfunction
assign ap_NS_fsm = _747_(28'hxxxxxxx, { 26'h0000000, _065_, 756'h000000400000080000010000002000000400000080000010000002000000400000080000010000002000000400000080000010000002000000400000080000010000002000000400000080000010000002000000400000080000000000001 }, { _271_, _298_, _297_, _296_, _295_, _294_, _293_, _292_, _291_, _290_, _289_, _288_, _287_, _286_, _285_, _284_, _283_, _282_, _281_, _280_, _279_, _278_, _277_, _276_, _275_, _274_, _273_, _272_ });
assign _272_ = ap_CS_fsm == 28'h8000000;
assign _273_ = ap_CS_fsm == 27'h4000000;
assign _274_ = ap_CS_fsm == 26'h2000000;
assign _275_ = ap_CS_fsm == 25'h1000000;
assign _276_ = ap_CS_fsm == 24'h800000;
assign _277_ = ap_CS_fsm == 23'h400000;
assign _278_ = ap_CS_fsm == 22'h200000;
assign _279_ = ap_CS_fsm == 21'h100000;
assign _280_ = ap_CS_fsm == 20'h80000;
assign _281_ = ap_CS_fsm == 19'h40000;
assign _282_ = ap_CS_fsm == 18'h20000;
assign _283_ = ap_CS_fsm == 17'h10000;
assign _284_ = ap_CS_fsm == 16'h8000;
assign _285_ = ap_CS_fsm == 15'h4000;
assign _286_ = ap_CS_fsm == 14'h2000;
assign _287_ = ap_CS_fsm == 13'h1000;
assign _288_ = ap_CS_fsm == 12'h800;
assign _289_ = ap_CS_fsm == 11'h400;
assign _290_ = ap_CS_fsm == 10'h200;
assign _291_ = ap_CS_fsm == 9'h100;
assign _292_ = ap_CS_fsm == 8'h80;
assign _293_ = ap_CS_fsm == 7'h40;
assign _294_ = ap_CS_fsm == 6'h20;
assign _295_ = ap_CS_fsm == 5'h10;
assign _296_ = ap_CS_fsm == 4'h8;
assign _297_ = ap_CS_fsm == 3'h4;
assign _298_ = ap_CS_fsm == 2'h2;
assign op_29_ap_vld = ap_CS_fsm[27] ? 1'h1 : 1'h0;
assign ap_idle = _070_ ? 1'h1 : 1'h0;
assign _058_ = _069_ ? grp_fu_917_p2[1:0] : trunc_ln1497_reg_1496;
assign _057_ = _068_ ? grp_fu_908_p2[1:0] : trunc_ln1497_1_reg_1501;
assign _055_ = _067_ ? grp_fu_854_p2 : sub_ln1497_reg_1423;
assign _044_ = ap_CS_fsm[20] ? grp_fu_946_p2[32:1] : ret_V_34_cast_reg_1489;
assign _042_ = ap_CS_fsm[20] ? grp_fu_946_p2 : ret_V_26_reg_1484;
assign _040_ = ap_CS_fsm[15] ? ret_V_24_fu_882_p3 : ret_V_24_reg_1418;
assign _045_ = ap_CS_fsm[9] ? grp_fu_629_p2[8:6] : ret_V_6_reg_1281;
assign _041_ = ap_CS_fsm[9] ? grp_fu_629_p2 : ret_V_25_reg_1276;
assign _061_ = ap_CS_fsm[9] ? grp_fu_609_p2[24:0] : trunc_ln851_1_reg_1271;
assign _049_ = ap_CS_fsm[9] ? grp_fu_609_p2[32:25] : ret_V_reg_1264;
assign _038_ = ap_CS_fsm[9] ? grp_fu_609_p2 : ret_V_23_reg_1259;
assign _033_ = _066_ ? grp_fu_682_p2 : ret_V_13_reg_1303;
assign _043_ = ap_CS_fsm[23] ? ret_V_27_fu_996_p3 : ret_V_27_reg_1516;
assign _031_ = ap_CS_fsm[23] ? r_fu_975_p3 : r_reg_1511;
assign _050_ = ap_CS_fsm[3] ? select_ln1193_fu_313_p3[8:6] : select_ln1193_reg_1103[8:6];
assign _029_ = ap_CS_fsm[3] ? grp_fu_281_p2[15:8] : p_Result_s_20_reg_1097;
assign _026_ = ap_CS_fsm[3] ? grp_fu_281_p2[7] : p_Result_12_reg_1091;
assign _025_ = ap_CS_fsm[3] ? grp_fu_281_p2[15] : p_Result_11_reg_1085;
assign _036_ = ap_CS_fsm[3] ? grp_fu_281_p2 : ret_V_21_reg_1079;
assign _060_ = ap_CS_fsm[5] ? grp_fu_365_p2[6:0] : trunc_ln790_reg_1157;
assign _028_ = ap_CS_fsm[5] ? grp_fu_365_p2[7] : p_Result_14_reg_1151;
assign _027_ = ap_CS_fsm[5] ? grp_fu_365_p2[8] : p_Result_13_reg_1145;
assign _037_ = ap_CS_fsm[5] ? grp_fu_365_p2 : ret_V_22_reg_1140;
assign _024_ = ap_CS_fsm[5] ? overflow_fu_379_p2 : overflow_reg_1134;
assign _018_ = ap_CS_fsm[2] ? add_ln731_reg_1053 : op_3_V_reg_1058[7:6];
assign _017_ = ap_CS_fsm[18] ? grp_fu_926_p2 : op_25_V_reg_1464;
assign _015_ = ap_CS_fsm[10] ? icmp_ln851_fu_672_p2 : icmp_ln851_reg_1288;
assign _014_ = ap_CS_fsm[11] ? icmp_ln851_3_fu_701_p2 : icmp_ln851_3_reg_1315;
assign _048_ = ap_CS_fsm[11] ? op_14[7:3] : ret_V_9_reg_1308;
assign _046_ = ap_CS_fsm[11] ? grp_fu_677_p2 : ret_V_7_reg_1298;
assign _052_ = ap_CS_fsm[8] ? select_ln69_fu_640_p3 : select_ln69_reg_1254;
assign _013_ = ap_CS_fsm[8] ? icmp_ln851_2_fu_635_p2 : icmp_ln851_2_reg_1249;
assign _056_ = ap_CS_fsm[13] ? ret_V_15_fu_803_p3[4] : tmp_13_reg_1373;
assign _035_ = ap_CS_fsm[13] ? ret_V_15_fu_803_p3 : ret_V_15_reg_1367;
assign _012_ = ap_CS_fsm[13] ? icmp_ln851_1_fu_781_p2 : icmp_ln851_1_reg_1362;
assign _063_ = ap_CS_fsm[7] ? op_8_V_fu_544_p3[5:0] : trunc_ln851_3_reg_1224;
assign _051_ = ap_CS_fsm[7] ? select_ln384_3_fu_559_p3 : select_ln384_3_reg_1219;
assign _020_ = ap_CS_fsm[7] ? op_8_V_fu_544_p3 : op_8_V_reg_1214;
assign _011_ = ap_CS_fsm[7] ? icmp_ln850_fu_500_p2 : icmp_ln850_reg_1209;
assign _010_ = ap_CS_fsm[6] ? icmp_ln790_fu_482_p2 : icmp_ln790_reg_1194;
assign _023_ = ap_CS_fsm[6] ? overflow_1_fu_477_p2 : overflow_1_reg_1188;
assign _022_ = ap_CS_fsm[6] ? or_ln384_fu_467_p2 : or_ln384_reg_1183;
assign _054_ = ap_CS_fsm[6] ? signbit_fu_433_p2 : signbit_reg_1178;
assign _064_ = ap_CS_fsm[6] ? or_ln1195_fu_416_p2[24:0] : trunc_ln851_reg_1173;
assign _021_ = ap_CS_fsm[6] ? or_ln1195_fu_416_p2 : or_ln1195_reg_1168;
assign _007_ = ap_CS_fsm[1] ? grp_fu_253_p2 : add_ln731_reg_1053;
assign _006_ = ap_CS_fsm[16] ? grp_fu_896_p2 : add_ln69_reg_1454;
assign _005_ = ap_CS_fsm[25] ? grp_fu_1023_p2 : add_ln69_5_reg_1541;
assign _004_ = ap_CS_fsm[25] ? grp_fu_1018_p2 : add_ln69_4_reg_1536;
assign _003_ = ap_CS_fsm[14] ? grp_fu_845_p2 : add_ln69_2_reg_1413;
assign _016_ = ap_CS_fsm[14] ? grp_fu_833_p2[28:25] : op_21_V_reg_1408;
assign _032_ = ap_CS_fsm[14] ? grp_fu_786_p2 : ret_V_10_reg_1398;
assign _002_ = ap_CS_fsm[12] ? grp_fu_717_p2 : add_ln69_1_reg_1357;
assign _053_ = ap_CS_fsm[12] ? select_ln850_7_fu_767_p3 : select_ln850_7_reg_1352;
assign _034_ = ap_CS_fsm[12] ? grp_fu_707_p2 : ret_V_14_reg_1347;
assign _062_ = ap_CS_fsm[12] ? grp_fu_494_p2[24:0] : trunc_ln851_2_reg_1342;
assign _039_ = ap_CS_fsm[12] ? grp_fu_494_p2[26:25] : ret_V_24_cast_reg_1335;
assign _030_ = ap_CS_fsm[12] ? grp_fu_494_p2 : r_V_reg_1330;
assign _047_ = ap_CS_fsm[12] ? ret_V_8_fu_734_p3 : ret_V_8_reg_1325;
assign _001_ = ap_CS_fsm[22] ? grp_fu_962_p2 : add_ln691_reg_1506;
assign _009_ = ap_CS_fsm[4] ? icmp_ln785_fu_357_p2 : icmp_ln785_reg_1124;
assign _000_ = ap_CS_fsm[4] ? Range1_all_ones_fu_352_p2 : Range1_all_ones_reg_1119;
assign _019_ = ap_CS_fsm[4] ? ret_V_20_fu_336_p2[9:6] : op_6_V_reg_1113;
assign _059_ = ap_CS_fsm[4] ? op_2[0] : trunc_ln728_reg_1108;
assign _008_ = ap_rst ? 28'h0000001 : ap_NS_fsm;
assign Range1_all_ones_fu_352_p2 = _075_ ? 1'h1 : 1'h0;
assign icmp_ln785_fu_357_p2 = _269_ ? 1'h1 : 1'h0;
assign icmp_ln790_fu_482_p2 = _076_ ? 1'h1 : 1'h0;
assign icmp_ln850_fu_500_p2 = _270_ ? 1'h1 : 1'h0;
assign icmp_ln851_1_fu_781_p2 = _077_ ? 1'h1 : 1'h0;
assign icmp_ln851_2_fu_635_p2 = _078_ ? 1'h1 : 1'h0;
assign icmp_ln851_3_fu_701_p2 = _079_ ? 1'h1 : 1'h0;
assign icmp_ln851_fu_672_p2 = _080_ ? 1'h1 : 1'h0;
assign op_8_V_fu_544_p3 = or_ln384_1_fu_539_p2 ? select_ln384_fu_532_p3 : ret_V_22_reg_1140[7:0];
assign r_fu_975_p3 = tmp_13_reg_1373 ? trunc_ln1497_reg_1496 : trunc_ln1497_1_reg_1501;
assign ret_V_15_fu_803_p3 = op_14[7] ? select_ln850_3_fu_798_p3 : ret_V_9_reg_1308;
assign ret_V_24_fu_882_p3 = r_V_reg_1330[35] ? select_ln850_2_fu_877_p3 : ret_V_24_cast_reg_1335;
assign ret_V_27_fu_996_p3 = ret_V_26_reg_1484[33] ? select_ln850_5_fu_990_p3 : ret_V_34_cast_reg_1489;
assign ret_V_8_fu_734_p3 = ret_V_23_reg_1259[32] ? select_ln850_fu_729_p3 : ret_V_reg_1264;
assign select_ln1193_fu_313_p3 = op_5 ? 9'h1c0 : 9'h000;
assign select_ln1498_fu_426_p3 = op_5 ? 32'd4261412864 : 32'd0;
assign select_ln384_2_fu_552_p3 = overflow_reg_1134 ? 2'h1 : 2'h3;
assign select_ln384_3_fu_559_p3 = or_ln384_reg_1183 ? select_ln384_2_fu_552_p3 : ret_V_21_reg_1079[7:6];
assign select_ln384_fu_532_p3 = overflow_1_reg_1188 ? 8'h7f : 8'h81;
assign select_ln69_fu_640_p3 = ret_V_19_fu_589_p2 ? 5'h1f : 5'h00;
assign select_ln850_2_fu_877_p3 = icmp_ln851_1_reg_1362 ? ret_V_24_cast_reg_1335 : ret_V_10_reg_1398;
assign select_ln850_3_fu_798_p3 = icmp_ln851_3_reg_1315 ? ret_V_9_reg_1308 : ret_V_14_reg_1347;
assign select_ln850_5_fu_990_p3 = op_16[0] ? add_ln691_reg_1506 : ret_V_34_cast_reg_1489;
assign select_ln850_6_fu_762_p3 = icmp_ln851_2_reg_1249 ? ret_V_6_reg_1281 : ret_V_13_reg_1303;
assign select_ln850_7_fu_767_p3 = ret_V_25_reg_1276[8] ? select_ln850_6_fu_762_p3 : ret_V_6_reg_1281;
assign select_ln850_fu_729_p3 = icmp_ln851_reg_1288 ? ret_V_reg_1264 : ret_V_7_reg_1298;
assign signbit_fu_433_p2 = _081_ ? 1'h1 : 1'h0;
assign ret_V_19_fu_589_p2 = or_ln1195_reg_1168[25] ^ and_ln353_fu_584_p2;
assign ret_V_20_fu_336_p2 = { op_3_V_reg_1058[7], op_3_V_reg_1058[7], op_3_V_reg_1058 } ^ { op_2, 6'h00 };
assign ap_CS_fsm_state1 = ap_CS_fsm[0];
assign ap_CS_fsm_state10 = ap_CS_fsm[9];
assign ap_CS_fsm_state11 = ap_CS_fsm[10];
assign ap_CS_fsm_state12 = ap_CS_fsm[11];
assign ap_CS_fsm_state13 = ap_CS_fsm[12];
assign ap_CS_fsm_state14 = ap_CS_fsm[13];
assign ap_CS_fsm_state15 = ap_CS_fsm[14];
assign ap_CS_fsm_state16 = ap_CS_fsm[15];
assign ap_CS_fsm_state17 = ap_CS_fsm[16];
assign ap_CS_fsm_state18 = ap_CS_fsm[17];
assign ap_CS_fsm_state19 = ap_CS_fsm[18];
assign ap_CS_fsm_state2 = ap_CS_fsm[1];
assign ap_CS_fsm_state20 = ap_CS_fsm[19];
assign ap_CS_fsm_state21 = ap_CS_fsm[20];
assign ap_CS_fsm_state22 = ap_CS_fsm[21];
assign ap_CS_fsm_state23 = ap_CS_fsm[22];
assign ap_CS_fsm_state24 = ap_CS_fsm[23];
assign ap_CS_fsm_state25 = ap_CS_fsm[24];
assign ap_CS_fsm_state26 = ap_CS_fsm[25];
assign ap_CS_fsm_state27 = ap_CS_fsm[26];
assign ap_CS_fsm_state28 = ap_CS_fsm[27];
assign ap_CS_fsm_state3 = ap_CS_fsm[2];
assign ap_CS_fsm_state4 = ap_CS_fsm[3];
assign ap_CS_fsm_state5 = ap_CS_fsm[4];
assign ap_CS_fsm_state6 = ap_CS_fsm[5];
assign ap_CS_fsm_state7 = ap_CS_fsm[6];
assign ap_CS_fsm_state8 = ap_CS_fsm[7];
assign ap_CS_fsm_state9 = ap_CS_fsm[8];
assign ap_done = op_29_ap_vld;
assign ap_ready = op_29_ap_vld;
assign conv_i188_fu_905_p1 = { ret_V_24_reg_1418[1], ret_V_24_reg_1418[1], ret_V_24_reg_1418[1], ret_V_24_reg_1418[1], ret_V_24_reg_1418[1], ret_V_24_reg_1418[1], ret_V_24_reg_1418[1], ret_V_24_reg_1418[1], ret_V_24_reg_1418[1], ret_V_24_reg_1418[1], ret_V_24_reg_1418[1], ret_V_24_reg_1418[1], ret_V_24_reg_1418[1], ret_V_24_reg_1418[1], ret_V_24_reg_1418[1], ret_V_24_reg_1418[1], ret_V_24_reg_1418[1], ret_V_24_reg_1418[1], ret_V_24_reg_1418[1], ret_V_24_reg_1418[1], ret_V_24_reg_1418[1], ret_V_24_reg_1418[1], ret_V_24_reg_1418[1], ret_V_24_reg_1418[1], ret_V_24_reg_1418[1], ret_V_24_reg_1418[1], ret_V_24_reg_1418[1], ret_V_24_reg_1418[1], ret_V_24_reg_1418[1], ret_V_24_reg_1418[1], ret_V_24_reg_1418 };
assign grp_fu_1018_p1 = { 16'h0000, r_reg_1511[1], r_reg_1511[1], r_reg_1511[1], r_reg_1511[1], r_reg_1511[1], r_reg_1511[1], r_reg_1511[1], r_reg_1511[1], r_reg_1511[1], r_reg_1511[1], r_reg_1511[1], r_reg_1511[1], r_reg_1511[1], r_reg_1511[1], r_reg_1511 };
assign grp_fu_1023_p0 = { op_18[3], op_18 };
assign grp_fu_1023_p1 = { op_17[1], op_17[1], op_17[1], op_17 };
assign grp_fu_1032_p0 = { add_ln69_5_reg_1541[4], add_ln69_5_reg_1541[4], add_ln69_5_reg_1541[4], add_ln69_5_reg_1541[4], add_ln69_5_reg_1541[4], add_ln69_5_reg_1541[4], add_ln69_5_reg_1541[4], add_ln69_5_reg_1541[4], add_ln69_5_reg_1541[4], add_ln69_5_reg_1541[4], add_ln69_5_reg_1541[4], add_ln69_5_reg_1541[4], add_ln69_5_reg_1541[4], add_ln69_5_reg_1541[4], add_ln69_5_reg_1541[4], add_ln69_5_reg_1541[4], add_ln69_5_reg_1541[4], add_ln69_5_reg_1541[4], add_ln69_5_reg_1541[4], add_ln69_5_reg_1541[4], add_ln69_5_reg_1541[4], add_ln69_5_reg_1541[4], add_ln69_5_reg_1541[4], add_ln69_5_reg_1541[4], add_ln69_5_reg_1541[4], add_ln69_5_reg_1541[4], add_ln69_5_reg_1541[4], add_ln69_5_reg_1541 };
assign grp_fu_253_p0 = op_1[1:0];
assign grp_fu_253_p1 = op_0[1:0];
assign grp_fu_281_p0 = { 2'h0, op_1, 6'h00 };
assign grp_fu_281_p1 = { add_ln731_reg_1053[1], add_ln731_reg_1053[1], add_ln731_reg_1053[1], add_ln731_reg_1053[1], add_ln731_reg_1053[1], add_ln731_reg_1053[1], add_ln731_reg_1053[1], add_ln731_reg_1053[1], add_ln731_reg_1053, 6'h00 };
assign grp_fu_365_p0 = { op_3_V_reg_1058[7], op_3_V_reg_1058 };
assign grp_fu_609_p0 = { op_4[31], op_4 };
assign grp_fu_609_p1 = { op_6_V_reg_1113[3], op_6_V_reg_1113[3], op_6_V_reg_1113[3], op_6_V_reg_1113[3], op_6_V_reg_1113, 25'h0000000 };
assign grp_fu_629_p0 = { select_ln384_3_reg_1219[1], select_ln384_3_reg_1219, 6'h00 };
assign grp_fu_629_p1 = { op_8_V_reg_1214[7], op_8_V_reg_1214 };
assign grp_fu_707_p0 = op_14[7:3];
assign grp_fu_717_p0 = { op_15[3], op_15 };
assign grp_fu_833_p0 = { select_ln850_7_reg_1352[2], select_ln850_7_reg_1352, 25'h0000000 };
assign grp_fu_833_p1 = { 3'h0, signbit_reg_1178, 25'h0000000 };
assign grp_fu_845_p0 = { add_ln69_1_reg_1357[4], add_ln69_1_reg_1357[4], add_ln69_1_reg_1357[4], add_ln69_1_reg_1357[4], add_ln69_1_reg_1357 };
assign grp_fu_845_p1 = { ret_V_8_reg_1325[7], ret_V_8_reg_1325 };
assign grp_fu_854_p1 = { ret_V_15_reg_1367[4], ret_V_15_reg_1367 };
assign grp_fu_896_p0 = { op_21_V_reg_1408[3], op_21_V_reg_1408[3], op_21_V_reg_1408[3], op_21_V_reg_1408[3], op_21_V_reg_1408[3], op_21_V_reg_1408[3], op_21_V_reg_1408[3], op_21_V_reg_1408[3], op_21_V_reg_1408[3], op_21_V_reg_1408[3], op_21_V_reg_1408[3], op_21_V_reg_1408[3], op_21_V_reg_1408[3], op_21_V_reg_1408 };
assign grp_fu_896_p1 = { op_13[15], op_13 };
assign grp_fu_908_p1 = { ret_V_15_reg_1367[4], ret_V_15_reg_1367[4], ret_V_15_reg_1367[4], ret_V_15_reg_1367[4], ret_V_15_reg_1367[4], ret_V_15_reg_1367[4], ret_V_15_reg_1367[4], ret_V_15_reg_1367[4], ret_V_15_reg_1367[4], ret_V_15_reg_1367[4], ret_V_15_reg_1367[4], ret_V_15_reg_1367[4], ret_V_15_reg_1367[4], ret_V_15_reg_1367[4], ret_V_15_reg_1367[4], ret_V_15_reg_1367[4], ret_V_15_reg_1367[4], ret_V_15_reg_1367[4], ret_V_15_reg_1367[4], ret_V_15_reg_1367[4], ret_V_15_reg_1367[4], ret_V_15_reg_1367[4], ret_V_15_reg_1367[4], ret_V_15_reg_1367[4], ret_V_15_reg_1367[4], ret_V_15_reg_1367[4], ret_V_15_reg_1367[4], ret_V_15_reg_1367 };
assign grp_fu_917_p1 = { sub_ln1497_reg_1423[5], sub_ln1497_reg_1423[5], sub_ln1497_reg_1423[5], sub_ln1497_reg_1423[5], sub_ln1497_reg_1423[5], sub_ln1497_reg_1423[5], sub_ln1497_reg_1423[5], sub_ln1497_reg_1423[5], sub_ln1497_reg_1423[5], sub_ln1497_reg_1423[5], sub_ln1497_reg_1423[5], sub_ln1497_reg_1423[5], sub_ln1497_reg_1423[5], sub_ln1497_reg_1423[5], sub_ln1497_reg_1423[5], sub_ln1497_reg_1423[5], sub_ln1497_reg_1423[5], sub_ln1497_reg_1423[5], sub_ln1497_reg_1423[5], sub_ln1497_reg_1423[5], sub_ln1497_reg_1423[5], sub_ln1497_reg_1423[5], sub_ln1497_reg_1423[5], sub_ln1497_reg_1423[5], sub_ln1497_reg_1423[5], sub_ln1497_reg_1423[5], sub_ln1497_reg_1423 };
assign grp_fu_926_p0 = { add_ln69_2_reg_1413[8], add_ln69_2_reg_1413[8], add_ln69_2_reg_1413[8], add_ln69_2_reg_1413[8], add_ln69_2_reg_1413[8], add_ln69_2_reg_1413[8], add_ln69_2_reg_1413[8], add_ln69_2_reg_1413[8], add_ln69_2_reg_1413 };
assign grp_fu_946_p0 = { op_25_V_reg_1464[16], op_25_V_reg_1464[16], op_25_V_reg_1464[16], op_25_V_reg_1464[16], op_25_V_reg_1464[16], op_25_V_reg_1464[16], op_25_V_reg_1464[16], op_25_V_reg_1464[16], op_25_V_reg_1464[16], op_25_V_reg_1464[16], op_25_V_reg_1464[16], op_25_V_reg_1464[16], op_25_V_reg_1464[16], op_25_V_reg_1464[16], op_25_V_reg_1464[16], op_25_V_reg_1464[16], op_25_V_reg_1464, 1'h0 };
assign grp_fu_946_p1 = { op_16[1], op_16[1], op_16[1], op_16[1], op_16[1], op_16[1], op_16[1], op_16[1], op_16[1], op_16[1], op_16[1], op_16[1], op_16[1], op_16[1], op_16[1], op_16[1], op_16[1], op_16[1], op_16[1], op_16[1], op_16[1], op_16[1], op_16[1], op_16[1], op_16[1], op_16[1], op_16[1], op_16[1], op_16[1], op_16[1], op_16[1], op_16[1], op_16 };
assign lhs_V_2_fu_615_p3 = { select_ln384_3_reg_1219, 6'h00 };
assign lhs_V_fu_266_p3 = { op_1, 6'h00 };
assign lhs_cast_fu_405_p3 = { trunc_ln728_reg_1108, 25'h0000000 };
assign lhs_fu_325_p3 = { op_2, 6'h00 };
assign op_29 = grp_fu_1032_p2;
assign op_3_V_fu_259_p3 = { add_ln731_reg_1053, 6'h00 };
assign op_9_V_fu_774_p3 = { signbit_reg_1178, 25'h0000000 };
assign p_Result_10_fu_980_p3 = ret_V_26_reg_1484[33];
assign p_Result_6_fu_722_p3 = ret_V_23_reg_1259[32];
assign p_Result_7_fu_870_p3 = r_V_reg_1330[35];
assign p_Result_8_fu_755_p3 = ret_V_25_reg_1276[8];
assign p_Result_9_fu_791_p3 = op_14[7];
assign p_Result_s_fu_577_p1 = op_4;
assign p_Result_s_fu_577_p3 = op_4[31];
assign p_Val2_2_fu_505_p4 = ret_V_21_reg_1079[7:6];
assign p_Val2_4_fu_514_p1 = ret_V_22_reg_1140[7:0];
assign rhs_1_fu_598_p3 = { op_6_V_reg_1113, 25'h0000000 };
assign rhs_3_fu_822_p3 = { select_ln850_7_reg_1352, 25'h0000000 };
assign select_ln1193_fu_313_p0 = op_5;
assign select_ln1498_fu_426_p0 = op_5;
assign sext_ln1196_fu_333_p1 = { op_3_V_reg_1058[7], op_3_V_reg_1058[7], op_3_V_reg_1058 };
assign sext_ln69_7_fu_1011_p1 = { r_reg_1511[1], r_reg_1511[1], r_reg_1511[1], r_reg_1511[1], r_reg_1511[1], r_reg_1511[1], r_reg_1511[1], r_reg_1511[1], r_reg_1511[1], r_reg_1511[1], r_reg_1511[1], r_reg_1511[1], r_reg_1511[1], r_reg_1511[1], r_reg_1511 };
assign sext_ln703_2_fu_595_p0 = op_4;
assign sext_ln703_4_fu_931_p0 = op_16;
assign signbit_fu_433_p1 = op_4;
assign tmp_1_fu_570_p3 = or_ln1195_reg_1168[25];
assign tmp_6_fu_439_p3 = ret_V_21_reg_1079[6];
assign tmp_fu_935_p3 = { op_25_V_reg_1464, 1'h0 };
assign trunc_ln1195_fu_412_p0 = op_4;
assign trunc_ln1195_fu_412_p1 = op_4[25:0];
assign trunc_ln1497_1_fu_971_p1 = grp_fu_908_p2[1:0];
assign trunc_ln1497_fu_967_p1 = grp_fu_917_p2[1:0];
assign trunc_ln728_fu_321_p1 = op_2[0];
assign trunc_ln790_fu_401_p1 = grp_fu_365_p2[6:0];
assign trunc_ln851_1_fu_658_p1 = grp_fu_609_p2[24:0];
assign trunc_ln851_2_fu_751_p1 = grp_fu_494_p2[24:0];
assign trunc_ln851_3_fu_566_p1 = op_8_V_fu_544_p3[5:0];
assign trunc_ln851_4_fu_697_p1 = op_14[2:0];
assign trunc_ln851_5_fu_987_p0 = op_16;
assign trunc_ln851_5_fu_987_p1 = op_16[0];
assign trunc_ln851_fu_422_p1 = or_ln1195_fu_416_p2[24:0];
assign \sub_9s_9ns_9_2_1_U3.top_sub_9s_9ns_9_2_1_Adder_2_U.ain_s0  = \sub_9s_9ns_9_2_1_U3.top_sub_9s_9ns_9_2_1_Adder_2_U.a ;
assign \sub_9s_9ns_9_2_1_U3.top_sub_9s_9ns_9_2_1_Adder_2_U.s  = { \sub_9s_9ns_9_2_1_U3.top_sub_9s_9ns_9_2_1_Adder_2_U.fas_s2 , \sub_9s_9ns_9_2_1_U3.top_sub_9s_9ns_9_2_1_Adder_2_U.sum_s1  };
assign \sub_9s_9ns_9_2_1_U3.top_sub_9s_9ns_9_2_1_Adder_2_U.u2.a  = \sub_9s_9ns_9_2_1_U3.top_sub_9s_9ns_9_2_1_Adder_2_U.ain_s1 ;
assign \sub_9s_9ns_9_2_1_U3.top_sub_9s_9ns_9_2_1_Adder_2_U.u2.b  = \sub_9s_9ns_9_2_1_U3.top_sub_9s_9ns_9_2_1_Adder_2_U.bin_s1 ;
assign \sub_9s_9ns_9_2_1_U3.top_sub_9s_9ns_9_2_1_Adder_2_U.u2.cin  = \sub_9s_9ns_9_2_1_U3.top_sub_9s_9ns_9_2_1_Adder_2_U.carry_s1 ;
assign \sub_9s_9ns_9_2_1_U3.top_sub_9s_9ns_9_2_1_Adder_2_U.facout_s2  = \sub_9s_9ns_9_2_1_U3.top_sub_9s_9ns_9_2_1_Adder_2_U.u2.cout ;
assign \sub_9s_9ns_9_2_1_U3.top_sub_9s_9ns_9_2_1_Adder_2_U.fas_s2  = \sub_9s_9ns_9_2_1_U3.top_sub_9s_9ns_9_2_1_Adder_2_U.u2.s ;
assign \sub_9s_9ns_9_2_1_U3.top_sub_9s_9ns_9_2_1_Adder_2_U.u1.a  = \sub_9s_9ns_9_2_1_U3.top_sub_9s_9ns_9_2_1_Adder_2_U.a [3:0];
assign \sub_9s_9ns_9_2_1_U3.top_sub_9s_9ns_9_2_1_Adder_2_U.u1.b  = \sub_9s_9ns_9_2_1_U3.top_sub_9s_9ns_9_2_1_Adder_2_U.bin_s0 [3:0];
assign \sub_9s_9ns_9_2_1_U3.top_sub_9s_9ns_9_2_1_Adder_2_U.u1.cin  = 1'h1;
assign \sub_9s_9ns_9_2_1_U3.top_sub_9s_9ns_9_2_1_Adder_2_U.facout_s1  = \sub_9s_9ns_9_2_1_U3.top_sub_9s_9ns_9_2_1_Adder_2_U.u1.cout ;
assign \sub_9s_9ns_9_2_1_U3.top_sub_9s_9ns_9_2_1_Adder_2_U.fas_s1  = \sub_9s_9ns_9_2_1_U3.top_sub_9s_9ns_9_2_1_Adder_2_U.u1.s ;
assign \sub_9s_9ns_9_2_1_U3.top_sub_9s_9ns_9_2_1_Adder_2_U.a  = \sub_9s_9ns_9_2_1_U3.din0 ;
assign \sub_9s_9ns_9_2_1_U3.top_sub_9s_9ns_9_2_1_Adder_2_U.b  = \sub_9s_9ns_9_2_1_U3.din1 ;
assign \sub_9s_9ns_9_2_1_U3.top_sub_9s_9ns_9_2_1_Adder_2_U.ce  = \sub_9s_9ns_9_2_1_U3.ce ;
assign \sub_9s_9ns_9_2_1_U3.top_sub_9s_9ns_9_2_1_Adder_2_U.clk  = \sub_9s_9ns_9_2_1_U3.clk ;
assign \sub_9s_9ns_9_2_1_U3.top_sub_9s_9ns_9_2_1_Adder_2_U.reset  = \sub_9s_9ns_9_2_1_U3.reset ;
assign \sub_9s_9ns_9_2_1_U3.dout  = \sub_9s_9ns_9_2_1_U3.top_sub_9s_9ns_9_2_1_Adder_2_U.s ;
assign \sub_9s_9ns_9_2_1_U3.ce  = 1'h1;
assign \sub_9s_9ns_9_2_1_U3.clk  = ap_clk;
assign \sub_9s_9ns_9_2_1_U3.din0  = { op_3_V_reg_1058[7], op_3_V_reg_1058 };
assign \sub_9s_9ns_9_2_1_U3.din1  = select_ln1193_reg_1103;
assign grp_fu_365_p2 = \sub_9s_9ns_9_2_1_U3.dout ;
assign \sub_9s_9ns_9_2_1_U3.reset  = ap_rst;
assign \sub_6ns_6s_6_2_1_U14.top_sub_6ns_6s_6_2_1_Adder_10_U.ain_s0  = \sub_6ns_6s_6_2_1_U14.top_sub_6ns_6s_6_2_1_Adder_10_U.a ;
assign \sub_6ns_6s_6_2_1_U14.top_sub_6ns_6s_6_2_1_Adder_10_U.s  = { \sub_6ns_6s_6_2_1_U14.top_sub_6ns_6s_6_2_1_Adder_10_U.fas_s2 , \sub_6ns_6s_6_2_1_U14.top_sub_6ns_6s_6_2_1_Adder_10_U.sum_s1  };
assign \sub_6ns_6s_6_2_1_U14.top_sub_6ns_6s_6_2_1_Adder_10_U.u2.a  = \sub_6ns_6s_6_2_1_U14.top_sub_6ns_6s_6_2_1_Adder_10_U.ain_s1 ;
assign \sub_6ns_6s_6_2_1_U14.top_sub_6ns_6s_6_2_1_Adder_10_U.u2.b  = \sub_6ns_6s_6_2_1_U14.top_sub_6ns_6s_6_2_1_Adder_10_U.bin_s1 ;
assign \sub_6ns_6s_6_2_1_U14.top_sub_6ns_6s_6_2_1_Adder_10_U.u2.cin  = \sub_6ns_6s_6_2_1_U14.top_sub_6ns_6s_6_2_1_Adder_10_U.carry_s1 ;
assign \sub_6ns_6s_6_2_1_U14.top_sub_6ns_6s_6_2_1_Adder_10_U.facout_s2  = \sub_6ns_6s_6_2_1_U14.top_sub_6ns_6s_6_2_1_Adder_10_U.u2.cout ;
assign \sub_6ns_6s_6_2_1_U14.top_sub_6ns_6s_6_2_1_Adder_10_U.fas_s2  = \sub_6ns_6s_6_2_1_U14.top_sub_6ns_6s_6_2_1_Adder_10_U.u2.s ;
assign \sub_6ns_6s_6_2_1_U14.top_sub_6ns_6s_6_2_1_Adder_10_U.u1.a  = \sub_6ns_6s_6_2_1_U14.top_sub_6ns_6s_6_2_1_Adder_10_U.a [2:0];
assign \sub_6ns_6s_6_2_1_U14.top_sub_6ns_6s_6_2_1_Adder_10_U.u1.b  = \sub_6ns_6s_6_2_1_U14.top_sub_6ns_6s_6_2_1_Adder_10_U.bin_s0 [2:0];
assign \sub_6ns_6s_6_2_1_U14.top_sub_6ns_6s_6_2_1_Adder_10_U.u1.cin  = 1'h1;
assign \sub_6ns_6s_6_2_1_U14.top_sub_6ns_6s_6_2_1_Adder_10_U.facout_s1  = \sub_6ns_6s_6_2_1_U14.top_sub_6ns_6s_6_2_1_Adder_10_U.u1.cout ;
assign \sub_6ns_6s_6_2_1_U14.top_sub_6ns_6s_6_2_1_Adder_10_U.fas_s1  = \sub_6ns_6s_6_2_1_U14.top_sub_6ns_6s_6_2_1_Adder_10_U.u1.s ;
assign \sub_6ns_6s_6_2_1_U14.top_sub_6ns_6s_6_2_1_Adder_10_U.a  = \sub_6ns_6s_6_2_1_U14.din0 ;
assign \sub_6ns_6s_6_2_1_U14.top_sub_6ns_6s_6_2_1_Adder_10_U.b  = \sub_6ns_6s_6_2_1_U14.din1 ;
assign \sub_6ns_6s_6_2_1_U14.top_sub_6ns_6s_6_2_1_Adder_10_U.ce  = \sub_6ns_6s_6_2_1_U14.ce ;
assign \sub_6ns_6s_6_2_1_U14.top_sub_6ns_6s_6_2_1_Adder_10_U.clk  = \sub_6ns_6s_6_2_1_U14.clk ;
assign \sub_6ns_6s_6_2_1_U14.top_sub_6ns_6s_6_2_1_Adder_10_U.reset  = \sub_6ns_6s_6_2_1_U14.reset ;
assign \sub_6ns_6s_6_2_1_U14.dout  = \sub_6ns_6s_6_2_1_U14.top_sub_6ns_6s_6_2_1_Adder_10_U.s ;
assign \sub_6ns_6s_6_2_1_U14.ce  = 1'h1;
assign \sub_6ns_6s_6_2_1_U14.clk  = ap_clk;
assign \sub_6ns_6s_6_2_1_U14.din0  = 6'h00;
assign \sub_6ns_6s_6_2_1_U14.din1  = { ret_V_15_reg_1367[4], ret_V_15_reg_1367 };
assign grp_fu_854_p2 = \sub_6ns_6s_6_2_1_U14.dout ;
assign \sub_6ns_6s_6_2_1_U14.reset  = ap_rst;
assign \sub_33s_33s_33_2_1_U5.top_sub_33s_33s_33_2_1_Adder_3_U.ain_s0  = \sub_33s_33s_33_2_1_U5.top_sub_33s_33s_33_2_1_Adder_3_U.a ;
assign \sub_33s_33s_33_2_1_U5.top_sub_33s_33s_33_2_1_Adder_3_U.s  = { \sub_33s_33s_33_2_1_U5.top_sub_33s_33s_33_2_1_Adder_3_U.fas_s2 , \sub_33s_33s_33_2_1_U5.top_sub_33s_33s_33_2_1_Adder_3_U.sum_s1  };
assign \sub_33s_33s_33_2_1_U5.top_sub_33s_33s_33_2_1_Adder_3_U.u2.a  = \sub_33s_33s_33_2_1_U5.top_sub_33s_33s_33_2_1_Adder_3_U.ain_s1 ;
assign \sub_33s_33s_33_2_1_U5.top_sub_33s_33s_33_2_1_Adder_3_U.u2.b  = \sub_33s_33s_33_2_1_U5.top_sub_33s_33s_33_2_1_Adder_3_U.bin_s1 ;
assign \sub_33s_33s_33_2_1_U5.top_sub_33s_33s_33_2_1_Adder_3_U.u2.cin  = \sub_33s_33s_33_2_1_U5.top_sub_33s_33s_33_2_1_Adder_3_U.carry_s1 ;
assign \sub_33s_33s_33_2_1_U5.top_sub_33s_33s_33_2_1_Adder_3_U.facout_s2  = \sub_33s_33s_33_2_1_U5.top_sub_33s_33s_33_2_1_Adder_3_U.u2.cout ;
assign \sub_33s_33s_33_2_1_U5.top_sub_33s_33s_33_2_1_Adder_3_U.fas_s2  = \sub_33s_33s_33_2_1_U5.top_sub_33s_33s_33_2_1_Adder_3_U.u2.s ;
assign \sub_33s_33s_33_2_1_U5.top_sub_33s_33s_33_2_1_Adder_3_U.u1.a  = \sub_33s_33s_33_2_1_U5.top_sub_33s_33s_33_2_1_Adder_3_U.a [15:0];
assign \sub_33s_33s_33_2_1_U5.top_sub_33s_33s_33_2_1_Adder_3_U.u1.b  = \sub_33s_33s_33_2_1_U5.top_sub_33s_33s_33_2_1_Adder_3_U.bin_s0 [15:0];
assign \sub_33s_33s_33_2_1_U5.top_sub_33s_33s_33_2_1_Adder_3_U.u1.cin  = 1'h1;
assign \sub_33s_33s_33_2_1_U5.top_sub_33s_33s_33_2_1_Adder_3_U.facout_s1  = \sub_33s_33s_33_2_1_U5.top_sub_33s_33s_33_2_1_Adder_3_U.u1.cout ;
assign \sub_33s_33s_33_2_1_U5.top_sub_33s_33s_33_2_1_Adder_3_U.fas_s1  = \sub_33s_33s_33_2_1_U5.top_sub_33s_33s_33_2_1_Adder_3_U.u1.s ;
assign \sub_33s_33s_33_2_1_U5.top_sub_33s_33s_33_2_1_Adder_3_U.a  = \sub_33s_33s_33_2_1_U5.din0 ;
assign \sub_33s_33s_33_2_1_U5.top_sub_33s_33s_33_2_1_Adder_3_U.b  = \sub_33s_33s_33_2_1_U5.din1 ;
assign \sub_33s_33s_33_2_1_U5.top_sub_33s_33s_33_2_1_Adder_3_U.ce  = \sub_33s_33s_33_2_1_U5.ce ;
assign \sub_33s_33s_33_2_1_U5.top_sub_33s_33s_33_2_1_Adder_3_U.clk  = \sub_33s_33s_33_2_1_U5.clk ;
assign \sub_33s_33s_33_2_1_U5.top_sub_33s_33s_33_2_1_Adder_3_U.reset  = \sub_33s_33s_33_2_1_U5.reset ;
assign \sub_33s_33s_33_2_1_U5.dout  = \sub_33s_33s_33_2_1_U5.top_sub_33s_33s_33_2_1_Adder_3_U.s ;
assign \sub_33s_33s_33_2_1_U5.ce  = 1'h1;
assign \sub_33s_33s_33_2_1_U5.clk  = ap_clk;
assign \sub_33s_33s_33_2_1_U5.din0  = { op_4[31], op_4 };
assign \sub_33s_33s_33_2_1_U5.din1  = { op_6_V_reg_1113[3], op_6_V_reg_1113[3], op_6_V_reg_1113[3], op_6_V_reg_1113[3], op_6_V_reg_1113, 25'h0000000 };
assign grp_fu_609_p2 = \sub_33s_33s_33_2_1_U5.dout ;
assign \sub_33s_33s_33_2_1_U5.reset  = ap_rst;
assign \sub_16ns_16s_16_2_1_U2.top_sub_16ns_16s_16_2_1_Adder_1_U.ain_s0  = \sub_16ns_16s_16_2_1_U2.top_sub_16ns_16s_16_2_1_Adder_1_U.a ;
assign \sub_16ns_16s_16_2_1_U2.top_sub_16ns_16s_16_2_1_Adder_1_U.s  = { \sub_16ns_16s_16_2_1_U2.top_sub_16ns_16s_16_2_1_Adder_1_U.fas_s2 , \sub_16ns_16s_16_2_1_U2.top_sub_16ns_16s_16_2_1_Adder_1_U.sum_s1  };
assign \sub_16ns_16s_16_2_1_U2.top_sub_16ns_16s_16_2_1_Adder_1_U.u2.a  = \sub_16ns_16s_16_2_1_U2.top_sub_16ns_16s_16_2_1_Adder_1_U.ain_s1 ;
assign \sub_16ns_16s_16_2_1_U2.top_sub_16ns_16s_16_2_1_Adder_1_U.u2.b  = \sub_16ns_16s_16_2_1_U2.top_sub_16ns_16s_16_2_1_Adder_1_U.bin_s1 ;
assign \sub_16ns_16s_16_2_1_U2.top_sub_16ns_16s_16_2_1_Adder_1_U.u2.cin  = \sub_16ns_16s_16_2_1_U2.top_sub_16ns_16s_16_2_1_Adder_1_U.carry_s1 ;
assign \sub_16ns_16s_16_2_1_U2.top_sub_16ns_16s_16_2_1_Adder_1_U.facout_s2  = \sub_16ns_16s_16_2_1_U2.top_sub_16ns_16s_16_2_1_Adder_1_U.u2.cout ;
assign \sub_16ns_16s_16_2_1_U2.top_sub_16ns_16s_16_2_1_Adder_1_U.fas_s2  = \sub_16ns_16s_16_2_1_U2.top_sub_16ns_16s_16_2_1_Adder_1_U.u2.s ;
assign \sub_16ns_16s_16_2_1_U2.top_sub_16ns_16s_16_2_1_Adder_1_U.u1.a  = \sub_16ns_16s_16_2_1_U2.top_sub_16ns_16s_16_2_1_Adder_1_U.a [7:0];
assign \sub_16ns_16s_16_2_1_U2.top_sub_16ns_16s_16_2_1_Adder_1_U.u1.b  = \sub_16ns_16s_16_2_1_U2.top_sub_16ns_16s_16_2_1_Adder_1_U.bin_s0 [7:0];
assign \sub_16ns_16s_16_2_1_U2.top_sub_16ns_16s_16_2_1_Adder_1_U.u1.cin  = 1'h1;
assign \sub_16ns_16s_16_2_1_U2.top_sub_16ns_16s_16_2_1_Adder_1_U.facout_s1  = \sub_16ns_16s_16_2_1_U2.top_sub_16ns_16s_16_2_1_Adder_1_U.u1.cout ;
assign \sub_16ns_16s_16_2_1_U2.top_sub_16ns_16s_16_2_1_Adder_1_U.fas_s1  = \sub_16ns_16s_16_2_1_U2.top_sub_16ns_16s_16_2_1_Adder_1_U.u1.s ;
assign \sub_16ns_16s_16_2_1_U2.top_sub_16ns_16s_16_2_1_Adder_1_U.a  = \sub_16ns_16s_16_2_1_U2.din0 ;
assign \sub_16ns_16s_16_2_1_U2.top_sub_16ns_16s_16_2_1_Adder_1_U.b  = \sub_16ns_16s_16_2_1_U2.din1 ;
assign \sub_16ns_16s_16_2_1_U2.top_sub_16ns_16s_16_2_1_Adder_1_U.ce  = \sub_16ns_16s_16_2_1_U2.ce ;
assign \sub_16ns_16s_16_2_1_U2.top_sub_16ns_16s_16_2_1_Adder_1_U.clk  = \sub_16ns_16s_16_2_1_U2.clk ;
assign \sub_16ns_16s_16_2_1_U2.top_sub_16ns_16s_16_2_1_Adder_1_U.reset  = \sub_16ns_16s_16_2_1_U2.reset ;
assign \sub_16ns_16s_16_2_1_U2.dout  = \sub_16ns_16s_16_2_1_U2.top_sub_16ns_16s_16_2_1_Adder_1_U.s ;
assign \sub_16ns_16s_16_2_1_U2.ce  = 1'h1;
assign \sub_16ns_16s_16_2_1_U2.clk  = ap_clk;
assign \sub_16ns_16s_16_2_1_U2.din0  = { 2'h0, op_1, 6'h00 };
assign \sub_16ns_16s_16_2_1_U2.din1  = { add_ln731_reg_1053[1], add_ln731_reg_1053[1], add_ln731_reg_1053[1], add_ln731_reg_1053[1], add_ln731_reg_1053[1], add_ln731_reg_1053[1], add_ln731_reg_1053[1], add_ln731_reg_1053[1], add_ln731_reg_1053, 6'h00 };
assign grp_fu_281_p2 = \sub_16ns_16s_16_2_1_U2.dout ;
assign \sub_16ns_16s_16_2_1_U2.reset  = ap_rst;
assign \shl_32s_32s_32_7_1_U17.din1_cast  = \shl_32s_32s_32_7_1_U17.din1 ;
assign \shl_32s_32s_32_7_1_U17.din1_mask  = 32'd31;
assign \shl_32s_32s_32_7_1_U17.ce  = 1'h1;
assign \shl_32s_32s_32_7_1_U17.clk  = ap_clk;
assign \shl_32s_32s_32_7_1_U17.din0  = { ret_V_24_reg_1418[1], ret_V_24_reg_1418[1], ret_V_24_reg_1418[1], ret_V_24_reg_1418[1], ret_V_24_reg_1418[1], ret_V_24_reg_1418[1], ret_V_24_reg_1418[1], ret_V_24_reg_1418[1], ret_V_24_reg_1418[1], ret_V_24_reg_1418[1], ret_V_24_reg_1418[1], ret_V_24_reg_1418[1], ret_V_24_reg_1418[1], ret_V_24_reg_1418[1], ret_V_24_reg_1418[1], ret_V_24_reg_1418[1], ret_V_24_reg_1418[1], ret_V_24_reg_1418[1], ret_V_24_reg_1418[1], ret_V_24_reg_1418[1], ret_V_24_reg_1418[1], ret_V_24_reg_1418[1], ret_V_24_reg_1418[1], ret_V_24_reg_1418[1], ret_V_24_reg_1418[1], ret_V_24_reg_1418[1], ret_V_24_reg_1418[1], ret_V_24_reg_1418[1], ret_V_24_reg_1418[1], ret_V_24_reg_1418[1], ret_V_24_reg_1418 };
assign \shl_32s_32s_32_7_1_U17.din1  = { sub_ln1497_reg_1423[5], sub_ln1497_reg_1423[5], sub_ln1497_reg_1423[5], sub_ln1497_reg_1423[5], sub_ln1497_reg_1423[5], sub_ln1497_reg_1423[5], sub_ln1497_reg_1423[5], sub_ln1497_reg_1423[5], sub_ln1497_reg_1423[5], sub_ln1497_reg_1423[5], sub_ln1497_reg_1423[5], sub_ln1497_reg_1423[5], sub_ln1497_reg_1423[5], sub_ln1497_reg_1423[5], sub_ln1497_reg_1423[5], sub_ln1497_reg_1423[5], sub_ln1497_reg_1423[5], sub_ln1497_reg_1423[5], sub_ln1497_reg_1423[5], sub_ln1497_reg_1423[5], sub_ln1497_reg_1423[5], sub_ln1497_reg_1423[5], sub_ln1497_reg_1423[5], sub_ln1497_reg_1423[5], sub_ln1497_reg_1423[5], sub_ln1497_reg_1423[5], sub_ln1497_reg_1423 };
assign grp_fu_917_p2 = \shl_32s_32s_32_7_1_U17.dout ;
assign \shl_32s_32s_32_7_1_U17.reset  = ap_rst;
assign \mul_32s_4s_36_7_1_U4.top_mul_32s_4s_36_7_1_Mul_DSP_0_U.p  = \mul_32s_4s_36_7_1_U4.top_mul_32s_4s_36_7_1_Mul_DSP_0_U.buff4 ;
assign \mul_32s_4s_36_7_1_U4.top_mul_32s_4s_36_7_1_Mul_DSP_0_U.a  = \mul_32s_4s_36_7_1_U4.din0 ;
assign \mul_32s_4s_36_7_1_U4.top_mul_32s_4s_36_7_1_Mul_DSP_0_U.b  = \mul_32s_4s_36_7_1_U4.din1 ;
assign \mul_32s_4s_36_7_1_U4.top_mul_32s_4s_36_7_1_Mul_DSP_0_U.ce  = \mul_32s_4s_36_7_1_U4.ce ;
assign \mul_32s_4s_36_7_1_U4.top_mul_32s_4s_36_7_1_Mul_DSP_0_U.clk  = \mul_32s_4s_36_7_1_U4.clk ;
assign \mul_32s_4s_36_7_1_U4.dout  = \mul_32s_4s_36_7_1_U4.top_mul_32s_4s_36_7_1_Mul_DSP_0_U.p ;
assign \mul_32s_4s_36_7_1_U4.ce  = 1'h1;
assign \mul_32s_4s_36_7_1_U4.clk  = ap_clk;
assign \mul_32s_4s_36_7_1_U4.din0  = op_4;
assign \mul_32s_4s_36_7_1_U4.din1  = op_6_V_reg_1113;
assign grp_fu_494_p2 = \mul_32s_4s_36_7_1_U4.dout ;
assign \mul_32s_4s_36_7_1_U4.reset  = ap_rst;
assign \ashr_32s_32s_32_7_1_U16.din1_cast  = \ashr_32s_32s_32_7_1_U16.din1 ;
assign \ashr_32s_32s_32_7_1_U16.din1_mask  = 32'd31;
assign \ashr_32s_32s_32_7_1_U16.ce  = 1'h1;
assign \ashr_32s_32s_32_7_1_U16.clk  = ap_clk;
assign \ashr_32s_32s_32_7_1_U16.din0  = { ret_V_24_reg_1418[1], ret_V_24_reg_1418[1], ret_V_24_reg_1418[1], ret_V_24_reg_1418[1], ret_V_24_reg_1418[1], ret_V_24_reg_1418[1], ret_V_24_reg_1418[1], ret_V_24_reg_1418[1], ret_V_24_reg_1418[1], ret_V_24_reg_1418[1], ret_V_24_reg_1418[1], ret_V_24_reg_1418[1], ret_V_24_reg_1418[1], ret_V_24_reg_1418[1], ret_V_24_reg_1418[1], ret_V_24_reg_1418[1], ret_V_24_reg_1418[1], ret_V_24_reg_1418[1], ret_V_24_reg_1418[1], ret_V_24_reg_1418[1], ret_V_24_reg_1418[1], ret_V_24_reg_1418[1], ret_V_24_reg_1418[1], ret_V_24_reg_1418[1], ret_V_24_reg_1418[1], ret_V_24_reg_1418[1], ret_V_24_reg_1418[1], ret_V_24_reg_1418[1], ret_V_24_reg_1418[1], ret_V_24_reg_1418[1], ret_V_24_reg_1418 };
assign \ashr_32s_32s_32_7_1_U16.din1  = { ret_V_15_reg_1367[4], ret_V_15_reg_1367[4], ret_V_15_reg_1367[4], ret_V_15_reg_1367[4], ret_V_15_reg_1367[4], ret_V_15_reg_1367[4], ret_V_15_reg_1367[4], ret_V_15_reg_1367[4], ret_V_15_reg_1367[4], ret_V_15_reg_1367[4], ret_V_15_reg_1367[4], ret_V_15_reg_1367[4], ret_V_15_reg_1367[4], ret_V_15_reg_1367[4], ret_V_15_reg_1367[4], ret_V_15_reg_1367[4], ret_V_15_reg_1367[4], ret_V_15_reg_1367[4], ret_V_15_reg_1367[4], ret_V_15_reg_1367[4], ret_V_15_reg_1367[4], ret_V_15_reg_1367[4], ret_V_15_reg_1367[4], ret_V_15_reg_1367[4], ret_V_15_reg_1367[4], ret_V_15_reg_1367[4], ret_V_15_reg_1367[4], ret_V_15_reg_1367 };
assign grp_fu_908_p2 = \ashr_32s_32s_32_7_1_U16.dout ;
assign \ashr_32s_32s_32_7_1_U16.reset  = ap_rst;
assign \add_9s_9s_9_2_1_U6.top_add_9s_9s_9_2_1_Adder_4_U.ain_s0  = \add_9s_9s_9_2_1_U6.top_add_9s_9s_9_2_1_Adder_4_U.a ;
assign \add_9s_9s_9_2_1_U6.top_add_9s_9s_9_2_1_Adder_4_U.bin_s0  = \add_9s_9s_9_2_1_U6.top_add_9s_9s_9_2_1_Adder_4_U.b ;
assign \add_9s_9s_9_2_1_U6.top_add_9s_9s_9_2_1_Adder_4_U.s  = { \add_9s_9s_9_2_1_U6.top_add_9s_9s_9_2_1_Adder_4_U.fas_s2 , \add_9s_9s_9_2_1_U6.top_add_9s_9s_9_2_1_Adder_4_U.sum_s1  };
assign \add_9s_9s_9_2_1_U6.top_add_9s_9s_9_2_1_Adder_4_U.u2.a  = \add_9s_9s_9_2_1_U6.top_add_9s_9s_9_2_1_Adder_4_U.ain_s1 ;
assign \add_9s_9s_9_2_1_U6.top_add_9s_9s_9_2_1_Adder_4_U.u2.b  = \add_9s_9s_9_2_1_U6.top_add_9s_9s_9_2_1_Adder_4_U.bin_s1 ;
assign \add_9s_9s_9_2_1_U6.top_add_9s_9s_9_2_1_Adder_4_U.u2.cin  = \add_9s_9s_9_2_1_U6.top_add_9s_9s_9_2_1_Adder_4_U.carry_s1 ;
assign \add_9s_9s_9_2_1_U6.top_add_9s_9s_9_2_1_Adder_4_U.facout_s2  = \add_9s_9s_9_2_1_U6.top_add_9s_9s_9_2_1_Adder_4_U.u2.cout ;
assign \add_9s_9s_9_2_1_U6.top_add_9s_9s_9_2_1_Adder_4_U.fas_s2  = \add_9s_9s_9_2_1_U6.top_add_9s_9s_9_2_1_Adder_4_U.u2.s ;
assign \add_9s_9s_9_2_1_U6.top_add_9s_9s_9_2_1_Adder_4_U.u1.a  = \add_9s_9s_9_2_1_U6.top_add_9s_9s_9_2_1_Adder_4_U.a [3:0];
assign \add_9s_9s_9_2_1_U6.top_add_9s_9s_9_2_1_Adder_4_U.u1.b  = \add_9s_9s_9_2_1_U6.top_add_9s_9s_9_2_1_Adder_4_U.b [3:0];
assign \add_9s_9s_9_2_1_U6.top_add_9s_9s_9_2_1_Adder_4_U.u1.cin  = 1'h0;
assign \add_9s_9s_9_2_1_U6.top_add_9s_9s_9_2_1_Adder_4_U.facout_s1  = \add_9s_9s_9_2_1_U6.top_add_9s_9s_9_2_1_Adder_4_U.u1.cout ;
assign \add_9s_9s_9_2_1_U6.top_add_9s_9s_9_2_1_Adder_4_U.fas_s1  = \add_9s_9s_9_2_1_U6.top_add_9s_9s_9_2_1_Adder_4_U.u1.s ;
assign \add_9s_9s_9_2_1_U6.top_add_9s_9s_9_2_1_Adder_4_U.a  = \add_9s_9s_9_2_1_U6.din0 ;
assign \add_9s_9s_9_2_1_U6.top_add_9s_9s_9_2_1_Adder_4_U.b  = \add_9s_9s_9_2_1_U6.din1 ;
assign \add_9s_9s_9_2_1_U6.top_add_9s_9s_9_2_1_Adder_4_U.ce  = \add_9s_9s_9_2_1_U6.ce ;
assign \add_9s_9s_9_2_1_U6.top_add_9s_9s_9_2_1_Adder_4_U.clk  = \add_9s_9s_9_2_1_U6.clk ;
assign \add_9s_9s_9_2_1_U6.top_add_9s_9s_9_2_1_Adder_4_U.reset  = \add_9s_9s_9_2_1_U6.reset ;
assign \add_9s_9s_9_2_1_U6.dout  = \add_9s_9s_9_2_1_U6.top_add_9s_9s_9_2_1_Adder_4_U.s ;
assign \add_9s_9s_9_2_1_U6.ce  = 1'h1;
assign \add_9s_9s_9_2_1_U6.clk  = ap_clk;
assign \add_9s_9s_9_2_1_U6.din0  = { select_ln384_3_reg_1219[1], select_ln384_3_reg_1219, 6'h00 };
assign \add_9s_9s_9_2_1_U6.din1  = { op_8_V_reg_1214[7], op_8_V_reg_1214 };
assign grp_fu_629_p2 = \add_9s_9s_9_2_1_U6.dout ;
assign \add_9s_9s_9_2_1_U6.reset  = ap_rst;
assign \add_9s_9s_9_2_1_U13.top_add_9s_9s_9_2_1_Adder_4_U.ain_s0  = \add_9s_9s_9_2_1_U13.top_add_9s_9s_9_2_1_Adder_4_U.a ;
assign \add_9s_9s_9_2_1_U13.top_add_9s_9s_9_2_1_Adder_4_U.bin_s0  = \add_9s_9s_9_2_1_U13.top_add_9s_9s_9_2_1_Adder_4_U.b ;
assign \add_9s_9s_9_2_1_U13.top_add_9s_9s_9_2_1_Adder_4_U.s  = { \add_9s_9s_9_2_1_U13.top_add_9s_9s_9_2_1_Adder_4_U.fas_s2 , \add_9s_9s_9_2_1_U13.top_add_9s_9s_9_2_1_Adder_4_U.sum_s1  };
assign \add_9s_9s_9_2_1_U13.top_add_9s_9s_9_2_1_Adder_4_U.u2.a  = \add_9s_9s_9_2_1_U13.top_add_9s_9s_9_2_1_Adder_4_U.ain_s1 ;
assign \add_9s_9s_9_2_1_U13.top_add_9s_9s_9_2_1_Adder_4_U.u2.b  = \add_9s_9s_9_2_1_U13.top_add_9s_9s_9_2_1_Adder_4_U.bin_s1 ;
assign \add_9s_9s_9_2_1_U13.top_add_9s_9s_9_2_1_Adder_4_U.u2.cin  = \add_9s_9s_9_2_1_U13.top_add_9s_9s_9_2_1_Adder_4_U.carry_s1 ;
assign \add_9s_9s_9_2_1_U13.top_add_9s_9s_9_2_1_Adder_4_U.facout_s2  = \add_9s_9s_9_2_1_U13.top_add_9s_9s_9_2_1_Adder_4_U.u2.cout ;
assign \add_9s_9s_9_2_1_U13.top_add_9s_9s_9_2_1_Adder_4_U.fas_s2  = \add_9s_9s_9_2_1_U13.top_add_9s_9s_9_2_1_Adder_4_U.u2.s ;
assign \add_9s_9s_9_2_1_U13.top_add_9s_9s_9_2_1_Adder_4_U.u1.a  = \add_9s_9s_9_2_1_U13.top_add_9s_9s_9_2_1_Adder_4_U.a [3:0];
assign \add_9s_9s_9_2_1_U13.top_add_9s_9s_9_2_1_Adder_4_U.u1.b  = \add_9s_9s_9_2_1_U13.top_add_9s_9s_9_2_1_Adder_4_U.b [3:0];
assign \add_9s_9s_9_2_1_U13.top_add_9s_9s_9_2_1_Adder_4_U.u1.cin  = 1'h0;
assign \add_9s_9s_9_2_1_U13.top_add_9s_9s_9_2_1_Adder_4_U.facout_s1  = \add_9s_9s_9_2_1_U13.top_add_9s_9s_9_2_1_Adder_4_U.u1.cout ;
assign \add_9s_9s_9_2_1_U13.top_add_9s_9s_9_2_1_Adder_4_U.fas_s1  = \add_9s_9s_9_2_1_U13.top_add_9s_9s_9_2_1_Adder_4_U.u1.s ;
assign \add_9s_9s_9_2_1_U13.top_add_9s_9s_9_2_1_Adder_4_U.a  = \add_9s_9s_9_2_1_U13.din0 ;
assign \add_9s_9s_9_2_1_U13.top_add_9s_9s_9_2_1_Adder_4_U.b  = \add_9s_9s_9_2_1_U13.din1 ;
assign \add_9s_9s_9_2_1_U13.top_add_9s_9s_9_2_1_Adder_4_U.ce  = \add_9s_9s_9_2_1_U13.ce ;
assign \add_9s_9s_9_2_1_U13.top_add_9s_9s_9_2_1_Adder_4_U.clk  = \add_9s_9s_9_2_1_U13.clk ;
assign \add_9s_9s_9_2_1_U13.top_add_9s_9s_9_2_1_Adder_4_U.reset  = \add_9s_9s_9_2_1_U13.reset ;
assign \add_9s_9s_9_2_1_U13.dout  = \add_9s_9s_9_2_1_U13.top_add_9s_9s_9_2_1_Adder_4_U.s ;
assign \add_9s_9s_9_2_1_U13.ce  = 1'h1;
assign \add_9s_9s_9_2_1_U13.clk  = ap_clk;
assign \add_9s_9s_9_2_1_U13.din0  = { add_ln69_1_reg_1357[4], add_ln69_1_reg_1357[4], add_ln69_1_reg_1357[4], add_ln69_1_reg_1357[4], add_ln69_1_reg_1357 };
assign \add_9s_9s_9_2_1_U13.din1  = { ret_V_8_reg_1325[7], ret_V_8_reg_1325 };
assign grp_fu_845_p2 = \add_9s_9s_9_2_1_U13.dout ;
assign \add_9s_9s_9_2_1_U13.reset  = ap_rst;
assign \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_5_U.ain_s0  = \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_5_U.a ;
assign \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_5_U.bin_s0  = \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_5_U.b ;
assign \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_5_U.s  = { \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_5_U.fas_s2 , \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_5_U.sum_s1  };
assign \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_5_U.u2.a  = \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_5_U.ain_s1 ;
assign \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_5_U.u2.b  = \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_5_U.bin_s1 ;
assign \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_5_U.u2.cin  = \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_5_U.carry_s1 ;
assign \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_5_U.facout_s2  = \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_5_U.u2.cout ;
assign \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_5_U.fas_s2  = \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_5_U.u2.s ;
assign \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_5_U.u1.a  = \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_5_U.a [3:0];
assign \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_5_U.u1.b  = \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_5_U.b [3:0];
assign \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_5_U.u1.cin  = 1'h0;
assign \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_5_U.facout_s1  = \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_5_U.u1.cout ;
assign \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_5_U.fas_s1  = \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_5_U.u1.s ;
assign \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_5_U.a  = \add_8ns_8ns_8_2_1_U7.din0 ;
assign \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_5_U.b  = \add_8ns_8ns_8_2_1_U7.din1 ;
assign \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_5_U.ce  = \add_8ns_8ns_8_2_1_U7.ce ;
assign \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_5_U.clk  = \add_8ns_8ns_8_2_1_U7.clk ;
assign \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_5_U.reset  = \add_8ns_8ns_8_2_1_U7.reset ;
assign \add_8ns_8ns_8_2_1_U7.dout  = \add_8ns_8ns_8_2_1_U7.top_add_8ns_8ns_8_2_1_Adder_5_U.s ;
assign \add_8ns_8ns_8_2_1_U7.ce  = 1'h1;
assign \add_8ns_8ns_8_2_1_U7.clk  = ap_clk;
assign \add_8ns_8ns_8_2_1_U7.din0  = ret_V_reg_1264;
assign \add_8ns_8ns_8_2_1_U7.din1  = 8'h01;
assign grp_fu_677_p2 = \add_8ns_8ns_8_2_1_U7.dout ;
assign \add_8ns_8ns_8_2_1_U7.reset  = ap_rst;
assign \add_5s_5s_5_2_1_U22.top_add_5s_5s_5_2_1_Adder_15_U.ain_s0  = \add_5s_5s_5_2_1_U22.top_add_5s_5s_5_2_1_Adder_15_U.a ;
assign \add_5s_5s_5_2_1_U22.top_add_5s_5s_5_2_1_Adder_15_U.bin_s0  = \add_5s_5s_5_2_1_U22.top_add_5s_5s_5_2_1_Adder_15_U.b ;
assign \add_5s_5s_5_2_1_U22.top_add_5s_5s_5_2_1_Adder_15_U.s  = { \add_5s_5s_5_2_1_U22.top_add_5s_5s_5_2_1_Adder_15_U.fas_s2 , \add_5s_5s_5_2_1_U22.top_add_5s_5s_5_2_1_Adder_15_U.sum_s1  };
assign \add_5s_5s_5_2_1_U22.top_add_5s_5s_5_2_1_Adder_15_U.u2.a  = \add_5s_5s_5_2_1_U22.top_add_5s_5s_5_2_1_Adder_15_U.ain_s1 ;
assign \add_5s_5s_5_2_1_U22.top_add_5s_5s_5_2_1_Adder_15_U.u2.b  = \add_5s_5s_5_2_1_U22.top_add_5s_5s_5_2_1_Adder_15_U.bin_s1 ;
assign \add_5s_5s_5_2_1_U22.top_add_5s_5s_5_2_1_Adder_15_U.u2.cin  = \add_5s_5s_5_2_1_U22.top_add_5s_5s_5_2_1_Adder_15_U.carry_s1 ;
assign \add_5s_5s_5_2_1_U22.top_add_5s_5s_5_2_1_Adder_15_U.facout_s2  = \add_5s_5s_5_2_1_U22.top_add_5s_5s_5_2_1_Adder_15_U.u2.cout ;
assign \add_5s_5s_5_2_1_U22.top_add_5s_5s_5_2_1_Adder_15_U.fas_s2  = \add_5s_5s_5_2_1_U22.top_add_5s_5s_5_2_1_Adder_15_U.u2.s ;
assign \add_5s_5s_5_2_1_U22.top_add_5s_5s_5_2_1_Adder_15_U.u1.a  = \add_5s_5s_5_2_1_U22.top_add_5s_5s_5_2_1_Adder_15_U.a [1:0];
assign \add_5s_5s_5_2_1_U22.top_add_5s_5s_5_2_1_Adder_15_U.u1.b  = \add_5s_5s_5_2_1_U22.top_add_5s_5s_5_2_1_Adder_15_U.b [1:0];
assign \add_5s_5s_5_2_1_U22.top_add_5s_5s_5_2_1_Adder_15_U.u1.cin  = 1'h0;
assign \add_5s_5s_5_2_1_U22.top_add_5s_5s_5_2_1_Adder_15_U.facout_s1  = \add_5s_5s_5_2_1_U22.top_add_5s_5s_5_2_1_Adder_15_U.u1.cout ;
assign \add_5s_5s_5_2_1_U22.top_add_5s_5s_5_2_1_Adder_15_U.fas_s1  = \add_5s_5s_5_2_1_U22.top_add_5s_5s_5_2_1_Adder_15_U.u1.s ;
assign \add_5s_5s_5_2_1_U22.top_add_5s_5s_5_2_1_Adder_15_U.a  = \add_5s_5s_5_2_1_U22.din0 ;
assign \add_5s_5s_5_2_1_U22.top_add_5s_5s_5_2_1_Adder_15_U.b  = \add_5s_5s_5_2_1_U22.din1 ;
assign \add_5s_5s_5_2_1_U22.top_add_5s_5s_5_2_1_Adder_15_U.ce  = \add_5s_5s_5_2_1_U22.ce ;
assign \add_5s_5s_5_2_1_U22.top_add_5s_5s_5_2_1_Adder_15_U.clk  = \add_5s_5s_5_2_1_U22.clk ;
assign \add_5s_5s_5_2_1_U22.top_add_5s_5s_5_2_1_Adder_15_U.reset  = \add_5s_5s_5_2_1_U22.reset ;
assign \add_5s_5s_5_2_1_U22.dout  = \add_5s_5s_5_2_1_U22.top_add_5s_5s_5_2_1_Adder_15_U.s ;
assign \add_5s_5s_5_2_1_U22.ce  = 1'h1;
assign \add_5s_5s_5_2_1_U22.clk  = ap_clk;
assign \add_5s_5s_5_2_1_U22.din0  = { op_18[3], op_18 };
assign \add_5s_5s_5_2_1_U22.din1  = { op_17[1], op_17[1], op_17[1], op_17 };
assign grp_fu_1023_p2 = \add_5s_5s_5_2_1_U22.dout ;
assign \add_5s_5s_5_2_1_U22.reset  = ap_rst;
assign \add_5s_5ns_5_2_1_U10.top_add_5s_5ns_5_2_1_Adder_8_U.ain_s0  = \add_5s_5ns_5_2_1_U10.top_add_5s_5ns_5_2_1_Adder_8_U.a ;
assign \add_5s_5ns_5_2_1_U10.top_add_5s_5ns_5_2_1_Adder_8_U.bin_s0  = \add_5s_5ns_5_2_1_U10.top_add_5s_5ns_5_2_1_Adder_8_U.b ;
assign \add_5s_5ns_5_2_1_U10.top_add_5s_5ns_5_2_1_Adder_8_U.s  = { \add_5s_5ns_5_2_1_U10.top_add_5s_5ns_5_2_1_Adder_8_U.fas_s2 , \add_5s_5ns_5_2_1_U10.top_add_5s_5ns_5_2_1_Adder_8_U.sum_s1  };
assign \add_5s_5ns_5_2_1_U10.top_add_5s_5ns_5_2_1_Adder_8_U.u2.a  = \add_5s_5ns_5_2_1_U10.top_add_5s_5ns_5_2_1_Adder_8_U.ain_s1 ;
assign \add_5s_5ns_5_2_1_U10.top_add_5s_5ns_5_2_1_Adder_8_U.u2.b  = \add_5s_5ns_5_2_1_U10.top_add_5s_5ns_5_2_1_Adder_8_U.bin_s1 ;
assign \add_5s_5ns_5_2_1_U10.top_add_5s_5ns_5_2_1_Adder_8_U.u2.cin  = \add_5s_5ns_5_2_1_U10.top_add_5s_5ns_5_2_1_Adder_8_U.carry_s1 ;
assign \add_5s_5ns_5_2_1_U10.top_add_5s_5ns_5_2_1_Adder_8_U.facout_s2  = \add_5s_5ns_5_2_1_U10.top_add_5s_5ns_5_2_1_Adder_8_U.u2.cout ;
assign \add_5s_5ns_5_2_1_U10.top_add_5s_5ns_5_2_1_Adder_8_U.fas_s2  = \add_5s_5ns_5_2_1_U10.top_add_5s_5ns_5_2_1_Adder_8_U.u2.s ;
assign \add_5s_5ns_5_2_1_U10.top_add_5s_5ns_5_2_1_Adder_8_U.u1.a  = \add_5s_5ns_5_2_1_U10.top_add_5s_5ns_5_2_1_Adder_8_U.a [1:0];
assign \add_5s_5ns_5_2_1_U10.top_add_5s_5ns_5_2_1_Adder_8_U.u1.b  = \add_5s_5ns_5_2_1_U10.top_add_5s_5ns_5_2_1_Adder_8_U.b [1:0];
assign \add_5s_5ns_5_2_1_U10.top_add_5s_5ns_5_2_1_Adder_8_U.u1.cin  = 1'h0;
assign \add_5s_5ns_5_2_1_U10.top_add_5s_5ns_5_2_1_Adder_8_U.facout_s1  = \add_5s_5ns_5_2_1_U10.top_add_5s_5ns_5_2_1_Adder_8_U.u1.cout ;
assign \add_5s_5ns_5_2_1_U10.top_add_5s_5ns_5_2_1_Adder_8_U.fas_s1  = \add_5s_5ns_5_2_1_U10.top_add_5s_5ns_5_2_1_Adder_8_U.u1.s ;
assign \add_5s_5ns_5_2_1_U10.top_add_5s_5ns_5_2_1_Adder_8_U.a  = \add_5s_5ns_5_2_1_U10.din0 ;
assign \add_5s_5ns_5_2_1_U10.top_add_5s_5ns_5_2_1_Adder_8_U.b  = \add_5s_5ns_5_2_1_U10.din1 ;
assign \add_5s_5ns_5_2_1_U10.top_add_5s_5ns_5_2_1_Adder_8_U.ce  = \add_5s_5ns_5_2_1_U10.ce ;
assign \add_5s_5ns_5_2_1_U10.top_add_5s_5ns_5_2_1_Adder_8_U.clk  = \add_5s_5ns_5_2_1_U10.clk ;
assign \add_5s_5ns_5_2_1_U10.top_add_5s_5ns_5_2_1_Adder_8_U.reset  = \add_5s_5ns_5_2_1_U10.reset ;
assign \add_5s_5ns_5_2_1_U10.dout  = \add_5s_5ns_5_2_1_U10.top_add_5s_5ns_5_2_1_Adder_8_U.s ;
assign \add_5s_5ns_5_2_1_U10.ce  = 1'h1;
assign \add_5s_5ns_5_2_1_U10.clk  = ap_clk;
assign \add_5s_5ns_5_2_1_U10.din0  = { op_15[3], op_15 };
assign \add_5s_5ns_5_2_1_U10.din1  = select_ln69_reg_1254;
assign grp_fu_717_p2 = \add_5s_5ns_5_2_1_U10.dout ;
assign \add_5s_5ns_5_2_1_U10.reset  = ap_rst;
assign \add_5ns_5ns_5_2_1_U9.top_add_5ns_5ns_5_2_1_Adder_7_U.ain_s0  = \add_5ns_5ns_5_2_1_U9.top_add_5ns_5ns_5_2_1_Adder_7_U.a ;
assign \add_5ns_5ns_5_2_1_U9.top_add_5ns_5ns_5_2_1_Adder_7_U.bin_s0  = \add_5ns_5ns_5_2_1_U9.top_add_5ns_5ns_5_2_1_Adder_7_U.b ;
assign \add_5ns_5ns_5_2_1_U9.top_add_5ns_5ns_5_2_1_Adder_7_U.s  = { \add_5ns_5ns_5_2_1_U9.top_add_5ns_5ns_5_2_1_Adder_7_U.fas_s2 , \add_5ns_5ns_5_2_1_U9.top_add_5ns_5ns_5_2_1_Adder_7_U.sum_s1  };
assign \add_5ns_5ns_5_2_1_U9.top_add_5ns_5ns_5_2_1_Adder_7_U.u2.a  = \add_5ns_5ns_5_2_1_U9.top_add_5ns_5ns_5_2_1_Adder_7_U.ain_s1 ;
assign \add_5ns_5ns_5_2_1_U9.top_add_5ns_5ns_5_2_1_Adder_7_U.u2.b  = \add_5ns_5ns_5_2_1_U9.top_add_5ns_5ns_5_2_1_Adder_7_U.bin_s1 ;
assign \add_5ns_5ns_5_2_1_U9.top_add_5ns_5ns_5_2_1_Adder_7_U.u2.cin  = \add_5ns_5ns_5_2_1_U9.top_add_5ns_5ns_5_2_1_Adder_7_U.carry_s1 ;
assign \add_5ns_5ns_5_2_1_U9.top_add_5ns_5ns_5_2_1_Adder_7_U.facout_s2  = \add_5ns_5ns_5_2_1_U9.top_add_5ns_5ns_5_2_1_Adder_7_U.u2.cout ;
assign \add_5ns_5ns_5_2_1_U9.top_add_5ns_5ns_5_2_1_Adder_7_U.fas_s2  = \add_5ns_5ns_5_2_1_U9.top_add_5ns_5ns_5_2_1_Adder_7_U.u2.s ;
assign \add_5ns_5ns_5_2_1_U9.top_add_5ns_5ns_5_2_1_Adder_7_U.u1.a  = \add_5ns_5ns_5_2_1_U9.top_add_5ns_5ns_5_2_1_Adder_7_U.a [1:0];
assign \add_5ns_5ns_5_2_1_U9.top_add_5ns_5ns_5_2_1_Adder_7_U.u1.b  = \add_5ns_5ns_5_2_1_U9.top_add_5ns_5ns_5_2_1_Adder_7_U.b [1:0];
assign \add_5ns_5ns_5_2_1_U9.top_add_5ns_5ns_5_2_1_Adder_7_U.u1.cin  = 1'h0;
assign \add_5ns_5ns_5_2_1_U9.top_add_5ns_5ns_5_2_1_Adder_7_U.facout_s1  = \add_5ns_5ns_5_2_1_U9.top_add_5ns_5ns_5_2_1_Adder_7_U.u1.cout ;
assign \add_5ns_5ns_5_2_1_U9.top_add_5ns_5ns_5_2_1_Adder_7_U.fas_s1  = \add_5ns_5ns_5_2_1_U9.top_add_5ns_5ns_5_2_1_Adder_7_U.u1.s ;
assign \add_5ns_5ns_5_2_1_U9.top_add_5ns_5ns_5_2_1_Adder_7_U.a  = \add_5ns_5ns_5_2_1_U9.din0 ;
assign \add_5ns_5ns_5_2_1_U9.top_add_5ns_5ns_5_2_1_Adder_7_U.b  = \add_5ns_5ns_5_2_1_U9.din1 ;
assign \add_5ns_5ns_5_2_1_U9.top_add_5ns_5ns_5_2_1_Adder_7_U.ce  = \add_5ns_5ns_5_2_1_U9.ce ;
assign \add_5ns_5ns_5_2_1_U9.top_add_5ns_5ns_5_2_1_Adder_7_U.clk  = \add_5ns_5ns_5_2_1_U9.clk ;
assign \add_5ns_5ns_5_2_1_U9.top_add_5ns_5ns_5_2_1_Adder_7_U.reset  = \add_5ns_5ns_5_2_1_U9.reset ;
assign \add_5ns_5ns_5_2_1_U9.dout  = \add_5ns_5ns_5_2_1_U9.top_add_5ns_5ns_5_2_1_Adder_7_U.s ;
assign \add_5ns_5ns_5_2_1_U9.ce  = 1'h1;
assign \add_5ns_5ns_5_2_1_U9.clk  = ap_clk;
assign \add_5ns_5ns_5_2_1_U9.din0  = op_14[7:3];
assign \add_5ns_5ns_5_2_1_U9.din1  = 5'h01;
assign grp_fu_707_p2 = \add_5ns_5ns_5_2_1_U9.dout ;
assign \add_5ns_5ns_5_2_1_U9.reset  = ap_rst;
assign \add_3ns_3ns_3_2_1_U8.top_add_3ns_3ns_3_2_1_Adder_6_U.ain_s0  = \add_3ns_3ns_3_2_1_U8.top_add_3ns_3ns_3_2_1_Adder_6_U.a ;
assign \add_3ns_3ns_3_2_1_U8.top_add_3ns_3ns_3_2_1_Adder_6_U.bin_s0  = \add_3ns_3ns_3_2_1_U8.top_add_3ns_3ns_3_2_1_Adder_6_U.b ;
assign \add_3ns_3ns_3_2_1_U8.top_add_3ns_3ns_3_2_1_Adder_6_U.s  = { \add_3ns_3ns_3_2_1_U8.top_add_3ns_3ns_3_2_1_Adder_6_U.fas_s2 , \add_3ns_3ns_3_2_1_U8.top_add_3ns_3ns_3_2_1_Adder_6_U.sum_s1  };
assign \add_3ns_3ns_3_2_1_U8.top_add_3ns_3ns_3_2_1_Adder_6_U.u2.a  = \add_3ns_3ns_3_2_1_U8.top_add_3ns_3ns_3_2_1_Adder_6_U.ain_s1 ;
assign \add_3ns_3ns_3_2_1_U8.top_add_3ns_3ns_3_2_1_Adder_6_U.u2.b  = \add_3ns_3ns_3_2_1_U8.top_add_3ns_3ns_3_2_1_Adder_6_U.bin_s1 ;
assign \add_3ns_3ns_3_2_1_U8.top_add_3ns_3ns_3_2_1_Adder_6_U.u2.cin  = \add_3ns_3ns_3_2_1_U8.top_add_3ns_3ns_3_2_1_Adder_6_U.carry_s1 ;
assign \add_3ns_3ns_3_2_1_U8.top_add_3ns_3ns_3_2_1_Adder_6_U.facout_s2  = \add_3ns_3ns_3_2_1_U8.top_add_3ns_3ns_3_2_1_Adder_6_U.u2.cout ;
assign \add_3ns_3ns_3_2_1_U8.top_add_3ns_3ns_3_2_1_Adder_6_U.fas_s2  = \add_3ns_3ns_3_2_1_U8.top_add_3ns_3ns_3_2_1_Adder_6_U.u2.s ;
assign \add_3ns_3ns_3_2_1_U8.top_add_3ns_3ns_3_2_1_Adder_6_U.u1.a  = \add_3ns_3ns_3_2_1_U8.top_add_3ns_3ns_3_2_1_Adder_6_U.a [0];
assign \add_3ns_3ns_3_2_1_U8.top_add_3ns_3ns_3_2_1_Adder_6_U.u1.b  = \add_3ns_3ns_3_2_1_U8.top_add_3ns_3ns_3_2_1_Adder_6_U.b [0];
assign \add_3ns_3ns_3_2_1_U8.top_add_3ns_3ns_3_2_1_Adder_6_U.u1.cin  = 1'h0;
assign \add_3ns_3ns_3_2_1_U8.top_add_3ns_3ns_3_2_1_Adder_6_U.facout_s1  = \add_3ns_3ns_3_2_1_U8.top_add_3ns_3ns_3_2_1_Adder_6_U.u1.cout ;
assign \add_3ns_3ns_3_2_1_U8.top_add_3ns_3ns_3_2_1_Adder_6_U.fas_s1  = \add_3ns_3ns_3_2_1_U8.top_add_3ns_3ns_3_2_1_Adder_6_U.u1.s ;
assign \add_3ns_3ns_3_2_1_U8.top_add_3ns_3ns_3_2_1_Adder_6_U.a  = \add_3ns_3ns_3_2_1_U8.din0 ;
assign \add_3ns_3ns_3_2_1_U8.top_add_3ns_3ns_3_2_1_Adder_6_U.b  = \add_3ns_3ns_3_2_1_U8.din1 ;
assign \add_3ns_3ns_3_2_1_U8.top_add_3ns_3ns_3_2_1_Adder_6_U.ce  = \add_3ns_3ns_3_2_1_U8.ce ;
assign \add_3ns_3ns_3_2_1_U8.top_add_3ns_3ns_3_2_1_Adder_6_U.clk  = \add_3ns_3ns_3_2_1_U8.clk ;
assign \add_3ns_3ns_3_2_1_U8.top_add_3ns_3ns_3_2_1_Adder_6_U.reset  = \add_3ns_3ns_3_2_1_U8.reset ;
assign \add_3ns_3ns_3_2_1_U8.dout  = \add_3ns_3ns_3_2_1_U8.top_add_3ns_3ns_3_2_1_Adder_6_U.s ;
assign \add_3ns_3ns_3_2_1_U8.ce  = 1'h1;
assign \add_3ns_3ns_3_2_1_U8.clk  = ap_clk;
assign \add_3ns_3ns_3_2_1_U8.din0  = ret_V_6_reg_1281;
assign \add_3ns_3ns_3_2_1_U8.din1  = 3'h1;
assign grp_fu_682_p2 = \add_3ns_3ns_3_2_1_U8.dout ;
assign \add_3ns_3ns_3_2_1_U8.reset  = ap_rst;
assign \add_34s_34s_34_2_1_U19.top_add_34s_34s_34_2_1_Adder_13_U.ain_s0  = \add_34s_34s_34_2_1_U19.top_add_34s_34s_34_2_1_Adder_13_U.a ;
assign \add_34s_34s_34_2_1_U19.top_add_34s_34s_34_2_1_Adder_13_U.bin_s0  = \add_34s_34s_34_2_1_U19.top_add_34s_34s_34_2_1_Adder_13_U.b ;
assign \add_34s_34s_34_2_1_U19.top_add_34s_34s_34_2_1_Adder_13_U.s  = { \add_34s_34s_34_2_1_U19.top_add_34s_34s_34_2_1_Adder_13_U.fas_s2 , \add_34s_34s_34_2_1_U19.top_add_34s_34s_34_2_1_Adder_13_U.sum_s1  };
assign \add_34s_34s_34_2_1_U19.top_add_34s_34s_34_2_1_Adder_13_U.u2.a  = \add_34s_34s_34_2_1_U19.top_add_34s_34s_34_2_1_Adder_13_U.ain_s1 ;
assign \add_34s_34s_34_2_1_U19.top_add_34s_34s_34_2_1_Adder_13_U.u2.b  = \add_34s_34s_34_2_1_U19.top_add_34s_34s_34_2_1_Adder_13_U.bin_s1 ;
assign \add_34s_34s_34_2_1_U19.top_add_34s_34s_34_2_1_Adder_13_U.u2.cin  = \add_34s_34s_34_2_1_U19.top_add_34s_34s_34_2_1_Adder_13_U.carry_s1 ;
assign \add_34s_34s_34_2_1_U19.top_add_34s_34s_34_2_1_Adder_13_U.facout_s2  = \add_34s_34s_34_2_1_U19.top_add_34s_34s_34_2_1_Adder_13_U.u2.cout ;
assign \add_34s_34s_34_2_1_U19.top_add_34s_34s_34_2_1_Adder_13_U.fas_s2  = \add_34s_34s_34_2_1_U19.top_add_34s_34s_34_2_1_Adder_13_U.u2.s ;
assign \add_34s_34s_34_2_1_U19.top_add_34s_34s_34_2_1_Adder_13_U.u1.a  = \add_34s_34s_34_2_1_U19.top_add_34s_34s_34_2_1_Adder_13_U.a [16:0];
assign \add_34s_34s_34_2_1_U19.top_add_34s_34s_34_2_1_Adder_13_U.u1.b  = \add_34s_34s_34_2_1_U19.top_add_34s_34s_34_2_1_Adder_13_U.b [16:0];
assign \add_34s_34s_34_2_1_U19.top_add_34s_34s_34_2_1_Adder_13_U.u1.cin  = 1'h0;
assign \add_34s_34s_34_2_1_U19.top_add_34s_34s_34_2_1_Adder_13_U.facout_s1  = \add_34s_34s_34_2_1_U19.top_add_34s_34s_34_2_1_Adder_13_U.u1.cout ;
assign \add_34s_34s_34_2_1_U19.top_add_34s_34s_34_2_1_Adder_13_U.fas_s1  = \add_34s_34s_34_2_1_U19.top_add_34s_34s_34_2_1_Adder_13_U.u1.s ;
assign \add_34s_34s_34_2_1_U19.top_add_34s_34s_34_2_1_Adder_13_U.a  = \add_34s_34s_34_2_1_U19.din0 ;
assign \add_34s_34s_34_2_1_U19.top_add_34s_34s_34_2_1_Adder_13_U.b  = \add_34s_34s_34_2_1_U19.din1 ;
assign \add_34s_34s_34_2_1_U19.top_add_34s_34s_34_2_1_Adder_13_U.ce  = \add_34s_34s_34_2_1_U19.ce ;
assign \add_34s_34s_34_2_1_U19.top_add_34s_34s_34_2_1_Adder_13_U.clk  = \add_34s_34s_34_2_1_U19.clk ;
assign \add_34s_34s_34_2_1_U19.top_add_34s_34s_34_2_1_Adder_13_U.reset  = \add_34s_34s_34_2_1_U19.reset ;
assign \add_34s_34s_34_2_1_U19.dout  = \add_34s_34s_34_2_1_U19.top_add_34s_34s_34_2_1_Adder_13_U.s ;
assign \add_34s_34s_34_2_1_U19.ce  = 1'h1;
assign \add_34s_34s_34_2_1_U19.clk  = ap_clk;
assign \add_34s_34s_34_2_1_U19.din0  = { op_25_V_reg_1464[16], op_25_V_reg_1464[16], op_25_V_reg_1464[16], op_25_V_reg_1464[16], op_25_V_reg_1464[16], op_25_V_reg_1464[16], op_25_V_reg_1464[16], op_25_V_reg_1464[16], op_25_V_reg_1464[16], op_25_V_reg_1464[16], op_25_V_reg_1464[16], op_25_V_reg_1464[16], op_25_V_reg_1464[16], op_25_V_reg_1464[16], op_25_V_reg_1464[16], op_25_V_reg_1464[16], op_25_V_reg_1464, 1'h0 };
assign \add_34s_34s_34_2_1_U19.din1  = { op_16[1], op_16[1], op_16[1], op_16[1], op_16[1], op_16[1], op_16[1], op_16[1], op_16[1], op_16[1], op_16[1], op_16[1], op_16[1], op_16[1], op_16[1], op_16[1], op_16[1], op_16[1], op_16[1], op_16[1], op_16[1], op_16[1], op_16[1], op_16[1], op_16[1], op_16[1], op_16[1], op_16[1], op_16[1], op_16[1], op_16[1], op_16[1], op_16 };
assign grp_fu_946_p2 = \add_34s_34s_34_2_1_U19.dout ;
assign \add_34s_34s_34_2_1_U19.reset  = ap_rst;
assign \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_16_U.ain_s0  = \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_16_U.a ;
assign \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_16_U.bin_s0  = \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_16_U.b ;
assign \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_16_U.s  = { \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_16_U.fas_s2 , \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_16_U.sum_s1  };
assign \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_16_U.u2.a  = \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_16_U.ain_s1 ;
assign \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_16_U.u2.b  = \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_16_U.bin_s1 ;
assign \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_16_U.u2.cin  = \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_16_U.carry_s1 ;
assign \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_16_U.facout_s2  = \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_16_U.u2.cout ;
assign \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_16_U.fas_s2  = \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_16_U.u2.s ;
assign \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_16_U.u1.a  = \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_16_U.a [15:0];
assign \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_16_U.u1.b  = \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_16_U.b [15:0];
assign \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_16_U.u1.cin  = 1'h0;
assign \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_16_U.facout_s1  = \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_16_U.u1.cout ;
assign \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_16_U.fas_s1  = \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_16_U.u1.s ;
assign \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_16_U.a  = \add_32s_32ns_32_2_1_U23.din0 ;
assign \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_16_U.b  = \add_32s_32ns_32_2_1_U23.din1 ;
assign \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_16_U.ce  = \add_32s_32ns_32_2_1_U23.ce ;
assign \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_16_U.clk  = \add_32s_32ns_32_2_1_U23.clk ;
assign \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_16_U.reset  = \add_32s_32ns_32_2_1_U23.reset ;
assign \add_32s_32ns_32_2_1_U23.dout  = \add_32s_32ns_32_2_1_U23.top_add_32s_32ns_32_2_1_Adder_16_U.s ;
assign \add_32s_32ns_32_2_1_U23.ce  = 1'h1;
assign \add_32s_32ns_32_2_1_U23.clk  = ap_clk;
assign \add_32s_32ns_32_2_1_U23.din0  = { add_ln69_5_reg_1541[4], add_ln69_5_reg_1541[4], add_ln69_5_reg_1541[4], add_ln69_5_reg_1541[4], add_ln69_5_reg_1541[4], add_ln69_5_reg_1541[4], add_ln69_5_reg_1541[4], add_ln69_5_reg_1541[4], add_ln69_5_reg_1541[4], add_ln69_5_reg_1541[4], add_ln69_5_reg_1541[4], add_ln69_5_reg_1541[4], add_ln69_5_reg_1541[4], add_ln69_5_reg_1541[4], add_ln69_5_reg_1541[4], add_ln69_5_reg_1541[4], add_ln69_5_reg_1541[4], add_ln69_5_reg_1541[4], add_ln69_5_reg_1541[4], add_ln69_5_reg_1541[4], add_ln69_5_reg_1541[4], add_ln69_5_reg_1541[4], add_ln69_5_reg_1541[4], add_ln69_5_reg_1541[4], add_ln69_5_reg_1541[4], add_ln69_5_reg_1541[4], add_ln69_5_reg_1541[4], add_ln69_5_reg_1541 };
assign \add_32s_32ns_32_2_1_U23.din1  = add_ln69_4_reg_1536;
assign grp_fu_1032_p2 = \add_32s_32ns_32_2_1_U23.dout ;
assign \add_32s_32ns_32_2_1_U23.reset  = ap_rst;
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_14_U.ain_s0  = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_14_U.a ;
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_14_U.bin_s0  = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_14_U.b ;
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_14_U.s  = { \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_14_U.fas_s2 , \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_14_U.sum_s1  };
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_14_U.u2.a  = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_14_U.ain_s1 ;
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_14_U.u2.b  = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_14_U.bin_s1 ;
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_14_U.u2.cin  = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_14_U.carry_s1 ;
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_14_U.facout_s2  = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_14_U.u2.cout ;
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_14_U.fas_s2  = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_14_U.u2.s ;
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_14_U.u1.a  = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_14_U.a [15:0];
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_14_U.u1.b  = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_14_U.b [15:0];
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_14_U.u1.cin  = 1'h0;
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_14_U.facout_s1  = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_14_U.u1.cout ;
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_14_U.fas_s1  = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_14_U.u1.s ;
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_14_U.a  = \add_32ns_32ns_32_2_1_U21.din0 ;
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_14_U.b  = \add_32ns_32ns_32_2_1_U21.din1 ;
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_14_U.ce  = \add_32ns_32ns_32_2_1_U21.ce ;
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_14_U.clk  = \add_32ns_32ns_32_2_1_U21.clk ;
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_14_U.reset  = \add_32ns_32ns_32_2_1_U21.reset ;
assign \add_32ns_32ns_32_2_1_U21.dout  = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_14_U.s ;
assign \add_32ns_32ns_32_2_1_U21.ce  = 1'h1;
assign \add_32ns_32ns_32_2_1_U21.clk  = ap_clk;
assign \add_32ns_32ns_32_2_1_U21.din0  = ret_V_27_reg_1516;
assign \add_32ns_32ns_32_2_1_U21.din1  = { 16'h0000, r_reg_1511[1], r_reg_1511[1], r_reg_1511[1], r_reg_1511[1], r_reg_1511[1], r_reg_1511[1], r_reg_1511[1], r_reg_1511[1], r_reg_1511[1], r_reg_1511[1], r_reg_1511[1], r_reg_1511[1], r_reg_1511[1], r_reg_1511[1], r_reg_1511 };
assign grp_fu_1018_p2 = \add_32ns_32ns_32_2_1_U21.dout ;
assign \add_32ns_32ns_32_2_1_U21.reset  = ap_rst;
assign \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_14_U.ain_s0  = \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_14_U.a ;
assign \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_14_U.bin_s0  = \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_14_U.b ;
assign \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_14_U.s  = { \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_14_U.fas_s2 , \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_14_U.sum_s1  };
assign \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_14_U.u2.a  = \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_14_U.ain_s1 ;
assign \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_14_U.u2.b  = \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_14_U.bin_s1 ;
assign \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_14_U.u2.cin  = \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_14_U.carry_s1 ;
assign \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_14_U.facout_s2  = \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_14_U.u2.cout ;
assign \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_14_U.fas_s2  = \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_14_U.u2.s ;
assign \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_14_U.u1.a  = \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_14_U.a [15:0];
assign \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_14_U.u1.b  = \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_14_U.b [15:0];
assign \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_14_U.u1.cin  = 1'h0;
assign \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_14_U.facout_s1  = \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_14_U.u1.cout ;
assign \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_14_U.fas_s1  = \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_14_U.u1.s ;
assign \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_14_U.a  = \add_32ns_32ns_32_2_1_U20.din0 ;
assign \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_14_U.b  = \add_32ns_32ns_32_2_1_U20.din1 ;
assign \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_14_U.ce  = \add_32ns_32ns_32_2_1_U20.ce ;
assign \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_14_U.clk  = \add_32ns_32ns_32_2_1_U20.clk ;
assign \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_14_U.reset  = \add_32ns_32ns_32_2_1_U20.reset ;
assign \add_32ns_32ns_32_2_1_U20.dout  = \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_14_U.s ;
assign \add_32ns_32ns_32_2_1_U20.ce  = 1'h1;
assign \add_32ns_32ns_32_2_1_U20.clk  = ap_clk;
assign \add_32ns_32ns_32_2_1_U20.din0  = ret_V_34_cast_reg_1489;
assign \add_32ns_32ns_32_2_1_U20.din1  = 32'd1;
assign grp_fu_962_p2 = \add_32ns_32ns_32_2_1_U20.dout ;
assign \add_32ns_32ns_32_2_1_U20.reset  = ap_rst;
assign \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_0_U.ain_s0  = \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_0_U.a ;
assign \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_0_U.bin_s0  = \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_0_U.b ;
assign \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_0_U.s  = { \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_0_U.fas_s2 , \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_0_U.sum_s1  };
assign \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_0_U.u2.a  = \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_0_U.ain_s1 ;
assign \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_0_U.u2.b  = \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_0_U.bin_s1 ;
assign \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_0_U.u2.cin  = \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_0_U.carry_s1 ;
assign \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_0_U.facout_s2  = \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_0_U.u2.cout ;
assign \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_0_U.fas_s2  = \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_0_U.u2.s ;
assign \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_0_U.u1.a  = \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_0_U.a [0];
assign \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_0_U.u1.b  = \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_0_U.b [0];
assign \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_0_U.u1.cin  = 1'h0;
assign \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_0_U.facout_s1  = \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_0_U.u1.cout ;
assign \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_0_U.fas_s1  = \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_0_U.u1.s ;
assign \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_0_U.a  = \add_2ns_2ns_2_2_1_U11.din0 ;
assign \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_0_U.b  = \add_2ns_2ns_2_2_1_U11.din1 ;
assign \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_0_U.ce  = \add_2ns_2ns_2_2_1_U11.ce ;
assign \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_0_U.clk  = \add_2ns_2ns_2_2_1_U11.clk ;
assign \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_0_U.reset  = \add_2ns_2ns_2_2_1_U11.reset ;
assign \add_2ns_2ns_2_2_1_U11.dout  = \add_2ns_2ns_2_2_1_U11.top_add_2ns_2ns_2_2_1_Adder_0_U.s ;
assign \add_2ns_2ns_2_2_1_U11.ce  = 1'h1;
assign \add_2ns_2ns_2_2_1_U11.clk  = ap_clk;
assign \add_2ns_2ns_2_2_1_U11.din0  = ret_V_24_cast_reg_1335;
assign \add_2ns_2ns_2_2_1_U11.din1  = 2'h1;
assign grp_fu_786_p2 = \add_2ns_2ns_2_2_1_U11.dout ;
assign \add_2ns_2ns_2_2_1_U11.reset  = ap_rst;
assign \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.ain_s0  = \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.a ;
assign \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.bin_s0  = \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.b ;
assign \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.s  = { \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.fas_s2 , \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.sum_s1  };
assign \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.u2.a  = \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.ain_s1 ;
assign \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.u2.b  = \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.bin_s1 ;
assign \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.u2.cin  = \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.carry_s1 ;
assign \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.facout_s2  = \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.u2.cout ;
assign \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.fas_s2  = \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.u2.s ;
assign \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.u1.a  = \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.a [0];
assign \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.u1.b  = \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.b [0];
assign \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.u1.cin  = 1'h0;
assign \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.facout_s1  = \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.u1.cout ;
assign \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.fas_s1  = \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.u1.s ;
assign \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.a  = \add_2ns_2ns_2_2_1_U1.din0 ;
assign \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.b  = \add_2ns_2ns_2_2_1_U1.din1 ;
assign \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.ce  = \add_2ns_2ns_2_2_1_U1.ce ;
assign \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.clk  = \add_2ns_2ns_2_2_1_U1.clk ;
assign \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.reset  = \add_2ns_2ns_2_2_1_U1.reset ;
assign \add_2ns_2ns_2_2_1_U1.dout  = \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.s ;
assign \add_2ns_2ns_2_2_1_U1.ce  = 1'h1;
assign \add_2ns_2ns_2_2_1_U1.clk  = ap_clk;
assign \add_2ns_2ns_2_2_1_U1.din0  = op_1[1:0];
assign \add_2ns_2ns_2_2_1_U1.din1  = op_0[1:0];
assign grp_fu_253_p2 = \add_2ns_2ns_2_2_1_U1.dout ;
assign \add_2ns_2ns_2_2_1_U1.reset  = ap_rst;
assign \add_29s_29ns_29_2_1_U12.top_add_29s_29ns_29_2_1_Adder_9_U.ain_s0  = \add_29s_29ns_29_2_1_U12.top_add_29s_29ns_29_2_1_Adder_9_U.a ;
assign \add_29s_29ns_29_2_1_U12.top_add_29s_29ns_29_2_1_Adder_9_U.bin_s0  = \add_29s_29ns_29_2_1_U12.top_add_29s_29ns_29_2_1_Adder_9_U.b ;
assign \add_29s_29ns_29_2_1_U12.top_add_29s_29ns_29_2_1_Adder_9_U.s  = { \add_29s_29ns_29_2_1_U12.top_add_29s_29ns_29_2_1_Adder_9_U.fas_s2 , \add_29s_29ns_29_2_1_U12.top_add_29s_29ns_29_2_1_Adder_9_U.sum_s1  };
assign \add_29s_29ns_29_2_1_U12.top_add_29s_29ns_29_2_1_Adder_9_U.u2.a  = \add_29s_29ns_29_2_1_U12.top_add_29s_29ns_29_2_1_Adder_9_U.ain_s1 ;
assign \add_29s_29ns_29_2_1_U12.top_add_29s_29ns_29_2_1_Adder_9_U.u2.b  = \add_29s_29ns_29_2_1_U12.top_add_29s_29ns_29_2_1_Adder_9_U.bin_s1 ;
assign \add_29s_29ns_29_2_1_U12.top_add_29s_29ns_29_2_1_Adder_9_U.u2.cin  = \add_29s_29ns_29_2_1_U12.top_add_29s_29ns_29_2_1_Adder_9_U.carry_s1 ;
assign \add_29s_29ns_29_2_1_U12.top_add_29s_29ns_29_2_1_Adder_9_U.facout_s2  = \add_29s_29ns_29_2_1_U12.top_add_29s_29ns_29_2_1_Adder_9_U.u2.cout ;
assign \add_29s_29ns_29_2_1_U12.top_add_29s_29ns_29_2_1_Adder_9_U.fas_s2  = \add_29s_29ns_29_2_1_U12.top_add_29s_29ns_29_2_1_Adder_9_U.u2.s ;
assign \add_29s_29ns_29_2_1_U12.top_add_29s_29ns_29_2_1_Adder_9_U.u1.a  = \add_29s_29ns_29_2_1_U12.top_add_29s_29ns_29_2_1_Adder_9_U.a [13:0];
assign \add_29s_29ns_29_2_1_U12.top_add_29s_29ns_29_2_1_Adder_9_U.u1.b  = \add_29s_29ns_29_2_1_U12.top_add_29s_29ns_29_2_1_Adder_9_U.b [13:0];
assign \add_29s_29ns_29_2_1_U12.top_add_29s_29ns_29_2_1_Adder_9_U.u1.cin  = 1'h0;
assign \add_29s_29ns_29_2_1_U12.top_add_29s_29ns_29_2_1_Adder_9_U.facout_s1  = \add_29s_29ns_29_2_1_U12.top_add_29s_29ns_29_2_1_Adder_9_U.u1.cout ;
assign \add_29s_29ns_29_2_1_U12.top_add_29s_29ns_29_2_1_Adder_9_U.fas_s1  = \add_29s_29ns_29_2_1_U12.top_add_29s_29ns_29_2_1_Adder_9_U.u1.s ;
assign \add_29s_29ns_29_2_1_U12.top_add_29s_29ns_29_2_1_Adder_9_U.a  = \add_29s_29ns_29_2_1_U12.din0 ;
assign \add_29s_29ns_29_2_1_U12.top_add_29s_29ns_29_2_1_Adder_9_U.b  = \add_29s_29ns_29_2_1_U12.din1 ;
assign \add_29s_29ns_29_2_1_U12.top_add_29s_29ns_29_2_1_Adder_9_U.ce  = \add_29s_29ns_29_2_1_U12.ce ;
assign \add_29s_29ns_29_2_1_U12.top_add_29s_29ns_29_2_1_Adder_9_U.clk  = \add_29s_29ns_29_2_1_U12.clk ;
assign \add_29s_29ns_29_2_1_U12.top_add_29s_29ns_29_2_1_Adder_9_U.reset  = \add_29s_29ns_29_2_1_U12.reset ;
assign \add_29s_29ns_29_2_1_U12.dout  = \add_29s_29ns_29_2_1_U12.top_add_29s_29ns_29_2_1_Adder_9_U.s ;
assign \add_29s_29ns_29_2_1_U12.ce  = 1'h1;
assign \add_29s_29ns_29_2_1_U12.clk  = ap_clk;
assign \add_29s_29ns_29_2_1_U12.din0  = { select_ln850_7_reg_1352[2], select_ln850_7_reg_1352, 25'h0000000 };
assign \add_29s_29ns_29_2_1_U12.din1  = { 3'h0, signbit_reg_1178, 25'h0000000 };
assign grp_fu_833_p2 = \add_29s_29ns_29_2_1_U12.dout ;
assign \add_29s_29ns_29_2_1_U12.reset  = ap_rst;
assign \add_17s_17s_17_2_1_U15.top_add_17s_17s_17_2_1_Adder_11_U.ain_s0  = \add_17s_17s_17_2_1_U15.top_add_17s_17s_17_2_1_Adder_11_U.a ;
assign \add_17s_17s_17_2_1_U15.top_add_17s_17s_17_2_1_Adder_11_U.bin_s0  = \add_17s_17s_17_2_1_U15.top_add_17s_17s_17_2_1_Adder_11_U.b ;
assign \add_17s_17s_17_2_1_U15.top_add_17s_17s_17_2_1_Adder_11_U.s  = { \add_17s_17s_17_2_1_U15.top_add_17s_17s_17_2_1_Adder_11_U.fas_s2 , \add_17s_17s_17_2_1_U15.top_add_17s_17s_17_2_1_Adder_11_U.sum_s1  };
assign \add_17s_17s_17_2_1_U15.top_add_17s_17s_17_2_1_Adder_11_U.u2.a  = \add_17s_17s_17_2_1_U15.top_add_17s_17s_17_2_1_Adder_11_U.ain_s1 ;
assign \add_17s_17s_17_2_1_U15.top_add_17s_17s_17_2_1_Adder_11_U.u2.b  = \add_17s_17s_17_2_1_U15.top_add_17s_17s_17_2_1_Adder_11_U.bin_s1 ;
assign \add_17s_17s_17_2_1_U15.top_add_17s_17s_17_2_1_Adder_11_U.u2.cin  = \add_17s_17s_17_2_1_U15.top_add_17s_17s_17_2_1_Adder_11_U.carry_s1 ;
assign \add_17s_17s_17_2_1_U15.top_add_17s_17s_17_2_1_Adder_11_U.facout_s2  = \add_17s_17s_17_2_1_U15.top_add_17s_17s_17_2_1_Adder_11_U.u2.cout ;
assign \add_17s_17s_17_2_1_U15.top_add_17s_17s_17_2_1_Adder_11_U.fas_s2  = \add_17s_17s_17_2_1_U15.top_add_17s_17s_17_2_1_Adder_11_U.u2.s ;
assign \add_17s_17s_17_2_1_U15.top_add_17s_17s_17_2_1_Adder_11_U.u1.a  = \add_17s_17s_17_2_1_U15.top_add_17s_17s_17_2_1_Adder_11_U.a [7:0];
assign \add_17s_17s_17_2_1_U15.top_add_17s_17s_17_2_1_Adder_11_U.u1.b  = \add_17s_17s_17_2_1_U15.top_add_17s_17s_17_2_1_Adder_11_U.b [7:0];
assign \add_17s_17s_17_2_1_U15.top_add_17s_17s_17_2_1_Adder_11_U.u1.cin  = 1'h0;
assign \add_17s_17s_17_2_1_U15.top_add_17s_17s_17_2_1_Adder_11_U.facout_s1  = \add_17s_17s_17_2_1_U15.top_add_17s_17s_17_2_1_Adder_11_U.u1.cout ;
assign \add_17s_17s_17_2_1_U15.top_add_17s_17s_17_2_1_Adder_11_U.fas_s1  = \add_17s_17s_17_2_1_U15.top_add_17s_17s_17_2_1_Adder_11_U.u1.s ;
assign \add_17s_17s_17_2_1_U15.top_add_17s_17s_17_2_1_Adder_11_U.a  = \add_17s_17s_17_2_1_U15.din0 ;
assign \add_17s_17s_17_2_1_U15.top_add_17s_17s_17_2_1_Adder_11_U.b  = \add_17s_17s_17_2_1_U15.din1 ;
assign \add_17s_17s_17_2_1_U15.top_add_17s_17s_17_2_1_Adder_11_U.ce  = \add_17s_17s_17_2_1_U15.ce ;
assign \add_17s_17s_17_2_1_U15.top_add_17s_17s_17_2_1_Adder_11_U.clk  = \add_17s_17s_17_2_1_U15.clk ;
assign \add_17s_17s_17_2_1_U15.top_add_17s_17s_17_2_1_Adder_11_U.reset  = \add_17s_17s_17_2_1_U15.reset ;
assign \add_17s_17s_17_2_1_U15.dout  = \add_17s_17s_17_2_1_U15.top_add_17s_17s_17_2_1_Adder_11_U.s ;
assign \add_17s_17s_17_2_1_U15.ce  = 1'h1;
assign \add_17s_17s_17_2_1_U15.clk  = ap_clk;
assign \add_17s_17s_17_2_1_U15.din0  = { op_21_V_reg_1408[3], op_21_V_reg_1408[3], op_21_V_reg_1408[3], op_21_V_reg_1408[3], op_21_V_reg_1408[3], op_21_V_reg_1408[3], op_21_V_reg_1408[3], op_21_V_reg_1408[3], op_21_V_reg_1408[3], op_21_V_reg_1408[3], op_21_V_reg_1408[3], op_21_V_reg_1408[3], op_21_V_reg_1408[3], op_21_V_reg_1408 };
assign \add_17s_17s_17_2_1_U15.din1  = { op_13[15], op_13 };
assign grp_fu_896_p2 = \add_17s_17s_17_2_1_U15.dout ;
assign \add_17s_17s_17_2_1_U15.reset  = ap_rst;
assign \add_17s_17ns_17_2_1_U18.top_add_17s_17ns_17_2_1_Adder_12_U.ain_s0  = \add_17s_17ns_17_2_1_U18.top_add_17s_17ns_17_2_1_Adder_12_U.a ;
assign \add_17s_17ns_17_2_1_U18.top_add_17s_17ns_17_2_1_Adder_12_U.bin_s0  = \add_17s_17ns_17_2_1_U18.top_add_17s_17ns_17_2_1_Adder_12_U.b ;
assign \add_17s_17ns_17_2_1_U18.top_add_17s_17ns_17_2_1_Adder_12_U.s  = { \add_17s_17ns_17_2_1_U18.top_add_17s_17ns_17_2_1_Adder_12_U.fas_s2 , \add_17s_17ns_17_2_1_U18.top_add_17s_17ns_17_2_1_Adder_12_U.sum_s1  };
assign \add_17s_17ns_17_2_1_U18.top_add_17s_17ns_17_2_1_Adder_12_U.u2.a  = \add_17s_17ns_17_2_1_U18.top_add_17s_17ns_17_2_1_Adder_12_U.ain_s1 ;
assign \add_17s_17ns_17_2_1_U18.top_add_17s_17ns_17_2_1_Adder_12_U.u2.b  = \add_17s_17ns_17_2_1_U18.top_add_17s_17ns_17_2_1_Adder_12_U.bin_s1 ;
assign \add_17s_17ns_17_2_1_U18.top_add_17s_17ns_17_2_1_Adder_12_U.u2.cin  = \add_17s_17ns_17_2_1_U18.top_add_17s_17ns_17_2_1_Adder_12_U.carry_s1 ;
assign \add_17s_17ns_17_2_1_U18.top_add_17s_17ns_17_2_1_Adder_12_U.facout_s2  = \add_17s_17ns_17_2_1_U18.top_add_17s_17ns_17_2_1_Adder_12_U.u2.cout ;
assign \add_17s_17ns_17_2_1_U18.top_add_17s_17ns_17_2_1_Adder_12_U.fas_s2  = \add_17s_17ns_17_2_1_U18.top_add_17s_17ns_17_2_1_Adder_12_U.u2.s ;
assign \add_17s_17ns_17_2_1_U18.top_add_17s_17ns_17_2_1_Adder_12_U.u1.a  = \add_17s_17ns_17_2_1_U18.top_add_17s_17ns_17_2_1_Adder_12_U.a [7:0];
assign \add_17s_17ns_17_2_1_U18.top_add_17s_17ns_17_2_1_Adder_12_U.u1.b  = \add_17s_17ns_17_2_1_U18.top_add_17s_17ns_17_2_1_Adder_12_U.b [7:0];
assign \add_17s_17ns_17_2_1_U18.top_add_17s_17ns_17_2_1_Adder_12_U.u1.cin  = 1'h0;
assign \add_17s_17ns_17_2_1_U18.top_add_17s_17ns_17_2_1_Adder_12_U.facout_s1  = \add_17s_17ns_17_2_1_U18.top_add_17s_17ns_17_2_1_Adder_12_U.u1.cout ;
assign \add_17s_17ns_17_2_1_U18.top_add_17s_17ns_17_2_1_Adder_12_U.fas_s1  = \add_17s_17ns_17_2_1_U18.top_add_17s_17ns_17_2_1_Adder_12_U.u1.s ;
assign \add_17s_17ns_17_2_1_U18.top_add_17s_17ns_17_2_1_Adder_12_U.a  = \add_17s_17ns_17_2_1_U18.din0 ;
assign \add_17s_17ns_17_2_1_U18.top_add_17s_17ns_17_2_1_Adder_12_U.b  = \add_17s_17ns_17_2_1_U18.din1 ;
assign \add_17s_17ns_17_2_1_U18.top_add_17s_17ns_17_2_1_Adder_12_U.ce  = \add_17s_17ns_17_2_1_U18.ce ;
assign \add_17s_17ns_17_2_1_U18.top_add_17s_17ns_17_2_1_Adder_12_U.clk  = \add_17s_17ns_17_2_1_U18.clk ;
assign \add_17s_17ns_17_2_1_U18.top_add_17s_17ns_17_2_1_Adder_12_U.reset  = \add_17s_17ns_17_2_1_U18.reset ;
assign \add_17s_17ns_17_2_1_U18.dout  = \add_17s_17ns_17_2_1_U18.top_add_17s_17ns_17_2_1_Adder_12_U.s ;
assign \add_17s_17ns_17_2_1_U18.ce  = 1'h1;
assign \add_17s_17ns_17_2_1_U18.clk  = ap_clk;
assign \add_17s_17ns_17_2_1_U18.din0  = { add_ln69_2_reg_1413[8], add_ln69_2_reg_1413[8], add_ln69_2_reg_1413[8], add_ln69_2_reg_1413[8], add_ln69_2_reg_1413[8], add_ln69_2_reg_1413[8], add_ln69_2_reg_1413[8], add_ln69_2_reg_1413[8], add_ln69_2_reg_1413 };
assign \add_17s_17ns_17_2_1_U18.din1  = add_ln69_reg_1454;
assign grp_fu_926_p2 = \add_17s_17ns_17_2_1_U18.dout ;
assign \add_17s_17ns_17_2_1_U18.reset  = ap_rst;
endmodule


// Machine B:
// Processed by function `add_clk_enable_signal` in `verilog_tricks.py`.
// Processed by function `remove_reset_signal` in `verilog_tricks.py`.
module top_B (
  ap_clk,
  ap_start,
  ap_done,
  ap_idle,
  ap_ready,
  op_0,
  op_1,
  op_2,
  op_4,
  op_5,
  op_13,
  op_14,
  op_15,
  op_16,
  op_17,
  op_18,
  op_29,
  op_29_ap_vld,
clk_enable
);
input clk_enable;


input ap_clk;
wire ap_rst;
assign ap_rst = op_29_ap_vld;
input ap_start;
input [7:0] op_0;
input [7:0] op_1;
input [15:0] op_13;
input [7:0] op_14;
input [3:0] op_15;
input [1:0] op_16;
input [1:0] op_17;
input [3:0] op_18;
input [3:0] op_2;
input [31:0] op_4;
input op_5;
output ap_done;
output ap_idle;
output ap_ready;
output [31:0] op_29;
output op_29_ap_vld;


reg Range1_all_ones_reg_1157;
reg [31:0] add_ln691_reg_1340;
reg [4:0] add_ln69_1_reg_1222;
reg [8:0] add_ln69_2_reg_1232;
reg [31:0] add_ln69_4_reg_1350;
reg [4:0] add_ln69_5_reg_1355;
reg [14:0] ap_CS_fsm = 15'h0001;
reg [31:0] conv_i188_reg_1302;
reg icmp_ln850_reg_1152;
reg icmp_ln851_1_reg_1280;
reg icmp_ln851_2_reg_1217;
reg icmp_ln851_3_reg_1270;
reg icmp_ln851_reg_1195;
reg [31:0] \mul_32s_4s_36_7_1_U1.top_mul_32s_4s_36_7_1_Multiplier_0_U.a_reg0 ;
reg [3:0] \mul_32s_4s_36_7_1_U1.top_mul_32s_4s_36_7_1_Multiplier_0_U.b_reg0 ;
reg [35:0] \mul_32s_4s_36_7_1_U1.top_mul_32s_4s_36_7_1_Multiplier_0_U.buff0 ;
reg [35:0] \mul_32s_4s_36_7_1_U1.top_mul_32s_4s_36_7_1_Multiplier_0_U.buff1 ;
reg [35:0] \mul_32s_4s_36_7_1_U1.top_mul_32s_4s_36_7_1_Multiplier_0_U.buff2 ;
reg [35:0] \mul_32s_4s_36_7_1_U1.top_mul_32s_4s_36_7_1_Multiplier_0_U.buff3 ;
reg [35:0] \mul_32s_4s_36_7_1_U1.top_mul_32s_4s_36_7_1_Multiplier_0_U.buff4 ;
reg [3:0] op_21_V_reg_1237;
reg [16:0] op_25_V_reg_1313;
reg [7:0] op_3_V_reg_1058;
reg [3:0] op_6_V_reg_1069;
reg [7:0] op_8_V_reg_1168;
reg [25:0] or_ln1195_reg_1081;
reg overflow_reg_1162;
reg p_Result_11_reg_1102;
reg p_Result_12_reg_1108;
reg p_Result_13_reg_1125;
reg p_Result_14_reg_1131;
reg [7:0] p_Result_s_20_reg_1114;
reg [35:0] r_V_reg_1247;
reg [2:0] ret_V_13_reg_1227;
reg [4:0] ret_V_14_reg_1275;
reg [4:0] ret_V_15_reg_1285;
reg [8:0] ret_V_22_reg_1120;
reg [32:0] ret_V_23_reg_1173;
reg [1:0] ret_V_24_cast_reg_1252;
reg [1:0] ret_V_24_reg_1292;
reg [8:0] ret_V_25_reg_1205;
reg [33:0] ret_V_26_reg_1328;
reg [31:0] ret_V_34_cast_reg_1333;
reg [2:0] ret_V_6_reg_1210;
reg [7:0] ret_V_7_reg_1200;
reg [4:0] ret_V_9_reg_1264;
reg [7:0] ret_V_reg_1178;
reg [15:0] sext_ln69_7_reg_1345;
reg [31:0] \shl_32s_32s_32_2_1_U2.din1_cast_array[0] ;
reg [31:0] \shl_32s_32s_32_2_1_U2.dout_array[0] ;
reg [31:0] shl_ln1497_reg_1323;
reg signbit_reg_1091;
reg [5:0] sub_ln1497_reg_1297;
reg trunc_ln728_reg_1064;
reg [6:0] trunc_ln790_reg_1137;
reg [24:0] trunc_ln851_1_reg_1185;
reg [24:0] trunc_ln851_2_reg_1259;
reg [5:0] trunc_ln851_3_reg_1190;
reg [24:0] trunc_ln851_reg_1086;
reg [9:0] _174_;
wire _000_;
wire [31:0] _001_;
wire [4:0] _002_;
wire [8:0] _003_;
wire [31:0] _004_;
wire [4:0] _005_;
wire [14:0] _006_;
wire [31:0] _007_;
wire _008_;
wire _009_;
wire _010_;
wire _011_;
wire _012_;
wire [3:0] _013_;
wire [16:0] _014_;
wire [1:0] _015_;
wire [3:0] _016_;
wire [7:0] _017_;
wire [25:0] _018_;
wire _019_;
wire _020_;
wire _021_;
wire _022_;
wire _023_;
wire [7:0] _024_;
wire [35:0] _025_;
wire [2:0] _026_;
wire [4:0] _027_;
wire [4:0] _028_;
wire [9:0] _029_;
wire [2:0] _030_;
wire [32:0] _031_;
wire [1:0] _032_;
wire [1:0] _033_;
wire [8:0] _034_;
wire [33:0] _035_;
wire [31:0] _036_;
wire [2:0] _037_;
wire [7:0] _038_;
wire [4:0] _039_;
wire [7:0] _040_;
wire [15:0] _041_;
wire [31:0] _042_;
wire _043_;
wire [5:0] _044_;
wire _045_;
wire _046_;
wire [24:0] _047_;
wire [24:0] _048_;
wire [5:0] _049_;
wire [24:0] _050_;
wire [1:0] _051_;
wire _052_;
wire _053_;
wire _054_;
wire _055_;
wire _056_;
wire _057_;
wire _058_;
wire _059_;
wire _060_;
wire _061_;
wire _062_;
wire _063_;
wire [31:0] _064_;
wire [3:0] _065_;
wire [35:0] _066_;
wire [35:0] _067_;
wire [35:0] _068_;
wire [35:0] _069_;
wire [35:0] _070_;
wire [31:0] _071_;
wire [31:0] _072_;
wire [31:0] _073_;
wire [31:0] _074_;
wire [31:0] _075_;
wire _076_;
wire _077_;
wire _078_;
wire _079_;
wire _080_;
wire _081_;
wire _082_;
wire _083_;
wire _084_;
wire _085_;
wire _086_;
wire _087_;
wire _088_;
wire _089_;
wire _090_;
wire _091_;
wire _092_;
wire Range1_all_ones_fu_435_p2;
wire [31:0] add_ln691_fu_989_p2;
wire [4:0] add_ln69_1_fu_695_p2;
wire [8:0] add_ln69_2_fu_732_p2;
wire [31:0] add_ln69_4_fu_1032_p2;
wire [4:0] add_ln69_5_fu_1038_p2;
wire [16:0] add_ln69_fu_913_p2;
wire [1:0] add_ln731_fu_253_p2;
wire and_ln353_fu_569_p2;
wire and_ln788_1_fu_601_p2;
wire and_ln788_fu_596_p2;
wire ap_CS_fsm_state1;
wire ap_CS_fsm_state10;
wire ap_CS_fsm_state11;
wire ap_CS_fsm_state12;
wire ap_CS_fsm_state13;
wire ap_CS_fsm_state14;
wire ap_CS_fsm_state15;
wire ap_CS_fsm_state2;
wire ap_CS_fsm_state3;
wire ap_CS_fsm_state4;
wire ap_CS_fsm_state5;
wire ap_CS_fsm_state6;
wire ap_CS_fsm_state8;
wire ap_CS_fsm_state9;
wire [14:0] ap_NS_fsm;
wire ap_clk;
wire ap_done;
wire ap_idle;
wire ap_ready;
wire ap_rst;
wire ap_start;
wire [31:0] ashr_ln1497_fu_969_p2;
wire [31:0] conv_i188_fu_894_p1;
wire [35:0] grp_fu_424_p2;
wire [31:0] grp_fu_900_p0;
wire [31:0] grp_fu_900_p1;
wire [31:0] grp_fu_900_p2;
wire icmp_ln785_fu_440_p2;
wire icmp_ln790_fu_479_p2;
wire icmp_ln850_fu_430_p2;
wire icmp_ln851_1_fu_836_p2;
wire icmp_ln851_2_fu_678_p2;
wire icmp_ln851_3_fu_824_p2;
wire icmp_ln851_fu_622_p2;
wire [7:0] lhs_V_2_fu_647_p3;
wire [13:0] lhs_V_fu_334_p3;
wire [25:0] lhs_cast_fu_299_p3;
wire [9:0] lhs_fu_271_p3;
wire \mul_32s_4s_36_7_1_U1.ce ;
wire \mul_32s_4s_36_7_1_U1.clk ;
wire [31:0] \mul_32s_4s_36_7_1_U1.din0 ;
wire [3:0] \mul_32s_4s_36_7_1_U1.din1 ;
wire [35:0] \mul_32s_4s_36_7_1_U1.dout ;
wire \mul_32s_4s_36_7_1_U1.reset ;
wire [31:0] \mul_32s_4s_36_7_1_U1.top_mul_32s_4s_36_7_1_Multiplier_0_U.a ;
wire [3:0] \mul_32s_4s_36_7_1_U1.top_mul_32s_4s_36_7_1_Multiplier_0_U.b ;
wire \mul_32s_4s_36_7_1_U1.top_mul_32s_4s_36_7_1_Multiplier_0_U.ce ;
wire \mul_32s_4s_36_7_1_U1.top_mul_32s_4s_36_7_1_Multiplier_0_U.clk ;
wire [35:0] \mul_32s_4s_36_7_1_U1.top_mul_32s_4s_36_7_1_Multiplier_0_U.p ;
wire [35:0] \mul_32s_4s_36_7_1_U1.top_mul_32s_4s_36_7_1_Multiplier_0_U.tmp_product ;
wire [7:0] op_0;
wire [7:0] op_1;
wire [15:0] op_13;
wire [7:0] op_14;
wire [3:0] op_15;
wire [1:0] op_16;
wire [1:0] op_17;
wire [3:0] op_18;
wire [3:0] op_2;
wire [16:0] op_25_V_fu_922_p2;
wire [31:0] op_29;
wire op_29_ap_vld;
wire [7:0] op_3_V_fu_259_p3;
wire [31:0] op_4;
wire op_5;
wire [7:0] op_8_V_fu_509_p3;
wire [25:0] op_9_V_fu_738_p3;
wire [25:0] or_ln1195_fu_310_p2;
wire or_ln384_1_fu_503_p2;
wire or_ln384_fu_617_p2;
wire or_ln785_fu_445_p2;
wire or_ln788_fu_484_p2;
wire overflow_1_fu_469_p2;
wire overflow_fu_455_p2;
wire p_Result_10_fu_998_p3;
wire p_Result_6_fu_701_p3;
wire p_Result_7_fu_860_p3;
wire p_Result_8_fu_745_p3;
wire p_Result_9_fu_841_p3;
wire [31:0] p_Result_s_fu_562_p1;
wire p_Result_s_fu_562_p3;
wire [1:0] p_Val2_2_fu_580_p4;
wire [7:0] p_Val2_4_fu_461_p1;
wire [28:0] p_Val2_9_fu_780_p2;
wire [1:0] r_fu_981_p3;
wire [1:0] ret_V_10_fu_867_p2;
wire [2:0] ret_V_13_fu_720_p2;
wire [4:0] ret_V_14_fu_830_p2;
wire [4:0] ret_V_15_fu_853_p3;
wire ret_V_19_fu_574_p2;
wire [9:0] ret_V_20_fu_283_p2;
wire [15:0] ret_V_21_fu_348_p2;
wire [15:0] ret_V_21_reg_1096;
wire [8:0] ret_V_22_fu_391_p2;
wire [32:0] ret_V_23_fu_531_p2;
wire [1:0] ret_V_24_fu_878_p3;
wire [8:0] ret_V_25_fu_662_p2;
wire [33:0] ret_V_26_fu_943_p2;
wire [31:0] ret_V_27_fu_1014_p3;
wire [7:0] ret_V_7_fu_627_p2;
wire [7:0] ret_V_8_fu_713_p3;
wire [4:0] ret_V_9_fu_810_p4;
wire [28:0] rhs_1_fu_520_p3;
wire [27:0] rhs_3_fu_768_p3;
wire select_ln1193_fu_383_p0;
wire [8:0] select_ln1193_fu_383_p3;
wire select_ln1498_fu_320_p0;
wire [31:0] select_ln1498_fu_320_p3;
wire [1:0] select_ln384_2_fu_632_p3;
wire [1:0] select_ln384_3_fu_639_p3;
wire [7:0] select_ln384_fu_495_p3;
wire [4:0] select_ln69_fu_683_p3;
wire [1:0] select_ln850_2_fu_872_p3;
wire [4:0] select_ln850_3_fu_848_p3;
wire [31:0] select_ln850_5_fu_1008_p3;
wire [2:0] select_ln850_6_fu_756_p3;
wire [2:0] select_ln850_7_fu_761_p3;
wire [7:0] select_ln850_fu_708_p3;
wire [28:0] sext_ln1192_1_fu_776_p1;
wire [33:0] sext_ln1192_2_fu_939_p1;
wire [8:0] sext_ln1192_fu_655_p1;
wire [32:0] sext_ln1193_fu_527_p1;
wire [9:0] sext_ln1196_fu_279_p1;
wire [5:0] sext_ln1497_fu_885_p1;
wire [16:0] sext_ln21_fu_906_p1;
wire [31:0] sext_ln545_fu_959_p1;
wire [16:0] sext_ln69_1_fu_909_p1;
wire [4:0] sext_ln69_2_fu_691_p1;
wire [8:0] sext_ln69_3_fu_729_p1;
wire [16:0] sext_ln69_4_fu_919_p1;
wire [4:0] sext_ln69_5_fu_1021_p1;
wire [4:0] sext_ln69_6_fu_1025_p1;
wire [15:0] sext_ln69_7_fu_994_p1;
wire [31:0] sext_ln69_8_fu_1044_p1;
wire [8:0] sext_ln69_fu_725_p1;
wire [8:0] sext_ln703_1_fu_380_p1;
wire [31:0] sext_ln703_2_fu_517_p0;
wire [32:0] sext_ln703_2_fu_517_p1;
wire [8:0] sext_ln703_3_fu_659_p1;
wire [1:0] sext_ln703_4_fu_928_p0;
wire [33:0] sext_ln703_4_fu_928_p1;
wire [15:0] sext_ln703_fu_345_p1;
wire \shl_32s_32s_32_2_1_U2.ce ;
wire \shl_32s_32s_32_2_1_U2.clk ;
wire [31:0] \shl_32s_32s_32_2_1_U2.din0 ;
wire [31:0] \shl_32s_32s_32_2_1_U2.din1 ;
wire [31:0] \shl_32s_32s_32_2_1_U2.din1_cast ;
wire [31:0] \shl_32s_32s_32_2_1_U2.din1_mask ;
wire [31:0] \shl_32s_32s_32_2_1_U2.dout ;
wire \shl_32s_32s_32_2_1_U2.reset ;
wire [31:0] signbit_fu_328_p1;
wire signbit_fu_328_p2;
wire [5:0] sub_ln1497_fu_888_p2;
wire tmp_13_fu_962_p3;
wire tmp_1_fu_555_p3;
wire tmp_6_fu_589_p3;
wire [17:0] tmp_fu_932_p3;
wire [31:0] trunc_ln1195_fu_306_p0;
wire [25:0] trunc_ln1195_fu_306_p1;
wire [1:0] trunc_ln1497_1_fu_977_p1;
wire [1:0] trunc_ln1497_fu_974_p1;
wire trunc_ln728_fu_267_p1;
wire [1:0] trunc_ln731_1_fu_249_p1;
wire [1:0] trunc_ln731_fu_245_p1;
wire [6:0] trunc_ln790_fu_413_p1;
wire [24:0] trunc_ln851_1_fu_547_p1;
wire [24:0] trunc_ln851_2_fu_806_p1;
wire [5:0] trunc_ln851_3_fu_551_p1;
wire [2:0] trunc_ln851_4_fu_820_p1;
wire [1:0] trunc_ln851_5_fu_1005_p0;
wire trunc_ln851_5_fu_1005_p1;
wire [24:0] trunc_ln851_fu_316_p1;
wire underflow_1_fu_490_p2;
wire underflow_fu_612_p2;
wire xor_ln785_1_fu_464_p2;
wire xor_ln785_fu_450_p2;
wire xor_ln786_fu_474_p2;
wire xor_ln788_fu_606_p2;
wire [28:0] zext_ln1192_fu_752_p1;
wire [15:0] zext_ln1193_fu_341_p1;
wire [31:0] zext_ln69_fu_1029_p1;


assign add_ln691_fu_989_p2 = ret_V_34_cast_reg_1333 + 1'h1;
assign add_ln69_1_fu_695_p2 = $signed(op_15) + $signed(select_ln69_fu_683_p3);
assign add_ln69_2_fu_732_p2 = $signed(add_ln69_1_reg_1222) + $signed(ret_V_8_fu_713_p3);
assign add_ln69_4_fu_1032_p2 = ret_V_27_fu_1014_p3 + sext_ln69_7_reg_1345;
assign add_ln69_5_fu_1038_p2 = $signed(op_18) + $signed(op_17);
assign add_ln69_fu_913_p2 = $signed(op_21_V_reg_1237) + $signed(op_13);
assign add_ln731_fu_253_p2 = op_1[1:0] + op_0[1:0];
assign op_25_V_fu_922_p2 = $signed(add_ln69_2_reg_1232) + $signed(add_ln69_fu_913_p2);
assign op_29 = $signed(add_ln69_5_reg_1355) + $signed(add_ln69_4_reg_1350);
assign p_Val2_9_fu_780_p2 = $signed({ select_ln850_7_fu_761_p3, 25'h0000000 }) + $signed({ 1'h0, signbit_reg_1091, 25'h0000000 });
assign ret_V_10_fu_867_p2 = ret_V_24_cast_reg_1252 + 1'h1;
assign ret_V_13_fu_720_p2 = ret_V_6_reg_1210 + 1'h1;
assign ret_V_14_fu_830_p2 = op_14[7:3] + 1'h1;
assign ret_V_25_fu_662_p2 = $signed({ select_ln384_3_fu_639_p3, 6'h00 }) + $signed(op_8_V_reg_1168);
assign { ret_V_26_fu_943_p2[33], ret_V_26_fu_943_p2[17:0] } = $signed({ op_25_V_reg_1313, 1'h0 }) + $signed(op_16);
assign ret_V_7_fu_627_p2 = ret_V_reg_1178 + 1'h1;
assign _052_ = ap_CS_fsm[4] & _055_;
assign _053_ = _056_ & ap_CS_fsm[0];
assign _054_ = ap_start & ap_CS_fsm[0];
assign and_ln353_fu_569_p2 = op_4[31] & icmp_ln850_reg_1152;
assign and_ln788_1_fu_601_p2 = p_Result_12_reg_1108 & and_ln788_fu_596_p2;
assign and_ln788_fu_596_p2 = ret_V_21_reg_1096[6] & Range1_all_ones_reg_1157;
assign overflow_1_fu_469_p2 = xor_ln785_1_fu_464_p2 & p_Result_14_reg_1131;
assign overflow_fu_455_p2 = xor_ln785_fu_450_p2 & or_ln785_fu_445_p2;
assign underflow_1_fu_490_p2 = p_Result_13_reg_1125 & or_ln788_fu_484_p2;
assign underflow_fu_612_p2 = xor_ln788_fu_606_p2 & p_Result_11_reg_1102;
assign xor_ln785_1_fu_464_p2 = ~ p_Result_13_reg_1125;
assign xor_ln786_fu_474_p2 = ~ p_Result_14_reg_1131;
assign xor_ln788_fu_606_p2 = ~ and_ln788_1_fu_601_p2;
assign xor_ln785_fu_450_p2 = ~ p_Result_11_reg_1102;
assign _055_ = ~ icmp_ln851_2_reg_1217;
assign _056_ = ~ ap_start;
assign _057_ = p_Result_s_20_reg_1114 == 8'hff;
assign _058_ = ! trunc_ln790_reg_1137;
assign _059_ = ! trunc_ln851_2_reg_1259;
assign _060_ = ! trunc_ln851_3_reg_1190;
assign _061_ = ! op_14[2:0];
assign _062_ = ! trunc_ln851_1_reg_1185;
assign _063_ = select_ln1498_fu_320_p3 == op_4;
assign \mul_32s_4s_36_7_1_U1.top_mul_32s_4s_36_7_1_Multiplier_0_U.tmp_product  = $signed(\mul_32s_4s_36_7_1_U1.top_mul_32s_4s_36_7_1_Multiplier_0_U.a_reg0 ) * $signed(\mul_32s_4s_36_7_1_U1.top_mul_32s_4s_36_7_1_Multiplier_0_U.b_reg0 );
always @(posedge \mul_32s_4s_36_7_1_U1.top_mul_32s_4s_36_7_1_Multiplier_0_U.clk )
\mul_32s_4s_36_7_1_U1.top_mul_32s_4s_36_7_1_Multiplier_0_U.a_reg0  <= _064_;
always @(posedge \mul_32s_4s_36_7_1_U1.top_mul_32s_4s_36_7_1_Multiplier_0_U.clk )
\mul_32s_4s_36_7_1_U1.top_mul_32s_4s_36_7_1_Multiplier_0_U.b_reg0  <= _065_;
always @(posedge \mul_32s_4s_36_7_1_U1.top_mul_32s_4s_36_7_1_Multiplier_0_U.clk )
\mul_32s_4s_36_7_1_U1.top_mul_32s_4s_36_7_1_Multiplier_0_U.buff0  <= _066_;
always @(posedge \mul_32s_4s_36_7_1_U1.top_mul_32s_4s_36_7_1_Multiplier_0_U.clk )
\mul_32s_4s_36_7_1_U1.top_mul_32s_4s_36_7_1_Multiplier_0_U.buff1  <= _067_;
always @(posedge \mul_32s_4s_36_7_1_U1.top_mul_32s_4s_36_7_1_Multiplier_0_U.clk )
\mul_32s_4s_36_7_1_U1.top_mul_32s_4s_36_7_1_Multiplier_0_U.buff2  <= _068_;
always @(posedge \mul_32s_4s_36_7_1_U1.top_mul_32s_4s_36_7_1_Multiplier_0_U.clk )
\mul_32s_4s_36_7_1_U1.top_mul_32s_4s_36_7_1_Multiplier_0_U.buff3  <= _069_;
always @(posedge \mul_32s_4s_36_7_1_U1.top_mul_32s_4s_36_7_1_Multiplier_0_U.clk )
\mul_32s_4s_36_7_1_U1.top_mul_32s_4s_36_7_1_Multiplier_0_U.buff4  <= _070_;
assign _070_ = \mul_32s_4s_36_7_1_U1.top_mul_32s_4s_36_7_1_Multiplier_0_U.ce  ? \mul_32s_4s_36_7_1_U1.top_mul_32s_4s_36_7_1_Multiplier_0_U.buff3  : \mul_32s_4s_36_7_1_U1.top_mul_32s_4s_36_7_1_Multiplier_0_U.buff4 ;
assign _069_ = \mul_32s_4s_36_7_1_U1.top_mul_32s_4s_36_7_1_Multiplier_0_U.ce  ? \mul_32s_4s_36_7_1_U1.top_mul_32s_4s_36_7_1_Multiplier_0_U.buff2  : \mul_32s_4s_36_7_1_U1.top_mul_32s_4s_36_7_1_Multiplier_0_U.buff3 ;
assign _068_ = \mul_32s_4s_36_7_1_U1.top_mul_32s_4s_36_7_1_Multiplier_0_U.ce  ? \mul_32s_4s_36_7_1_U1.top_mul_32s_4s_36_7_1_Multiplier_0_U.buff1  : \mul_32s_4s_36_7_1_U1.top_mul_32s_4s_36_7_1_Multiplier_0_U.buff2 ;
assign _067_ = \mul_32s_4s_36_7_1_U1.top_mul_32s_4s_36_7_1_Multiplier_0_U.ce  ? \mul_32s_4s_36_7_1_U1.top_mul_32s_4s_36_7_1_Multiplier_0_U.buff0  : \mul_32s_4s_36_7_1_U1.top_mul_32s_4s_36_7_1_Multiplier_0_U.buff1 ;
assign _066_ = \mul_32s_4s_36_7_1_U1.top_mul_32s_4s_36_7_1_Multiplier_0_U.ce  ? \mul_32s_4s_36_7_1_U1.top_mul_32s_4s_36_7_1_Multiplier_0_U.tmp_product  : \mul_32s_4s_36_7_1_U1.top_mul_32s_4s_36_7_1_Multiplier_0_U.buff0 ;
assign _065_ = \mul_32s_4s_36_7_1_U1.top_mul_32s_4s_36_7_1_Multiplier_0_U.ce  ? \mul_32s_4s_36_7_1_U1.top_mul_32s_4s_36_7_1_Multiplier_0_U.b  : \mul_32s_4s_36_7_1_U1.top_mul_32s_4s_36_7_1_Multiplier_0_U.b_reg0 ;
assign _064_ = \mul_32s_4s_36_7_1_U1.top_mul_32s_4s_36_7_1_Multiplier_0_U.ce  ? \mul_32s_4s_36_7_1_U1.top_mul_32s_4s_36_7_1_Multiplier_0_U.a  : \mul_32s_4s_36_7_1_U1.top_mul_32s_4s_36_7_1_Multiplier_0_U.a_reg0 ;
always @(posedge \shl_32s_32s_32_2_1_U2.clk )
\shl_32s_32s_32_2_1_U2.dout_array[0]  <= _072_;
always @(posedge \shl_32s_32s_32_2_1_U2.clk )
\shl_32s_32s_32_2_1_U2.din1_cast_array[0]  <= _071_;
assign _073_ = \shl_32s_32s_32_2_1_U2.ce  ? \shl_32s_32s_32_2_1_U2.din1  : \shl_32s_32s_32_2_1_U2.din1_cast_array[0] ;
assign _071_ = \shl_32s_32s_32_2_1_U2.reset  ? 32'd0 : _073_;
assign _074_ = \shl_32s_32s_32_2_1_U2.ce  ? _075_ : \shl_32s_32s_32_2_1_U2.dout_array[0] ;
assign _072_ = \shl_32s_32s_32_2_1_U2.reset  ? 32'd0 : _074_;
assign _075_ = \shl_32s_32s_32_2_1_U2.din0  << { \shl_32s_32s_32_2_1_U2.din1 [31:16], 16'h0000 };
assign \shl_32s_32s_32_2_1_U2.dout  = \shl_32s_32s_32_2_1_U2.dout_array[0]  << \shl_32s_32s_32_2_1_U2.din1_cast_array[0] [15:0];
assign _076_ = | p_Result_s_20_reg_1114;
assign _077_ = | trunc_ln851_reg_1086;
assign or_ln1195_fu_310_p2 = op_4[25:0] | { trunc_ln728_reg_1064, 25'h0000000 };
assign or_ln384_1_fu_503_p2 = underflow_1_fu_490_p2 | overflow_1_fu_469_p2;
assign or_ln384_fu_617_p2 = underflow_fu_612_p2 | overflow_reg_1162;
assign or_ln785_fu_445_p2 = p_Result_12_reg_1108 | icmp_ln785_fu_440_p2;
assign or_ln788_fu_484_p2 = xor_ln786_fu_474_p2 | icmp_ln790_fu_479_p2;
always @(posedge ap_clk)
op_3_V_reg_1058[5:0] <= 6'h00;
always @(posedge ap_clk)
ret_V_22_reg_1120[5:0] <= 6'h00;
always @(posedge ap_clk)
trunc_ln790_reg_1137[5:0] <= 6'h00;
always @(posedge ap_clk)
shl_ln1497_reg_1323 <= _042_;
always @(posedge ap_clk)
ret_V_26_reg_1328 <= _035_;
always @(posedge ap_clk)
ret_V_34_cast_reg_1333 <= _036_;
always @(posedge ap_clk)
ret_V_24_reg_1292 <= _033_;
always @(posedge ap_clk)
sub_ln1497_reg_1297 <= _044_;
always @(posedge ap_clk)
ret_V_13_reg_1227 <= _026_;
always @(posedge ap_clk)
or_ln1195_reg_1081 <= _018_;
always @(posedge ap_clk)
trunc_ln851_reg_1086 <= _050_;
always @(posedge ap_clk)
signbit_reg_1091 <= _043_;
always @(posedge ap_clk)
_174_ <= _029_;
assign ret_V_21_reg_1096[15:6] = _174_;
always @(posedge ap_clk)
p_Result_11_reg_1102 <= _020_;
always @(posedge ap_clk)
p_Result_12_reg_1108 <= _021_;
always @(posedge ap_clk)
p_Result_s_20_reg_1114 <= _024_;
always @(posedge ap_clk)
ret_V_22_reg_1120[8:6] <= _030_;
always @(posedge ap_clk)
p_Result_13_reg_1125 <= _022_;
always @(posedge ap_clk)
p_Result_14_reg_1131 <= _023_;
always @(posedge ap_clk)
trunc_ln790_reg_1137[6] <= _046_;
always @(posedge ap_clk)
op_3_V_reg_1058[7:6] <= _015_;
always @(posedge ap_clk)
trunc_ln728_reg_1064 <= _045_;
always @(posedge ap_clk)
op_6_V_reg_1069 <= _016_;
always @(posedge ap_clk)
op_21_V_reg_1237 <= _013_;
always @(posedge ap_clk)
r_V_reg_1247 <= _025_;
always @(posedge ap_clk)
ret_V_24_cast_reg_1252 <= _032_;
always @(posedge ap_clk)
trunc_ln851_2_reg_1259 <= _048_;
always @(posedge ap_clk)
ret_V_9_reg_1264 <= _039_;
always @(posedge ap_clk)
icmp_ln851_3_reg_1270 <= _011_;
always @(posedge ap_clk)
ret_V_14_reg_1275 <= _027_;
always @(posedge ap_clk)
icmp_ln851_1_reg_1280 <= _009_;
always @(posedge ap_clk)
ret_V_15_reg_1285 <= _028_;
always @(posedge ap_clk)
conv_i188_reg_1302 <= _007_;
always @(posedge ap_clk)
op_25_V_reg_1313 <= _014_;
always @(posedge ap_clk)
add_ln69_4_reg_1350 <= _004_;
always @(posedge ap_clk)
add_ln69_5_reg_1355 <= _005_;
always @(posedge ap_clk)
add_ln69_2_reg_1232 <= _003_;
always @(posedge ap_clk)
icmp_ln851_reg_1195 <= _012_;
always @(posedge ap_clk)
ret_V_7_reg_1200 <= _038_;
always @(posedge ap_clk)
ret_V_25_reg_1205 <= _034_;
always @(posedge ap_clk)
ret_V_6_reg_1210 <= _037_;
always @(posedge ap_clk)
icmp_ln851_2_reg_1217 <= _010_;
always @(posedge ap_clk)
add_ln69_1_reg_1222 <= _002_;
always @(posedge ap_clk)
add_ln691_reg_1340 <= _001_;
always @(posedge ap_clk)
sext_ln69_7_reg_1345 <= _041_;
always @(posedge ap_clk)
icmp_ln850_reg_1152 <= _008_;
always @(posedge ap_clk)
Range1_all_ones_reg_1157 <= _000_;
always @(posedge ap_clk)
overflow_reg_1162 <= _019_;
always @(posedge ap_clk)
op_8_V_reg_1168 <= _017_;
always @(posedge ap_clk)
ret_V_23_reg_1173 <= _031_;
always @(posedge ap_clk)
ret_V_reg_1178 <= _040_;
always @(posedge ap_clk)
trunc_ln851_1_reg_1185 <= _047_;
always @(posedge ap_clk)
trunc_ln851_3_reg_1190 <= _049_;
always @(posedge ap_clk)
ap_CS_fsm <= _006_;
assign _051_ = _054_ ? 2'h2 : 2'h1;
assign _078_ = ap_CS_fsm == 1'h1;
function [14:0] _218_;
input [14:0] a;
input [224:0] b;
input [14:0] s;
case (s)
15'b000000000000001:
_218_ = b[14:0];
15'b000000000000010:
_218_ = b[29:15];
15'b000000000000100:
_218_ = b[44:30];
15'b000000000001000:
_218_ = b[59:45];
15'b000000000010000:
_218_ = b[74:60];
15'b000000000100000:
_218_ = b[89:75];
15'b000000001000000:
_218_ = b[104:90];
15'b000000010000000:
_218_ = b[119:105];
15'b000000100000000:
_218_ = b[134:120];
15'b000001000000000:
_218_ = b[149:135];
15'b000010000000000:
_218_ = b[164:150];
15'b000100000000000:
_218_ = b[179:165];
15'b001000000000000:
_218_ = b[194:180];
15'b010000000000000:
_218_ = b[209:195];
15'b100000000000000:
_218_ = b[224:210];
15'b000000000000000:
_218_ = a;
default:
_218_ = 15'bx;
endcase
endfunction
assign ap_NS_fsm = _218_(15'hxxxx, { 13'h0000, _051_, 210'h00020008002000800200080020008002000800200080020000001 }, { _078_, _092_, _091_, _090_, _089_, _088_, _087_, _086_, _085_, _084_, _083_, _082_, _081_, _080_, _079_ });
assign _079_ = ap_CS_fsm == 15'h4000;
assign _080_ = ap_CS_fsm == 14'h2000;
assign _081_ = ap_CS_fsm == 13'h1000;
assign _082_ = ap_CS_fsm == 12'h800;
assign _083_ = ap_CS_fsm == 11'h400;
assign _084_ = ap_CS_fsm == 10'h200;
assign _085_ = ap_CS_fsm == 9'h100;
assign _086_ = ap_CS_fsm == 8'h80;
assign _087_ = ap_CS_fsm == 7'h40;
assign _088_ = ap_CS_fsm == 6'h20;
assign _089_ = ap_CS_fsm == 5'h10;
assign _090_ = ap_CS_fsm == 4'h8;
assign _091_ = ap_CS_fsm == 3'h4;
assign _092_ = ap_CS_fsm == 2'h2;
assign op_29_ap_vld = ap_CS_fsm[14] ? 1'h1 : 1'h0;
assign ap_idle = _053_ ? 1'h1 : 1'h0;
assign _036_ = ap_CS_fsm[11] ? { ret_V_26_fu_943_p2[33], ret_V_26_fu_943_p2[33], ret_V_26_fu_943_p2[33], ret_V_26_fu_943_p2[33], ret_V_26_fu_943_p2[33], ret_V_26_fu_943_p2[33], ret_V_26_fu_943_p2[33], ret_V_26_fu_943_p2[33], ret_V_26_fu_943_p2[33], ret_V_26_fu_943_p2[33], ret_V_26_fu_943_p2[33], ret_V_26_fu_943_p2[33], ret_V_26_fu_943_p2[33], ret_V_26_fu_943_p2[33], ret_V_26_fu_943_p2[33], ret_V_26_fu_943_p2[17:1] } : ret_V_34_cast_reg_1333;
assign _035_ = ap_CS_fsm[11] ? { ret_V_26_fu_943_p2[33], ret_V_26_fu_943_p2[33], ret_V_26_fu_943_p2[33], ret_V_26_fu_943_p2[33], ret_V_26_fu_943_p2[33], ret_V_26_fu_943_p2[33], ret_V_26_fu_943_p2[33], ret_V_26_fu_943_p2[33], ret_V_26_fu_943_p2[33], ret_V_26_fu_943_p2[33], ret_V_26_fu_943_p2[33], ret_V_26_fu_943_p2[33], ret_V_26_fu_943_p2[33], ret_V_26_fu_943_p2[33], ret_V_26_fu_943_p2[33], ret_V_26_fu_943_p2[33], ret_V_26_fu_943_p2[17:0] } : ret_V_26_reg_1328;
assign _042_ = ap_CS_fsm[11] ? grp_fu_900_p2 : shl_ln1497_reg_1323;
assign _044_ = ap_CS_fsm[9] ? sub_ln1497_fu_888_p2 : sub_ln1497_reg_1297;
assign _033_ = ap_CS_fsm[9] ? ret_V_24_fu_878_p3 : ret_V_24_reg_1292;
assign _026_ = _052_ ? ret_V_13_fu_720_p2 : ret_V_13_reg_1227;
assign _046_ = ap_CS_fsm[1] ? ret_V_22_fu_391_p2[6] : trunc_ln790_reg_1137[6];
assign _023_ = ap_CS_fsm[1] ? ret_V_22_fu_391_p2[7] : p_Result_14_reg_1131;
assign _022_ = ap_CS_fsm[1] ? ret_V_22_fu_391_p2[8] : p_Result_13_reg_1125;
assign _030_ = ap_CS_fsm[1] ? ret_V_22_fu_391_p2[8:6] : ret_V_22_reg_1120[8:6];
assign _024_ = ap_CS_fsm[1] ? ret_V_21_fu_348_p2[15:8] : p_Result_s_20_reg_1114;
assign _021_ = ap_CS_fsm[1] ? ret_V_21_fu_348_p2[7] : p_Result_12_reg_1108;
assign _020_ = ap_CS_fsm[1] ? ret_V_21_fu_348_p2[15] : p_Result_11_reg_1102;
assign _029_ = ap_CS_fsm[1] ? ret_V_21_fu_348_p2[15:6] : ret_V_21_reg_1096[15:6];
assign _043_ = ap_CS_fsm[1] ? signbit_fu_328_p2 : signbit_reg_1091;
assign _050_ = ap_CS_fsm[1] ? or_ln1195_fu_310_p2[24:0] : trunc_ln851_reg_1086;
assign _018_ = ap_CS_fsm[1] ? or_ln1195_fu_310_p2 : or_ln1195_reg_1081;
assign _016_ = ap_CS_fsm[0] ? ret_V_20_fu_283_p2[9:6] : op_6_V_reg_1069;
assign _045_ = ap_CS_fsm[0] ? op_2[0] : trunc_ln728_reg_1064;
assign _015_ = ap_CS_fsm[0] ? add_ln731_fu_253_p2 : op_3_V_reg_1058[7:6];
assign _013_ = ap_CS_fsm[5] ? p_Val2_9_fu_780_p2[28:25] : op_21_V_reg_1237;
assign _027_ = ap_CS_fsm[7] ? ret_V_14_fu_830_p2 : ret_V_14_reg_1275;
assign _011_ = ap_CS_fsm[7] ? icmp_ln851_3_fu_824_p2 : icmp_ln851_3_reg_1270;
assign _039_ = ap_CS_fsm[7] ? op_14[7:3] : ret_V_9_reg_1264;
assign _048_ = ap_CS_fsm[7] ? grp_fu_424_p2[24:0] : trunc_ln851_2_reg_1259;
assign _032_ = ap_CS_fsm[7] ? grp_fu_424_p2[26:25] : ret_V_24_cast_reg_1252;
assign _025_ = ap_CS_fsm[7] ? grp_fu_424_p2 : r_V_reg_1247;
assign _028_ = ap_CS_fsm[8] ? ret_V_15_fu_853_p3 : ret_V_15_reg_1285;
assign _009_ = ap_CS_fsm[8] ? icmp_ln851_1_fu_836_p2 : icmp_ln851_1_reg_1280;
assign _014_ = ap_CS_fsm[10] ? op_25_V_fu_922_p2 : op_25_V_reg_1313;
assign _007_ = ap_CS_fsm[10] ? { ret_V_24_reg_1292[1], ret_V_24_reg_1292[1], ret_V_24_reg_1292[1], ret_V_24_reg_1292[1], ret_V_24_reg_1292[1], ret_V_24_reg_1292[1], ret_V_24_reg_1292[1], ret_V_24_reg_1292[1], ret_V_24_reg_1292[1], ret_V_24_reg_1292[1], ret_V_24_reg_1292[1], ret_V_24_reg_1292[1], ret_V_24_reg_1292[1], ret_V_24_reg_1292[1], ret_V_24_reg_1292[1], ret_V_24_reg_1292[1], ret_V_24_reg_1292[1], ret_V_24_reg_1292[1], ret_V_24_reg_1292[1], ret_V_24_reg_1292[1], ret_V_24_reg_1292[1], ret_V_24_reg_1292[1], ret_V_24_reg_1292[1], ret_V_24_reg_1292[1], ret_V_24_reg_1292[1], ret_V_24_reg_1292[1], ret_V_24_reg_1292[1], ret_V_24_reg_1292[1], ret_V_24_reg_1292[1], ret_V_24_reg_1292[1], ret_V_24_reg_1292 } : conv_i188_reg_1302;
assign _005_ = ap_CS_fsm[13] ? add_ln69_5_fu_1038_p2 : add_ln69_5_reg_1355;
assign _004_ = ap_CS_fsm[13] ? add_ln69_4_fu_1032_p2 : add_ln69_4_reg_1350;
assign _003_ = ap_CS_fsm[4] ? add_ln69_2_fu_732_p2 : add_ln69_2_reg_1232;
assign _002_ = ap_CS_fsm[3] ? add_ln69_1_fu_695_p2 : add_ln69_1_reg_1222;
assign _010_ = ap_CS_fsm[3] ? icmp_ln851_2_fu_678_p2 : icmp_ln851_2_reg_1217;
assign _037_ = ap_CS_fsm[3] ? ret_V_25_fu_662_p2[8:6] : ret_V_6_reg_1210;
assign _034_ = ap_CS_fsm[3] ? ret_V_25_fu_662_p2 : ret_V_25_reg_1205;
assign _038_ = ap_CS_fsm[3] ? ret_V_7_fu_627_p2 : ret_V_7_reg_1200;
assign _012_ = ap_CS_fsm[3] ? icmp_ln851_fu_622_p2 : icmp_ln851_reg_1195;
assign _041_ = ap_CS_fsm[12] ? { r_fu_981_p3[1], r_fu_981_p3[1], r_fu_981_p3[1], r_fu_981_p3[1], r_fu_981_p3[1], r_fu_981_p3[1], r_fu_981_p3[1], r_fu_981_p3[1], r_fu_981_p3[1], r_fu_981_p3[1], r_fu_981_p3[1], r_fu_981_p3[1], r_fu_981_p3[1], r_fu_981_p3[1], r_fu_981_p3 } : sext_ln69_7_reg_1345;
assign _001_ = ap_CS_fsm[12] ? add_ln691_fu_989_p2 : add_ln691_reg_1340;
assign _049_ = ap_CS_fsm[2] ? op_8_V_fu_509_p3[5:0] : trunc_ln851_3_reg_1190;
assign _047_ = ap_CS_fsm[2] ? ret_V_23_fu_531_p2[24:0] : trunc_ln851_1_reg_1185;
assign _040_ = ap_CS_fsm[2] ? ret_V_23_fu_531_p2[32:25] : ret_V_reg_1178;
assign _031_ = ap_CS_fsm[2] ? ret_V_23_fu_531_p2 : ret_V_23_reg_1173;
assign _017_ = ap_CS_fsm[2] ? op_8_V_fu_509_p3 : op_8_V_reg_1168;
assign _019_ = ap_CS_fsm[2] ? overflow_fu_455_p2 : overflow_reg_1162;
assign _000_ = ap_CS_fsm[2] ? Range1_all_ones_fu_435_p2 : Range1_all_ones_reg_1157;
assign _008_ = ap_CS_fsm[2] ? icmp_ln850_fu_430_p2 : icmp_ln850_reg_1152;
assign _006_ = ap_rst ? 15'h0001 : ap_NS_fsm;
assign trunc_ln1497_1_fu_977_p1 = $signed(conv_i188_reg_1302) >>> { ret_V_15_reg_1285[4], ret_V_15_reg_1285[4], ret_V_15_reg_1285[4], ret_V_15_reg_1285[4], ret_V_15_reg_1285[4], ret_V_15_reg_1285[4], ret_V_15_reg_1285[4], ret_V_15_reg_1285[4], ret_V_15_reg_1285[4], ret_V_15_reg_1285[4], ret_V_15_reg_1285[4], ret_V_15_reg_1285[4], ret_V_15_reg_1285[4], ret_V_15_reg_1285[4], ret_V_15_reg_1285[4], ret_V_15_reg_1285[4], ret_V_15_reg_1285[4], ret_V_15_reg_1285[4], ret_V_15_reg_1285[4], ret_V_15_reg_1285[4], ret_V_15_reg_1285[4], ret_V_15_reg_1285[4], ret_V_15_reg_1285[4], ret_V_15_reg_1285[4], ret_V_15_reg_1285[4], ret_V_15_reg_1285[4], ret_V_15_reg_1285[4], ret_V_15_reg_1285 };
assign ret_V_21_fu_348_p2 = $signed({ 1'h0, op_1, 6'h00 }) - $signed(op_3_V_reg_1058);
assign ret_V_22_fu_391_p2 = $signed(op_3_V_reg_1058) - $signed(select_ln1193_fu_383_p3);
assign ret_V_23_fu_531_p2 = $signed(op_4) - $signed({ op_6_V_reg_1069, 25'h0000000 });
assign sub_ln1497_fu_888_p2 = $signed(1'h0) - $signed(ret_V_15_reg_1285);
assign Range1_all_ones_fu_435_p2 = _057_ ? 1'h1 : 1'h0;
assign icmp_ln785_fu_440_p2 = _076_ ? 1'h1 : 1'h0;
assign icmp_ln790_fu_479_p2 = _058_ ? 1'h1 : 1'h0;
assign icmp_ln850_fu_430_p2 = _077_ ? 1'h1 : 1'h0;
assign icmp_ln851_1_fu_836_p2 = _059_ ? 1'h1 : 1'h0;
assign icmp_ln851_2_fu_678_p2 = _060_ ? 1'h1 : 1'h0;
assign icmp_ln851_3_fu_824_p2 = _061_ ? 1'h1 : 1'h0;
assign icmp_ln851_fu_622_p2 = _062_ ? 1'h1 : 1'h0;
assign op_8_V_fu_509_p3 = or_ln384_1_fu_503_p2 ? select_ln384_fu_495_p3 : ret_V_22_reg_1120[7:0];
assign r_fu_981_p3 = ret_V_15_reg_1285[4] ? shl_ln1497_reg_1323[1:0] : trunc_ln1497_1_fu_977_p1;
assign ret_V_15_fu_853_p3 = op_14[7] ? select_ln850_3_fu_848_p3 : ret_V_9_reg_1264;
assign ret_V_24_fu_878_p3 = r_V_reg_1247[35] ? select_ln850_2_fu_872_p3 : ret_V_24_cast_reg_1252;
assign ret_V_27_fu_1014_p3 = ret_V_26_reg_1328[33] ? select_ln850_5_fu_1008_p3 : ret_V_34_cast_reg_1333;
assign ret_V_8_fu_713_p3 = ret_V_23_reg_1173[32] ? select_ln850_fu_708_p3 : ret_V_reg_1178;
assign select_ln1193_fu_383_p3 = op_5 ? 9'h1c0 : 9'h000;
assign select_ln1498_fu_320_p3 = op_5 ? 32'd4261412864 : 32'd0;
assign select_ln384_2_fu_632_p3 = overflow_reg_1162 ? 2'h1 : 2'h3;
assign select_ln384_3_fu_639_p3 = or_ln384_fu_617_p2 ? select_ln384_2_fu_632_p3 : ret_V_21_reg_1096[7:6];
assign select_ln384_fu_495_p3 = overflow_1_fu_469_p2 ? 8'h7f : 8'h81;
assign select_ln69_fu_683_p3 = ret_V_19_fu_574_p2 ? 5'h1f : 5'h00;
assign select_ln850_2_fu_872_p3 = icmp_ln851_1_reg_1280 ? ret_V_24_cast_reg_1252 : ret_V_10_fu_867_p2;
assign select_ln850_3_fu_848_p3 = icmp_ln851_3_reg_1270 ? ret_V_9_reg_1264 : ret_V_14_reg_1275;
assign select_ln850_5_fu_1008_p3 = op_16[0] ? add_ln691_reg_1340 : ret_V_34_cast_reg_1333;
assign select_ln850_6_fu_756_p3 = icmp_ln851_2_reg_1217 ? ret_V_6_reg_1210 : ret_V_13_reg_1227;
assign select_ln850_7_fu_761_p3 = ret_V_25_reg_1205[8] ? select_ln850_6_fu_756_p3 : ret_V_6_reg_1210;
assign select_ln850_fu_708_p3 = icmp_ln851_reg_1195 ? ret_V_reg_1178 : ret_V_7_reg_1200;
assign signbit_fu_328_p2 = _063_ ? 1'h1 : 1'h0;
assign ret_V_19_fu_574_p2 = or_ln1195_reg_1081[25] ^ and_ln353_fu_569_p2;
assign ret_V_20_fu_283_p2 = { add_ln731_fu_253_p2[1], add_ln731_fu_253_p2[1], add_ln731_fu_253_p2, 6'h00 } ^ { op_2, 6'h00 };
assign ap_CS_fsm_state1 = ap_CS_fsm[0];
assign ap_CS_fsm_state10 = ap_CS_fsm[9];
assign ap_CS_fsm_state11 = ap_CS_fsm[10];
assign ap_CS_fsm_state12 = ap_CS_fsm[11];
assign ap_CS_fsm_state13 = ap_CS_fsm[12];
assign ap_CS_fsm_state14 = ap_CS_fsm[13];
assign ap_CS_fsm_state15 = ap_CS_fsm[14];
assign ap_CS_fsm_state2 = ap_CS_fsm[1];
assign ap_CS_fsm_state3 = ap_CS_fsm[2];
assign ap_CS_fsm_state4 = ap_CS_fsm[3];
assign ap_CS_fsm_state5 = ap_CS_fsm[4];
assign ap_CS_fsm_state6 = ap_CS_fsm[5];
assign ap_CS_fsm_state8 = ap_CS_fsm[7];
assign ap_CS_fsm_state9 = ap_CS_fsm[8];
assign ap_done = op_29_ap_vld;
assign ap_ready = op_29_ap_vld;
assign ashr_ln1497_fu_969_p2[1:0] = trunc_ln1497_1_fu_977_p1;
assign conv_i188_fu_894_p1 = { ret_V_24_reg_1292[1], ret_V_24_reg_1292[1], ret_V_24_reg_1292[1], ret_V_24_reg_1292[1], ret_V_24_reg_1292[1], ret_V_24_reg_1292[1], ret_V_24_reg_1292[1], ret_V_24_reg_1292[1], ret_V_24_reg_1292[1], ret_V_24_reg_1292[1], ret_V_24_reg_1292[1], ret_V_24_reg_1292[1], ret_V_24_reg_1292[1], ret_V_24_reg_1292[1], ret_V_24_reg_1292[1], ret_V_24_reg_1292[1], ret_V_24_reg_1292[1], ret_V_24_reg_1292[1], ret_V_24_reg_1292[1], ret_V_24_reg_1292[1], ret_V_24_reg_1292[1], ret_V_24_reg_1292[1], ret_V_24_reg_1292[1], ret_V_24_reg_1292[1], ret_V_24_reg_1292[1], ret_V_24_reg_1292[1], ret_V_24_reg_1292[1], ret_V_24_reg_1292[1], ret_V_24_reg_1292[1], ret_V_24_reg_1292[1], ret_V_24_reg_1292 };
assign grp_fu_900_p0 = { ret_V_24_reg_1292[1], ret_V_24_reg_1292[1], ret_V_24_reg_1292[1], ret_V_24_reg_1292[1], ret_V_24_reg_1292[1], ret_V_24_reg_1292[1], ret_V_24_reg_1292[1], ret_V_24_reg_1292[1], ret_V_24_reg_1292[1], ret_V_24_reg_1292[1], ret_V_24_reg_1292[1], ret_V_24_reg_1292[1], ret_V_24_reg_1292[1], ret_V_24_reg_1292[1], ret_V_24_reg_1292[1], ret_V_24_reg_1292[1], ret_V_24_reg_1292[1], ret_V_24_reg_1292[1], ret_V_24_reg_1292[1], ret_V_24_reg_1292[1], ret_V_24_reg_1292[1], ret_V_24_reg_1292[1], ret_V_24_reg_1292[1], ret_V_24_reg_1292[1], ret_V_24_reg_1292[1], ret_V_24_reg_1292[1], ret_V_24_reg_1292[1], ret_V_24_reg_1292[1], ret_V_24_reg_1292[1], ret_V_24_reg_1292[1], ret_V_24_reg_1292 };
assign grp_fu_900_p1 = { sub_ln1497_reg_1297[5], sub_ln1497_reg_1297[5], sub_ln1497_reg_1297[5], sub_ln1497_reg_1297[5], sub_ln1497_reg_1297[5], sub_ln1497_reg_1297[5], sub_ln1497_reg_1297[5], sub_ln1497_reg_1297[5], sub_ln1497_reg_1297[5], sub_ln1497_reg_1297[5], sub_ln1497_reg_1297[5], sub_ln1497_reg_1297[5], sub_ln1497_reg_1297[5], sub_ln1497_reg_1297[5], sub_ln1497_reg_1297[5], sub_ln1497_reg_1297[5], sub_ln1497_reg_1297[5], sub_ln1497_reg_1297[5], sub_ln1497_reg_1297[5], sub_ln1497_reg_1297[5], sub_ln1497_reg_1297[5], sub_ln1497_reg_1297[5], sub_ln1497_reg_1297[5], sub_ln1497_reg_1297[5], sub_ln1497_reg_1297[5], sub_ln1497_reg_1297[5], sub_ln1497_reg_1297 };
assign lhs_V_2_fu_647_p3 = { select_ln384_3_fu_639_p3, 6'h00 };
assign lhs_V_fu_334_p3 = { op_1, 6'h00 };
assign lhs_cast_fu_299_p3 = { trunc_ln728_reg_1064, 25'h0000000 };
assign lhs_fu_271_p3 = { op_2, 6'h00 };
assign op_3_V_fu_259_p3 = { add_ln731_fu_253_p2, 6'h00 };
assign op_9_V_fu_738_p3 = { signbit_reg_1091, 25'h0000000 };
assign p_Result_10_fu_998_p3 = ret_V_26_reg_1328[33];
assign p_Result_6_fu_701_p3 = ret_V_23_reg_1173[32];
assign p_Result_7_fu_860_p3 = r_V_reg_1247[35];
assign p_Result_8_fu_745_p3 = ret_V_25_reg_1205[8];
assign p_Result_9_fu_841_p3 = op_14[7];
assign p_Result_s_fu_562_p1 = op_4;
assign p_Result_s_fu_562_p3 = op_4[31];
assign p_Val2_2_fu_580_p4 = ret_V_21_reg_1096[7:6];
assign p_Val2_4_fu_461_p1 = ret_V_22_reg_1120[7:0];
assign ret_V_26_fu_943_p2[32:18] = { ret_V_26_fu_943_p2[33], ret_V_26_fu_943_p2[33], ret_V_26_fu_943_p2[33], ret_V_26_fu_943_p2[33], ret_V_26_fu_943_p2[33], ret_V_26_fu_943_p2[33], ret_V_26_fu_943_p2[33], ret_V_26_fu_943_p2[33], ret_V_26_fu_943_p2[33], ret_V_26_fu_943_p2[33], ret_V_26_fu_943_p2[33], ret_V_26_fu_943_p2[33], ret_V_26_fu_943_p2[33], ret_V_26_fu_943_p2[33], ret_V_26_fu_943_p2[33] };
assign ret_V_9_fu_810_p4 = op_14[7:3];
assign rhs_1_fu_520_p3 = { op_6_V_reg_1069, 25'h0000000 };
assign rhs_3_fu_768_p3 = { select_ln850_7_fu_761_p3, 25'h0000000 };
assign select_ln1193_fu_383_p0 = op_5;
assign select_ln1498_fu_320_p0 = op_5;
assign sext_ln1192_1_fu_776_p1 = { select_ln850_7_fu_761_p3[2], select_ln850_7_fu_761_p3, 25'h0000000 };
assign sext_ln1192_2_fu_939_p1 = { op_25_V_reg_1313[16], op_25_V_reg_1313[16], op_25_V_reg_1313[16], op_25_V_reg_1313[16], op_25_V_reg_1313[16], op_25_V_reg_1313[16], op_25_V_reg_1313[16], op_25_V_reg_1313[16], op_25_V_reg_1313[16], op_25_V_reg_1313[16], op_25_V_reg_1313[16], op_25_V_reg_1313[16], op_25_V_reg_1313[16], op_25_V_reg_1313[16], op_25_V_reg_1313[16], op_25_V_reg_1313[16], op_25_V_reg_1313, 1'h0 };
assign sext_ln1192_fu_655_p1 = { select_ln384_3_fu_639_p3[1], select_ln384_3_fu_639_p3, 6'h00 };
assign sext_ln1193_fu_527_p1 = { op_6_V_reg_1069[3], op_6_V_reg_1069[3], op_6_V_reg_1069[3], op_6_V_reg_1069[3], op_6_V_reg_1069, 25'h0000000 };
assign sext_ln1196_fu_279_p1 = { add_ln731_fu_253_p2[1], add_ln731_fu_253_p2[1], add_ln731_fu_253_p2, 6'h00 };
assign sext_ln1497_fu_885_p1 = { ret_V_15_reg_1285[4], ret_V_15_reg_1285 };
assign sext_ln21_fu_906_p1 = { op_21_V_reg_1237[3], op_21_V_reg_1237[3], op_21_V_reg_1237[3], op_21_V_reg_1237[3], op_21_V_reg_1237[3], op_21_V_reg_1237[3], op_21_V_reg_1237[3], op_21_V_reg_1237[3], op_21_V_reg_1237[3], op_21_V_reg_1237[3], op_21_V_reg_1237[3], op_21_V_reg_1237[3], op_21_V_reg_1237[3], op_21_V_reg_1237 };
assign sext_ln545_fu_959_p1 = { ret_V_15_reg_1285[4], ret_V_15_reg_1285[4], ret_V_15_reg_1285[4], ret_V_15_reg_1285[4], ret_V_15_reg_1285[4], ret_V_15_reg_1285[4], ret_V_15_reg_1285[4], ret_V_15_reg_1285[4], ret_V_15_reg_1285[4], ret_V_15_reg_1285[4], ret_V_15_reg_1285[4], ret_V_15_reg_1285[4], ret_V_15_reg_1285[4], ret_V_15_reg_1285[4], ret_V_15_reg_1285[4], ret_V_15_reg_1285[4], ret_V_15_reg_1285[4], ret_V_15_reg_1285[4], ret_V_15_reg_1285[4], ret_V_15_reg_1285[4], ret_V_15_reg_1285[4], ret_V_15_reg_1285[4], ret_V_15_reg_1285[4], ret_V_15_reg_1285[4], ret_V_15_reg_1285[4], ret_V_15_reg_1285[4], ret_V_15_reg_1285[4], ret_V_15_reg_1285 };
assign sext_ln69_1_fu_909_p1 = { op_13[15], op_13 };
assign sext_ln69_2_fu_691_p1 = { op_15[3], op_15 };
assign sext_ln69_3_fu_729_p1 = { add_ln69_1_reg_1222[4], add_ln69_1_reg_1222[4], add_ln69_1_reg_1222[4], add_ln69_1_reg_1222[4], add_ln69_1_reg_1222 };
assign sext_ln69_4_fu_919_p1 = { add_ln69_2_reg_1232[8], add_ln69_2_reg_1232[8], add_ln69_2_reg_1232[8], add_ln69_2_reg_1232[8], add_ln69_2_reg_1232[8], add_ln69_2_reg_1232[8], add_ln69_2_reg_1232[8], add_ln69_2_reg_1232[8], add_ln69_2_reg_1232 };
assign sext_ln69_5_fu_1021_p1 = { op_17[1], op_17[1], op_17[1], op_17 };
assign sext_ln69_6_fu_1025_p1 = { op_18[3], op_18 };
assign sext_ln69_7_fu_994_p1 = { r_fu_981_p3[1], r_fu_981_p3[1], r_fu_981_p3[1], r_fu_981_p3[1], r_fu_981_p3[1], r_fu_981_p3[1], r_fu_981_p3[1], r_fu_981_p3[1], r_fu_981_p3[1], r_fu_981_p3[1], r_fu_981_p3[1], r_fu_981_p3[1], r_fu_981_p3[1], r_fu_981_p3[1], r_fu_981_p3 };
assign sext_ln69_8_fu_1044_p1 = { add_ln69_5_reg_1355[4], add_ln69_5_reg_1355[4], add_ln69_5_reg_1355[4], add_ln69_5_reg_1355[4], add_ln69_5_reg_1355[4], add_ln69_5_reg_1355[4], add_ln69_5_reg_1355[4], add_ln69_5_reg_1355[4], add_ln69_5_reg_1355[4], add_ln69_5_reg_1355[4], add_ln69_5_reg_1355[4], add_ln69_5_reg_1355[4], add_ln69_5_reg_1355[4], add_ln69_5_reg_1355[4], add_ln69_5_reg_1355[4], add_ln69_5_reg_1355[4], add_ln69_5_reg_1355[4], add_ln69_5_reg_1355[4], add_ln69_5_reg_1355[4], add_ln69_5_reg_1355[4], add_ln69_5_reg_1355[4], add_ln69_5_reg_1355[4], add_ln69_5_reg_1355[4], add_ln69_5_reg_1355[4], add_ln69_5_reg_1355[4], add_ln69_5_reg_1355[4], add_ln69_5_reg_1355[4], add_ln69_5_reg_1355 };
assign sext_ln69_fu_725_p1 = { ret_V_8_fu_713_p3[7], ret_V_8_fu_713_p3 };
assign sext_ln703_1_fu_380_p1 = { op_3_V_reg_1058[7], op_3_V_reg_1058 };
assign sext_ln703_2_fu_517_p0 = op_4;
assign sext_ln703_2_fu_517_p1 = { op_4[31], op_4 };
assign sext_ln703_3_fu_659_p1 = { op_8_V_reg_1168[7], op_8_V_reg_1168 };
assign sext_ln703_4_fu_928_p0 = op_16;
assign sext_ln703_4_fu_928_p1 = { op_16[1], op_16[1], op_16[1], op_16[1], op_16[1], op_16[1], op_16[1], op_16[1], op_16[1], op_16[1], op_16[1], op_16[1], op_16[1], op_16[1], op_16[1], op_16[1], op_16[1], op_16[1], op_16[1], op_16[1], op_16[1], op_16[1], op_16[1], op_16[1], op_16[1], op_16[1], op_16[1], op_16[1], op_16[1], op_16[1], op_16[1], op_16[1], op_16 };
assign sext_ln703_fu_345_p1 = { op_3_V_reg_1058[7], op_3_V_reg_1058[7], op_3_V_reg_1058[7], op_3_V_reg_1058[7], op_3_V_reg_1058[7], op_3_V_reg_1058[7], op_3_V_reg_1058[7], op_3_V_reg_1058[7], op_3_V_reg_1058 };
assign signbit_fu_328_p1 = op_4;
assign tmp_13_fu_962_p3 = ret_V_15_reg_1285[4];
assign tmp_1_fu_555_p3 = or_ln1195_reg_1081[25];
assign tmp_6_fu_589_p3 = ret_V_21_reg_1096[6];
assign tmp_fu_932_p3 = { op_25_V_reg_1313, 1'h0 };
assign trunc_ln1195_fu_306_p0 = op_4;
assign trunc_ln1195_fu_306_p1 = op_4[25:0];
assign trunc_ln1497_fu_974_p1 = shl_ln1497_reg_1323[1:0];
assign trunc_ln728_fu_267_p1 = op_2[0];
assign trunc_ln731_1_fu_249_p1 = op_1[1:0];
assign trunc_ln731_fu_245_p1 = op_0[1:0];
assign trunc_ln790_fu_413_p1 = ret_V_22_fu_391_p2[6:0];
assign trunc_ln851_1_fu_547_p1 = ret_V_23_fu_531_p2[24:0];
assign trunc_ln851_2_fu_806_p1 = grp_fu_424_p2[24:0];
assign trunc_ln851_3_fu_551_p1 = op_8_V_fu_509_p3[5:0];
assign trunc_ln851_4_fu_820_p1 = op_14[2:0];
assign trunc_ln851_5_fu_1005_p0 = op_16;
assign trunc_ln851_5_fu_1005_p1 = op_16[0];
assign trunc_ln851_fu_316_p1 = or_ln1195_fu_310_p2[24:0];
assign zext_ln1192_fu_752_p1 = { 3'h0, signbit_reg_1091, 25'h0000000 };
assign zext_ln1193_fu_341_p1 = { 2'h0, op_1, 6'h00 };
assign zext_ln69_fu_1029_p1 = { 16'h0000, sext_ln69_7_reg_1345 };
assign \shl_32s_32s_32_2_1_U2.din1_cast  = \shl_32s_32s_32_2_1_U2.din1 ;
assign \shl_32s_32s_32_2_1_U2.din1_mask  = 32'd65535;
assign \shl_32s_32s_32_2_1_U2.ce  = 1'h1;
assign \shl_32s_32s_32_2_1_U2.clk  = ap_clk;
assign \shl_32s_32s_32_2_1_U2.din0  = { ret_V_24_reg_1292[1], ret_V_24_reg_1292[1], ret_V_24_reg_1292[1], ret_V_24_reg_1292[1], ret_V_24_reg_1292[1], ret_V_24_reg_1292[1], ret_V_24_reg_1292[1], ret_V_24_reg_1292[1], ret_V_24_reg_1292[1], ret_V_24_reg_1292[1], ret_V_24_reg_1292[1], ret_V_24_reg_1292[1], ret_V_24_reg_1292[1], ret_V_24_reg_1292[1], ret_V_24_reg_1292[1], ret_V_24_reg_1292[1], ret_V_24_reg_1292[1], ret_V_24_reg_1292[1], ret_V_24_reg_1292[1], ret_V_24_reg_1292[1], ret_V_24_reg_1292[1], ret_V_24_reg_1292[1], ret_V_24_reg_1292[1], ret_V_24_reg_1292[1], ret_V_24_reg_1292[1], ret_V_24_reg_1292[1], ret_V_24_reg_1292[1], ret_V_24_reg_1292[1], ret_V_24_reg_1292[1], ret_V_24_reg_1292[1], ret_V_24_reg_1292 };
assign \shl_32s_32s_32_2_1_U2.din1  = { sub_ln1497_reg_1297[5], sub_ln1497_reg_1297[5], sub_ln1497_reg_1297[5], sub_ln1497_reg_1297[5], sub_ln1497_reg_1297[5], sub_ln1497_reg_1297[5], sub_ln1497_reg_1297[5], sub_ln1497_reg_1297[5], sub_ln1497_reg_1297[5], sub_ln1497_reg_1297[5], sub_ln1497_reg_1297[5], sub_ln1497_reg_1297[5], sub_ln1497_reg_1297[5], sub_ln1497_reg_1297[5], sub_ln1497_reg_1297[5], sub_ln1497_reg_1297[5], sub_ln1497_reg_1297[5], sub_ln1497_reg_1297[5], sub_ln1497_reg_1297[5], sub_ln1497_reg_1297[5], sub_ln1497_reg_1297[5], sub_ln1497_reg_1297[5], sub_ln1497_reg_1297[5], sub_ln1497_reg_1297[5], sub_ln1497_reg_1297[5], sub_ln1497_reg_1297[5], sub_ln1497_reg_1297 };
assign grp_fu_900_p2 = \shl_32s_32s_32_2_1_U2.dout ;
assign \shl_32s_32s_32_2_1_U2.reset  = ap_rst;
assign \mul_32s_4s_36_7_1_U1.top_mul_32s_4s_36_7_1_Multiplier_0_U.p  = \mul_32s_4s_36_7_1_U1.top_mul_32s_4s_36_7_1_Multiplier_0_U.buff4 ;
assign \mul_32s_4s_36_7_1_U1.top_mul_32s_4s_36_7_1_Multiplier_0_U.a  = \mul_32s_4s_36_7_1_U1.din0 ;
assign \mul_32s_4s_36_7_1_U1.top_mul_32s_4s_36_7_1_Multiplier_0_U.b  = \mul_32s_4s_36_7_1_U1.din1 ;
assign \mul_32s_4s_36_7_1_U1.top_mul_32s_4s_36_7_1_Multiplier_0_U.ce  = \mul_32s_4s_36_7_1_U1.ce ;
assign \mul_32s_4s_36_7_1_U1.top_mul_32s_4s_36_7_1_Multiplier_0_U.clk  = \mul_32s_4s_36_7_1_U1.clk ;
assign \mul_32s_4s_36_7_1_U1.dout  = \mul_32s_4s_36_7_1_U1.top_mul_32s_4s_36_7_1_Multiplier_0_U.p ;
assign \mul_32s_4s_36_7_1_U1.ce  = 1'h1;
assign \mul_32s_4s_36_7_1_U1.clk  = ap_clk;
assign \mul_32s_4s_36_7_1_U1.din0  = op_4;
assign \mul_32s_4s_36_7_1_U1.din1  = op_6_V_reg_1069;
assign grp_fu_424_p2 = \mul_32s_4s_36_7_1_U1.dout ;
assign \mul_32s_4s_36_7_1_U1.reset  = ap_rst;
endmodule


// Product machine:
module top_A_times_top_B (ap_start, op_0, op_1, op_13, op_14, op_15, op_16, op_17, op_18, op_2, op_4, op_5, ap_clk, unsafe_signal);
input ap_start;
input [7:0] op_0;
input [7:0] op_1;
input [15:0] op_13;
input [7:0] op_14;
input [3:0] op_15;
input [1:0] op_16;
input [1:0] op_17;
input [3:0] op_18;
input [3:0] op_2;
input [31:0] op_4;
input op_5;
input ap_clk;
output unsafe_signal;
reg _setup;
initial _setup = 1'b0;
always @ (posedge ap_clk) _setup <= 1'b1;
reg ap_start_internal;
always @ (posedge ap_clk) if (!_setup) ap_start_internal <= ap_start;
reg [7:0] op_0_internal;
always @ (posedge ap_clk) if (!_setup) op_0_internal <= op_0;
reg [7:0] op_1_internal;
always @ (posedge ap_clk) if (!_setup) op_1_internal <= op_1;
reg [15:0] op_13_internal;
always @ (posedge ap_clk) if (!_setup) op_13_internal <= op_13;
reg [7:0] op_14_internal;
always @ (posedge ap_clk) if (!_setup) op_14_internal <= op_14;
reg [3:0] op_15_internal;
always @ (posedge ap_clk) if (!_setup) op_15_internal <= op_15;
reg [1:0] op_16_internal;
always @ (posedge ap_clk) if (!_setup) op_16_internal <= op_16;
reg [1:0] op_17_internal;
always @ (posedge ap_clk) if (!_setup) op_17_internal <= op_17;
reg [3:0] op_18_internal;
always @ (posedge ap_clk) if (!_setup) op_18_internal <= op_18;
reg [3:0] op_2_internal;
always @ (posedge ap_clk) if (!_setup) op_2_internal <= op_2;
reg [31:0] op_4_internal;
always @ (posedge ap_clk) if (!_setup) op_4_internal <= op_4;
reg op_5_internal;
always @ (posedge ap_clk) if (!_setup) op_5_internal <= op_5;
wire ap_done_A;
wire ap_done_B;
wire ap_done_eq;
assign ap_done_eq = ap_done_A == ap_done_B;
wire ap_idle_A;
wire ap_idle_B;
wire ap_idle_eq;
assign ap_idle_eq = ap_idle_A == ap_idle_B;
wire ap_ready_A;
wire ap_ready_B;
wire ap_ready_eq;
assign ap_ready_eq = ap_ready_A == ap_ready_B;
wire [31:0] op_29_A;
wire [31:0] op_29_B;
wire op_29_eq;
assign op_29_eq = op_29_A == op_29_B;
wire op_29_ap_vld_A;
wire op_29_ap_vld_B;
wire clk_enable_A;
wire clk_enable_B;
assign clk_enable_A = _setup & (~op_29_ap_vld_A | op_29_ap_vld_B);
assign clk_enable_B = _setup;
wire divergent;
assign divergent = ~(ap_done_eq & ap_idle_eq & ap_ready_eq & op_29_eq);
assign unsafe_signal = op_29_ap_vld_A & op_29_ap_vld_B & divergent;
top_A instance_A (
    .ap_clk(ap_clk),
    .clk_enable(clk_enable_A),
    .ap_start(ap_start_internal),
    .op_0(op_0_internal),
    .op_1(op_1_internal),
    .op_13(op_13_internal),
    .op_14(op_14_internal),
    .op_15(op_15_internal),
    .op_16(op_16_internal),
    .op_17(op_17_internal),
    .op_18(op_18_internal),
    .op_2(op_2_internal),
    .op_4(op_4_internal),
    .op_5(op_5_internal),
    .ap_done(ap_done_A),
    .ap_idle(ap_idle_A),
    .ap_ready(ap_ready_A),
    .op_29(op_29_A),
    .op_29_ap_vld(op_29_ap_vld_A)
);
top_B instance_B (
    .ap_clk(ap_clk),
    .clk_enable(clk_enable_B),
    .ap_start(ap_start_internal),
    .op_0(op_0_internal),
    .op_1(op_1_internal),
    .op_13(op_13_internal),
    .op_14(op_14_internal),
    .op_15(op_15_internal),
    .op_16(op_16_internal),
    .op_17(op_17_internal),
    .op_18(op_18_internal),
    .op_2(op_2_internal),
    .op_4(op_4_internal),
    .op_5(op_5_internal),
    .ap_done(ap_done_B),
    .ap_idle(ap_idle_B),
    .ap_ready(ap_ready_B),
    .op_29(op_29_B),
    .op_29_ap_vld(op_29_ap_vld_B)
);
endmodule
