// Processed by function `construct_kairos` in `verilog_tricks.py`.
// Machine A:
// Processed by function `add_clk_enable_signal` in `verilog_tricks.py`.
// Processed by function `remove_reset_signal` in `verilog_tricks.py`.
module top_A (
  ap_clk,
  ap_start,
  ap_done,
  ap_idle,
  ap_ready,
  op_0,
  op_4,
  op_5,
  op_6,
  op_10,
  op_14,
  op_15,
  op_16,
  op_17,
  op_18,
  op_29,
  op_29_ap_vld,
clk_enable
);
input clk_enable;


input ap_clk;
wire ap_rst;
assign ap_rst = op_29_ap_vld;
input ap_start;
input op_0;
input op_10;
input [3:0] op_14;
input [7:0] op_15;
input [1:0] op_16;
input [7:0] op_17;
input op_18;
input [1:0] op_4;
input [3:0] op_5;
input [1:0] op_6;
output ap_done;
output ap_idle;
output ap_ready;
output [31:0] op_29;
output op_29_ap_vld;


reg [4:0] \add_10ns_10ns_10_2_1_U10.top_add_10ns_10ns_10_2_1_Adder_7_U.ain_s1 ;
reg [4:0] \add_10ns_10ns_10_2_1_U10.top_add_10ns_10ns_10_2_1_Adder_7_U.bin_s1 ;
reg \add_10ns_10ns_10_2_1_U10.top_add_10ns_10ns_10_2_1_Adder_7_U.carry_s1 ;
reg [4:0] \add_10ns_10ns_10_2_1_U10.top_add_10ns_10ns_10_2_1_Adder_7_U.sum_s1 ;
reg [5:0] \add_11s_11s_11_2_1_U12.top_add_11s_11s_11_2_1_Adder_9_U.ain_s1 ;
reg [5:0] \add_11s_11s_11_2_1_U12.top_add_11s_11s_11_2_1_Adder_9_U.bin_s1 ;
reg \add_11s_11s_11_2_1_U12.top_add_11s_11s_11_2_1_Adder_9_U.carry_s1 ;
reg [4:0] \add_11s_11s_11_2_1_U12.top_add_11s_11s_11_2_1_Adder_9_U.sum_s1 ;
reg [5:0] \add_12ns_12s_12_2_1_U8.top_add_12ns_12s_12_2_1_Adder_5_U.ain_s1 ;
reg [5:0] \add_12ns_12s_12_2_1_U8.top_add_12ns_12s_12_2_1_Adder_5_U.bin_s1 ;
reg \add_12ns_12s_12_2_1_U8.top_add_12ns_12s_12_2_1_Adder_5_U.carry_s1 ;
reg [5:0] \add_12ns_12s_12_2_1_U8.top_add_12ns_12s_12_2_1_Adder_5_U.sum_s1 ;
reg \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.ain_s1 ;
reg \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.bin_s1 ;
reg \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.carry_s1 ;
reg \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.sum_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.ain_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.bin_s1 ;
reg \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.carry_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.sum_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.ain_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.bin_s1 ;
reg \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.carry_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.sum_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_11_U.ain_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_11_U.bin_s1 ;
reg \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_11_U.carry_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_11_U.sum_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.ain_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.bin_s1 ;
reg \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.carry_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.sum_s1 ;
reg [15:0] \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_12_U.ain_s1 ;
reg [15:0] \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_12_U.bin_s1 ;
reg \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_12_U.carry_s1 ;
reg [15:0] \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_12_U.sum_s1 ;
reg [15:0] \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_16_U.ain_s1 ;
reg [15:0] \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_16_U.bin_s1 ;
reg \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_16_U.carry_s1 ;
reg [15:0] \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_16_U.sum_s1 ;
reg [17:0] \add_36s_36s_36_2_1_U19.top_add_36s_36s_36_2_1_Adder_14_U.ain_s1 ;
reg [17:0] \add_36s_36s_36_2_1_U19.top_add_36s_36s_36_2_1_Adder_14_U.bin_s1 ;
reg \add_36s_36s_36_2_1_U19.top_add_36s_36s_36_2_1_Adder_14_U.carry_s1 ;
reg [17:0] \add_36s_36s_36_2_1_U19.top_add_36s_36s_36_2_1_Adder_14_U.sum_s1 ;
reg [18:0] \add_37s_37s_37_2_1_U13.top_add_37s_37s_37_2_1_Adder_10_U.ain_s1 ;
reg [18:0] \add_37s_37s_37_2_1_U13.top_add_37s_37s_37_2_1_Adder_10_U.bin_s1 ;
reg \add_37s_37s_37_2_1_U13.top_add_37s_37s_37_2_1_Adder_10_U.carry_s1 ;
reg [17:0] \add_37s_37s_37_2_1_U13.top_add_37s_37s_37_2_1_Adder_10_U.sum_s1 ;
reg [18:0] \add_38s_38s_38_2_1_U16.top_add_38s_38s_38_2_1_Adder_13_U.ain_s1 ;
reg [18:0] \add_38s_38s_38_2_1_U16.top_add_38s_38s_38_2_1_Adder_13_U.bin_s1 ;
reg \add_38s_38s_38_2_1_U16.top_add_38s_38s_38_2_1_Adder_13_U.carry_s1 ;
reg [18:0] \add_38s_38s_38_2_1_U16.top_add_38s_38s_38_2_1_Adder_13_U.sum_s1 ;
reg [1:0] \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_3_U.ain_s1 ;
reg [1:0] \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_3_U.bin_s1 ;
reg \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_3_U.carry_s1 ;
reg \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_3_U.sum_s1 ;
reg [1:0] \add_3s_3ns_3_2_1_U7.top_add_3s_3ns_3_2_1_Adder_4_U.ain_s1 ;
reg [1:0] \add_3s_3ns_3_2_1_U7.top_add_3s_3ns_3_2_1_Adder_4_U.bin_s1 ;
reg \add_3s_3ns_3_2_1_U7.top_add_3s_3ns_3_2_1_Adder_4_U.carry_s1 ;
reg \add_3s_3ns_3_2_1_U7.top_add_3s_3ns_3_2_1_Adder_4_U.sum_s1 ;
reg [1:0] \add_4s_4ns_4_2_1_U11.top_add_4s_4ns_4_2_1_Adder_8_U.ain_s1 ;
reg [1:0] \add_4s_4ns_4_2_1_U11.top_add_4s_4ns_4_2_1_Adder_8_U.bin_s1 ;
reg \add_4s_4ns_4_2_1_U11.top_add_4s_4ns_4_2_1_Adder_8_U.carry_s1 ;
reg [1:0] \add_4s_4ns_4_2_1_U11.top_add_4s_4ns_4_2_1_Adder_8_U.sum_s1 ;
reg [2:0] \add_6ns_6s_6_2_1_U9.top_add_6ns_6s_6_2_1_Adder_6_U.ain_s1 ;
reg [2:0] \add_6ns_6s_6_2_1_U9.top_add_6ns_6s_6_2_1_Adder_6_U.bin_s1 ;
reg \add_6ns_6s_6_2_1_U9.top_add_6ns_6s_6_2_1_Adder_6_U.carry_s1 ;
reg [2:0] \add_6ns_6s_6_2_1_U9.top_add_6ns_6s_6_2_1_Adder_6_U.sum_s1 ;
reg [4:0] \add_9ns_9ns_9_2_1_U21.top_add_9ns_9ns_9_2_1_Adder_15_U.ain_s1 ;
reg [4:0] \add_9ns_9ns_9_2_1_U21.top_add_9ns_9ns_9_2_1_Adder_15_U.bin_s1 ;
reg \add_9ns_9ns_9_2_1_U21.top_add_9ns_9ns_9_2_1_Adder_15_U.carry_s1 ;
reg [3:0] \add_9ns_9ns_9_2_1_U21.top_add_9ns_9ns_9_2_1_Adder_15_U.sum_s1 ;
reg [31:0] add_ln691_1_reg_1605;
reg [31:0] add_ln691_2_reg_1652;
reg [31:0] add_ln691_3_reg_1704;
reg [3:0] add_ln691_reg_1523;
reg [8:0] add_ln69_reg_1719;
reg and_ln786_1_reg_1492;
reg and_ln786_reg_1347;
reg [42:0] ap_CS_fsm = 43'h00000000001;
reg icmp_ln768_reg_1291;
reg icmp_ln786_reg_1296;
reg icmp_ln851_1_reg_1217;
reg icmp_ln851_2_reg_1179;
reg icmp_ln851_3_reg_1419;
reg icmp_ln851_4_reg_1588;
reg icmp_ln851_5_reg_1635;
reg icmp_ln851_6_reg_1682;
reg icmp_ln851_reg_1276;
reg [3:0] \mul_4s_2s_6_7_1_U1.top_mul_4s_2s_6_7_1_Mul_DSP_0_U.a_reg0 ;
reg [1:0] \mul_4s_2s_6_7_1_U1.top_mul_4s_2s_6_7_1_Mul_DSP_0_U.b_reg0 ;
reg [5:0] \mul_4s_2s_6_7_1_U1.top_mul_4s_2s_6_7_1_Mul_DSP_0_U.buff0 ;
reg [5:0] \mul_4s_2s_6_7_1_U1.top_mul_4s_2s_6_7_1_Mul_DSP_0_U.buff1 ;
reg [5:0] \mul_4s_2s_6_7_1_U1.top_mul_4s_2s_6_7_1_Mul_DSP_0_U.buff2 ;
reg [5:0] \mul_4s_2s_6_7_1_U1.top_mul_4s_2s_6_7_1_Mul_DSP_0_U.buff3 ;
reg [5:0] \mul_4s_2s_6_7_1_U1.top_mul_4s_2s_6_7_1_Mul_DSP_0_U.buff4 ;
reg [3:0] op_11_V_reg_1389;
reg [7:0] op_13_V_reg_1563;
reg [10:0] op_22_V_reg_1568;
reg [31:0] op_24_V_reg_1620;
reg [31:0] op_26_V_reg_1667;
reg [1:0] or_ln1195_reg_1286;
reg or_ln340_1_reg_1517;
reg or_ln340_reg_1341;
reg or_ln785_1_reg_1480;
reg or_ln785_reg_1312;
reg or_ln786_reg_1335;
reg p_Result_16_reg_1251;
reg p_Result_17_reg_1263;
reg p_Result_19_reg_1441;
reg p_Result_20_reg_1457;
reg [1:0] p_Result_s_18_reg_1270;
reg [3:0] p_Val2_5_reg_1358;
reg [7:0] p_Val2_8_reg_1449;
reg [19:0] r_V_1_reg_1436;
reg [5:0] r_V_reg_1189;
reg [9:0] ret_V_10_reg_1528;
reg [4:0] ret_V_20_reg_1222;
reg [2:0] ret_V_21_reg_1329;
reg [1:0] ret_V_22_reg_1281;
reg [2:0] ret_V_23_reg_1384;
reg [11:0] ret_V_24_reg_1424;
reg [4:0] ret_V_25_reg_1244;
reg [5:0] ret_V_26_reg_1470;
reg [3:0] ret_V_27_reg_1543;
reg [36:0] ret_V_28_reg_1593;
reg [31:0] ret_V_29_cast_reg_1598;
reg [31:0] ret_V_29_reg_1610;
reg [2:0] ret_V_2_reg_1302;
reg [37:0] ret_V_30_reg_1640;
reg [31:0] ret_V_31_cast_reg_1645;
reg [31:0] ret_V_31_reg_1657;
reg [35:0] ret_V_32_reg_1687;
reg [31:0] ret_V_33_cast_reg_1692;
reg [31:0] ret_V_33_reg_1714;
reg [1:0] ret_V_3_cast_reg_1194;
reg [1:0] ret_V_4_reg_1239;
reg [9:0] ret_V_8_reg_1429;
reg [9:0] ret_V_9_reg_1506;
reg [2:0] ret_V_reg_1227;
reg sel_tmp11_reg_1369;
reg sel_tmp24_reg_1538;
reg [7:0] select_ln340_1_reg_1533;
reg [3:0] select_ln340_reg_1364;
reg [8:0] select_ln69_reg_1699;
reg [2:0] select_ln703_reg_1353;
reg [7:0] select_ln785_1_reg_1548;
reg [3:0] select_ln785_reg_1379;
reg [3:0] sext_ln850_reg_1499;
reg [1:0] \shl_20s_2ns_20_7_1_U6.din1_cast_array[0] ;
reg [1:0] \shl_20s_2ns_20_7_1_U6.din1_cast_array[1] ;
reg [1:0] \shl_20s_2ns_20_7_1_U6.din1_cast_array[2] ;
reg [1:0] \shl_20s_2ns_20_7_1_U6.din1_cast_array[3] ;
reg [1:0] \shl_20s_2ns_20_7_1_U6.din1_cast_array[4] ;
reg [1:0] \shl_20s_2ns_20_7_1_U6.din1_cast_array[5] ;
reg [19:0] \shl_20s_2ns_20_7_1_U6.dout_array[0] ;
reg [19:0] \shl_20s_2ns_20_7_1_U6.dout_array[1] ;
reg [19:0] \shl_20s_2ns_20_7_1_U6.dout_array[2] ;
reg [19:0] \shl_20s_2ns_20_7_1_U6.dout_array[3] ;
reg [19:0] \shl_20s_2ns_20_7_1_U6.dout_array[4] ;
reg [19:0] \shl_20s_2ns_20_7_1_U6.dout_array[5] ;
reg [2:0] \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.ain_s1 ;
reg [2:0] \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.bin_s1 ;
reg \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.carry_s1 ;
reg [1:0] \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.sum_s1 ;
reg [2:0] \sub_5s_5s_5_2_1_U2.top_sub_5s_5s_5_2_1_Adder_0_U.ain_s1 ;
reg [2:0] \sub_5s_5s_5_2_1_U2.top_sub_5s_5s_5_2_1_Adder_0_U.bin_s1 ;
reg \sub_5s_5s_5_2_1_U2.top_sub_5s_5s_5_2_1_Adder_0_U.carry_s1 ;
reg [1:0] \sub_5s_5s_5_2_1_U2.top_sub_5s_5s_5_2_1_Adder_0_U.sum_s1 ;
reg tmp_12_reg_1463;
reg [2:0] tmp_3_reg_1475;
reg tmp_reg_1184;
reg [2:0] trunc_ln731_reg_1258;
reg [2:0] trunc_ln851_1_reg_1201;
reg [2:0] trunc_ln851_3_reg_1394;
reg [3:0] trunc_ln851_4_reg_1573;
reg [1:0] trunc_ln851_reg_1234;
reg xor_ln785_1_reg_1486;
reg xor_ln785_reg_1318;
reg xor_ln786_2_reg_1511;
wire [31:0] _000_;
wire [31:0] _001_;
wire [31:0] _002_;
wire [3:0] _003_;
wire [8:0] _004_;
wire _005_;
wire _006_;
wire [42:0] _007_;
wire _008_;
wire _009_;
wire _010_;
wire _011_;
wire _012_;
wire _013_;
wire _014_;
wire _015_;
wire _016_;
wire [3:0] _017_;
wire [7:0] _018_;
wire [10:0] _019_;
wire [31:0] _020_;
wire [31:0] _021_;
wire [1:0] _022_;
wire _023_;
wire _024_;
wire _025_;
wire _026_;
wire _027_;
wire _028_;
wire _029_;
wire _030_;
wire _031_;
wire [1:0] _032_;
wire [2:0] _033_;
wire [7:0] _034_;
wire [19:0] _035_;
wire [5:0] _036_;
wire [9:0] _037_;
wire [4:0] _038_;
wire [2:0] _039_;
wire [1:0] _040_;
wire [2:0] _041_;
wire [11:0] _042_;
wire [4:0] _043_;
wire [5:0] _044_;
wire [3:0] _045_;
wire [36:0] _046_;
wire [31:0] _047_;
wire [31:0] _048_;
wire [2:0] _049_;
wire [37:0] _050_;
wire [31:0] _051_;
wire [31:0] _052_;
wire [35:0] _053_;
wire [31:0] _054_;
wire [31:0] _055_;
wire [1:0] _056_;
wire [1:0] _057_;
wire [9:0] _058_;
wire [9:0] _059_;
wire [2:0] _060_;
wire _061_;
wire _062_;
wire [7:0] _063_;
wire [3:0] _064_;
wire [8:0] _065_;
wire [2:0] _066_;
wire [7:0] _067_;
wire [3:0] _068_;
wire [3:0] _069_;
wire _070_;
wire [2:0] _071_;
wire _072_;
wire [2:0] _073_;
wire [2:0] _074_;
wire [2:0] _075_;
wire [3:0] _076_;
wire [1:0] _077_;
wire _078_;
wire _079_;
wire _080_;
wire [1:0] _081_;
wire _082_;
wire _083_;
wire _084_;
wire _085_;
wire _086_;
wire _087_;
wire _088_;
wire _089_;
wire _090_;
wire _091_;
wire _092_;
wire _093_;
wire _094_;
wire _095_;
wire _096_;
wire _097_;
wire [4:0] _098_;
wire [4:0] _099_;
wire _100_;
wire [4:0] _101_;
wire [5:0] _102_;
wire [5:0] _103_;
wire [5:0] _104_;
wire [5:0] _105_;
wire _106_;
wire [4:0] _107_;
wire [5:0] _108_;
wire [6:0] _109_;
wire [5:0] _110_;
wire [5:0] _111_;
wire _112_;
wire [5:0] _113_;
wire [6:0] _114_;
wire [6:0] _115_;
wire _116_;
wire _117_;
wire _118_;
wire _119_;
wire [1:0] _120_;
wire [1:0] _121_;
wire [15:0] _122_;
wire [15:0] _123_;
wire _124_;
wire [15:0] _125_;
wire [16:0] _126_;
wire [16:0] _127_;
wire [15:0] _128_;
wire [15:0] _129_;
wire _130_;
wire [15:0] _131_;
wire [16:0] _132_;
wire [16:0] _133_;
wire [15:0] _134_;
wire [15:0] _135_;
wire _136_;
wire [15:0] _137_;
wire [16:0] _138_;
wire [16:0] _139_;
wire [15:0] _140_;
wire [15:0] _141_;
wire _142_;
wire [15:0] _143_;
wire [16:0] _144_;
wire [16:0] _145_;
wire [15:0] _146_;
wire [15:0] _147_;
wire _148_;
wire [15:0] _149_;
wire [16:0] _150_;
wire [16:0] _151_;
wire [15:0] _152_;
wire [15:0] _153_;
wire _154_;
wire [15:0] _155_;
wire [16:0] _156_;
wire [16:0] _157_;
wire [17:0] _158_;
wire [17:0] _159_;
wire _160_;
wire [17:0] _161_;
wire [18:0] _162_;
wire [18:0] _163_;
wire [18:0] _164_;
wire [18:0] _165_;
wire _166_;
wire [17:0] _167_;
wire [18:0] _168_;
wire [19:0] _169_;
wire [18:0] _170_;
wire [18:0] _171_;
wire _172_;
wire [18:0] _173_;
wire [19:0] _174_;
wire [19:0] _175_;
wire [1:0] _176_;
wire [1:0] _177_;
wire _178_;
wire _179_;
wire [1:0] _180_;
wire [2:0] _181_;
wire [1:0] _182_;
wire [1:0] _183_;
wire _184_;
wire _185_;
wire [1:0] _186_;
wire [2:0] _187_;
wire [1:0] _188_;
wire [1:0] _189_;
wire _190_;
wire [1:0] _191_;
wire [2:0] _192_;
wire [2:0] _193_;
wire [2:0] _194_;
wire [2:0] _195_;
wire _196_;
wire [2:0] _197_;
wire [3:0] _198_;
wire [3:0] _199_;
wire [4:0] _200_;
wire [4:0] _201_;
wire _202_;
wire [3:0] _203_;
wire [4:0] _204_;
wire [5:0] _205_;
wire [3:0] _206_;
wire [1:0] _207_;
wire [5:0] _208_;
wire [5:0] _209_;
wire [5:0] _210_;
wire [5:0] _211_;
wire [5:0] _212_;
wire [1:0] _213_;
wire [1:0] _214_;
wire [1:0] _215_;
wire [1:0] _216_;
wire [1:0] _217_;
wire [1:0] _218_;
wire [19:0] _219_;
wire [19:0] _220_;
wire [19:0] _221_;
wire [19:0] _222_;
wire [19:0] _223_;
wire [19:0] _224_;
wire [1:0] _225_;
wire [19:0] _226_;
wire [1:0] _227_;
wire [19:0] _228_;
wire [1:0] _229_;
wire [19:0] _230_;
wire [1:0] _231_;
wire [19:0] _232_;
wire [1:0] _233_;
wire [19:0] _234_;
wire [1:0] _235_;
wire [19:0] _236_;
wire [19:0] _237_;
wire [2:0] _238_;
wire [2:0] _239_;
wire _240_;
wire [1:0] _241_;
wire [2:0] _242_;
wire [3:0] _243_;
wire [2:0] _244_;
wire [2:0] _245_;
wire _246_;
wire [1:0] _247_;
wire [2:0] _248_;
wire [3:0] _249_;
wire _250_;
wire _251_;
wire _252_;
wire _253_;
wire _254_;
wire _255_;
wire _256_;
wire _257_;
wire _258_;
wire _259_;
wire _260_;
wire _261_;
wire _262_;
wire _263_;
wire _264_;
wire _265_;
wire _266_;
wire _267_;
wire _268_;
wire _269_;
wire _270_;
wire _271_;
wire _272_;
wire _273_;
wire _274_;
wire _275_;
wire _276_;
wire _277_;
wire _278_;
wire _279_;
wire _280_;
wire _281_;
wire _282_;
wire _283_;
wire _284_;
wire _285_;
wire _286_;
wire _287_;
wire _288_;
wire _289_;
wire _290_;
wire _291_;
wire _292_;
wire _293_;
wire _294_;
wire _295_;
wire _296_;
wire _297_;
wire _298_;
wire \add_10ns_10ns_10_2_1_U10.ce ;
wire \add_10ns_10ns_10_2_1_U10.clk ;
wire [9:0] \add_10ns_10ns_10_2_1_U10.din0 ;
wire [9:0] \add_10ns_10ns_10_2_1_U10.din1 ;
wire [9:0] \add_10ns_10ns_10_2_1_U10.dout ;
wire \add_10ns_10ns_10_2_1_U10.reset ;
wire [9:0] \add_10ns_10ns_10_2_1_U10.top_add_10ns_10ns_10_2_1_Adder_7_U.a ;
wire [9:0] \add_10ns_10ns_10_2_1_U10.top_add_10ns_10ns_10_2_1_Adder_7_U.ain_s0 ;
wire [9:0] \add_10ns_10ns_10_2_1_U10.top_add_10ns_10ns_10_2_1_Adder_7_U.b ;
wire [9:0] \add_10ns_10ns_10_2_1_U10.top_add_10ns_10ns_10_2_1_Adder_7_U.bin_s0 ;
wire \add_10ns_10ns_10_2_1_U10.top_add_10ns_10ns_10_2_1_Adder_7_U.ce ;
wire \add_10ns_10ns_10_2_1_U10.top_add_10ns_10ns_10_2_1_Adder_7_U.clk ;
wire \add_10ns_10ns_10_2_1_U10.top_add_10ns_10ns_10_2_1_Adder_7_U.facout_s1 ;
wire \add_10ns_10ns_10_2_1_U10.top_add_10ns_10ns_10_2_1_Adder_7_U.facout_s2 ;
wire [4:0] \add_10ns_10ns_10_2_1_U10.top_add_10ns_10ns_10_2_1_Adder_7_U.fas_s1 ;
wire [4:0] \add_10ns_10ns_10_2_1_U10.top_add_10ns_10ns_10_2_1_Adder_7_U.fas_s2 ;
wire \add_10ns_10ns_10_2_1_U10.top_add_10ns_10ns_10_2_1_Adder_7_U.reset ;
wire [9:0] \add_10ns_10ns_10_2_1_U10.top_add_10ns_10ns_10_2_1_Adder_7_U.s ;
wire [4:0] \add_10ns_10ns_10_2_1_U10.top_add_10ns_10ns_10_2_1_Adder_7_U.u1.a ;
wire [4:0] \add_10ns_10ns_10_2_1_U10.top_add_10ns_10ns_10_2_1_Adder_7_U.u1.b ;
wire \add_10ns_10ns_10_2_1_U10.top_add_10ns_10ns_10_2_1_Adder_7_U.u1.cin ;
wire \add_10ns_10ns_10_2_1_U10.top_add_10ns_10ns_10_2_1_Adder_7_U.u1.cout ;
wire [4:0] \add_10ns_10ns_10_2_1_U10.top_add_10ns_10ns_10_2_1_Adder_7_U.u1.s ;
wire [4:0] \add_10ns_10ns_10_2_1_U10.top_add_10ns_10ns_10_2_1_Adder_7_U.u2.a ;
wire [4:0] \add_10ns_10ns_10_2_1_U10.top_add_10ns_10ns_10_2_1_Adder_7_U.u2.b ;
wire \add_10ns_10ns_10_2_1_U10.top_add_10ns_10ns_10_2_1_Adder_7_U.u2.cin ;
wire \add_10ns_10ns_10_2_1_U10.top_add_10ns_10ns_10_2_1_Adder_7_U.u2.cout ;
wire [4:0] \add_10ns_10ns_10_2_1_U10.top_add_10ns_10ns_10_2_1_Adder_7_U.u2.s ;
wire \add_11s_11s_11_2_1_U12.ce ;
wire \add_11s_11s_11_2_1_U12.clk ;
wire [10:0] \add_11s_11s_11_2_1_U12.din0 ;
wire [10:0] \add_11s_11s_11_2_1_U12.din1 ;
wire [10:0] \add_11s_11s_11_2_1_U12.dout ;
wire \add_11s_11s_11_2_1_U12.reset ;
wire [10:0] \add_11s_11s_11_2_1_U12.top_add_11s_11s_11_2_1_Adder_9_U.a ;
wire [10:0] \add_11s_11s_11_2_1_U12.top_add_11s_11s_11_2_1_Adder_9_U.ain_s0 ;
wire [10:0] \add_11s_11s_11_2_1_U12.top_add_11s_11s_11_2_1_Adder_9_U.b ;
wire [10:0] \add_11s_11s_11_2_1_U12.top_add_11s_11s_11_2_1_Adder_9_U.bin_s0 ;
wire \add_11s_11s_11_2_1_U12.top_add_11s_11s_11_2_1_Adder_9_U.ce ;
wire \add_11s_11s_11_2_1_U12.top_add_11s_11s_11_2_1_Adder_9_U.clk ;
wire \add_11s_11s_11_2_1_U12.top_add_11s_11s_11_2_1_Adder_9_U.facout_s1 ;
wire \add_11s_11s_11_2_1_U12.top_add_11s_11s_11_2_1_Adder_9_U.facout_s2 ;
wire [4:0] \add_11s_11s_11_2_1_U12.top_add_11s_11s_11_2_1_Adder_9_U.fas_s1 ;
wire [5:0] \add_11s_11s_11_2_1_U12.top_add_11s_11s_11_2_1_Adder_9_U.fas_s2 ;
wire \add_11s_11s_11_2_1_U12.top_add_11s_11s_11_2_1_Adder_9_U.reset ;
wire [10:0] \add_11s_11s_11_2_1_U12.top_add_11s_11s_11_2_1_Adder_9_U.s ;
wire [4:0] \add_11s_11s_11_2_1_U12.top_add_11s_11s_11_2_1_Adder_9_U.u1.a ;
wire [4:0] \add_11s_11s_11_2_1_U12.top_add_11s_11s_11_2_1_Adder_9_U.u1.b ;
wire \add_11s_11s_11_2_1_U12.top_add_11s_11s_11_2_1_Adder_9_U.u1.cin ;
wire \add_11s_11s_11_2_1_U12.top_add_11s_11s_11_2_1_Adder_9_U.u1.cout ;
wire [4:0] \add_11s_11s_11_2_1_U12.top_add_11s_11s_11_2_1_Adder_9_U.u1.s ;
wire [5:0] \add_11s_11s_11_2_1_U12.top_add_11s_11s_11_2_1_Adder_9_U.u2.a ;
wire [5:0] \add_11s_11s_11_2_1_U12.top_add_11s_11s_11_2_1_Adder_9_U.u2.b ;
wire \add_11s_11s_11_2_1_U12.top_add_11s_11s_11_2_1_Adder_9_U.u2.cin ;
wire \add_11s_11s_11_2_1_U12.top_add_11s_11s_11_2_1_Adder_9_U.u2.cout ;
wire [5:0] \add_11s_11s_11_2_1_U12.top_add_11s_11s_11_2_1_Adder_9_U.u2.s ;
wire \add_12ns_12s_12_2_1_U8.ce ;
wire \add_12ns_12s_12_2_1_U8.clk ;
wire [11:0] \add_12ns_12s_12_2_1_U8.din0 ;
wire [11:0] \add_12ns_12s_12_2_1_U8.din1 ;
wire [11:0] \add_12ns_12s_12_2_1_U8.dout ;
wire \add_12ns_12s_12_2_1_U8.reset ;
wire [11:0] \add_12ns_12s_12_2_1_U8.top_add_12ns_12s_12_2_1_Adder_5_U.a ;
wire [11:0] \add_12ns_12s_12_2_1_U8.top_add_12ns_12s_12_2_1_Adder_5_U.ain_s0 ;
wire [11:0] \add_12ns_12s_12_2_1_U8.top_add_12ns_12s_12_2_1_Adder_5_U.b ;
wire [11:0] \add_12ns_12s_12_2_1_U8.top_add_12ns_12s_12_2_1_Adder_5_U.bin_s0 ;
wire \add_12ns_12s_12_2_1_U8.top_add_12ns_12s_12_2_1_Adder_5_U.ce ;
wire \add_12ns_12s_12_2_1_U8.top_add_12ns_12s_12_2_1_Adder_5_U.clk ;
wire \add_12ns_12s_12_2_1_U8.top_add_12ns_12s_12_2_1_Adder_5_U.facout_s1 ;
wire \add_12ns_12s_12_2_1_U8.top_add_12ns_12s_12_2_1_Adder_5_U.facout_s2 ;
wire [5:0] \add_12ns_12s_12_2_1_U8.top_add_12ns_12s_12_2_1_Adder_5_U.fas_s1 ;
wire [5:0] \add_12ns_12s_12_2_1_U8.top_add_12ns_12s_12_2_1_Adder_5_U.fas_s2 ;
wire \add_12ns_12s_12_2_1_U8.top_add_12ns_12s_12_2_1_Adder_5_U.reset ;
wire [11:0] \add_12ns_12s_12_2_1_U8.top_add_12ns_12s_12_2_1_Adder_5_U.s ;
wire [5:0] \add_12ns_12s_12_2_1_U8.top_add_12ns_12s_12_2_1_Adder_5_U.u1.a ;
wire [5:0] \add_12ns_12s_12_2_1_U8.top_add_12ns_12s_12_2_1_Adder_5_U.u1.b ;
wire \add_12ns_12s_12_2_1_U8.top_add_12ns_12s_12_2_1_Adder_5_U.u1.cin ;
wire \add_12ns_12s_12_2_1_U8.top_add_12ns_12s_12_2_1_Adder_5_U.u1.cout ;
wire [5:0] \add_12ns_12s_12_2_1_U8.top_add_12ns_12s_12_2_1_Adder_5_U.u1.s ;
wire [5:0] \add_12ns_12s_12_2_1_U8.top_add_12ns_12s_12_2_1_Adder_5_U.u2.a ;
wire [5:0] \add_12ns_12s_12_2_1_U8.top_add_12ns_12s_12_2_1_Adder_5_U.u2.b ;
wire \add_12ns_12s_12_2_1_U8.top_add_12ns_12s_12_2_1_Adder_5_U.u2.cin ;
wire \add_12ns_12s_12_2_1_U8.top_add_12ns_12s_12_2_1_Adder_5_U.u2.cout ;
wire [5:0] \add_12ns_12s_12_2_1_U8.top_add_12ns_12s_12_2_1_Adder_5_U.u2.s ;
wire \add_2ns_2ns_2_2_1_U3.ce ;
wire \add_2ns_2ns_2_2_1_U3.clk ;
wire [1:0] \add_2ns_2ns_2_2_1_U3.din0 ;
wire [1:0] \add_2ns_2ns_2_2_1_U3.din1 ;
wire [1:0] \add_2ns_2ns_2_2_1_U3.dout ;
wire \add_2ns_2ns_2_2_1_U3.reset ;
wire [1:0] \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.a ;
wire [1:0] \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.ain_s0 ;
wire [1:0] \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.b ;
wire [1:0] \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.bin_s0 ;
wire \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.ce ;
wire \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.clk ;
wire \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.facout_s1 ;
wire \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.facout_s2 ;
wire \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.fas_s1 ;
wire \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.fas_s2 ;
wire \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.reset ;
wire [1:0] \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.s ;
wire \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.a ;
wire \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.b ;
wire \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.cin ;
wire \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.cout ;
wire \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.s ;
wire \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.a ;
wire \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.b ;
wire \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.cin ;
wire \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.cout ;
wire \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.s ;
wire \add_32ns_32ns_32_2_1_U14.ce ;
wire \add_32ns_32ns_32_2_1_U14.clk ;
wire [31:0] \add_32ns_32ns_32_2_1_U14.din0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U14.din1 ;
wire [31:0] \add_32ns_32ns_32_2_1_U14.dout ;
wire \add_32ns_32ns_32_2_1_U14.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.a ;
wire [31:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.ain_s0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.b ;
wire [31:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.bin_s0 ;
wire \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.ce ;
wire \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.clk ;
wire \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.facout_s1 ;
wire \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.facout_s2 ;
wire [15:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.fas_s1 ;
wire [15:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.fas_s2 ;
wire \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.b ;
wire \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.cin ;
wire \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.b ;
wire \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.cin ;
wire \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.s ;
wire \add_32ns_32ns_32_2_1_U17.ce ;
wire \add_32ns_32ns_32_2_1_U17.clk ;
wire [31:0] \add_32ns_32ns_32_2_1_U17.din0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U17.din1 ;
wire [31:0] \add_32ns_32ns_32_2_1_U17.dout ;
wire \add_32ns_32ns_32_2_1_U17.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.a ;
wire [31:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.ain_s0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.b ;
wire [31:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.bin_s0 ;
wire \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.ce ;
wire \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.clk ;
wire \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.facout_s1 ;
wire \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.facout_s2 ;
wire [15:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.fas_s1 ;
wire [15:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.fas_s2 ;
wire \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.b ;
wire \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.cin ;
wire \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.b ;
wire \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.cin ;
wire \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.s ;
wire \add_32ns_32ns_32_2_1_U18.ce ;
wire \add_32ns_32ns_32_2_1_U18.clk ;
wire [31:0] \add_32ns_32ns_32_2_1_U18.din0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U18.din1 ;
wire [31:0] \add_32ns_32ns_32_2_1_U18.dout ;
wire \add_32ns_32ns_32_2_1_U18.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_11_U.a ;
wire [31:0] \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_11_U.ain_s0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_11_U.b ;
wire [31:0] \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_11_U.bin_s0 ;
wire \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_11_U.ce ;
wire \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_11_U.clk ;
wire \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_11_U.facout_s1 ;
wire \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_11_U.facout_s2 ;
wire [15:0] \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_11_U.fas_s1 ;
wire [15:0] \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_11_U.fas_s2 ;
wire \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_11_U.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_11_U.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.b ;
wire \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.cin ;
wire \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.b ;
wire \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.cin ;
wire \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.s ;
wire \add_32ns_32ns_32_2_1_U20.ce ;
wire \add_32ns_32ns_32_2_1_U20.clk ;
wire [31:0] \add_32ns_32ns_32_2_1_U20.din0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U20.din1 ;
wire [31:0] \add_32ns_32ns_32_2_1_U20.dout ;
wire \add_32ns_32ns_32_2_1_U20.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.a ;
wire [31:0] \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.ain_s0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.b ;
wire [31:0] \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.bin_s0 ;
wire \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.ce ;
wire \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.clk ;
wire \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.facout_s1 ;
wire \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.facout_s2 ;
wire [15:0] \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.fas_s1 ;
wire [15:0] \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.fas_s2 ;
wire \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.b ;
wire \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.cin ;
wire \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.b ;
wire \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.cin ;
wire \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.s ;
wire \add_32ns_32s_32_2_1_U15.ce ;
wire \add_32ns_32s_32_2_1_U15.clk ;
wire [31:0] \add_32ns_32s_32_2_1_U15.din0 ;
wire [31:0] \add_32ns_32s_32_2_1_U15.din1 ;
wire [31:0] \add_32ns_32s_32_2_1_U15.dout ;
wire \add_32ns_32s_32_2_1_U15.reset ;
wire [31:0] \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_12_U.a ;
wire [31:0] \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_12_U.ain_s0 ;
wire [31:0] \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_12_U.b ;
wire [31:0] \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_12_U.bin_s0 ;
wire \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_12_U.ce ;
wire \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_12_U.clk ;
wire \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_12_U.facout_s1 ;
wire \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_12_U.facout_s2 ;
wire [15:0] \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_12_U.fas_s1 ;
wire [15:0] \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_12_U.fas_s2 ;
wire \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_12_U.reset ;
wire [31:0] \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_12_U.s ;
wire [15:0] \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_12_U.u1.a ;
wire [15:0] \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_12_U.u1.b ;
wire \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_12_U.u1.cin ;
wire \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_12_U.u1.cout ;
wire [15:0] \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_12_U.u1.s ;
wire [15:0] \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_12_U.u2.a ;
wire [15:0] \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_12_U.u2.b ;
wire \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_12_U.u2.cin ;
wire \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_12_U.u2.cout ;
wire [15:0] \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_12_U.u2.s ;
wire \add_32s_32ns_32_2_1_U22.ce ;
wire \add_32s_32ns_32_2_1_U22.clk ;
wire [31:0] \add_32s_32ns_32_2_1_U22.din0 ;
wire [31:0] \add_32s_32ns_32_2_1_U22.din1 ;
wire [31:0] \add_32s_32ns_32_2_1_U22.dout ;
wire \add_32s_32ns_32_2_1_U22.reset ;
wire [31:0] \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_16_U.a ;
wire [31:0] \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_16_U.ain_s0 ;
wire [31:0] \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_16_U.b ;
wire [31:0] \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_16_U.bin_s0 ;
wire \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_16_U.ce ;
wire \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_16_U.clk ;
wire \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_16_U.facout_s1 ;
wire \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_16_U.facout_s2 ;
wire [15:0] \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_16_U.fas_s1 ;
wire [15:0] \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_16_U.fas_s2 ;
wire \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_16_U.reset ;
wire [31:0] \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_16_U.s ;
wire [15:0] \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_16_U.u1.a ;
wire [15:0] \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_16_U.u1.b ;
wire \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_16_U.u1.cin ;
wire \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_16_U.u1.cout ;
wire [15:0] \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_16_U.u1.s ;
wire [15:0] \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_16_U.u2.a ;
wire [15:0] \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_16_U.u2.b ;
wire \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_16_U.u2.cin ;
wire \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_16_U.u2.cout ;
wire [15:0] \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_16_U.u2.s ;
wire \add_36s_36s_36_2_1_U19.ce ;
wire \add_36s_36s_36_2_1_U19.clk ;
wire [35:0] \add_36s_36s_36_2_1_U19.din0 ;
wire [35:0] \add_36s_36s_36_2_1_U19.din1 ;
wire [35:0] \add_36s_36s_36_2_1_U19.dout ;
wire \add_36s_36s_36_2_1_U19.reset ;
wire [35:0] \add_36s_36s_36_2_1_U19.top_add_36s_36s_36_2_1_Adder_14_U.a ;
wire [35:0] \add_36s_36s_36_2_1_U19.top_add_36s_36s_36_2_1_Adder_14_U.ain_s0 ;
wire [35:0] \add_36s_36s_36_2_1_U19.top_add_36s_36s_36_2_1_Adder_14_U.b ;
wire [35:0] \add_36s_36s_36_2_1_U19.top_add_36s_36s_36_2_1_Adder_14_U.bin_s0 ;
wire \add_36s_36s_36_2_1_U19.top_add_36s_36s_36_2_1_Adder_14_U.ce ;
wire \add_36s_36s_36_2_1_U19.top_add_36s_36s_36_2_1_Adder_14_U.clk ;
wire \add_36s_36s_36_2_1_U19.top_add_36s_36s_36_2_1_Adder_14_U.facout_s1 ;
wire \add_36s_36s_36_2_1_U19.top_add_36s_36s_36_2_1_Adder_14_U.facout_s2 ;
wire [17:0] \add_36s_36s_36_2_1_U19.top_add_36s_36s_36_2_1_Adder_14_U.fas_s1 ;
wire [17:0] \add_36s_36s_36_2_1_U19.top_add_36s_36s_36_2_1_Adder_14_U.fas_s2 ;
wire \add_36s_36s_36_2_1_U19.top_add_36s_36s_36_2_1_Adder_14_U.reset ;
wire [35:0] \add_36s_36s_36_2_1_U19.top_add_36s_36s_36_2_1_Adder_14_U.s ;
wire [17:0] \add_36s_36s_36_2_1_U19.top_add_36s_36s_36_2_1_Adder_14_U.u1.a ;
wire [17:0] \add_36s_36s_36_2_1_U19.top_add_36s_36s_36_2_1_Adder_14_U.u1.b ;
wire \add_36s_36s_36_2_1_U19.top_add_36s_36s_36_2_1_Adder_14_U.u1.cin ;
wire \add_36s_36s_36_2_1_U19.top_add_36s_36s_36_2_1_Adder_14_U.u1.cout ;
wire [17:0] \add_36s_36s_36_2_1_U19.top_add_36s_36s_36_2_1_Adder_14_U.u1.s ;
wire [17:0] \add_36s_36s_36_2_1_U19.top_add_36s_36s_36_2_1_Adder_14_U.u2.a ;
wire [17:0] \add_36s_36s_36_2_1_U19.top_add_36s_36s_36_2_1_Adder_14_U.u2.b ;
wire \add_36s_36s_36_2_1_U19.top_add_36s_36s_36_2_1_Adder_14_U.u2.cin ;
wire \add_36s_36s_36_2_1_U19.top_add_36s_36s_36_2_1_Adder_14_U.u2.cout ;
wire [17:0] \add_36s_36s_36_2_1_U19.top_add_36s_36s_36_2_1_Adder_14_U.u2.s ;
wire \add_37s_37s_37_2_1_U13.ce ;
wire \add_37s_37s_37_2_1_U13.clk ;
wire [36:0] \add_37s_37s_37_2_1_U13.din0 ;
wire [36:0] \add_37s_37s_37_2_1_U13.din1 ;
wire [36:0] \add_37s_37s_37_2_1_U13.dout ;
wire \add_37s_37s_37_2_1_U13.reset ;
wire [36:0] \add_37s_37s_37_2_1_U13.top_add_37s_37s_37_2_1_Adder_10_U.a ;
wire [36:0] \add_37s_37s_37_2_1_U13.top_add_37s_37s_37_2_1_Adder_10_U.ain_s0 ;
wire [36:0] \add_37s_37s_37_2_1_U13.top_add_37s_37s_37_2_1_Adder_10_U.b ;
wire [36:0] \add_37s_37s_37_2_1_U13.top_add_37s_37s_37_2_1_Adder_10_U.bin_s0 ;
wire \add_37s_37s_37_2_1_U13.top_add_37s_37s_37_2_1_Adder_10_U.ce ;
wire \add_37s_37s_37_2_1_U13.top_add_37s_37s_37_2_1_Adder_10_U.clk ;
wire \add_37s_37s_37_2_1_U13.top_add_37s_37s_37_2_1_Adder_10_U.facout_s1 ;
wire \add_37s_37s_37_2_1_U13.top_add_37s_37s_37_2_1_Adder_10_U.facout_s2 ;
wire [17:0] \add_37s_37s_37_2_1_U13.top_add_37s_37s_37_2_1_Adder_10_U.fas_s1 ;
wire [18:0] \add_37s_37s_37_2_1_U13.top_add_37s_37s_37_2_1_Adder_10_U.fas_s2 ;
wire \add_37s_37s_37_2_1_U13.top_add_37s_37s_37_2_1_Adder_10_U.reset ;
wire [36:0] \add_37s_37s_37_2_1_U13.top_add_37s_37s_37_2_1_Adder_10_U.s ;
wire [17:0] \add_37s_37s_37_2_1_U13.top_add_37s_37s_37_2_1_Adder_10_U.u1.a ;
wire [17:0] \add_37s_37s_37_2_1_U13.top_add_37s_37s_37_2_1_Adder_10_U.u1.b ;
wire \add_37s_37s_37_2_1_U13.top_add_37s_37s_37_2_1_Adder_10_U.u1.cin ;
wire \add_37s_37s_37_2_1_U13.top_add_37s_37s_37_2_1_Adder_10_U.u1.cout ;
wire [17:0] \add_37s_37s_37_2_1_U13.top_add_37s_37s_37_2_1_Adder_10_U.u1.s ;
wire [18:0] \add_37s_37s_37_2_1_U13.top_add_37s_37s_37_2_1_Adder_10_U.u2.a ;
wire [18:0] \add_37s_37s_37_2_1_U13.top_add_37s_37s_37_2_1_Adder_10_U.u2.b ;
wire \add_37s_37s_37_2_1_U13.top_add_37s_37s_37_2_1_Adder_10_U.u2.cin ;
wire \add_37s_37s_37_2_1_U13.top_add_37s_37s_37_2_1_Adder_10_U.u2.cout ;
wire [18:0] \add_37s_37s_37_2_1_U13.top_add_37s_37s_37_2_1_Adder_10_U.u2.s ;
wire \add_38s_38s_38_2_1_U16.ce ;
wire \add_38s_38s_38_2_1_U16.clk ;
wire [37:0] \add_38s_38s_38_2_1_U16.din0 ;
wire [37:0] \add_38s_38s_38_2_1_U16.din1 ;
wire [37:0] \add_38s_38s_38_2_1_U16.dout ;
wire \add_38s_38s_38_2_1_U16.reset ;
wire [37:0] \add_38s_38s_38_2_1_U16.top_add_38s_38s_38_2_1_Adder_13_U.a ;
wire [37:0] \add_38s_38s_38_2_1_U16.top_add_38s_38s_38_2_1_Adder_13_U.ain_s0 ;
wire [37:0] \add_38s_38s_38_2_1_U16.top_add_38s_38s_38_2_1_Adder_13_U.b ;
wire [37:0] \add_38s_38s_38_2_1_U16.top_add_38s_38s_38_2_1_Adder_13_U.bin_s0 ;
wire \add_38s_38s_38_2_1_U16.top_add_38s_38s_38_2_1_Adder_13_U.ce ;
wire \add_38s_38s_38_2_1_U16.top_add_38s_38s_38_2_1_Adder_13_U.clk ;
wire \add_38s_38s_38_2_1_U16.top_add_38s_38s_38_2_1_Adder_13_U.facout_s1 ;
wire \add_38s_38s_38_2_1_U16.top_add_38s_38s_38_2_1_Adder_13_U.facout_s2 ;
wire [18:0] \add_38s_38s_38_2_1_U16.top_add_38s_38s_38_2_1_Adder_13_U.fas_s1 ;
wire [18:0] \add_38s_38s_38_2_1_U16.top_add_38s_38s_38_2_1_Adder_13_U.fas_s2 ;
wire \add_38s_38s_38_2_1_U16.top_add_38s_38s_38_2_1_Adder_13_U.reset ;
wire [37:0] \add_38s_38s_38_2_1_U16.top_add_38s_38s_38_2_1_Adder_13_U.s ;
wire [18:0] \add_38s_38s_38_2_1_U16.top_add_38s_38s_38_2_1_Adder_13_U.u1.a ;
wire [18:0] \add_38s_38s_38_2_1_U16.top_add_38s_38s_38_2_1_Adder_13_U.u1.b ;
wire \add_38s_38s_38_2_1_U16.top_add_38s_38s_38_2_1_Adder_13_U.u1.cin ;
wire \add_38s_38s_38_2_1_U16.top_add_38s_38s_38_2_1_Adder_13_U.u1.cout ;
wire [18:0] \add_38s_38s_38_2_1_U16.top_add_38s_38s_38_2_1_Adder_13_U.u1.s ;
wire [18:0] \add_38s_38s_38_2_1_U16.top_add_38s_38s_38_2_1_Adder_13_U.u2.a ;
wire [18:0] \add_38s_38s_38_2_1_U16.top_add_38s_38s_38_2_1_Adder_13_U.u2.b ;
wire \add_38s_38s_38_2_1_U16.top_add_38s_38s_38_2_1_Adder_13_U.u2.cin ;
wire \add_38s_38s_38_2_1_U16.top_add_38s_38s_38_2_1_Adder_13_U.u2.cout ;
wire [18:0] \add_38s_38s_38_2_1_U16.top_add_38s_38s_38_2_1_Adder_13_U.u2.s ;
wire \add_3ns_3ns_3_2_1_U5.ce ;
wire \add_3ns_3ns_3_2_1_U5.clk ;
wire [2:0] \add_3ns_3ns_3_2_1_U5.din0 ;
wire [2:0] \add_3ns_3ns_3_2_1_U5.din1 ;
wire [2:0] \add_3ns_3ns_3_2_1_U5.dout ;
wire \add_3ns_3ns_3_2_1_U5.reset ;
wire [2:0] \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_3_U.a ;
wire [2:0] \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_3_U.ain_s0 ;
wire [2:0] \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_3_U.b ;
wire [2:0] \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_3_U.bin_s0 ;
wire \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_3_U.ce ;
wire \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_3_U.clk ;
wire \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_3_U.facout_s1 ;
wire \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_3_U.facout_s2 ;
wire \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_3_U.fas_s1 ;
wire [1:0] \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_3_U.fas_s2 ;
wire \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_3_U.reset ;
wire [2:0] \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_3_U.s ;
wire \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_3_U.u1.a ;
wire \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_3_U.u1.b ;
wire \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_3_U.u1.cin ;
wire \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_3_U.u1.cout ;
wire \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_3_U.u1.s ;
wire [1:0] \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_3_U.u2.a ;
wire [1:0] \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_3_U.u2.b ;
wire \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_3_U.u2.cin ;
wire \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_3_U.u2.cout ;
wire [1:0] \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_3_U.u2.s ;
wire \add_3s_3ns_3_2_1_U7.ce ;
wire \add_3s_3ns_3_2_1_U7.clk ;
wire [2:0] \add_3s_3ns_3_2_1_U7.din0 ;
wire [2:0] \add_3s_3ns_3_2_1_U7.din1 ;
wire [2:0] \add_3s_3ns_3_2_1_U7.dout ;
wire \add_3s_3ns_3_2_1_U7.reset ;
wire [2:0] \add_3s_3ns_3_2_1_U7.top_add_3s_3ns_3_2_1_Adder_4_U.a ;
wire [2:0] \add_3s_3ns_3_2_1_U7.top_add_3s_3ns_3_2_1_Adder_4_U.ain_s0 ;
wire [2:0] \add_3s_3ns_3_2_1_U7.top_add_3s_3ns_3_2_1_Adder_4_U.b ;
wire [2:0] \add_3s_3ns_3_2_1_U7.top_add_3s_3ns_3_2_1_Adder_4_U.bin_s0 ;
wire \add_3s_3ns_3_2_1_U7.top_add_3s_3ns_3_2_1_Adder_4_U.ce ;
wire \add_3s_3ns_3_2_1_U7.top_add_3s_3ns_3_2_1_Adder_4_U.clk ;
wire \add_3s_3ns_3_2_1_U7.top_add_3s_3ns_3_2_1_Adder_4_U.facout_s1 ;
wire \add_3s_3ns_3_2_1_U7.top_add_3s_3ns_3_2_1_Adder_4_U.facout_s2 ;
wire \add_3s_3ns_3_2_1_U7.top_add_3s_3ns_3_2_1_Adder_4_U.fas_s1 ;
wire [1:0] \add_3s_3ns_3_2_1_U7.top_add_3s_3ns_3_2_1_Adder_4_U.fas_s2 ;
wire \add_3s_3ns_3_2_1_U7.top_add_3s_3ns_3_2_1_Adder_4_U.reset ;
wire [2:0] \add_3s_3ns_3_2_1_U7.top_add_3s_3ns_3_2_1_Adder_4_U.s ;
wire \add_3s_3ns_3_2_1_U7.top_add_3s_3ns_3_2_1_Adder_4_U.u1.a ;
wire \add_3s_3ns_3_2_1_U7.top_add_3s_3ns_3_2_1_Adder_4_U.u1.b ;
wire \add_3s_3ns_3_2_1_U7.top_add_3s_3ns_3_2_1_Adder_4_U.u1.cin ;
wire \add_3s_3ns_3_2_1_U7.top_add_3s_3ns_3_2_1_Adder_4_U.u1.cout ;
wire \add_3s_3ns_3_2_1_U7.top_add_3s_3ns_3_2_1_Adder_4_U.u1.s ;
wire [1:0] \add_3s_3ns_3_2_1_U7.top_add_3s_3ns_3_2_1_Adder_4_U.u2.a ;
wire [1:0] \add_3s_3ns_3_2_1_U7.top_add_3s_3ns_3_2_1_Adder_4_U.u2.b ;
wire \add_3s_3ns_3_2_1_U7.top_add_3s_3ns_3_2_1_Adder_4_U.u2.cin ;
wire \add_3s_3ns_3_2_1_U7.top_add_3s_3ns_3_2_1_Adder_4_U.u2.cout ;
wire [1:0] \add_3s_3ns_3_2_1_U7.top_add_3s_3ns_3_2_1_Adder_4_U.u2.s ;
wire \add_4s_4ns_4_2_1_U11.ce ;
wire \add_4s_4ns_4_2_1_U11.clk ;
wire [3:0] \add_4s_4ns_4_2_1_U11.din0 ;
wire [3:0] \add_4s_4ns_4_2_1_U11.din1 ;
wire [3:0] \add_4s_4ns_4_2_1_U11.dout ;
wire \add_4s_4ns_4_2_1_U11.reset ;
wire [3:0] \add_4s_4ns_4_2_1_U11.top_add_4s_4ns_4_2_1_Adder_8_U.a ;
wire [3:0] \add_4s_4ns_4_2_1_U11.top_add_4s_4ns_4_2_1_Adder_8_U.ain_s0 ;
wire [3:0] \add_4s_4ns_4_2_1_U11.top_add_4s_4ns_4_2_1_Adder_8_U.b ;
wire [3:0] \add_4s_4ns_4_2_1_U11.top_add_4s_4ns_4_2_1_Adder_8_U.bin_s0 ;
wire \add_4s_4ns_4_2_1_U11.top_add_4s_4ns_4_2_1_Adder_8_U.ce ;
wire \add_4s_4ns_4_2_1_U11.top_add_4s_4ns_4_2_1_Adder_8_U.clk ;
wire \add_4s_4ns_4_2_1_U11.top_add_4s_4ns_4_2_1_Adder_8_U.facout_s1 ;
wire \add_4s_4ns_4_2_1_U11.top_add_4s_4ns_4_2_1_Adder_8_U.facout_s2 ;
wire [1:0] \add_4s_4ns_4_2_1_U11.top_add_4s_4ns_4_2_1_Adder_8_U.fas_s1 ;
wire [1:0] \add_4s_4ns_4_2_1_U11.top_add_4s_4ns_4_2_1_Adder_8_U.fas_s2 ;
wire \add_4s_4ns_4_2_1_U11.top_add_4s_4ns_4_2_1_Adder_8_U.reset ;
wire [3:0] \add_4s_4ns_4_2_1_U11.top_add_4s_4ns_4_2_1_Adder_8_U.s ;
wire [1:0] \add_4s_4ns_4_2_1_U11.top_add_4s_4ns_4_2_1_Adder_8_U.u1.a ;
wire [1:0] \add_4s_4ns_4_2_1_U11.top_add_4s_4ns_4_2_1_Adder_8_U.u1.b ;
wire \add_4s_4ns_4_2_1_U11.top_add_4s_4ns_4_2_1_Adder_8_U.u1.cin ;
wire \add_4s_4ns_4_2_1_U11.top_add_4s_4ns_4_2_1_Adder_8_U.u1.cout ;
wire [1:0] \add_4s_4ns_4_2_1_U11.top_add_4s_4ns_4_2_1_Adder_8_U.u1.s ;
wire [1:0] \add_4s_4ns_4_2_1_U11.top_add_4s_4ns_4_2_1_Adder_8_U.u2.a ;
wire [1:0] \add_4s_4ns_4_2_1_U11.top_add_4s_4ns_4_2_1_Adder_8_U.u2.b ;
wire \add_4s_4ns_4_2_1_U11.top_add_4s_4ns_4_2_1_Adder_8_U.u2.cin ;
wire \add_4s_4ns_4_2_1_U11.top_add_4s_4ns_4_2_1_Adder_8_U.u2.cout ;
wire [1:0] \add_4s_4ns_4_2_1_U11.top_add_4s_4ns_4_2_1_Adder_8_U.u2.s ;
wire \add_6ns_6s_6_2_1_U9.ce ;
wire \add_6ns_6s_6_2_1_U9.clk ;
wire [5:0] \add_6ns_6s_6_2_1_U9.din0 ;
wire [5:0] \add_6ns_6s_6_2_1_U9.din1 ;
wire [5:0] \add_6ns_6s_6_2_1_U9.dout ;
wire \add_6ns_6s_6_2_1_U9.reset ;
wire [5:0] \add_6ns_6s_6_2_1_U9.top_add_6ns_6s_6_2_1_Adder_6_U.a ;
wire [5:0] \add_6ns_6s_6_2_1_U9.top_add_6ns_6s_6_2_1_Adder_6_U.ain_s0 ;
wire [5:0] \add_6ns_6s_6_2_1_U9.top_add_6ns_6s_6_2_1_Adder_6_U.b ;
wire [5:0] \add_6ns_6s_6_2_1_U9.top_add_6ns_6s_6_2_1_Adder_6_U.bin_s0 ;
wire \add_6ns_6s_6_2_1_U9.top_add_6ns_6s_6_2_1_Adder_6_U.ce ;
wire \add_6ns_6s_6_2_1_U9.top_add_6ns_6s_6_2_1_Adder_6_U.clk ;
wire \add_6ns_6s_6_2_1_U9.top_add_6ns_6s_6_2_1_Adder_6_U.facout_s1 ;
wire \add_6ns_6s_6_2_1_U9.top_add_6ns_6s_6_2_1_Adder_6_U.facout_s2 ;
wire [2:0] \add_6ns_6s_6_2_1_U9.top_add_6ns_6s_6_2_1_Adder_6_U.fas_s1 ;
wire [2:0] \add_6ns_6s_6_2_1_U9.top_add_6ns_6s_6_2_1_Adder_6_U.fas_s2 ;
wire \add_6ns_6s_6_2_1_U9.top_add_6ns_6s_6_2_1_Adder_6_U.reset ;
wire [5:0] \add_6ns_6s_6_2_1_U9.top_add_6ns_6s_6_2_1_Adder_6_U.s ;
wire [2:0] \add_6ns_6s_6_2_1_U9.top_add_6ns_6s_6_2_1_Adder_6_U.u1.a ;
wire [2:0] \add_6ns_6s_6_2_1_U9.top_add_6ns_6s_6_2_1_Adder_6_U.u1.b ;
wire \add_6ns_6s_6_2_1_U9.top_add_6ns_6s_6_2_1_Adder_6_U.u1.cin ;
wire \add_6ns_6s_6_2_1_U9.top_add_6ns_6s_6_2_1_Adder_6_U.u1.cout ;
wire [2:0] \add_6ns_6s_6_2_1_U9.top_add_6ns_6s_6_2_1_Adder_6_U.u1.s ;
wire [2:0] \add_6ns_6s_6_2_1_U9.top_add_6ns_6s_6_2_1_Adder_6_U.u2.a ;
wire [2:0] \add_6ns_6s_6_2_1_U9.top_add_6ns_6s_6_2_1_Adder_6_U.u2.b ;
wire \add_6ns_6s_6_2_1_U9.top_add_6ns_6s_6_2_1_Adder_6_U.u2.cin ;
wire \add_6ns_6s_6_2_1_U9.top_add_6ns_6s_6_2_1_Adder_6_U.u2.cout ;
wire [2:0] \add_6ns_6s_6_2_1_U9.top_add_6ns_6s_6_2_1_Adder_6_U.u2.s ;
wire \add_9ns_9ns_9_2_1_U21.ce ;
wire \add_9ns_9ns_9_2_1_U21.clk ;
wire [8:0] \add_9ns_9ns_9_2_1_U21.din0 ;
wire [8:0] \add_9ns_9ns_9_2_1_U21.din1 ;
wire [8:0] \add_9ns_9ns_9_2_1_U21.dout ;
wire \add_9ns_9ns_9_2_1_U21.reset ;
wire [8:0] \add_9ns_9ns_9_2_1_U21.top_add_9ns_9ns_9_2_1_Adder_15_U.a ;
wire [8:0] \add_9ns_9ns_9_2_1_U21.top_add_9ns_9ns_9_2_1_Adder_15_U.ain_s0 ;
wire [8:0] \add_9ns_9ns_9_2_1_U21.top_add_9ns_9ns_9_2_1_Adder_15_U.b ;
wire [8:0] \add_9ns_9ns_9_2_1_U21.top_add_9ns_9ns_9_2_1_Adder_15_U.bin_s0 ;
wire \add_9ns_9ns_9_2_1_U21.top_add_9ns_9ns_9_2_1_Adder_15_U.ce ;
wire \add_9ns_9ns_9_2_1_U21.top_add_9ns_9ns_9_2_1_Adder_15_U.clk ;
wire \add_9ns_9ns_9_2_1_U21.top_add_9ns_9ns_9_2_1_Adder_15_U.facout_s1 ;
wire \add_9ns_9ns_9_2_1_U21.top_add_9ns_9ns_9_2_1_Adder_15_U.facout_s2 ;
wire [3:0] \add_9ns_9ns_9_2_1_U21.top_add_9ns_9ns_9_2_1_Adder_15_U.fas_s1 ;
wire [4:0] \add_9ns_9ns_9_2_1_U21.top_add_9ns_9ns_9_2_1_Adder_15_U.fas_s2 ;
wire \add_9ns_9ns_9_2_1_U21.top_add_9ns_9ns_9_2_1_Adder_15_U.reset ;
wire [8:0] \add_9ns_9ns_9_2_1_U21.top_add_9ns_9ns_9_2_1_Adder_15_U.s ;
wire [3:0] \add_9ns_9ns_9_2_1_U21.top_add_9ns_9ns_9_2_1_Adder_15_U.u1.a ;
wire [3:0] \add_9ns_9ns_9_2_1_U21.top_add_9ns_9ns_9_2_1_Adder_15_U.u1.b ;
wire \add_9ns_9ns_9_2_1_U21.top_add_9ns_9ns_9_2_1_Adder_15_U.u1.cin ;
wire \add_9ns_9ns_9_2_1_U21.top_add_9ns_9ns_9_2_1_Adder_15_U.u1.cout ;
wire [3:0] \add_9ns_9ns_9_2_1_U21.top_add_9ns_9ns_9_2_1_Adder_15_U.u1.s ;
wire [4:0] \add_9ns_9ns_9_2_1_U21.top_add_9ns_9ns_9_2_1_Adder_15_U.u2.a ;
wire [4:0] \add_9ns_9ns_9_2_1_U21.top_add_9ns_9ns_9_2_1_Adder_15_U.u2.b ;
wire \add_9ns_9ns_9_2_1_U21.top_add_9ns_9ns_9_2_1_Adder_15_U.u2.cin ;
wire \add_9ns_9ns_9_2_1_U21.top_add_9ns_9ns_9_2_1_Adder_15_U.u2.cout ;
wire [4:0] \add_9ns_9ns_9_2_1_U21.top_add_9ns_9ns_9_2_1_Adder_15_U.u2.s ;
wire and_ln340_1_fu_573_p2;
wire and_ln340_2_fu_828_p2;
wire and_ln340_3_fu_840_p2;
wire and_ln340_fu_560_p2;
wire and_ln785_1_fu_577_p2;
wire and_ln785_3_fu_889_p2;
wire and_ln785_4_fu_844_p2;
wire and_ln785_fu_612_p2;
wire and_ln786_1_fu_745_p2;
wire and_ln786_fu_486_p2;
wire ap_CS_fsm_state1;
wire ap_CS_fsm_state10;
wire ap_CS_fsm_state11;
wire ap_CS_fsm_state12;
wire ap_CS_fsm_state13;
wire ap_CS_fsm_state14;
wire ap_CS_fsm_state15;
wire ap_CS_fsm_state16;
wire ap_CS_fsm_state17;
wire ap_CS_fsm_state18;
wire ap_CS_fsm_state19;
wire ap_CS_fsm_state20;
wire ap_CS_fsm_state21;
wire ap_CS_fsm_state22;
wire ap_CS_fsm_state23;
wire ap_CS_fsm_state24;
wire ap_CS_fsm_state25;
wire ap_CS_fsm_state26;
wire ap_CS_fsm_state27;
wire ap_CS_fsm_state28;
wire ap_CS_fsm_state29;
wire ap_CS_fsm_state30;
wire ap_CS_fsm_state31;
wire ap_CS_fsm_state32;
wire ap_CS_fsm_state33;
wire ap_CS_fsm_state34;
wire ap_CS_fsm_state35;
wire ap_CS_fsm_state36;
wire ap_CS_fsm_state37;
wire ap_CS_fsm_state38;
wire ap_CS_fsm_state39;
wire ap_CS_fsm_state40;
wire ap_CS_fsm_state41;
wire ap_CS_fsm_state42;
wire ap_CS_fsm_state43;
wire ap_CS_fsm_state7;
wire ap_CS_fsm_state8;
wire ap_CS_fsm_state9;
wire [42:0] ap_NS_fsm;
wire ap_clk;
wire ap_done;
wire ap_idle;
wire ap_ready;
wire ap_rst;
wire ap_start;
wire [37:0] grp_fu_1004_p0;
wire [37:0] grp_fu_1004_p1;
wire [37:0] grp_fu_1004_p2;
wire [31:0] grp_fu_1030_p2;
wire [31:0] grp_fu_1058_p1;
wire [31:0] grp_fu_1058_p2;
wire [35:0] grp_fu_1078_p0;
wire [35:0] grp_fu_1078_p1;
wire [35:0] grp_fu_1078_p2;
wire [31:0] grp_fu_1104_p2;
wire [8:0] grp_fu_1124_p0;
wire [8:0] grp_fu_1124_p2;
wire [31:0] grp_fu_1151_p0;
wire [31:0] grp_fu_1151_p2;
wire [5:0] grp_fu_237_p2;
wire [4:0] grp_fu_289_p0;
wire [4:0] grp_fu_289_p2;
wire [1:0] grp_fu_300_p2;
wire [4:0] grp_fu_305_p2;
wire [2:0] grp_fu_360_p2;
wire [19:0] grp_fu_437_p0;
wire [19:0] grp_fu_437_p1;
wire [19:0] grp_fu_437_p2;
wire [2:0] grp_fu_597_p0;
wire [2:0] grp_fu_597_p2;
wire [11:0] grp_fu_650_p0;
wire [11:0] grp_fu_650_p1;
wire [11:0] grp_fu_650_p2;
wire [5:0] grp_fu_666_p0;
wire [5:0] grp_fu_666_p1;
wire [5:0] grp_fu_666_p2;
wire [9:0] grp_fu_731_p2;
wire [3:0] grp_fu_752_p0;
wire [3:0] grp_fu_752_p2;
wire [10:0] grp_fu_906_p0;
wire [10:0] grp_fu_906_p1;
wire [10:0] grp_fu_906_p2;
wire [36:0] grp_fu_935_p0;
wire [36:0] grp_fu_935_p1;
wire [36:0] grp_fu_935_p2;
wire [31:0] grp_fu_956_p2;
wire [31:0] grp_fu_984_p1;
wire [31:0] grp_fu_984_p2;
wire icmp_ln768_fu_403_p2;
wire icmp_ln786_fu_408_p2;
wire icmp_ln851_1_fu_295_p2;
wire icmp_ln851_2_fu_247_p2;
wire icmp_ln851_3_fu_672_p2;
wire icmp_ln851_4_fu_941_p2;
wire icmp_ln851_5_fu_1014_p2;
wire icmp_ln851_6_fu_1088_p2;
wire icmp_ln851_fu_355_p2;
wire [1:0] lhs_V_fu_390_p3;
wire [1:0] lhs_fu_275_p1;
wire [2:0] lhs_fu_275_p3;
wire \mul_4s_2s_6_7_1_U1.ce ;
wire \mul_4s_2s_6_7_1_U1.clk ;
wire [3:0] \mul_4s_2s_6_7_1_U1.din0 ;
wire [1:0] \mul_4s_2s_6_7_1_U1.din1 ;
wire [5:0] \mul_4s_2s_6_7_1_U1.dout ;
wire \mul_4s_2s_6_7_1_U1.reset ;
wire [3:0] \mul_4s_2s_6_7_1_U1.top_mul_4s_2s_6_7_1_Mul_DSP_0_U.a ;
wire [1:0] \mul_4s_2s_6_7_1_U1.top_mul_4s_2s_6_7_1_Mul_DSP_0_U.b ;
wire \mul_4s_2s_6_7_1_U1.top_mul_4s_2s_6_7_1_Mul_DSP_0_U.ce ;
wire \mul_4s_2s_6_7_1_U1.top_mul_4s_2s_6_7_1_Mul_DSP_0_U.clk ;
wire [5:0] \mul_4s_2s_6_7_1_U1.top_mul_4s_2s_6_7_1_Mul_DSP_0_U.p ;
wire [5:0] \mul_4s_2s_6_7_1_U1.top_mul_4s_2s_6_7_1_Mul_DSP_0_U.tmp_product ;
wire op_0;
wire op_10;
wire [3:0] op_11_V_fu_623_p3;
wire [7:0] op_13_V_fu_912_p3;
wire [3:0] op_14;
wire [7:0] op_15;
wire [1:0] op_16;
wire [7:0] op_17;
wire op_18;
wire [31:0] op_29;
wire op_29_ap_vld;
wire [1:0] op_4;
wire [3:0] op_5;
wire [1:0] op_6;
wire [16:0] op_7_V_fu_413_p4;
wire [1:0] or_ln1195_fu_398_p1;
wire [1:0] or_ln1195_fu_398_p2;
wire or_ln340_1_fu_767_p2;
wire or_ln340_fu_476_p2;
wire or_ln785_1_fu_736_p2;
wire or_ln785_2_fu_607_p2;
wire or_ln785_3_fu_581_p2;
wire or_ln785_4_fu_884_p2;
wire or_ln785_5_fu_848_p2;
wire or_ln785_fu_425_p2;
wire or_ln786_fu_471_p2;
wire overflow_1_fu_758_p2;
wire overflow_fu_462_p2;
wire [7:0] p_Result_11_fu_814_p4;
wire p_Result_12_fu_860_p3;
wire p_Result_13_fu_961_p3;
wire p_Result_14_fu_1035_p3;
wire p_Result_15_fu_1129_p3;
wire p_Result_18_fu_506_p3;
wire p_Result_1_fu_365_p3;
wire p_Result_3_fu_772_p3;
wire [3:0] p_Result_7_fu_545_p4;
wire p_Result_s_fu_443_p3;
wire [3:0] p_Val2_5_fu_499_p3;
wire [2:0] p_Val2_6_fu_539_p2;
wire [7:0] p_Val2_9_fu_809_p2;
wire [9:0] ret_V_10_fu_784_p3;
wire [2:0] ret_V_21_fu_455_p3;
wire [1:0] ret_V_22_fu_377_p3;
wire [3:0] ret_V_27_fu_872_p3;
wire [31:0] ret_V_29_fu_973_p3;
wire [31:0] ret_V_31_fu_1047_p3;
wire [31:0] ret_V_33_fu_1141_p3;
wire [4:0] rhs_1_fu_635_p3;
wire [36:0] rhs_5_fu_993_p3;
wire [34:0] rhs_7_fu_1067_p3;
wire sel_tmp11_fu_587_p2;
wire sel_tmp24_fu_854_p2;
wire [7:0] select_ln340_1_fu_833_p3;
wire [3:0] select_ln340_fu_565_p3;
wire [8:0] select_ln69_fu_1109_p3;
wire [2:0] select_ln703_fu_491_p3;
wire [7:0] select_ln785_1_fu_894_p3;
wire [3:0] select_ln785_fu_617_p3;
wire [1:0] select_ln850_1_fu_372_p3;
wire [9:0] select_ln850_2_fu_779_p3;
wire [3:0] select_ln850_3_fu_867_p3;
wire [31:0] select_ln850_4_fu_968_p3;
wire [31:0] select_ln850_5_fu_1042_p3;
wire [31:0] select_ln850_6_fu_1136_p3;
wire [2:0] select_ln850_fu_450_p3;
wire [9:0] sext_ln1192_fu_642_p1;
wire [3:0] sext_ln1193_fu_286_p0;
wire [4:0] sext_ln1193_fu_286_p1;
wire [7:0] sext_ln69_2_fu_1117_p1;
wire [3:0] sext_ln703_1_fu_632_p0;
wire [7:0] sext_ln703_3_fu_989_p0;
wire [7:0] sext_ln703_4_fu_1063_p0;
wire [3:0] sext_ln850_fu_749_p1;
wire \shl_20s_2ns_20_7_1_U6.ce ;
wire \shl_20s_2ns_20_7_1_U6.clk ;
wire [19:0] \shl_20s_2ns_20_7_1_U6.din0 ;
wire [19:0] \shl_20s_2ns_20_7_1_U6.din1 ;
wire [1:0] \shl_20s_2ns_20_7_1_U6.din1_cast ;
wire [1:0] \shl_20s_2ns_20_7_1_U6.din1_mask ;
wire [19:0] \shl_20s_2ns_20_7_1_U6.dout ;
wire \shl_20s_2ns_20_7_1_U6.reset ;
wire \sub_5ns_5s_5_2_1_U4.ce ;
wire \sub_5ns_5s_5_2_1_U4.clk ;
wire [4:0] \sub_5ns_5s_5_2_1_U4.din0 ;
wire [4:0] \sub_5ns_5s_5_2_1_U4.din1 ;
wire [4:0] \sub_5ns_5s_5_2_1_U4.dout ;
wire \sub_5ns_5s_5_2_1_U4.reset ;
wire [4:0] \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.a ;
wire [4:0] \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.ain_s0 ;
wire [4:0] \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.b ;
wire [4:0] \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.bin_s0 ;
wire \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.ce ;
wire \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.clk ;
wire \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.facout_s1 ;
wire \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.facout_s2 ;
wire [1:0] \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.fas_s1 ;
wire [2:0] \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.fas_s2 ;
wire \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.reset ;
wire [4:0] \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.s ;
wire [1:0] \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.u1.a ;
wire [1:0] \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.u1.b ;
wire \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.u1.cin ;
wire \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.u1.cout ;
wire [1:0] \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.u1.s ;
wire [2:0] \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.u2.a ;
wire [2:0] \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.u2.b ;
wire \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.u2.cin ;
wire \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.u2.cout ;
wire [2:0] \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.u2.s ;
wire \sub_5s_5s_5_2_1_U2.ce ;
wire \sub_5s_5s_5_2_1_U2.clk ;
wire [4:0] \sub_5s_5s_5_2_1_U2.din0 ;
wire [4:0] \sub_5s_5s_5_2_1_U2.din1 ;
wire [4:0] \sub_5s_5s_5_2_1_U2.dout ;
wire \sub_5s_5s_5_2_1_U2.reset ;
wire [4:0] \sub_5s_5s_5_2_1_U2.top_sub_5s_5s_5_2_1_Adder_0_U.a ;
wire [4:0] \sub_5s_5s_5_2_1_U2.top_sub_5s_5s_5_2_1_Adder_0_U.ain_s0 ;
wire [4:0] \sub_5s_5s_5_2_1_U2.top_sub_5s_5s_5_2_1_Adder_0_U.b ;
wire [4:0] \sub_5s_5s_5_2_1_U2.top_sub_5s_5s_5_2_1_Adder_0_U.bin_s0 ;
wire \sub_5s_5s_5_2_1_U2.top_sub_5s_5s_5_2_1_Adder_0_U.ce ;
wire \sub_5s_5s_5_2_1_U2.top_sub_5s_5s_5_2_1_Adder_0_U.clk ;
wire \sub_5s_5s_5_2_1_U2.top_sub_5s_5s_5_2_1_Adder_0_U.facout_s1 ;
wire \sub_5s_5s_5_2_1_U2.top_sub_5s_5s_5_2_1_Adder_0_U.facout_s2 ;
wire [1:0] \sub_5s_5s_5_2_1_U2.top_sub_5s_5s_5_2_1_Adder_0_U.fas_s1 ;
wire [2:0] \sub_5s_5s_5_2_1_U2.top_sub_5s_5s_5_2_1_Adder_0_U.fas_s2 ;
wire \sub_5s_5s_5_2_1_U2.top_sub_5s_5s_5_2_1_Adder_0_U.reset ;
wire [4:0] \sub_5s_5s_5_2_1_U2.top_sub_5s_5s_5_2_1_Adder_0_U.s ;
wire [1:0] \sub_5s_5s_5_2_1_U2.top_sub_5s_5s_5_2_1_Adder_0_U.u1.a ;
wire [1:0] \sub_5s_5s_5_2_1_U2.top_sub_5s_5s_5_2_1_Adder_0_U.u1.b ;
wire \sub_5s_5s_5_2_1_U2.top_sub_5s_5s_5_2_1_Adder_0_U.u1.cin ;
wire \sub_5s_5s_5_2_1_U2.top_sub_5s_5s_5_2_1_Adder_0_U.u1.cout ;
wire [1:0] \sub_5s_5s_5_2_1_U2.top_sub_5s_5s_5_2_1_Adder_0_U.u1.s ;
wire [2:0] \sub_5s_5s_5_2_1_U2.top_sub_5s_5s_5_2_1_Adder_0_U.u2.a ;
wire [2:0] \sub_5s_5s_5_2_1_U2.top_sub_5s_5s_5_2_1_Adder_0_U.u2.b ;
wire \sub_5s_5s_5_2_1_U2.top_sub_5s_5s_5_2_1_Adder_0_U.u2.cin ;
wire \sub_5s_5s_5_2_1_U2.top_sub_5s_5s_5_2_1_Adder_0_U.u2.cout ;
wire [2:0] \sub_5s_5s_5_2_1_U2.top_sub_5s_5s_5_2_1_Adder_0_U.u2.s ;
wire tmp_13_fu_791_p3;
wire [14:0] tmp_16_fu_924_p3;
wire tmp_7_fu_513_p3;
wire tmp_8_fu_520_p3;
wire [1:0] tmp_fu_253_p1;
wire [2:0] trunc_ln731_fu_333_p1;
wire [2:0] trunc_ln851_1_fu_271_p1;
wire [3:0] trunc_ln851_2_fu_243_p0;
wire [1:0] trunc_ln851_2_fu_243_p1;
wire [2:0] trunc_ln851_3_fu_628_p1;
wire [3:0] trunc_ln851_4_fu_917_p1;
wire [7:0] trunc_ln851_5_fu_1010_p0;
wire [4:0] trunc_ln851_5_fu_1010_p1;
wire [7:0] trunc_ln851_6_fu_1084_p0;
wire [2:0] trunc_ln851_6_fu_1084_p1;
wire [1:0] trunc_ln851_fu_321_p1;
wire xor_ln1499_fu_384_p2;
wire xor_ln340_1_fu_823_p2;
wire xor_ln340_fu_555_p2;
wire xor_ln365_1_fu_533_p2;
wire xor_ln365_2_fu_798_p2;
wire xor_ln365_3_fu_803_p2;
wire xor_ln365_fu_527_p2;
wire xor_ln785_1_fu_740_p2;
wire xor_ln785_2_fu_602_p2;
wire xor_ln785_3_fu_879_p2;
wire xor_ln785_fu_429_p2;
wire xor_ln786_1_fu_481_p2;
wire xor_ln786_2_fu_762_p2;
wire xor_ln786_fu_466_p2;


assign _082_ = icmp_ln851_4_reg_1588 & ap_CS_fsm[25];
assign _083_ = icmp_ln851_5_reg_1635 & ap_CS_fsm[32];
assign _084_ = icmp_ln851_6_reg_1682 & ap_CS_fsm[39];
assign _085_ = icmp_ln851_3_reg_1419 & ap_CS_fsm[18];
assign _086_ = _091_ & ap_CS_fsm[18];
assign _087_ = _092_ & ap_CS_fsm[20];
assign _088_ = ap_CS_fsm[13] & _093_;
assign _089_ = _094_ & ap_CS_fsm[0];
assign _090_ = ap_start & ap_CS_fsm[0];
assign and_ln340_1_fu_573_p2 = or_ln786_reg_1335 & or_ln340_reg_1341;
assign and_ln340_2_fu_828_p2 = xor_ln786_2_reg_1511 & xor_ln340_1_fu_823_p2;
assign and_ln340_3_fu_840_p2 = xor_ln786_2_reg_1511 & or_ln340_1_reg_1517;
assign and_ln340_fu_560_p2 = xor_ln340_fu_555_p2 & or_ln786_reg_1335;
assign and_ln785_1_fu_577_p2 = xor_ln785_reg_1318 & and_ln786_reg_1347;
assign and_ln785_3_fu_889_p2 = or_ln785_4_fu_884_p2 & and_ln786_1_reg_1492;
assign and_ln785_4_fu_844_p2 = xor_ln785_1_reg_1486 & and_ln786_1_reg_1492;
assign and_ln785_fu_612_p2 = or_ln785_2_fu_607_p2 & and_ln786_reg_1347;
assign and_ln786_1_fu_745_p2 = tmp_12_reg_1463 & p_Result_20_reg_1457;
assign and_ln786_fu_486_p2 = xor_ln786_1_fu_481_p2 & p_Result_17_reg_1263;
assign overflow_1_fu_758_p2 = xor_ln785_1_reg_1486 & or_ln785_1_reg_1480;
assign overflow_fu_462_p2 = xor_ln785_reg_1318 & or_ln785_reg_1312;
assign sel_tmp11_fu_587_p2 = xor_ln365_1_fu_533_p2 & or_ln785_3_fu_581_p2;
assign sel_tmp24_fu_854_p2 = xor_ln365_3_fu_803_p2 & or_ln785_5_fu_848_p2;
assign xor_ln786_fu_466_p2 = ~ p_Result_17_reg_1263;
assign xor_ln365_1_fu_533_p2 = ~ xor_ln365_fu_527_p2;
assign xor_ln365_3_fu_803_p2 = ~ xor_ln365_2_fu_798_p2;
assign xor_ln785_1_fu_740_p2 = ~ p_Result_19_reg_1441;
assign xor_ln785_fu_429_p2 = ~ p_Result_16_reg_1251;
assign xor_ln786_2_fu_762_p2 = ~ and_ln786_1_reg_1492;
assign xor_ln340_1_fu_823_p2 = ~ or_ln340_1_reg_1517;
assign xor_ln340_fu_555_p2 = ~ or_ln340_reg_1341;
assign xor_ln785_3_fu_879_p2 = ~ or_ln785_1_reg_1480;
assign xor_ln785_2_fu_602_p2 = ~ or_ln785_reg_1312;
assign xor_ln786_1_fu_481_p2 = ~ icmp_ln786_reg_1296;
assign xor_ln1499_fu_384_p2 = ~ op_0;
assign p_Val2_6_fu_539_p2 = ~ { trunc_ln731_reg_1258[1:0], 1'h0 };
assign p_Val2_9_fu_809_p2[6:0] = ~ p_Val2_8_reg_1449[6:0];
assign _091_ = ~ icmp_ln851_2_reg_1179;
assign _092_ = ~ sel_tmp24_reg_1538;
assign _093_ = ~ sel_tmp11_reg_1369;
assign _094_ = ~ ap_start;
assign _095_ = ! trunc_ln851_1_reg_1201;
assign _096_ = ! op_5[1:0];
assign _097_ = ! trunc_ln851_reg_1234;
always @(posedge \add_10ns_10ns_10_2_1_U10.top_add_10ns_10ns_10_2_1_Adder_7_U.clk )
\add_10ns_10ns_10_2_1_U10.top_add_10ns_10ns_10_2_1_Adder_7_U.bin_s1  <= _099_;
always @(posedge \add_10ns_10ns_10_2_1_U10.top_add_10ns_10ns_10_2_1_Adder_7_U.clk )
\add_10ns_10ns_10_2_1_U10.top_add_10ns_10ns_10_2_1_Adder_7_U.ain_s1  <= _098_;
always @(posedge \add_10ns_10ns_10_2_1_U10.top_add_10ns_10ns_10_2_1_Adder_7_U.clk )
\add_10ns_10ns_10_2_1_U10.top_add_10ns_10ns_10_2_1_Adder_7_U.sum_s1  <= _101_;
always @(posedge \add_10ns_10ns_10_2_1_U10.top_add_10ns_10ns_10_2_1_Adder_7_U.clk )
\add_10ns_10ns_10_2_1_U10.top_add_10ns_10ns_10_2_1_Adder_7_U.carry_s1  <= _100_;
assign _099_ = \add_10ns_10ns_10_2_1_U10.top_add_10ns_10ns_10_2_1_Adder_7_U.ce  ? \add_10ns_10ns_10_2_1_U10.top_add_10ns_10ns_10_2_1_Adder_7_U.b [9:5] : \add_10ns_10ns_10_2_1_U10.top_add_10ns_10ns_10_2_1_Adder_7_U.bin_s1 ;
assign _098_ = \add_10ns_10ns_10_2_1_U10.top_add_10ns_10ns_10_2_1_Adder_7_U.ce  ? \add_10ns_10ns_10_2_1_U10.top_add_10ns_10ns_10_2_1_Adder_7_U.a [9:5] : \add_10ns_10ns_10_2_1_U10.top_add_10ns_10ns_10_2_1_Adder_7_U.ain_s1 ;
assign _100_ = \add_10ns_10ns_10_2_1_U10.top_add_10ns_10ns_10_2_1_Adder_7_U.ce  ? \add_10ns_10ns_10_2_1_U10.top_add_10ns_10ns_10_2_1_Adder_7_U.facout_s1  : \add_10ns_10ns_10_2_1_U10.top_add_10ns_10ns_10_2_1_Adder_7_U.carry_s1 ;
assign _101_ = \add_10ns_10ns_10_2_1_U10.top_add_10ns_10ns_10_2_1_Adder_7_U.ce  ? \add_10ns_10ns_10_2_1_U10.top_add_10ns_10ns_10_2_1_Adder_7_U.fas_s1  : \add_10ns_10ns_10_2_1_U10.top_add_10ns_10ns_10_2_1_Adder_7_U.sum_s1 ;
assign _102_ = \add_10ns_10ns_10_2_1_U10.top_add_10ns_10ns_10_2_1_Adder_7_U.u1.a  + \add_10ns_10ns_10_2_1_U10.top_add_10ns_10ns_10_2_1_Adder_7_U.u1.b ;
assign { \add_10ns_10ns_10_2_1_U10.top_add_10ns_10ns_10_2_1_Adder_7_U.u1.cout , \add_10ns_10ns_10_2_1_U10.top_add_10ns_10ns_10_2_1_Adder_7_U.u1.s  } = _102_ + \add_10ns_10ns_10_2_1_U10.top_add_10ns_10ns_10_2_1_Adder_7_U.u1.cin ;
assign _103_ = \add_10ns_10ns_10_2_1_U10.top_add_10ns_10ns_10_2_1_Adder_7_U.u2.a  + \add_10ns_10ns_10_2_1_U10.top_add_10ns_10ns_10_2_1_Adder_7_U.u2.b ;
assign { \add_10ns_10ns_10_2_1_U10.top_add_10ns_10ns_10_2_1_Adder_7_U.u2.cout , \add_10ns_10ns_10_2_1_U10.top_add_10ns_10ns_10_2_1_Adder_7_U.u2.s  } = _103_ + \add_10ns_10ns_10_2_1_U10.top_add_10ns_10ns_10_2_1_Adder_7_U.u2.cin ;
always @(posedge \add_11s_11s_11_2_1_U12.top_add_11s_11s_11_2_1_Adder_9_U.clk )
\add_11s_11s_11_2_1_U12.top_add_11s_11s_11_2_1_Adder_9_U.bin_s1  <= _105_;
always @(posedge \add_11s_11s_11_2_1_U12.top_add_11s_11s_11_2_1_Adder_9_U.clk )
\add_11s_11s_11_2_1_U12.top_add_11s_11s_11_2_1_Adder_9_U.ain_s1  <= _104_;
always @(posedge \add_11s_11s_11_2_1_U12.top_add_11s_11s_11_2_1_Adder_9_U.clk )
\add_11s_11s_11_2_1_U12.top_add_11s_11s_11_2_1_Adder_9_U.sum_s1  <= _107_;
always @(posedge \add_11s_11s_11_2_1_U12.top_add_11s_11s_11_2_1_Adder_9_U.clk )
\add_11s_11s_11_2_1_U12.top_add_11s_11s_11_2_1_Adder_9_U.carry_s1  <= _106_;
assign _105_ = \add_11s_11s_11_2_1_U12.top_add_11s_11s_11_2_1_Adder_9_U.ce  ? \add_11s_11s_11_2_1_U12.top_add_11s_11s_11_2_1_Adder_9_U.b [10:5] : \add_11s_11s_11_2_1_U12.top_add_11s_11s_11_2_1_Adder_9_U.bin_s1 ;
assign _104_ = \add_11s_11s_11_2_1_U12.top_add_11s_11s_11_2_1_Adder_9_U.ce  ? \add_11s_11s_11_2_1_U12.top_add_11s_11s_11_2_1_Adder_9_U.a [10:5] : \add_11s_11s_11_2_1_U12.top_add_11s_11s_11_2_1_Adder_9_U.ain_s1 ;
assign _106_ = \add_11s_11s_11_2_1_U12.top_add_11s_11s_11_2_1_Adder_9_U.ce  ? \add_11s_11s_11_2_1_U12.top_add_11s_11s_11_2_1_Adder_9_U.facout_s1  : \add_11s_11s_11_2_1_U12.top_add_11s_11s_11_2_1_Adder_9_U.carry_s1 ;
assign _107_ = \add_11s_11s_11_2_1_U12.top_add_11s_11s_11_2_1_Adder_9_U.ce  ? \add_11s_11s_11_2_1_U12.top_add_11s_11s_11_2_1_Adder_9_U.fas_s1  : \add_11s_11s_11_2_1_U12.top_add_11s_11s_11_2_1_Adder_9_U.sum_s1 ;
assign _108_ = \add_11s_11s_11_2_1_U12.top_add_11s_11s_11_2_1_Adder_9_U.u1.a  + \add_11s_11s_11_2_1_U12.top_add_11s_11s_11_2_1_Adder_9_U.u1.b ;
assign { \add_11s_11s_11_2_1_U12.top_add_11s_11s_11_2_1_Adder_9_U.u1.cout , \add_11s_11s_11_2_1_U12.top_add_11s_11s_11_2_1_Adder_9_U.u1.s  } = _108_ + \add_11s_11s_11_2_1_U12.top_add_11s_11s_11_2_1_Adder_9_U.u1.cin ;
assign _109_ = \add_11s_11s_11_2_1_U12.top_add_11s_11s_11_2_1_Adder_9_U.u2.a  + \add_11s_11s_11_2_1_U12.top_add_11s_11s_11_2_1_Adder_9_U.u2.b ;
assign { \add_11s_11s_11_2_1_U12.top_add_11s_11s_11_2_1_Adder_9_U.u2.cout , \add_11s_11s_11_2_1_U12.top_add_11s_11s_11_2_1_Adder_9_U.u2.s  } = _109_ + \add_11s_11s_11_2_1_U12.top_add_11s_11s_11_2_1_Adder_9_U.u2.cin ;
always @(posedge \add_12ns_12s_12_2_1_U8.top_add_12ns_12s_12_2_1_Adder_5_U.clk )
\add_12ns_12s_12_2_1_U8.top_add_12ns_12s_12_2_1_Adder_5_U.bin_s1  <= _111_;
always @(posedge \add_12ns_12s_12_2_1_U8.top_add_12ns_12s_12_2_1_Adder_5_U.clk )
\add_12ns_12s_12_2_1_U8.top_add_12ns_12s_12_2_1_Adder_5_U.ain_s1  <= _110_;
always @(posedge \add_12ns_12s_12_2_1_U8.top_add_12ns_12s_12_2_1_Adder_5_U.clk )
\add_12ns_12s_12_2_1_U8.top_add_12ns_12s_12_2_1_Adder_5_U.sum_s1  <= _113_;
always @(posedge \add_12ns_12s_12_2_1_U8.top_add_12ns_12s_12_2_1_Adder_5_U.clk )
\add_12ns_12s_12_2_1_U8.top_add_12ns_12s_12_2_1_Adder_5_U.carry_s1  <= _112_;
assign _111_ = \add_12ns_12s_12_2_1_U8.top_add_12ns_12s_12_2_1_Adder_5_U.ce  ? \add_12ns_12s_12_2_1_U8.top_add_12ns_12s_12_2_1_Adder_5_U.b [11:6] : \add_12ns_12s_12_2_1_U8.top_add_12ns_12s_12_2_1_Adder_5_U.bin_s1 ;
assign _110_ = \add_12ns_12s_12_2_1_U8.top_add_12ns_12s_12_2_1_Adder_5_U.ce  ? \add_12ns_12s_12_2_1_U8.top_add_12ns_12s_12_2_1_Adder_5_U.a [11:6] : \add_12ns_12s_12_2_1_U8.top_add_12ns_12s_12_2_1_Adder_5_U.ain_s1 ;
assign _112_ = \add_12ns_12s_12_2_1_U8.top_add_12ns_12s_12_2_1_Adder_5_U.ce  ? \add_12ns_12s_12_2_1_U8.top_add_12ns_12s_12_2_1_Adder_5_U.facout_s1  : \add_12ns_12s_12_2_1_U8.top_add_12ns_12s_12_2_1_Adder_5_U.carry_s1 ;
assign _113_ = \add_12ns_12s_12_2_1_U8.top_add_12ns_12s_12_2_1_Adder_5_U.ce  ? \add_12ns_12s_12_2_1_U8.top_add_12ns_12s_12_2_1_Adder_5_U.fas_s1  : \add_12ns_12s_12_2_1_U8.top_add_12ns_12s_12_2_1_Adder_5_U.sum_s1 ;
assign _114_ = \add_12ns_12s_12_2_1_U8.top_add_12ns_12s_12_2_1_Adder_5_U.u1.a  + \add_12ns_12s_12_2_1_U8.top_add_12ns_12s_12_2_1_Adder_5_U.u1.b ;
assign { \add_12ns_12s_12_2_1_U8.top_add_12ns_12s_12_2_1_Adder_5_U.u1.cout , \add_12ns_12s_12_2_1_U8.top_add_12ns_12s_12_2_1_Adder_5_U.u1.s  } = _114_ + \add_12ns_12s_12_2_1_U8.top_add_12ns_12s_12_2_1_Adder_5_U.u1.cin ;
assign _115_ = \add_12ns_12s_12_2_1_U8.top_add_12ns_12s_12_2_1_Adder_5_U.u2.a  + \add_12ns_12s_12_2_1_U8.top_add_12ns_12s_12_2_1_Adder_5_U.u2.b ;
assign { \add_12ns_12s_12_2_1_U8.top_add_12ns_12s_12_2_1_Adder_5_U.u2.cout , \add_12ns_12s_12_2_1_U8.top_add_12ns_12s_12_2_1_Adder_5_U.u2.s  } = _115_ + \add_12ns_12s_12_2_1_U8.top_add_12ns_12s_12_2_1_Adder_5_U.u2.cin ;
always @(posedge \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.clk )
\add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.bin_s1  <= _117_;
always @(posedge \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.clk )
\add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.ain_s1  <= _116_;
always @(posedge \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.clk )
\add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.sum_s1  <= _119_;
always @(posedge \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.clk )
\add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.carry_s1  <= _118_;
assign _117_ = \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.ce  ? \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.b [1] : \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.bin_s1 ;
assign _116_ = \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.ce  ? \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.a [1] : \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.ain_s1 ;
assign _118_ = \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.ce  ? \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.facout_s1  : \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.carry_s1 ;
assign _119_ = \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.ce  ? \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.fas_s1  : \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.sum_s1 ;
assign _120_ = \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.a  + \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.b ;
assign { \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.cout , \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.s  } = _120_ + \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.cin ;
assign _121_ = \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.a  + \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.b ;
assign { \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.cout , \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.s  } = _121_ + \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.cin ;
always @(posedge \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.clk )
\add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.bin_s1  <= _123_;
always @(posedge \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.clk )
\add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.ain_s1  <= _122_;
always @(posedge \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.clk )
\add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.sum_s1  <= _125_;
always @(posedge \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.clk )
\add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.carry_s1  <= _124_;
assign _123_ = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.ce  ? \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.b [31:16] : \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.bin_s1 ;
assign _122_ = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.ce  ? \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.a [31:16] : \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.ain_s1 ;
assign _124_ = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.ce  ? \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.facout_s1  : \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.carry_s1 ;
assign _125_ = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.ce  ? \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.fas_s1  : \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.sum_s1 ;
assign _126_ = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.a  + \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.b ;
assign { \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.cout , \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.s  } = _126_ + \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.cin ;
assign _127_ = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.a  + \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.b ;
assign { \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.cout , \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.s  } = _127_ + \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.cin ;
always @(posedge \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.clk )
\add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.bin_s1  <= _129_;
always @(posedge \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.clk )
\add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.ain_s1  <= _128_;
always @(posedge \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.clk )
\add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.sum_s1  <= _131_;
always @(posedge \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.clk )
\add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.carry_s1  <= _130_;
assign _129_ = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.ce  ? \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.b [31:16] : \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.bin_s1 ;
assign _128_ = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.ce  ? \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.a [31:16] : \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.ain_s1 ;
assign _130_ = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.ce  ? \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.facout_s1  : \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.carry_s1 ;
assign _131_ = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.ce  ? \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.fas_s1  : \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.sum_s1 ;
assign _132_ = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.a  + \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.b ;
assign { \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.cout , \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.s  } = _132_ + \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.cin ;
assign _133_ = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.a  + \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.b ;
assign { \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.cout , \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.s  } = _133_ + \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.cin ;
always @(posedge \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_11_U.clk )
\add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_11_U.bin_s1  <= _135_;
always @(posedge \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_11_U.clk )
\add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_11_U.ain_s1  <= _134_;
always @(posedge \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_11_U.clk )
\add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_11_U.sum_s1  <= _137_;
always @(posedge \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_11_U.clk )
\add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_11_U.carry_s1  <= _136_;
assign _135_ = \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_11_U.ce  ? \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_11_U.b [31:16] : \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_11_U.bin_s1 ;
assign _134_ = \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_11_U.ce  ? \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_11_U.a [31:16] : \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_11_U.ain_s1 ;
assign _136_ = \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_11_U.ce  ? \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_11_U.facout_s1  : \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_11_U.carry_s1 ;
assign _137_ = \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_11_U.ce  ? \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_11_U.fas_s1  : \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_11_U.sum_s1 ;
assign _138_ = \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.a  + \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.b ;
assign { \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.cout , \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.s  } = _138_ + \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.cin ;
assign _139_ = \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.a  + \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.b ;
assign { \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.cout , \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.s  } = _139_ + \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.cin ;
always @(posedge \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.clk )
\add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.bin_s1  <= _141_;
always @(posedge \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.clk )
\add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.ain_s1  <= _140_;
always @(posedge \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.clk )
\add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.sum_s1  <= _143_;
always @(posedge \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.clk )
\add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.carry_s1  <= _142_;
assign _141_ = \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.ce  ? \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.b [31:16] : \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.bin_s1 ;
assign _140_ = \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.ce  ? \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.a [31:16] : \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.ain_s1 ;
assign _142_ = \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.ce  ? \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.facout_s1  : \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.carry_s1 ;
assign _143_ = \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.ce  ? \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.fas_s1  : \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.sum_s1 ;
assign _144_ = \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.a  + \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.b ;
assign { \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.cout , \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.s  } = _144_ + \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.cin ;
assign _145_ = \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.a  + \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.b ;
assign { \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.cout , \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.s  } = _145_ + \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.cin ;
always @(posedge \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_12_U.clk )
\add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_12_U.bin_s1  <= _147_;
always @(posedge \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_12_U.clk )
\add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_12_U.ain_s1  <= _146_;
always @(posedge \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_12_U.clk )
\add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_12_U.sum_s1  <= _149_;
always @(posedge \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_12_U.clk )
\add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_12_U.carry_s1  <= _148_;
assign _147_ = \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_12_U.ce  ? \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_12_U.b [31:16] : \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_12_U.bin_s1 ;
assign _146_ = \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_12_U.ce  ? \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_12_U.a [31:16] : \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_12_U.ain_s1 ;
assign _148_ = \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_12_U.ce  ? \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_12_U.facout_s1  : \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_12_U.carry_s1 ;
assign _149_ = \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_12_U.ce  ? \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_12_U.fas_s1  : \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_12_U.sum_s1 ;
assign _150_ = \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_12_U.u1.a  + \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_12_U.u1.b ;
assign { \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_12_U.u1.cout , \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_12_U.u1.s  } = _150_ + \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_12_U.u1.cin ;
assign _151_ = \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_12_U.u2.a  + \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_12_U.u2.b ;
assign { \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_12_U.u2.cout , \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_12_U.u2.s  } = _151_ + \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_12_U.u2.cin ;
always @(posedge \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_16_U.clk )
\add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_16_U.bin_s1  <= _153_;
always @(posedge \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_16_U.clk )
\add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_16_U.ain_s1  <= _152_;
always @(posedge \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_16_U.clk )
\add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_16_U.sum_s1  <= _155_;
always @(posedge \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_16_U.clk )
\add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_16_U.carry_s1  <= _154_;
assign _153_ = \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_16_U.ce  ? \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_16_U.b [31:16] : \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_16_U.bin_s1 ;
assign _152_ = \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_16_U.ce  ? \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_16_U.a [31:16] : \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_16_U.ain_s1 ;
assign _154_ = \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_16_U.ce  ? \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_16_U.facout_s1  : \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_16_U.carry_s1 ;
assign _155_ = \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_16_U.ce  ? \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_16_U.fas_s1  : \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_16_U.sum_s1 ;
assign _156_ = \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_16_U.u1.a  + \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_16_U.u1.b ;
assign { \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_16_U.u1.cout , \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_16_U.u1.s  } = _156_ + \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_16_U.u1.cin ;
assign _157_ = \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_16_U.u2.a  + \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_16_U.u2.b ;
assign { \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_16_U.u2.cout , \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_16_U.u2.s  } = _157_ + \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_16_U.u2.cin ;
always @(posedge \add_36s_36s_36_2_1_U19.top_add_36s_36s_36_2_1_Adder_14_U.clk )
\add_36s_36s_36_2_1_U19.top_add_36s_36s_36_2_1_Adder_14_U.bin_s1  <= _159_;
always @(posedge \add_36s_36s_36_2_1_U19.top_add_36s_36s_36_2_1_Adder_14_U.clk )
\add_36s_36s_36_2_1_U19.top_add_36s_36s_36_2_1_Adder_14_U.ain_s1  <= _158_;
always @(posedge \add_36s_36s_36_2_1_U19.top_add_36s_36s_36_2_1_Adder_14_U.clk )
\add_36s_36s_36_2_1_U19.top_add_36s_36s_36_2_1_Adder_14_U.sum_s1  <= _161_;
always @(posedge \add_36s_36s_36_2_1_U19.top_add_36s_36s_36_2_1_Adder_14_U.clk )
\add_36s_36s_36_2_1_U19.top_add_36s_36s_36_2_1_Adder_14_U.carry_s1  <= _160_;
assign _159_ = \add_36s_36s_36_2_1_U19.top_add_36s_36s_36_2_1_Adder_14_U.ce  ? \add_36s_36s_36_2_1_U19.top_add_36s_36s_36_2_1_Adder_14_U.b [35:18] : \add_36s_36s_36_2_1_U19.top_add_36s_36s_36_2_1_Adder_14_U.bin_s1 ;
assign _158_ = \add_36s_36s_36_2_1_U19.top_add_36s_36s_36_2_1_Adder_14_U.ce  ? \add_36s_36s_36_2_1_U19.top_add_36s_36s_36_2_1_Adder_14_U.a [35:18] : \add_36s_36s_36_2_1_U19.top_add_36s_36s_36_2_1_Adder_14_U.ain_s1 ;
assign _160_ = \add_36s_36s_36_2_1_U19.top_add_36s_36s_36_2_1_Adder_14_U.ce  ? \add_36s_36s_36_2_1_U19.top_add_36s_36s_36_2_1_Adder_14_U.facout_s1  : \add_36s_36s_36_2_1_U19.top_add_36s_36s_36_2_1_Adder_14_U.carry_s1 ;
assign _161_ = \add_36s_36s_36_2_1_U19.top_add_36s_36s_36_2_1_Adder_14_U.ce  ? \add_36s_36s_36_2_1_U19.top_add_36s_36s_36_2_1_Adder_14_U.fas_s1  : \add_36s_36s_36_2_1_U19.top_add_36s_36s_36_2_1_Adder_14_U.sum_s1 ;
assign _162_ = \add_36s_36s_36_2_1_U19.top_add_36s_36s_36_2_1_Adder_14_U.u1.a  + \add_36s_36s_36_2_1_U19.top_add_36s_36s_36_2_1_Adder_14_U.u1.b ;
assign { \add_36s_36s_36_2_1_U19.top_add_36s_36s_36_2_1_Adder_14_U.u1.cout , \add_36s_36s_36_2_1_U19.top_add_36s_36s_36_2_1_Adder_14_U.u1.s  } = _162_ + \add_36s_36s_36_2_1_U19.top_add_36s_36s_36_2_1_Adder_14_U.u1.cin ;
assign _163_ = \add_36s_36s_36_2_1_U19.top_add_36s_36s_36_2_1_Adder_14_U.u2.a  + \add_36s_36s_36_2_1_U19.top_add_36s_36s_36_2_1_Adder_14_U.u2.b ;
assign { \add_36s_36s_36_2_1_U19.top_add_36s_36s_36_2_1_Adder_14_U.u2.cout , \add_36s_36s_36_2_1_U19.top_add_36s_36s_36_2_1_Adder_14_U.u2.s  } = _163_ + \add_36s_36s_36_2_1_U19.top_add_36s_36s_36_2_1_Adder_14_U.u2.cin ;
always @(posedge \add_37s_37s_37_2_1_U13.top_add_37s_37s_37_2_1_Adder_10_U.clk )
\add_37s_37s_37_2_1_U13.top_add_37s_37s_37_2_1_Adder_10_U.bin_s1  <= _165_;
always @(posedge \add_37s_37s_37_2_1_U13.top_add_37s_37s_37_2_1_Adder_10_U.clk )
\add_37s_37s_37_2_1_U13.top_add_37s_37s_37_2_1_Adder_10_U.ain_s1  <= _164_;
always @(posedge \add_37s_37s_37_2_1_U13.top_add_37s_37s_37_2_1_Adder_10_U.clk )
\add_37s_37s_37_2_1_U13.top_add_37s_37s_37_2_1_Adder_10_U.sum_s1  <= _167_;
always @(posedge \add_37s_37s_37_2_1_U13.top_add_37s_37s_37_2_1_Adder_10_U.clk )
\add_37s_37s_37_2_1_U13.top_add_37s_37s_37_2_1_Adder_10_U.carry_s1  <= _166_;
assign _165_ = \add_37s_37s_37_2_1_U13.top_add_37s_37s_37_2_1_Adder_10_U.ce  ? \add_37s_37s_37_2_1_U13.top_add_37s_37s_37_2_1_Adder_10_U.b [36:18] : \add_37s_37s_37_2_1_U13.top_add_37s_37s_37_2_1_Adder_10_U.bin_s1 ;
assign _164_ = \add_37s_37s_37_2_1_U13.top_add_37s_37s_37_2_1_Adder_10_U.ce  ? \add_37s_37s_37_2_1_U13.top_add_37s_37s_37_2_1_Adder_10_U.a [36:18] : \add_37s_37s_37_2_1_U13.top_add_37s_37s_37_2_1_Adder_10_U.ain_s1 ;
assign _166_ = \add_37s_37s_37_2_1_U13.top_add_37s_37s_37_2_1_Adder_10_U.ce  ? \add_37s_37s_37_2_1_U13.top_add_37s_37s_37_2_1_Adder_10_U.facout_s1  : \add_37s_37s_37_2_1_U13.top_add_37s_37s_37_2_1_Adder_10_U.carry_s1 ;
assign _167_ = \add_37s_37s_37_2_1_U13.top_add_37s_37s_37_2_1_Adder_10_U.ce  ? \add_37s_37s_37_2_1_U13.top_add_37s_37s_37_2_1_Adder_10_U.fas_s1  : \add_37s_37s_37_2_1_U13.top_add_37s_37s_37_2_1_Adder_10_U.sum_s1 ;
assign _168_ = \add_37s_37s_37_2_1_U13.top_add_37s_37s_37_2_1_Adder_10_U.u1.a  + \add_37s_37s_37_2_1_U13.top_add_37s_37s_37_2_1_Adder_10_U.u1.b ;
assign { \add_37s_37s_37_2_1_U13.top_add_37s_37s_37_2_1_Adder_10_U.u1.cout , \add_37s_37s_37_2_1_U13.top_add_37s_37s_37_2_1_Adder_10_U.u1.s  } = _168_ + \add_37s_37s_37_2_1_U13.top_add_37s_37s_37_2_1_Adder_10_U.u1.cin ;
assign _169_ = \add_37s_37s_37_2_1_U13.top_add_37s_37s_37_2_1_Adder_10_U.u2.a  + \add_37s_37s_37_2_1_U13.top_add_37s_37s_37_2_1_Adder_10_U.u2.b ;
assign { \add_37s_37s_37_2_1_U13.top_add_37s_37s_37_2_1_Adder_10_U.u2.cout , \add_37s_37s_37_2_1_U13.top_add_37s_37s_37_2_1_Adder_10_U.u2.s  } = _169_ + \add_37s_37s_37_2_1_U13.top_add_37s_37s_37_2_1_Adder_10_U.u2.cin ;
always @(posedge \add_38s_38s_38_2_1_U16.top_add_38s_38s_38_2_1_Adder_13_U.clk )
\add_38s_38s_38_2_1_U16.top_add_38s_38s_38_2_1_Adder_13_U.bin_s1  <= _171_;
always @(posedge \add_38s_38s_38_2_1_U16.top_add_38s_38s_38_2_1_Adder_13_U.clk )
\add_38s_38s_38_2_1_U16.top_add_38s_38s_38_2_1_Adder_13_U.ain_s1  <= _170_;
always @(posedge \add_38s_38s_38_2_1_U16.top_add_38s_38s_38_2_1_Adder_13_U.clk )
\add_38s_38s_38_2_1_U16.top_add_38s_38s_38_2_1_Adder_13_U.sum_s1  <= _173_;
always @(posedge \add_38s_38s_38_2_1_U16.top_add_38s_38s_38_2_1_Adder_13_U.clk )
\add_38s_38s_38_2_1_U16.top_add_38s_38s_38_2_1_Adder_13_U.carry_s1  <= _172_;
assign _171_ = \add_38s_38s_38_2_1_U16.top_add_38s_38s_38_2_1_Adder_13_U.ce  ? \add_38s_38s_38_2_1_U16.top_add_38s_38s_38_2_1_Adder_13_U.b [37:19] : \add_38s_38s_38_2_1_U16.top_add_38s_38s_38_2_1_Adder_13_U.bin_s1 ;
assign _170_ = \add_38s_38s_38_2_1_U16.top_add_38s_38s_38_2_1_Adder_13_U.ce  ? \add_38s_38s_38_2_1_U16.top_add_38s_38s_38_2_1_Adder_13_U.a [37:19] : \add_38s_38s_38_2_1_U16.top_add_38s_38s_38_2_1_Adder_13_U.ain_s1 ;
assign _172_ = \add_38s_38s_38_2_1_U16.top_add_38s_38s_38_2_1_Adder_13_U.ce  ? \add_38s_38s_38_2_1_U16.top_add_38s_38s_38_2_1_Adder_13_U.facout_s1  : \add_38s_38s_38_2_1_U16.top_add_38s_38s_38_2_1_Adder_13_U.carry_s1 ;
assign _173_ = \add_38s_38s_38_2_1_U16.top_add_38s_38s_38_2_1_Adder_13_U.ce  ? \add_38s_38s_38_2_1_U16.top_add_38s_38s_38_2_1_Adder_13_U.fas_s1  : \add_38s_38s_38_2_1_U16.top_add_38s_38s_38_2_1_Adder_13_U.sum_s1 ;
assign _174_ = \add_38s_38s_38_2_1_U16.top_add_38s_38s_38_2_1_Adder_13_U.u1.a  + \add_38s_38s_38_2_1_U16.top_add_38s_38s_38_2_1_Adder_13_U.u1.b ;
assign { \add_38s_38s_38_2_1_U16.top_add_38s_38s_38_2_1_Adder_13_U.u1.cout , \add_38s_38s_38_2_1_U16.top_add_38s_38s_38_2_1_Adder_13_U.u1.s  } = _174_ + \add_38s_38s_38_2_1_U16.top_add_38s_38s_38_2_1_Adder_13_U.u1.cin ;
assign _175_ = \add_38s_38s_38_2_1_U16.top_add_38s_38s_38_2_1_Adder_13_U.u2.a  + \add_38s_38s_38_2_1_U16.top_add_38s_38s_38_2_1_Adder_13_U.u2.b ;
assign { \add_38s_38s_38_2_1_U16.top_add_38s_38s_38_2_1_Adder_13_U.u2.cout , \add_38s_38s_38_2_1_U16.top_add_38s_38s_38_2_1_Adder_13_U.u2.s  } = _175_ + \add_38s_38s_38_2_1_U16.top_add_38s_38s_38_2_1_Adder_13_U.u2.cin ;
always @(posedge \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_3_U.clk )
\add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_3_U.bin_s1  <= _177_;
always @(posedge \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_3_U.clk )
\add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_3_U.ain_s1  <= _176_;
always @(posedge \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_3_U.clk )
\add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_3_U.sum_s1  <= _179_;
always @(posedge \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_3_U.clk )
\add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_3_U.carry_s1  <= _178_;
assign _177_ = \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_3_U.ce  ? \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_3_U.b [2:1] : \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_3_U.bin_s1 ;
assign _176_ = \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_3_U.ce  ? \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_3_U.a [2:1] : \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_3_U.ain_s1 ;
assign _178_ = \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_3_U.ce  ? \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_3_U.facout_s1  : \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_3_U.carry_s1 ;
assign _179_ = \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_3_U.ce  ? \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_3_U.fas_s1  : \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_3_U.sum_s1 ;
assign _180_ = \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_3_U.u1.a  + \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_3_U.u1.b ;
assign { \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_3_U.u1.cout , \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_3_U.u1.s  } = _180_ + \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_3_U.u1.cin ;
assign _181_ = \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_3_U.u2.a  + \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_3_U.u2.b ;
assign { \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_3_U.u2.cout , \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_3_U.u2.s  } = _181_ + \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_3_U.u2.cin ;
always @(posedge \add_3s_3ns_3_2_1_U7.top_add_3s_3ns_3_2_1_Adder_4_U.clk )
\add_3s_3ns_3_2_1_U7.top_add_3s_3ns_3_2_1_Adder_4_U.bin_s1  <= _183_;
always @(posedge \add_3s_3ns_3_2_1_U7.top_add_3s_3ns_3_2_1_Adder_4_U.clk )
\add_3s_3ns_3_2_1_U7.top_add_3s_3ns_3_2_1_Adder_4_U.ain_s1  <= _182_;
always @(posedge \add_3s_3ns_3_2_1_U7.top_add_3s_3ns_3_2_1_Adder_4_U.clk )
\add_3s_3ns_3_2_1_U7.top_add_3s_3ns_3_2_1_Adder_4_U.sum_s1  <= _185_;
always @(posedge \add_3s_3ns_3_2_1_U7.top_add_3s_3ns_3_2_1_Adder_4_U.clk )
\add_3s_3ns_3_2_1_U7.top_add_3s_3ns_3_2_1_Adder_4_U.carry_s1  <= _184_;
assign _183_ = \add_3s_3ns_3_2_1_U7.top_add_3s_3ns_3_2_1_Adder_4_U.ce  ? \add_3s_3ns_3_2_1_U7.top_add_3s_3ns_3_2_1_Adder_4_U.b [2:1] : \add_3s_3ns_3_2_1_U7.top_add_3s_3ns_3_2_1_Adder_4_U.bin_s1 ;
assign _182_ = \add_3s_3ns_3_2_1_U7.top_add_3s_3ns_3_2_1_Adder_4_U.ce  ? \add_3s_3ns_3_2_1_U7.top_add_3s_3ns_3_2_1_Adder_4_U.a [2:1] : \add_3s_3ns_3_2_1_U7.top_add_3s_3ns_3_2_1_Adder_4_U.ain_s1 ;
assign _184_ = \add_3s_3ns_3_2_1_U7.top_add_3s_3ns_3_2_1_Adder_4_U.ce  ? \add_3s_3ns_3_2_1_U7.top_add_3s_3ns_3_2_1_Adder_4_U.facout_s1  : \add_3s_3ns_3_2_1_U7.top_add_3s_3ns_3_2_1_Adder_4_U.carry_s1 ;
assign _185_ = \add_3s_3ns_3_2_1_U7.top_add_3s_3ns_3_2_1_Adder_4_U.ce  ? \add_3s_3ns_3_2_1_U7.top_add_3s_3ns_3_2_1_Adder_4_U.fas_s1  : \add_3s_3ns_3_2_1_U7.top_add_3s_3ns_3_2_1_Adder_4_U.sum_s1 ;
assign _186_ = \add_3s_3ns_3_2_1_U7.top_add_3s_3ns_3_2_1_Adder_4_U.u1.a  + \add_3s_3ns_3_2_1_U7.top_add_3s_3ns_3_2_1_Adder_4_U.u1.b ;
assign { \add_3s_3ns_3_2_1_U7.top_add_3s_3ns_3_2_1_Adder_4_U.u1.cout , \add_3s_3ns_3_2_1_U7.top_add_3s_3ns_3_2_1_Adder_4_U.u1.s  } = _186_ + \add_3s_3ns_3_2_1_U7.top_add_3s_3ns_3_2_1_Adder_4_U.u1.cin ;
assign _187_ = \add_3s_3ns_3_2_1_U7.top_add_3s_3ns_3_2_1_Adder_4_U.u2.a  + \add_3s_3ns_3_2_1_U7.top_add_3s_3ns_3_2_1_Adder_4_U.u2.b ;
assign { \add_3s_3ns_3_2_1_U7.top_add_3s_3ns_3_2_1_Adder_4_U.u2.cout , \add_3s_3ns_3_2_1_U7.top_add_3s_3ns_3_2_1_Adder_4_U.u2.s  } = _187_ + \add_3s_3ns_3_2_1_U7.top_add_3s_3ns_3_2_1_Adder_4_U.u2.cin ;
always @(posedge \add_4s_4ns_4_2_1_U11.top_add_4s_4ns_4_2_1_Adder_8_U.clk )
\add_4s_4ns_4_2_1_U11.top_add_4s_4ns_4_2_1_Adder_8_U.bin_s1  <= _189_;
always @(posedge \add_4s_4ns_4_2_1_U11.top_add_4s_4ns_4_2_1_Adder_8_U.clk )
\add_4s_4ns_4_2_1_U11.top_add_4s_4ns_4_2_1_Adder_8_U.ain_s1  <= _188_;
always @(posedge \add_4s_4ns_4_2_1_U11.top_add_4s_4ns_4_2_1_Adder_8_U.clk )
\add_4s_4ns_4_2_1_U11.top_add_4s_4ns_4_2_1_Adder_8_U.sum_s1  <= _191_;
always @(posedge \add_4s_4ns_4_2_1_U11.top_add_4s_4ns_4_2_1_Adder_8_U.clk )
\add_4s_4ns_4_2_1_U11.top_add_4s_4ns_4_2_1_Adder_8_U.carry_s1  <= _190_;
assign _189_ = \add_4s_4ns_4_2_1_U11.top_add_4s_4ns_4_2_1_Adder_8_U.ce  ? \add_4s_4ns_4_2_1_U11.top_add_4s_4ns_4_2_1_Adder_8_U.b [3:2] : \add_4s_4ns_4_2_1_U11.top_add_4s_4ns_4_2_1_Adder_8_U.bin_s1 ;
assign _188_ = \add_4s_4ns_4_2_1_U11.top_add_4s_4ns_4_2_1_Adder_8_U.ce  ? \add_4s_4ns_4_2_1_U11.top_add_4s_4ns_4_2_1_Adder_8_U.a [3:2] : \add_4s_4ns_4_2_1_U11.top_add_4s_4ns_4_2_1_Adder_8_U.ain_s1 ;
assign _190_ = \add_4s_4ns_4_2_1_U11.top_add_4s_4ns_4_2_1_Adder_8_U.ce  ? \add_4s_4ns_4_2_1_U11.top_add_4s_4ns_4_2_1_Adder_8_U.facout_s1  : \add_4s_4ns_4_2_1_U11.top_add_4s_4ns_4_2_1_Adder_8_U.carry_s1 ;
assign _191_ = \add_4s_4ns_4_2_1_U11.top_add_4s_4ns_4_2_1_Adder_8_U.ce  ? \add_4s_4ns_4_2_1_U11.top_add_4s_4ns_4_2_1_Adder_8_U.fas_s1  : \add_4s_4ns_4_2_1_U11.top_add_4s_4ns_4_2_1_Adder_8_U.sum_s1 ;
assign _192_ = \add_4s_4ns_4_2_1_U11.top_add_4s_4ns_4_2_1_Adder_8_U.u1.a  + \add_4s_4ns_4_2_1_U11.top_add_4s_4ns_4_2_1_Adder_8_U.u1.b ;
assign { \add_4s_4ns_4_2_1_U11.top_add_4s_4ns_4_2_1_Adder_8_U.u1.cout , \add_4s_4ns_4_2_1_U11.top_add_4s_4ns_4_2_1_Adder_8_U.u1.s  } = _192_ + \add_4s_4ns_4_2_1_U11.top_add_4s_4ns_4_2_1_Adder_8_U.u1.cin ;
assign _193_ = \add_4s_4ns_4_2_1_U11.top_add_4s_4ns_4_2_1_Adder_8_U.u2.a  + \add_4s_4ns_4_2_1_U11.top_add_4s_4ns_4_2_1_Adder_8_U.u2.b ;
assign { \add_4s_4ns_4_2_1_U11.top_add_4s_4ns_4_2_1_Adder_8_U.u2.cout , \add_4s_4ns_4_2_1_U11.top_add_4s_4ns_4_2_1_Adder_8_U.u2.s  } = _193_ + \add_4s_4ns_4_2_1_U11.top_add_4s_4ns_4_2_1_Adder_8_U.u2.cin ;
always @(posedge \add_6ns_6s_6_2_1_U9.top_add_6ns_6s_6_2_1_Adder_6_U.clk )
\add_6ns_6s_6_2_1_U9.top_add_6ns_6s_6_2_1_Adder_6_U.bin_s1  <= _195_;
always @(posedge \add_6ns_6s_6_2_1_U9.top_add_6ns_6s_6_2_1_Adder_6_U.clk )
\add_6ns_6s_6_2_1_U9.top_add_6ns_6s_6_2_1_Adder_6_U.ain_s1  <= _194_;
always @(posedge \add_6ns_6s_6_2_1_U9.top_add_6ns_6s_6_2_1_Adder_6_U.clk )
\add_6ns_6s_6_2_1_U9.top_add_6ns_6s_6_2_1_Adder_6_U.sum_s1  <= _197_;
always @(posedge \add_6ns_6s_6_2_1_U9.top_add_6ns_6s_6_2_1_Adder_6_U.clk )
\add_6ns_6s_6_2_1_U9.top_add_6ns_6s_6_2_1_Adder_6_U.carry_s1  <= _196_;
assign _195_ = \add_6ns_6s_6_2_1_U9.top_add_6ns_6s_6_2_1_Adder_6_U.ce  ? \add_6ns_6s_6_2_1_U9.top_add_6ns_6s_6_2_1_Adder_6_U.b [5:3] : \add_6ns_6s_6_2_1_U9.top_add_6ns_6s_6_2_1_Adder_6_U.bin_s1 ;
assign _194_ = \add_6ns_6s_6_2_1_U9.top_add_6ns_6s_6_2_1_Adder_6_U.ce  ? \add_6ns_6s_6_2_1_U9.top_add_6ns_6s_6_2_1_Adder_6_U.a [5:3] : \add_6ns_6s_6_2_1_U9.top_add_6ns_6s_6_2_1_Adder_6_U.ain_s1 ;
assign _196_ = \add_6ns_6s_6_2_1_U9.top_add_6ns_6s_6_2_1_Adder_6_U.ce  ? \add_6ns_6s_6_2_1_U9.top_add_6ns_6s_6_2_1_Adder_6_U.facout_s1  : \add_6ns_6s_6_2_1_U9.top_add_6ns_6s_6_2_1_Adder_6_U.carry_s1 ;
assign _197_ = \add_6ns_6s_6_2_1_U9.top_add_6ns_6s_6_2_1_Adder_6_U.ce  ? \add_6ns_6s_6_2_1_U9.top_add_6ns_6s_6_2_1_Adder_6_U.fas_s1  : \add_6ns_6s_6_2_1_U9.top_add_6ns_6s_6_2_1_Adder_6_U.sum_s1 ;
assign _198_ = \add_6ns_6s_6_2_1_U9.top_add_6ns_6s_6_2_1_Adder_6_U.u1.a  + \add_6ns_6s_6_2_1_U9.top_add_6ns_6s_6_2_1_Adder_6_U.u1.b ;
assign { \add_6ns_6s_6_2_1_U9.top_add_6ns_6s_6_2_1_Adder_6_U.u1.cout , \add_6ns_6s_6_2_1_U9.top_add_6ns_6s_6_2_1_Adder_6_U.u1.s  } = _198_ + \add_6ns_6s_6_2_1_U9.top_add_6ns_6s_6_2_1_Adder_6_U.u1.cin ;
assign _199_ = \add_6ns_6s_6_2_1_U9.top_add_6ns_6s_6_2_1_Adder_6_U.u2.a  + \add_6ns_6s_6_2_1_U9.top_add_6ns_6s_6_2_1_Adder_6_U.u2.b ;
assign { \add_6ns_6s_6_2_1_U9.top_add_6ns_6s_6_2_1_Adder_6_U.u2.cout , \add_6ns_6s_6_2_1_U9.top_add_6ns_6s_6_2_1_Adder_6_U.u2.s  } = _199_ + \add_6ns_6s_6_2_1_U9.top_add_6ns_6s_6_2_1_Adder_6_U.u2.cin ;
always @(posedge \add_9ns_9ns_9_2_1_U21.top_add_9ns_9ns_9_2_1_Adder_15_U.clk )
\add_9ns_9ns_9_2_1_U21.top_add_9ns_9ns_9_2_1_Adder_15_U.bin_s1  <= _201_;
always @(posedge \add_9ns_9ns_9_2_1_U21.top_add_9ns_9ns_9_2_1_Adder_15_U.clk )
\add_9ns_9ns_9_2_1_U21.top_add_9ns_9ns_9_2_1_Adder_15_U.ain_s1  <= _200_;
always @(posedge \add_9ns_9ns_9_2_1_U21.top_add_9ns_9ns_9_2_1_Adder_15_U.clk )
\add_9ns_9ns_9_2_1_U21.top_add_9ns_9ns_9_2_1_Adder_15_U.sum_s1  <= _203_;
always @(posedge \add_9ns_9ns_9_2_1_U21.top_add_9ns_9ns_9_2_1_Adder_15_U.clk )
\add_9ns_9ns_9_2_1_U21.top_add_9ns_9ns_9_2_1_Adder_15_U.carry_s1  <= _202_;
assign _201_ = \add_9ns_9ns_9_2_1_U21.top_add_9ns_9ns_9_2_1_Adder_15_U.ce  ? \add_9ns_9ns_9_2_1_U21.top_add_9ns_9ns_9_2_1_Adder_15_U.b [8:4] : \add_9ns_9ns_9_2_1_U21.top_add_9ns_9ns_9_2_1_Adder_15_U.bin_s1 ;
assign _200_ = \add_9ns_9ns_9_2_1_U21.top_add_9ns_9ns_9_2_1_Adder_15_U.ce  ? \add_9ns_9ns_9_2_1_U21.top_add_9ns_9ns_9_2_1_Adder_15_U.a [8:4] : \add_9ns_9ns_9_2_1_U21.top_add_9ns_9ns_9_2_1_Adder_15_U.ain_s1 ;
assign _202_ = \add_9ns_9ns_9_2_1_U21.top_add_9ns_9ns_9_2_1_Adder_15_U.ce  ? \add_9ns_9ns_9_2_1_U21.top_add_9ns_9ns_9_2_1_Adder_15_U.facout_s1  : \add_9ns_9ns_9_2_1_U21.top_add_9ns_9ns_9_2_1_Adder_15_U.carry_s1 ;
assign _203_ = \add_9ns_9ns_9_2_1_U21.top_add_9ns_9ns_9_2_1_Adder_15_U.ce  ? \add_9ns_9ns_9_2_1_U21.top_add_9ns_9ns_9_2_1_Adder_15_U.fas_s1  : \add_9ns_9ns_9_2_1_U21.top_add_9ns_9ns_9_2_1_Adder_15_U.sum_s1 ;
assign _204_ = \add_9ns_9ns_9_2_1_U21.top_add_9ns_9ns_9_2_1_Adder_15_U.u1.a  + \add_9ns_9ns_9_2_1_U21.top_add_9ns_9ns_9_2_1_Adder_15_U.u1.b ;
assign { \add_9ns_9ns_9_2_1_U21.top_add_9ns_9ns_9_2_1_Adder_15_U.u1.cout , \add_9ns_9ns_9_2_1_U21.top_add_9ns_9ns_9_2_1_Adder_15_U.u1.s  } = _204_ + \add_9ns_9ns_9_2_1_U21.top_add_9ns_9ns_9_2_1_Adder_15_U.u1.cin ;
assign _205_ = \add_9ns_9ns_9_2_1_U21.top_add_9ns_9ns_9_2_1_Adder_15_U.u2.a  + \add_9ns_9ns_9_2_1_U21.top_add_9ns_9ns_9_2_1_Adder_15_U.u2.b ;
assign { \add_9ns_9ns_9_2_1_U21.top_add_9ns_9ns_9_2_1_Adder_15_U.u2.cout , \add_9ns_9ns_9_2_1_U21.top_add_9ns_9ns_9_2_1_Adder_15_U.u2.s  } = _205_ + \add_9ns_9ns_9_2_1_U21.top_add_9ns_9ns_9_2_1_Adder_15_U.u2.cin ;
assign \mul_4s_2s_6_7_1_U1.top_mul_4s_2s_6_7_1_Mul_DSP_0_U.tmp_product  = $signed(\mul_4s_2s_6_7_1_U1.top_mul_4s_2s_6_7_1_Mul_DSP_0_U.a_reg0 ) * $signed(\mul_4s_2s_6_7_1_U1.top_mul_4s_2s_6_7_1_Mul_DSP_0_U.b_reg0 );
always @(posedge \mul_4s_2s_6_7_1_U1.top_mul_4s_2s_6_7_1_Mul_DSP_0_U.clk )
\mul_4s_2s_6_7_1_U1.top_mul_4s_2s_6_7_1_Mul_DSP_0_U.a_reg0  <= _206_;
always @(posedge \mul_4s_2s_6_7_1_U1.top_mul_4s_2s_6_7_1_Mul_DSP_0_U.clk )
\mul_4s_2s_6_7_1_U1.top_mul_4s_2s_6_7_1_Mul_DSP_0_U.b_reg0  <= _207_;
always @(posedge \mul_4s_2s_6_7_1_U1.top_mul_4s_2s_6_7_1_Mul_DSP_0_U.clk )
\mul_4s_2s_6_7_1_U1.top_mul_4s_2s_6_7_1_Mul_DSP_0_U.buff0  <= _208_;
always @(posedge \mul_4s_2s_6_7_1_U1.top_mul_4s_2s_6_7_1_Mul_DSP_0_U.clk )
\mul_4s_2s_6_7_1_U1.top_mul_4s_2s_6_7_1_Mul_DSP_0_U.buff1  <= _209_;
always @(posedge \mul_4s_2s_6_7_1_U1.top_mul_4s_2s_6_7_1_Mul_DSP_0_U.clk )
\mul_4s_2s_6_7_1_U1.top_mul_4s_2s_6_7_1_Mul_DSP_0_U.buff2  <= _210_;
always @(posedge \mul_4s_2s_6_7_1_U1.top_mul_4s_2s_6_7_1_Mul_DSP_0_U.clk )
\mul_4s_2s_6_7_1_U1.top_mul_4s_2s_6_7_1_Mul_DSP_0_U.buff3  <= _211_;
always @(posedge \mul_4s_2s_6_7_1_U1.top_mul_4s_2s_6_7_1_Mul_DSP_0_U.clk )
\mul_4s_2s_6_7_1_U1.top_mul_4s_2s_6_7_1_Mul_DSP_0_U.buff4  <= _212_;
assign _212_ = \mul_4s_2s_6_7_1_U1.top_mul_4s_2s_6_7_1_Mul_DSP_0_U.ce  ? \mul_4s_2s_6_7_1_U1.top_mul_4s_2s_6_7_1_Mul_DSP_0_U.buff3  : \mul_4s_2s_6_7_1_U1.top_mul_4s_2s_6_7_1_Mul_DSP_0_U.buff4 ;
assign _211_ = \mul_4s_2s_6_7_1_U1.top_mul_4s_2s_6_7_1_Mul_DSP_0_U.ce  ? \mul_4s_2s_6_7_1_U1.top_mul_4s_2s_6_7_1_Mul_DSP_0_U.buff2  : \mul_4s_2s_6_7_1_U1.top_mul_4s_2s_6_7_1_Mul_DSP_0_U.buff3 ;
assign _210_ = \mul_4s_2s_6_7_1_U1.top_mul_4s_2s_6_7_1_Mul_DSP_0_U.ce  ? \mul_4s_2s_6_7_1_U1.top_mul_4s_2s_6_7_1_Mul_DSP_0_U.buff1  : \mul_4s_2s_6_7_1_U1.top_mul_4s_2s_6_7_1_Mul_DSP_0_U.buff2 ;
assign _209_ = \mul_4s_2s_6_7_1_U1.top_mul_4s_2s_6_7_1_Mul_DSP_0_U.ce  ? \mul_4s_2s_6_7_1_U1.top_mul_4s_2s_6_7_1_Mul_DSP_0_U.buff0  : \mul_4s_2s_6_7_1_U1.top_mul_4s_2s_6_7_1_Mul_DSP_0_U.buff1 ;
assign _208_ = \mul_4s_2s_6_7_1_U1.top_mul_4s_2s_6_7_1_Mul_DSP_0_U.ce  ? \mul_4s_2s_6_7_1_U1.top_mul_4s_2s_6_7_1_Mul_DSP_0_U.tmp_product  : \mul_4s_2s_6_7_1_U1.top_mul_4s_2s_6_7_1_Mul_DSP_0_U.buff0 ;
assign _207_ = \mul_4s_2s_6_7_1_U1.top_mul_4s_2s_6_7_1_Mul_DSP_0_U.ce  ? \mul_4s_2s_6_7_1_U1.top_mul_4s_2s_6_7_1_Mul_DSP_0_U.b  : \mul_4s_2s_6_7_1_U1.top_mul_4s_2s_6_7_1_Mul_DSP_0_U.b_reg0 ;
assign _206_ = \mul_4s_2s_6_7_1_U1.top_mul_4s_2s_6_7_1_Mul_DSP_0_U.ce  ? \mul_4s_2s_6_7_1_U1.top_mul_4s_2s_6_7_1_Mul_DSP_0_U.a  : \mul_4s_2s_6_7_1_U1.top_mul_4s_2s_6_7_1_Mul_DSP_0_U.a_reg0 ;
always @(posedge \shl_20s_2ns_20_7_1_U6.clk )
\shl_20s_2ns_20_7_1_U6.dout_array[5]  <= _224_;
always @(posedge \shl_20s_2ns_20_7_1_U6.clk )
\shl_20s_2ns_20_7_1_U6.din1_cast_array[5]  <= _218_;
always @(posedge \shl_20s_2ns_20_7_1_U6.clk )
\shl_20s_2ns_20_7_1_U6.dout_array[4]  <= _223_;
always @(posedge \shl_20s_2ns_20_7_1_U6.clk )
\shl_20s_2ns_20_7_1_U6.din1_cast_array[4]  <= _217_;
always @(posedge \shl_20s_2ns_20_7_1_U6.clk )
\shl_20s_2ns_20_7_1_U6.dout_array[3]  <= _222_;
always @(posedge \shl_20s_2ns_20_7_1_U6.clk )
\shl_20s_2ns_20_7_1_U6.din1_cast_array[3]  <= _216_;
always @(posedge \shl_20s_2ns_20_7_1_U6.clk )
\shl_20s_2ns_20_7_1_U6.dout_array[2]  <= _221_;
always @(posedge \shl_20s_2ns_20_7_1_U6.clk )
\shl_20s_2ns_20_7_1_U6.din1_cast_array[2]  <= _215_;
always @(posedge \shl_20s_2ns_20_7_1_U6.clk )
\shl_20s_2ns_20_7_1_U6.dout_array[1]  <= _220_;
always @(posedge \shl_20s_2ns_20_7_1_U6.clk )
\shl_20s_2ns_20_7_1_U6.din1_cast_array[1]  <= _214_;
always @(posedge \shl_20s_2ns_20_7_1_U6.clk )
\shl_20s_2ns_20_7_1_U6.dout_array[0]  <= _219_;
always @(posedge \shl_20s_2ns_20_7_1_U6.clk )
\shl_20s_2ns_20_7_1_U6.din1_cast_array[0]  <= _213_;
assign _225_ = \shl_20s_2ns_20_7_1_U6.ce  ? \shl_20s_2ns_20_7_1_U6.din1_cast_array[4]  : \shl_20s_2ns_20_7_1_U6.din1_cast_array[5] ;
assign _218_ = \shl_20s_2ns_20_7_1_U6.reset  ? 2'h0 : _225_;
assign _226_ = \shl_20s_2ns_20_7_1_U6.ce  ? _237_ : \shl_20s_2ns_20_7_1_U6.dout_array[5] ;
assign _224_ = \shl_20s_2ns_20_7_1_U6.reset  ? 20'h00000 : _226_;
assign _227_ = \shl_20s_2ns_20_7_1_U6.ce  ? \shl_20s_2ns_20_7_1_U6.din1_cast_array[3]  : \shl_20s_2ns_20_7_1_U6.din1_cast_array[4] ;
assign _217_ = \shl_20s_2ns_20_7_1_U6.reset  ? 2'h0 : _227_;
assign _228_ = \shl_20s_2ns_20_7_1_U6.ce  ? \shl_20s_2ns_20_7_1_U6.dout_array[3]  : \shl_20s_2ns_20_7_1_U6.dout_array[4] ;
assign _223_ = \shl_20s_2ns_20_7_1_U6.reset  ? 20'h00000 : _228_;
assign _229_ = \shl_20s_2ns_20_7_1_U6.ce  ? \shl_20s_2ns_20_7_1_U6.din1_cast_array[2]  : \shl_20s_2ns_20_7_1_U6.din1_cast_array[3] ;
assign _216_ = \shl_20s_2ns_20_7_1_U6.reset  ? 2'h0 : _229_;
assign _230_ = \shl_20s_2ns_20_7_1_U6.ce  ? \shl_20s_2ns_20_7_1_U6.dout_array[2]  : \shl_20s_2ns_20_7_1_U6.dout_array[3] ;
assign _222_ = \shl_20s_2ns_20_7_1_U6.reset  ? 20'h00000 : _230_;
assign _231_ = \shl_20s_2ns_20_7_1_U6.ce  ? \shl_20s_2ns_20_7_1_U6.din1_cast_array[1]  : \shl_20s_2ns_20_7_1_U6.din1_cast_array[2] ;
assign _215_ = \shl_20s_2ns_20_7_1_U6.reset  ? 2'h0 : _231_;
assign _232_ = \shl_20s_2ns_20_7_1_U6.ce  ? \shl_20s_2ns_20_7_1_U6.dout_array[1]  : \shl_20s_2ns_20_7_1_U6.dout_array[2] ;
assign _221_ = \shl_20s_2ns_20_7_1_U6.reset  ? 20'h00000 : _232_;
assign _233_ = \shl_20s_2ns_20_7_1_U6.ce  ? \shl_20s_2ns_20_7_1_U6.din1_cast_array[0]  : \shl_20s_2ns_20_7_1_U6.din1_cast_array[1] ;
assign _214_ = \shl_20s_2ns_20_7_1_U6.reset  ? 2'h0 : _233_;
assign _234_ = \shl_20s_2ns_20_7_1_U6.ce  ? \shl_20s_2ns_20_7_1_U6.dout_array[0]  : \shl_20s_2ns_20_7_1_U6.dout_array[1] ;
assign _220_ = \shl_20s_2ns_20_7_1_U6.reset  ? 20'h00000 : _234_;
assign _235_ = \shl_20s_2ns_20_7_1_U6.ce  ? \shl_20s_2ns_20_7_1_U6.din1 [1:0] : \shl_20s_2ns_20_7_1_U6.din1_cast_array[0] ;
assign _213_ = \shl_20s_2ns_20_7_1_U6.reset  ? 2'h0 : _235_;
assign _236_ = \shl_20s_2ns_20_7_1_U6.ce  ? \shl_20s_2ns_20_7_1_U6.din0  : \shl_20s_2ns_20_7_1_U6.dout_array[0] ;
assign _219_ = \shl_20s_2ns_20_7_1_U6.reset  ? 20'h00000 : _236_;
assign _237_ = \shl_20s_2ns_20_7_1_U6.dout_array[4]  << { \shl_20s_2ns_20_7_1_U6.din1_cast_array[4] [1], 1'h0 };
assign \shl_20s_2ns_20_7_1_U6.dout  = \shl_20s_2ns_20_7_1_U6.dout_array[5]  << \shl_20s_2ns_20_7_1_U6.din1_cast_array[5] [0];
assign \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.bin_s0  = ~ \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.b ;
always @(posedge \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.clk )
\sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.bin_s1  <= _239_;
always @(posedge \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.clk )
\sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.ain_s1  <= _238_;
always @(posedge \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.clk )
\sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.sum_s1  <= _241_;
always @(posedge \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.clk )
\sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.carry_s1  <= _240_;
assign _239_ = \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.ce  ? \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.bin_s0 [4:2] : \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.bin_s1 ;
assign _238_ = \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.ce  ? \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.a [4:2] : \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.ain_s1 ;
assign _240_ = \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.ce  ? \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.facout_s1  : \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.carry_s1 ;
assign _241_ = \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.ce  ? \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.fas_s1  : \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.sum_s1 ;
assign _242_ = \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.u1.a  + \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.u1.b ;
assign { \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.u1.cout , \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.u1.s  } = _242_ + \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.u1.cin ;
assign _243_ = \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.u2.a  + \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.u2.b ;
assign { \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.u2.cout , \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.u2.s  } = _243_ + \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.u2.cin ;
assign \sub_5s_5s_5_2_1_U2.top_sub_5s_5s_5_2_1_Adder_0_U.bin_s0  = ~ \sub_5s_5s_5_2_1_U2.top_sub_5s_5s_5_2_1_Adder_0_U.b ;
always @(posedge \sub_5s_5s_5_2_1_U2.top_sub_5s_5s_5_2_1_Adder_0_U.clk )
\sub_5s_5s_5_2_1_U2.top_sub_5s_5s_5_2_1_Adder_0_U.bin_s1  <= _245_;
always @(posedge \sub_5s_5s_5_2_1_U2.top_sub_5s_5s_5_2_1_Adder_0_U.clk )
\sub_5s_5s_5_2_1_U2.top_sub_5s_5s_5_2_1_Adder_0_U.ain_s1  <= _244_;
always @(posedge \sub_5s_5s_5_2_1_U2.top_sub_5s_5s_5_2_1_Adder_0_U.clk )
\sub_5s_5s_5_2_1_U2.top_sub_5s_5s_5_2_1_Adder_0_U.sum_s1  <= _247_;
always @(posedge \sub_5s_5s_5_2_1_U2.top_sub_5s_5s_5_2_1_Adder_0_U.clk )
\sub_5s_5s_5_2_1_U2.top_sub_5s_5s_5_2_1_Adder_0_U.carry_s1  <= _246_;
assign _245_ = \sub_5s_5s_5_2_1_U2.top_sub_5s_5s_5_2_1_Adder_0_U.ce  ? \sub_5s_5s_5_2_1_U2.top_sub_5s_5s_5_2_1_Adder_0_U.bin_s0 [4:2] : \sub_5s_5s_5_2_1_U2.top_sub_5s_5s_5_2_1_Adder_0_U.bin_s1 ;
assign _244_ = \sub_5s_5s_5_2_1_U2.top_sub_5s_5s_5_2_1_Adder_0_U.ce  ? \sub_5s_5s_5_2_1_U2.top_sub_5s_5s_5_2_1_Adder_0_U.a [4:2] : \sub_5s_5s_5_2_1_U2.top_sub_5s_5s_5_2_1_Adder_0_U.ain_s1 ;
assign _246_ = \sub_5s_5s_5_2_1_U2.top_sub_5s_5s_5_2_1_Adder_0_U.ce  ? \sub_5s_5s_5_2_1_U2.top_sub_5s_5s_5_2_1_Adder_0_U.facout_s1  : \sub_5s_5s_5_2_1_U2.top_sub_5s_5s_5_2_1_Adder_0_U.carry_s1 ;
assign _247_ = \sub_5s_5s_5_2_1_U2.top_sub_5s_5s_5_2_1_Adder_0_U.ce  ? \sub_5s_5s_5_2_1_U2.top_sub_5s_5s_5_2_1_Adder_0_U.fas_s1  : \sub_5s_5s_5_2_1_U2.top_sub_5s_5s_5_2_1_Adder_0_U.sum_s1 ;
assign _248_ = \sub_5s_5s_5_2_1_U2.top_sub_5s_5s_5_2_1_Adder_0_U.u1.a  + \sub_5s_5s_5_2_1_U2.top_sub_5s_5s_5_2_1_Adder_0_U.u1.b ;
assign { \sub_5s_5s_5_2_1_U2.top_sub_5s_5s_5_2_1_Adder_0_U.u1.cout , \sub_5s_5s_5_2_1_U2.top_sub_5s_5s_5_2_1_Adder_0_U.u1.s  } = _248_ + \sub_5s_5s_5_2_1_U2.top_sub_5s_5s_5_2_1_Adder_0_U.u1.cin ;
assign _249_ = \sub_5s_5s_5_2_1_U2.top_sub_5s_5s_5_2_1_Adder_0_U.u2.a  + \sub_5s_5s_5_2_1_U2.top_sub_5s_5s_5_2_1_Adder_0_U.u2.b ;
assign { \sub_5s_5s_5_2_1_U2.top_sub_5s_5s_5_2_1_Adder_0_U.u2.cout , \sub_5s_5s_5_2_1_U2.top_sub_5s_5s_5_2_1_Adder_0_U.u2.s  } = _249_ + \sub_5s_5s_5_2_1_U2.top_sub_5s_5s_5_2_1_Adder_0_U.u2.cin ;
assign _250_ = | p_Result_s_18_reg_1270;
assign _251_ = p_Result_s_18_reg_1270 != 2'h3;
assign _252_ = | trunc_ln851_3_reg_1394;
assign _253_ = | trunc_ln851_4_reg_1573;
assign _254_ = | op_15[4:0];
assign _255_ = | op_17[2:0];
assign or_ln1195_fu_398_p2 = op_4 | { xor_ln1499_fu_384_p2, 1'h0 };
assign or_ln340_1_fu_767_p2 = p_Result_19_reg_1441 | overflow_1_fu_758_p2;
assign or_ln340_fu_476_p2 = p_Result_16_reg_1251 | overflow_fu_462_p2;
assign or_ln785_1_fu_736_p2 = tmp_12_reg_1463 | p_Result_20_reg_1457;
assign or_ln785_2_fu_607_p2 = xor_ln785_2_fu_602_p2 | p_Result_16_reg_1251;
assign or_ln785_3_fu_581_p2 = and_ln785_1_fu_577_p2 | and_ln340_1_fu_573_p2;
assign or_ln785_4_fu_884_p2 = xor_ln785_3_fu_879_p2 | p_Result_19_reg_1441;
assign or_ln785_5_fu_848_p2 = and_ln785_4_fu_844_p2 | and_ln340_3_fu_840_p2;
assign or_ln785_fu_425_p2 = p_Result_17_reg_1263 | icmp_ln768_reg_1291;
assign or_ln786_fu_471_p2 = xor_ln786_fu_466_p2 | icmp_ln786_reg_1296;
always @(posedge ap_clk)
p_Val2_5_reg_1358[0] <= 1'h0;
always @(posedge ap_clk)
select_ln785_reg_1379 <= _068_;
always @(posedge ap_clk)
select_ln785_1_reg_1548 <= _067_;
always @(posedge ap_clk)
select_ln69_reg_1699 <= _065_;
always @(posedge ap_clk)
ret_V_9_reg_1506 <= _059_;
always @(posedge ap_clk)
ret_V_32_reg_1687 <= _053_;
always @(posedge ap_clk)
ret_V_33_cast_reg_1692 <= _054_;
always @(posedge ap_clk)
ret_V_31_reg_1657 <= _052_;
always @(posedge ap_clk)
ret_V_30_reg_1640 <= _050_;
always @(posedge ap_clk)
ret_V_31_cast_reg_1645 <= _051_;
always @(posedge ap_clk)
ret_V_29_reg_1610 <= _048_;
always @(posedge ap_clk)
ret_V_28_reg_1593 <= _046_;
always @(posedge ap_clk)
ret_V_29_cast_reg_1598 <= _047_;
always @(posedge ap_clk)
ret_V_10_reg_1528 <= _037_;
always @(posedge ap_clk)
select_ln340_1_reg_1533 <= _063_;
always @(posedge ap_clk)
sel_tmp24_reg_1538 <= _062_;
always @(posedge ap_clk)
ret_V_27_reg_1543 <= _045_;
always @(posedge ap_clk)
r_V_reg_1189 <= _036_;
always @(posedge ap_clk)
ret_V_3_cast_reg_1194 <= _056_;
always @(posedge ap_clk)
trunc_ln851_1_reg_1201 <= _074_;
always @(posedge ap_clk)
select_ln703_reg_1353 <= _066_;
always @(posedge ap_clk)
p_Val2_5_reg_1358[3:1] <= _033_;
always @(posedge ap_clk)
select_ln340_reg_1364 <= _064_;
always @(posedge ap_clk)
sel_tmp11_reg_1369 <= _061_;
always @(posedge ap_clk)
ret_V_24_reg_1424 <= _042_;
always @(posedge ap_clk)
ret_V_8_reg_1429 <= _058_;
always @(posedge ap_clk)
r_V_1_reg_1436 <= _035_;
always @(posedge ap_clk)
p_Result_19_reg_1441 <= _030_;
always @(posedge ap_clk)
p_Val2_8_reg_1449 <= _034_;
always @(posedge ap_clk)
p_Result_20_reg_1457 <= _031_;
always @(posedge ap_clk)
tmp_12_reg_1463 <= _070_;
always @(posedge ap_clk)
ret_V_26_reg_1470 <= _044_;
always @(posedge ap_clk)
tmp_3_reg_1475 <= _071_;
always @(posedge ap_clk)
ret_V_20_reg_1222 <= _038_;
always @(posedge ap_clk)
ret_V_reg_1227 <= _060_;
always @(posedge ap_clk)
trunc_ln851_reg_1234 <= _077_;
always @(posedge ap_clk)
ret_V_4_reg_1239 <= _057_;
always @(posedge ap_clk)
ret_V_25_reg_1244 <= _043_;
always @(posedge ap_clk)
p_Result_16_reg_1251 <= _028_;
always @(posedge ap_clk)
trunc_ln731_reg_1258 <= _073_;
always @(posedge ap_clk)
p_Result_17_reg_1263 <= _029_;
always @(posedge ap_clk)
p_Result_s_18_reg_1270 <= _032_;
always @(posedge ap_clk)
ret_V_2_reg_1302 <= _049_;
always @(posedge ap_clk)
or_ln785_reg_1312 <= _026_;
always @(posedge ap_clk)
xor_ln785_reg_1318 <= _079_;
always @(posedge ap_clk)
xor_ln786_2_reg_1511 <= _080_;
always @(posedge ap_clk)
or_ln340_1_reg_1517 <= _023_;
always @(posedge ap_clk)
op_26_V_reg_1667 <= _021_;
always @(posedge ap_clk)
op_24_V_reg_1620 <= _020_;
always @(posedge ap_clk)
op_13_V_reg_1563 <= _018_;
always @(posedge ap_clk)
op_22_V_reg_1568 <= _019_;
always @(posedge ap_clk)
trunc_ln851_4_reg_1573 <= _076_;
always @(posedge ap_clk)
ret_V_23_reg_1384 <= _041_;
always @(posedge ap_clk)
op_11_V_reg_1389 <= _017_;
always @(posedge ap_clk)
trunc_ln851_3_reg_1394 <= _075_;
always @(posedge ap_clk)
icmp_ln851_6_reg_1682 <= _015_;
always @(posedge ap_clk)
icmp_ln851_5_reg_1635 <= _014_;
always @(posedge ap_clk)
icmp_ln851_4_reg_1588 <= _013_;
always @(posedge ap_clk)
icmp_ln851_3_reg_1419 <= _012_;
always @(posedge ap_clk)
icmp_ln851_2_reg_1179 <= _011_;
always @(posedge ap_clk)
tmp_reg_1184 <= _072_;
always @(posedge ap_clk)
icmp_ln851_1_reg_1217 <= _010_;
always @(posedge ap_clk)
icmp_ln851_reg_1276 <= _016_;
always @(posedge ap_clk)
ret_V_22_reg_1281 <= _040_;
always @(posedge ap_clk)
or_ln1195_reg_1286 <= _022_;
always @(posedge ap_clk)
icmp_ln768_reg_1291 <= _008_;
always @(posedge ap_clk)
icmp_ln786_reg_1296 <= _009_;
always @(posedge ap_clk)
ret_V_21_reg_1329 <= _039_;
always @(posedge ap_clk)
or_ln786_reg_1335 <= _027_;
always @(posedge ap_clk)
or_ln340_reg_1341 <= _024_;
always @(posedge ap_clk)
and_ln786_reg_1347 <= _006_;
always @(posedge ap_clk)
or_ln785_1_reg_1480 <= _025_;
always @(posedge ap_clk)
xor_ln785_1_reg_1486 <= _078_;
always @(posedge ap_clk)
and_ln786_1_reg_1492 <= _005_;
always @(posedge ap_clk)
sext_ln850_reg_1499 <= _069_;
always @(posedge ap_clk)
ret_V_33_reg_1714 <= _055_;
always @(posedge ap_clk)
add_ln69_reg_1719 <= _004_;
always @(posedge ap_clk)
add_ln691_reg_1523 <= _003_;
always @(posedge ap_clk)
add_ln691_3_reg_1704 <= _002_;
always @(posedge ap_clk)
add_ln691_2_reg_1652 <= _001_;
always @(posedge ap_clk)
add_ln691_1_reg_1605 <= _000_;
always @(posedge ap_clk)
ap_CS_fsm <= _007_;
assign _081_ = _090_ ? 2'h2 : 2'h1;
assign _256_ = ap_CS_fsm == 1'h1;
function [42:0] _738_;
input [42:0] a;
input [1848:0] b;
input [42:0] s;
case (s)
43'b0000000000000000000000000000000000000000001:
_738_ = b[42:0];
43'b0000000000000000000000000000000000000000010:
_738_ = b[85:43];
43'b0000000000000000000000000000000000000000100:
_738_ = b[128:86];
43'b0000000000000000000000000000000000000001000:
_738_ = b[171:129];
43'b0000000000000000000000000000000000000010000:
_738_ = b[214:172];
43'b0000000000000000000000000000000000000100000:
_738_ = b[257:215];
43'b0000000000000000000000000000000000001000000:
_738_ = b[300:258];
43'b0000000000000000000000000000000000010000000:
_738_ = b[343:301];
43'b0000000000000000000000000000000000100000000:
_738_ = b[386:344];
43'b0000000000000000000000000000000001000000000:
_738_ = b[429:387];
43'b0000000000000000000000000000000010000000000:
_738_ = b[472:430];
43'b0000000000000000000000000000000100000000000:
_738_ = b[515:473];
43'b0000000000000000000000000000001000000000000:
_738_ = b[558:516];
43'b0000000000000000000000000000010000000000000:
_738_ = b[601:559];
43'b0000000000000000000000000000100000000000000:
_738_ = b[644:602];
43'b0000000000000000000000000001000000000000000:
_738_ = b[687:645];
43'b0000000000000000000000000010000000000000000:
_738_ = b[730:688];
43'b0000000000000000000000000100000000000000000:
_738_ = b[773:731];
43'b0000000000000000000000001000000000000000000:
_738_ = b[816:774];
43'b0000000000000000000000010000000000000000000:
_738_ = b[859:817];
43'b0000000000000000000000100000000000000000000:
_738_ = b[902:860];
43'b0000000000000000000001000000000000000000000:
_738_ = b[945:903];
43'b0000000000000000000010000000000000000000000:
_738_ = b[988:946];
43'b0000000000000000000100000000000000000000000:
_738_ = b[1031:989];
43'b0000000000000000001000000000000000000000000:
_738_ = b[1074:1032];
43'b0000000000000000010000000000000000000000000:
_738_ = b[1117:1075];
43'b0000000000000000100000000000000000000000000:
_738_ = b[1160:1118];
43'b0000000000000001000000000000000000000000000:
_738_ = b[1203:1161];
43'b0000000000000010000000000000000000000000000:
_738_ = b[1246:1204];
43'b0000000000000100000000000000000000000000000:
_738_ = b[1289:1247];
43'b0000000000001000000000000000000000000000000:
_738_ = b[1332:1290];
43'b0000000000010000000000000000000000000000000:
_738_ = b[1375:1333];
43'b0000000000100000000000000000000000000000000:
_738_ = b[1418:1376];
43'b0000000001000000000000000000000000000000000:
_738_ = b[1461:1419];
43'b0000000010000000000000000000000000000000000:
_738_ = b[1504:1462];
43'b0000000100000000000000000000000000000000000:
_738_ = b[1547:1505];
43'b0000001000000000000000000000000000000000000:
_738_ = b[1590:1548];
43'b0000010000000000000000000000000000000000000:
_738_ = b[1633:1591];
43'b0000100000000000000000000000000000000000000:
_738_ = b[1676:1634];
43'b0001000000000000000000000000000000000000000:
_738_ = b[1719:1677];
43'b0010000000000000000000000000000000000000000:
_738_ = b[1762:1720];
43'b0100000000000000000000000000000000000000000:
_738_ = b[1805:1763];
43'b1000000000000000000000000000000000000000000:
_738_ = b[1848:1806];
43'b0000000000000000000000000000000000000000000:
_738_ = a;
default:
_738_ = 43'bx;
endcase
endfunction
assign ap_NS_fsm = _738_(43'hxxxxxxxxxxx, { 41'h00000000000, _081_, 1806'h00000000002000000000080000000002000000000080000000002000000000080000000002000000000080000000002000000000080000000002000000000080000000002000000000080000000002000000000080000000002000000000080000000002000000000080000000002000000000080000000002000000000080000000002000000000080000000002000000000080000000002000000000080000000002000000000080000000002000000000080000000002000000000080000000002000000000080000000002000000000080000000002000000000000000000001 }, { _256_, _298_, _297_, _296_, _295_, _294_, _293_, _292_, _291_, _290_, _289_, _288_, _287_, _286_, _285_, _284_, _283_, _282_, _281_, _280_, _279_, _278_, _277_, _276_, _275_, _274_, _273_, _272_, _271_, _270_, _269_, _268_, _267_, _266_, _265_, _264_, _263_, _262_, _261_, _260_, _259_, _258_, _257_ });
assign _257_ = ap_CS_fsm == 43'h40000000000;
assign _258_ = ap_CS_fsm == 42'h20000000000;
assign _259_ = ap_CS_fsm == 41'h10000000000;
assign _260_ = ap_CS_fsm == 40'h8000000000;
assign _261_ = ap_CS_fsm == 39'h4000000000;
assign _262_ = ap_CS_fsm == 38'h2000000000;
assign _263_ = ap_CS_fsm == 37'h1000000000;
assign _264_ = ap_CS_fsm == 36'h800000000;
assign _265_ = ap_CS_fsm == 35'h400000000;
assign _266_ = ap_CS_fsm == 34'h200000000;
assign _267_ = ap_CS_fsm == 33'h100000000;
assign _268_ = ap_CS_fsm == 32'd2147483648;
assign _269_ = ap_CS_fsm == 31'h40000000;
assign _270_ = ap_CS_fsm == 30'h20000000;
assign _271_ = ap_CS_fsm == 29'h10000000;
assign _272_ = ap_CS_fsm == 28'h8000000;
assign _273_ = ap_CS_fsm == 27'h4000000;
assign _274_ = ap_CS_fsm == 26'h2000000;
assign _275_ = ap_CS_fsm == 25'h1000000;
assign _276_ = ap_CS_fsm == 24'h800000;
assign _277_ = ap_CS_fsm == 23'h400000;
assign _278_ = ap_CS_fsm == 22'h200000;
assign _279_ = ap_CS_fsm == 21'h100000;
assign _280_ = ap_CS_fsm == 20'h80000;
assign _281_ = ap_CS_fsm == 19'h40000;
assign _282_ = ap_CS_fsm == 18'h20000;
assign _283_ = ap_CS_fsm == 17'h10000;
assign _284_ = ap_CS_fsm == 16'h8000;
assign _285_ = ap_CS_fsm == 15'h4000;
assign _286_ = ap_CS_fsm == 14'h2000;
assign _287_ = ap_CS_fsm == 13'h1000;
assign _288_ = ap_CS_fsm == 12'h800;
assign _289_ = ap_CS_fsm == 11'h400;
assign _290_ = ap_CS_fsm == 10'h200;
assign _291_ = ap_CS_fsm == 9'h100;
assign _292_ = ap_CS_fsm == 8'h80;
assign _293_ = ap_CS_fsm == 7'h40;
assign _294_ = ap_CS_fsm == 6'h20;
assign _295_ = ap_CS_fsm == 5'h10;
assign _296_ = ap_CS_fsm == 4'h8;
assign _297_ = ap_CS_fsm == 3'h4;
assign _298_ = ap_CS_fsm == 2'h2;
assign op_29_ap_vld = ap_CS_fsm[42] ? 1'h1 : 1'h0;
assign ap_idle = _089_ ? 1'h1 : 1'h0;
assign _068_ = _088_ ? select_ln785_fu_617_p3 : select_ln785_reg_1379;
assign _067_ = _087_ ? select_ln785_1_fu_894_p3 : select_ln785_1_reg_1548;
assign _065_ = ap_CS_fsm[38] ? select_ln69_fu_1109_p3 : select_ln69_reg_1699;
assign _059_ = _086_ ? grp_fu_731_p2 : ret_V_9_reg_1506;
assign _054_ = ap_CS_fsm[37] ? grp_fu_1078_p2[34:3] : ret_V_33_cast_reg_1692;
assign _053_ = ap_CS_fsm[37] ? grp_fu_1078_p2 : ret_V_32_reg_1687;
assign _052_ = ap_CS_fsm[33] ? ret_V_31_fu_1047_p3 : ret_V_31_reg_1657;
assign _051_ = ap_CS_fsm[30] ? grp_fu_1004_p2[36:5] : ret_V_31_cast_reg_1645;
assign _050_ = ap_CS_fsm[30] ? grp_fu_1004_p2 : ret_V_30_reg_1640;
assign _048_ = ap_CS_fsm[26] ? ret_V_29_fu_973_p3 : ret_V_29_reg_1610;
assign _047_ = ap_CS_fsm[23] ? grp_fu_935_p2[35:4] : ret_V_29_cast_reg_1598;
assign _046_ = ap_CS_fsm[23] ? grp_fu_935_p2 : ret_V_28_reg_1593;
assign _045_ = ap_CS_fsm[19] ? ret_V_27_fu_872_p3 : ret_V_27_reg_1543;
assign _062_ = ap_CS_fsm[19] ? sel_tmp24_fu_854_p2 : sel_tmp24_reg_1538;
assign _063_ = ap_CS_fsm[19] ? select_ln340_1_fu_833_p3 : select_ln340_1_reg_1533;
assign _037_ = ap_CS_fsm[19] ? ret_V_10_fu_784_p3 : ret_V_10_reg_1528;
assign _074_ = ap_CS_fsm[6] ? grp_fu_237_p2[2:0] : trunc_ln851_1_reg_1201;
assign _056_ = ap_CS_fsm[6] ? grp_fu_237_p2[4:3] : ret_V_3_cast_reg_1194;
assign _036_ = ap_CS_fsm[6] ? grp_fu_237_p2 : r_V_reg_1189;
assign _061_ = ap_CS_fsm[12] ? sel_tmp11_fu_587_p2 : sel_tmp11_reg_1369;
assign _064_ = ap_CS_fsm[12] ? select_ln340_fu_565_p3 : select_ln340_reg_1364;
assign _033_ = ap_CS_fsm[12] ? trunc_ln731_reg_1258 : p_Val2_5_reg_1358[3:1];
assign _066_ = ap_CS_fsm[12] ? select_ln703_fu_491_p3 : select_ln703_reg_1353;
assign _071_ = ap_CS_fsm[16] ? grp_fu_666_p2[5:3] : tmp_3_reg_1475;
assign _044_ = ap_CS_fsm[16] ? grp_fu_666_p2 : ret_V_26_reg_1470;
assign _070_ = ap_CS_fsm[16] ? grp_fu_437_p2[19] : tmp_12_reg_1463;
assign _031_ = ap_CS_fsm[16] ? grp_fu_437_p2[18] : p_Result_20_reg_1457;
assign _034_ = ap_CS_fsm[16] ? grp_fu_437_p2[18:11] : p_Val2_8_reg_1449;
assign _030_ = ap_CS_fsm[16] ? grp_fu_437_p2[19] : p_Result_19_reg_1441;
assign _035_ = ap_CS_fsm[16] ? grp_fu_437_p2 : r_V_1_reg_1436;
assign _058_ = ap_CS_fsm[16] ? grp_fu_650_p2[11:2] : ret_V_8_reg_1429;
assign _042_ = ap_CS_fsm[16] ? grp_fu_650_p2 : ret_V_24_reg_1424;
assign _032_ = ap_CS_fsm[8] ? grp_fu_305_p2[4:3] : p_Result_s_18_reg_1270;
assign _029_ = ap_CS_fsm[8] ? grp_fu_305_p2[2] : p_Result_17_reg_1263;
assign _073_ = ap_CS_fsm[8] ? grp_fu_305_p2[2:0] : trunc_ln731_reg_1258;
assign _028_ = ap_CS_fsm[8] ? grp_fu_305_p2[4] : p_Result_16_reg_1251;
assign _043_ = ap_CS_fsm[8] ? grp_fu_305_p2 : ret_V_25_reg_1244;
assign _057_ = ap_CS_fsm[8] ? grp_fu_300_p2 : ret_V_4_reg_1239;
assign _077_ = ap_CS_fsm[8] ? grp_fu_289_p2[1:0] : trunc_ln851_reg_1234;
assign _060_ = ap_CS_fsm[8] ? grp_fu_289_p2[4:2] : ret_V_reg_1227;
assign _038_ = ap_CS_fsm[8] ? grp_fu_289_p2 : ret_V_20_reg_1222;
assign _079_ = ap_CS_fsm[10] ? xor_ln785_fu_429_p2 : xor_ln785_reg_1318;
assign _026_ = ap_CS_fsm[10] ? or_ln785_fu_425_p2 : or_ln785_reg_1312;
assign _049_ = ap_CS_fsm[10] ? grp_fu_360_p2 : ret_V_2_reg_1302;
assign _023_ = ap_CS_fsm[18] ? or_ln340_1_fu_767_p2 : or_ln340_1_reg_1517;
assign _080_ = ap_CS_fsm[18] ? xor_ln786_2_fu_762_p2 : xor_ln786_2_reg_1511;
assign _021_ = ap_CS_fsm[35] ? grp_fu_1058_p2 : op_26_V_reg_1667;
assign _020_ = ap_CS_fsm[28] ? grp_fu_984_p2 : op_24_V_reg_1620;
assign _076_ = ap_CS_fsm[21] ? op_13_V_fu_912_p3[3:0] : trunc_ln851_4_reg_1573;
assign _019_ = ap_CS_fsm[21] ? grp_fu_906_p2 : op_22_V_reg_1568;
assign _018_ = ap_CS_fsm[21] ? op_13_V_fu_912_p3 : op_13_V_reg_1563;
assign _075_ = ap_CS_fsm[14] ? op_11_V_fu_623_p3[2:0] : trunc_ln851_3_reg_1394;
assign _017_ = ap_CS_fsm[14] ? op_11_V_fu_623_p3 : op_11_V_reg_1389;
assign _041_ = ap_CS_fsm[14] ? grp_fu_597_p2 : ret_V_23_reg_1384;
assign _015_ = ap_CS_fsm[36] ? icmp_ln851_6_fu_1088_p2 : icmp_ln851_6_reg_1682;
assign _014_ = ap_CS_fsm[29] ? icmp_ln851_5_fu_1014_p2 : icmp_ln851_5_reg_1635;
assign _013_ = ap_CS_fsm[22] ? icmp_ln851_4_fu_941_p2 : icmp_ln851_4_reg_1588;
assign _012_ = ap_CS_fsm[15] ? icmp_ln851_3_fu_672_p2 : icmp_ln851_3_reg_1419;
assign _072_ = ap_CS_fsm[0] ? op_4[1] : tmp_reg_1184;
assign _011_ = ap_CS_fsm[0] ? icmp_ln851_2_fu_247_p2 : icmp_ln851_2_reg_1179;
assign _010_ = ap_CS_fsm[7] ? icmp_ln851_1_fu_295_p2 : icmp_ln851_1_reg_1217;
assign _009_ = ap_CS_fsm[9] ? icmp_ln786_fu_408_p2 : icmp_ln786_reg_1296;
assign _008_ = ap_CS_fsm[9] ? icmp_ln768_fu_403_p2 : icmp_ln768_reg_1291;
assign _022_ = ap_CS_fsm[9] ? or_ln1195_fu_398_p2 : or_ln1195_reg_1286;
assign _040_ = ap_CS_fsm[9] ? ret_V_22_fu_377_p3 : ret_V_22_reg_1281;
assign _016_ = ap_CS_fsm[9] ? icmp_ln851_fu_355_p2 : icmp_ln851_reg_1276;
assign _006_ = ap_CS_fsm[11] ? and_ln786_fu_486_p2 : and_ln786_reg_1347;
assign _024_ = ap_CS_fsm[11] ? or_ln340_fu_476_p2 : or_ln340_reg_1341;
assign _027_ = ap_CS_fsm[11] ? or_ln786_fu_471_p2 : or_ln786_reg_1335;
assign _039_ = ap_CS_fsm[11] ? ret_V_21_fu_455_p3 : ret_V_21_reg_1329;
assign _069_ = ap_CS_fsm[17] ? { tmp_3_reg_1475[2], tmp_3_reg_1475 } : sext_ln850_reg_1499;
assign _005_ = ap_CS_fsm[17] ? and_ln786_1_fu_745_p2 : and_ln786_1_reg_1492;
assign _078_ = ap_CS_fsm[17] ? xor_ln785_1_fu_740_p2 : xor_ln785_1_reg_1486;
assign _025_ = ap_CS_fsm[17] ? or_ln785_1_fu_736_p2 : or_ln785_1_reg_1480;
assign _004_ = ap_CS_fsm[40] ? grp_fu_1124_p2 : add_ln69_reg_1719;
assign _055_ = ap_CS_fsm[40] ? ret_V_33_fu_1141_p3 : ret_V_33_reg_1714;
assign _003_ = _085_ ? grp_fu_752_p2 : add_ln691_reg_1523;
assign _002_ = _084_ ? grp_fu_1104_p2 : add_ln691_3_reg_1704;
assign _001_ = _083_ ? grp_fu_1030_p2 : add_ln691_2_reg_1652;
assign _000_ = _082_ ? grp_fu_956_p2 : add_ln691_1_reg_1605;
assign _007_ = ap_rst ? 43'h00000000001 : ap_NS_fsm;
assign icmp_ln768_fu_403_p2 = _250_ ? 1'h1 : 1'h0;
assign icmp_ln786_fu_408_p2 = _251_ ? 1'h1 : 1'h0;
assign icmp_ln851_1_fu_295_p2 = _095_ ? 1'h1 : 1'h0;
assign icmp_ln851_2_fu_247_p2 = _096_ ? 1'h1 : 1'h0;
assign icmp_ln851_3_fu_672_p2 = _252_ ? 1'h1 : 1'h0;
assign icmp_ln851_4_fu_941_p2 = _253_ ? 1'h1 : 1'h0;
assign icmp_ln851_5_fu_1014_p2 = _254_ ? 1'h1 : 1'h0;
assign icmp_ln851_6_fu_1088_p2 = _255_ ? 1'h1 : 1'h0;
assign icmp_ln851_fu_355_p2 = _097_ ? 1'h1 : 1'h0;
assign op_11_V_fu_623_p3 = sel_tmp11_reg_1369 ? p_Val2_5_reg_1358 : select_ln785_reg_1379;
assign op_13_V_fu_912_p3 = sel_tmp24_reg_1538 ? p_Val2_8_reg_1449 : select_ln785_1_reg_1548;
assign ret_V_10_fu_784_p3 = ret_V_24_reg_1424[11] ? select_ln850_2_fu_779_p3 : ret_V_8_reg_1429;
assign ret_V_21_fu_455_p3 = ret_V_20_reg_1222[4] ? select_ln850_fu_450_p3 : ret_V_reg_1227;
assign ret_V_22_fu_377_p3 = r_V_reg_1189[5] ? select_ln850_1_fu_372_p3 : ret_V_3_cast_reg_1194;
assign ret_V_27_fu_872_p3 = ret_V_26_reg_1470[5] ? select_ln850_3_fu_867_p3 : sext_ln850_reg_1499;
assign ret_V_29_fu_973_p3 = ret_V_28_reg_1593[36] ? select_ln850_4_fu_968_p3 : ret_V_29_cast_reg_1598;
assign ret_V_31_fu_1047_p3 = ret_V_30_reg_1640[37] ? select_ln850_5_fu_1042_p3 : ret_V_31_cast_reg_1645;
assign ret_V_33_fu_1141_p3 = ret_V_32_reg_1687[35] ? select_ln850_6_fu_1136_p3 : ret_V_33_cast_reg_1692;
assign select_ln340_1_fu_833_p3 = and_ln340_2_fu_828_p2 ? p_Val2_8_reg_1449 : { p_Result_19_reg_1441, p_Val2_9_fu_809_p2[6:0] };
assign select_ln340_fu_565_p3 = and_ln340_fu_560_p2 ? { trunc_ln731_reg_1258, 1'h0 } : { ret_V_25_reg_1244[3], p_Val2_6_fu_539_p2 };
assign select_ln69_fu_1109_p3 = op_18 ? 9'h1ff : 9'h000;
assign select_ln703_fu_491_p3 = op_10 ? 3'h7 : 3'h0;
assign select_ln785_1_fu_894_p3 = and_ln785_3_fu_889_p2 ? p_Val2_8_reg_1449 : select_ln340_1_reg_1533;
assign select_ln785_fu_617_p3 = and_ln785_fu_612_p2 ? p_Val2_5_reg_1358 : select_ln340_reg_1364;
assign select_ln850_1_fu_372_p3 = icmp_ln851_1_reg_1217 ? ret_V_3_cast_reg_1194 : ret_V_4_reg_1239;
assign select_ln850_2_fu_779_p3 = icmp_ln851_2_reg_1179 ? ret_V_8_reg_1429 : ret_V_9_reg_1506;
assign select_ln850_3_fu_867_p3 = icmp_ln851_3_reg_1419 ? add_ln691_reg_1523 : sext_ln850_reg_1499;
assign select_ln850_4_fu_968_p3 = icmp_ln851_4_reg_1588 ? add_ln691_1_reg_1605 : ret_V_29_cast_reg_1598;
assign select_ln850_5_fu_1042_p3 = icmp_ln851_5_reg_1635 ? add_ln691_2_reg_1652 : ret_V_31_cast_reg_1645;
assign select_ln850_6_fu_1136_p3 = icmp_ln851_6_reg_1682 ? add_ln691_3_reg_1704 : ret_V_33_cast_reg_1692;
assign select_ln850_fu_450_p3 = icmp_ln851_reg_1276 ? ret_V_reg_1227 : ret_V_2_reg_1302;
assign xor_ln365_2_fu_798_p2 = r_V_1_reg_1436[18] ^ tmp_12_reg_1463;
assign xor_ln365_fu_527_p2 = ret_V_25_reg_1244[2] ^ ret_V_25_reg_1244[3];
assign ap_CS_fsm_state1 = ap_CS_fsm[0];
assign ap_CS_fsm_state10 = ap_CS_fsm[9];
assign ap_CS_fsm_state11 = ap_CS_fsm[10];
assign ap_CS_fsm_state12 = ap_CS_fsm[11];
assign ap_CS_fsm_state13 = ap_CS_fsm[12];
assign ap_CS_fsm_state14 = ap_CS_fsm[13];
assign ap_CS_fsm_state15 = ap_CS_fsm[14];
assign ap_CS_fsm_state16 = ap_CS_fsm[15];
assign ap_CS_fsm_state17 = ap_CS_fsm[16];
assign ap_CS_fsm_state18 = ap_CS_fsm[17];
assign ap_CS_fsm_state19 = ap_CS_fsm[18];
assign ap_CS_fsm_state20 = ap_CS_fsm[19];
assign ap_CS_fsm_state21 = ap_CS_fsm[20];
assign ap_CS_fsm_state22 = ap_CS_fsm[21];
assign ap_CS_fsm_state23 = ap_CS_fsm[22];
assign ap_CS_fsm_state24 = ap_CS_fsm[23];
assign ap_CS_fsm_state25 = ap_CS_fsm[24];
assign ap_CS_fsm_state26 = ap_CS_fsm[25];
assign ap_CS_fsm_state27 = ap_CS_fsm[26];
assign ap_CS_fsm_state28 = ap_CS_fsm[27];
assign ap_CS_fsm_state29 = ap_CS_fsm[28];
assign ap_CS_fsm_state30 = ap_CS_fsm[29];
assign ap_CS_fsm_state31 = ap_CS_fsm[30];
assign ap_CS_fsm_state32 = ap_CS_fsm[31];
assign ap_CS_fsm_state33 = ap_CS_fsm[32];
assign ap_CS_fsm_state34 = ap_CS_fsm[33];
assign ap_CS_fsm_state35 = ap_CS_fsm[34];
assign ap_CS_fsm_state36 = ap_CS_fsm[35];
assign ap_CS_fsm_state37 = ap_CS_fsm[36];
assign ap_CS_fsm_state38 = ap_CS_fsm[37];
assign ap_CS_fsm_state39 = ap_CS_fsm[38];
assign ap_CS_fsm_state40 = ap_CS_fsm[39];
assign ap_CS_fsm_state41 = ap_CS_fsm[40];
assign ap_CS_fsm_state42 = ap_CS_fsm[41];
assign ap_CS_fsm_state43 = ap_CS_fsm[42];
assign ap_CS_fsm_state7 = ap_CS_fsm[6];
assign ap_CS_fsm_state8 = ap_CS_fsm[7];
assign ap_CS_fsm_state9 = ap_CS_fsm[8];
assign ap_done = op_29_ap_vld;
assign ap_ready = op_29_ap_vld;
assign grp_fu_1004_p0 = { op_24_V_reg_1620[31], op_24_V_reg_1620, 5'h00 };
assign grp_fu_1004_p1 = { op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15 };
assign grp_fu_1058_p1 = { 30'h00000000, op_16 };
assign grp_fu_1078_p0 = { op_26_V_reg_1667[31], op_26_V_reg_1667, 3'h0 };
assign grp_fu_1078_p1 = { op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17 };
assign grp_fu_1124_p0 = { 1'h0, ret_V_21_reg_1329[2], ret_V_21_reg_1329[2], ret_V_21_reg_1329[2], ret_V_21_reg_1329[2], ret_V_21_reg_1329[2], ret_V_21_reg_1329 };
assign grp_fu_1151_p0 = { add_ln69_reg_1719[8], add_ln69_reg_1719[8], add_ln69_reg_1719[8], add_ln69_reg_1719[8], add_ln69_reg_1719[8], add_ln69_reg_1719[8], add_ln69_reg_1719[8], add_ln69_reg_1719[8], add_ln69_reg_1719[8], add_ln69_reg_1719[8], add_ln69_reg_1719[8], add_ln69_reg_1719[8], add_ln69_reg_1719[8], add_ln69_reg_1719[8], add_ln69_reg_1719[8], add_ln69_reg_1719[8], add_ln69_reg_1719[8], add_ln69_reg_1719[8], add_ln69_reg_1719[8], add_ln69_reg_1719[8], add_ln69_reg_1719[8], add_ln69_reg_1719[8], add_ln69_reg_1719[8], add_ln69_reg_1719 };
assign grp_fu_289_p0 = { op_4[1], op_4[1], op_4, 1'h0 };
assign grp_fu_437_p0 = { tmp_reg_1184, tmp_reg_1184, tmp_reg_1184, tmp_reg_1184, or_ln1195_reg_1286, 14'h0000 };
assign grp_fu_437_p1 = { 18'h00000, ret_V_22_reg_1281 };
assign grp_fu_597_p0 = { op_6[1], op_6 };
assign grp_fu_650_p0 = { 2'h0, ret_V_21_reg_1329[2], ret_V_21_reg_1329[2], ret_V_21_reg_1329[2], ret_V_21_reg_1329[2], ret_V_21_reg_1329[2], ret_V_21_reg_1329, 2'h0 };
assign grp_fu_650_p1 = { op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5 };
assign grp_fu_666_p0 = { ret_V_23_reg_1384, 3'h0 };
assign grp_fu_666_p1 = { op_11_V_reg_1389[3], op_11_V_reg_1389[3], op_11_V_reg_1389 };
assign grp_fu_752_p0 = { tmp_3_reg_1475[2], tmp_3_reg_1475 };
assign grp_fu_906_p0 = { ret_V_27_reg_1543[3], ret_V_27_reg_1543[3], ret_V_27_reg_1543[3], ret_V_27_reg_1543[3], ret_V_27_reg_1543[3], ret_V_27_reg_1543[3], ret_V_27_reg_1543[3], ret_V_27_reg_1543 };
assign grp_fu_906_p1 = { ret_V_10_reg_1528[9], ret_V_10_reg_1528 };
assign grp_fu_935_p0 = { op_22_V_reg_1568[10], op_22_V_reg_1568[10], op_22_V_reg_1568[10], op_22_V_reg_1568[10], op_22_V_reg_1568[10], op_22_V_reg_1568[10], op_22_V_reg_1568[10], op_22_V_reg_1568[10], op_22_V_reg_1568[10], op_22_V_reg_1568[10], op_22_V_reg_1568[10], op_22_V_reg_1568[10], op_22_V_reg_1568[10], op_22_V_reg_1568[10], op_22_V_reg_1568[10], op_22_V_reg_1568[10], op_22_V_reg_1568[10], op_22_V_reg_1568[10], op_22_V_reg_1568[10], op_22_V_reg_1568[10], op_22_V_reg_1568[10], op_22_V_reg_1568[10], op_22_V_reg_1568, 4'h0 };
assign grp_fu_935_p1 = { op_13_V_reg_1563[7], op_13_V_reg_1563[7], op_13_V_reg_1563[7], op_13_V_reg_1563[7], op_13_V_reg_1563[7], op_13_V_reg_1563[7], op_13_V_reg_1563[7], op_13_V_reg_1563[7], op_13_V_reg_1563[7], op_13_V_reg_1563[7], op_13_V_reg_1563[7], op_13_V_reg_1563[7], op_13_V_reg_1563[7], op_13_V_reg_1563[7], op_13_V_reg_1563[7], op_13_V_reg_1563[7], op_13_V_reg_1563[7], op_13_V_reg_1563[7], op_13_V_reg_1563[7], op_13_V_reg_1563[7], op_13_V_reg_1563[7], op_13_V_reg_1563[7], op_13_V_reg_1563[7], op_13_V_reg_1563[7], op_13_V_reg_1563[7], op_13_V_reg_1563[7], op_13_V_reg_1563[7], op_13_V_reg_1563[7], op_13_V_reg_1563[7], op_13_V_reg_1563 };
assign grp_fu_984_p1 = { op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14 };
assign lhs_V_fu_390_p3 = { xor_ln1499_fu_384_p2, 1'h0 };
assign lhs_fu_275_p1 = op_4;
assign lhs_fu_275_p3 = { op_4, 1'h0 };
assign op_29 = grp_fu_1151_p2;
assign op_7_V_fu_413_p4 = { tmp_reg_1184, or_ln1195_reg_1286, 14'h0000 };
assign or_ln1195_fu_398_p1 = op_4;
assign p_Result_11_fu_814_p4 = { p_Result_19_reg_1441, p_Val2_9_fu_809_p2[6:0] };
assign p_Result_12_fu_860_p3 = ret_V_26_reg_1470[5];
assign p_Result_13_fu_961_p3 = ret_V_28_reg_1593[36];
assign p_Result_14_fu_1035_p3 = ret_V_30_reg_1640[37];
assign p_Result_15_fu_1129_p3 = ret_V_32_reg_1687[35];
assign p_Result_18_fu_506_p3 = ret_V_25_reg_1244[3];
assign p_Result_1_fu_365_p3 = r_V_reg_1189[5];
assign p_Result_3_fu_772_p3 = ret_V_24_reg_1424[11];
assign p_Result_7_fu_545_p4 = { ret_V_25_reg_1244[3], p_Val2_6_fu_539_p2 };
assign p_Result_s_fu_443_p3 = ret_V_20_reg_1222[4];
assign p_Val2_5_fu_499_p3 = { trunc_ln731_reg_1258, 1'h0 };
assign rhs_1_fu_635_p3 = { ret_V_21_reg_1329, 2'h0 };
assign rhs_5_fu_993_p3 = { op_24_V_reg_1620, 5'h00 };
assign rhs_7_fu_1067_p3 = { op_26_V_reg_1667, 3'h0 };
assign sext_ln1192_fu_642_p1 = { ret_V_21_reg_1329[2], ret_V_21_reg_1329[2], ret_V_21_reg_1329[2], ret_V_21_reg_1329[2], ret_V_21_reg_1329[2], ret_V_21_reg_1329, 2'h0 };
assign sext_ln1193_fu_286_p0 = op_5;
assign sext_ln1193_fu_286_p1 = { op_5[3], op_5 };
assign sext_ln69_2_fu_1117_p1 = { ret_V_21_reg_1329[2], ret_V_21_reg_1329[2], ret_V_21_reg_1329[2], ret_V_21_reg_1329[2], ret_V_21_reg_1329[2], ret_V_21_reg_1329 };
assign sext_ln703_1_fu_632_p0 = op_5;
assign sext_ln703_3_fu_989_p0 = op_15;
assign sext_ln703_4_fu_1063_p0 = op_17;
assign sext_ln850_fu_749_p1 = { tmp_3_reg_1475[2], tmp_3_reg_1475 };
assign tmp_13_fu_791_p3 = r_V_1_reg_1436[18];
assign tmp_16_fu_924_p3 = { op_22_V_reg_1568, 4'h0 };
assign tmp_7_fu_513_p3 = ret_V_25_reg_1244[3];
assign tmp_8_fu_520_p3 = ret_V_25_reg_1244[2];
assign tmp_fu_253_p1 = op_4;
assign trunc_ln731_fu_333_p1 = grp_fu_305_p2[2:0];
assign trunc_ln851_1_fu_271_p1 = grp_fu_237_p2[2:0];
assign trunc_ln851_2_fu_243_p0 = op_5;
assign trunc_ln851_2_fu_243_p1 = op_5[1:0];
assign trunc_ln851_3_fu_628_p1 = op_11_V_fu_623_p3[2:0];
assign trunc_ln851_4_fu_917_p1 = op_13_V_fu_912_p3[3:0];
assign trunc_ln851_5_fu_1010_p0 = op_15;
assign trunc_ln851_5_fu_1010_p1 = op_15[4:0];
assign trunc_ln851_6_fu_1084_p0 = op_17;
assign trunc_ln851_6_fu_1084_p1 = op_17[2:0];
assign trunc_ln851_fu_321_p1 = grp_fu_289_p2[1:0];
assign \sub_5s_5s_5_2_1_U2.top_sub_5s_5s_5_2_1_Adder_0_U.ain_s0  = \sub_5s_5s_5_2_1_U2.top_sub_5s_5s_5_2_1_Adder_0_U.a ;
assign \sub_5s_5s_5_2_1_U2.top_sub_5s_5s_5_2_1_Adder_0_U.s  = { \sub_5s_5s_5_2_1_U2.top_sub_5s_5s_5_2_1_Adder_0_U.fas_s2 , \sub_5s_5s_5_2_1_U2.top_sub_5s_5s_5_2_1_Adder_0_U.sum_s1  };
assign \sub_5s_5s_5_2_1_U2.top_sub_5s_5s_5_2_1_Adder_0_U.u2.a  = \sub_5s_5s_5_2_1_U2.top_sub_5s_5s_5_2_1_Adder_0_U.ain_s1 ;
assign \sub_5s_5s_5_2_1_U2.top_sub_5s_5s_5_2_1_Adder_0_U.u2.b  = \sub_5s_5s_5_2_1_U2.top_sub_5s_5s_5_2_1_Adder_0_U.bin_s1 ;
assign \sub_5s_5s_5_2_1_U2.top_sub_5s_5s_5_2_1_Adder_0_U.u2.cin  = \sub_5s_5s_5_2_1_U2.top_sub_5s_5s_5_2_1_Adder_0_U.carry_s1 ;
assign \sub_5s_5s_5_2_1_U2.top_sub_5s_5s_5_2_1_Adder_0_U.facout_s2  = \sub_5s_5s_5_2_1_U2.top_sub_5s_5s_5_2_1_Adder_0_U.u2.cout ;
assign \sub_5s_5s_5_2_1_U2.top_sub_5s_5s_5_2_1_Adder_0_U.fas_s2  = \sub_5s_5s_5_2_1_U2.top_sub_5s_5s_5_2_1_Adder_0_U.u2.s ;
assign \sub_5s_5s_5_2_1_U2.top_sub_5s_5s_5_2_1_Adder_0_U.u1.a  = \sub_5s_5s_5_2_1_U2.top_sub_5s_5s_5_2_1_Adder_0_U.a [1:0];
assign \sub_5s_5s_5_2_1_U2.top_sub_5s_5s_5_2_1_Adder_0_U.u1.b  = \sub_5s_5s_5_2_1_U2.top_sub_5s_5s_5_2_1_Adder_0_U.bin_s0 [1:0];
assign \sub_5s_5s_5_2_1_U2.top_sub_5s_5s_5_2_1_Adder_0_U.u1.cin  = 1'h1;
assign \sub_5s_5s_5_2_1_U2.top_sub_5s_5s_5_2_1_Adder_0_U.facout_s1  = \sub_5s_5s_5_2_1_U2.top_sub_5s_5s_5_2_1_Adder_0_U.u1.cout ;
assign \sub_5s_5s_5_2_1_U2.top_sub_5s_5s_5_2_1_Adder_0_U.fas_s1  = \sub_5s_5s_5_2_1_U2.top_sub_5s_5s_5_2_1_Adder_0_U.u1.s ;
assign \sub_5s_5s_5_2_1_U2.top_sub_5s_5s_5_2_1_Adder_0_U.a  = \sub_5s_5s_5_2_1_U2.din0 ;
assign \sub_5s_5s_5_2_1_U2.top_sub_5s_5s_5_2_1_Adder_0_U.b  = \sub_5s_5s_5_2_1_U2.din1 ;
assign \sub_5s_5s_5_2_1_U2.top_sub_5s_5s_5_2_1_Adder_0_U.ce  = \sub_5s_5s_5_2_1_U2.ce ;
assign \sub_5s_5s_5_2_1_U2.top_sub_5s_5s_5_2_1_Adder_0_U.clk  = \sub_5s_5s_5_2_1_U2.clk ;
assign \sub_5s_5s_5_2_1_U2.top_sub_5s_5s_5_2_1_Adder_0_U.reset  = \sub_5s_5s_5_2_1_U2.reset ;
assign \sub_5s_5s_5_2_1_U2.dout  = \sub_5s_5s_5_2_1_U2.top_sub_5s_5s_5_2_1_Adder_0_U.s ;
assign \sub_5s_5s_5_2_1_U2.ce  = 1'h1;
assign \sub_5s_5s_5_2_1_U2.clk  = ap_clk;
assign \sub_5s_5s_5_2_1_U2.din0  = { op_4[1], op_4[1], op_4, 1'h0 };
assign \sub_5s_5s_5_2_1_U2.din1  = { op_5[3], op_5 };
assign grp_fu_289_p2 = \sub_5s_5s_5_2_1_U2.dout ;
assign \sub_5s_5s_5_2_1_U2.reset  = ap_rst;
assign \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.ain_s0  = \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.a ;
assign \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.s  = { \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.fas_s2 , \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.sum_s1  };
assign \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.u2.a  = \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.ain_s1 ;
assign \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.u2.b  = \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.bin_s1 ;
assign \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.u2.cin  = \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.carry_s1 ;
assign \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.facout_s2  = \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.u2.cout ;
assign \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.fas_s2  = \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.u2.s ;
assign \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.u1.a  = \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.a [1:0];
assign \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.u1.b  = \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.bin_s0 [1:0];
assign \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.u1.cin  = 1'h1;
assign \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.facout_s1  = \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.u1.cout ;
assign \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.fas_s1  = \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.u1.s ;
assign \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.a  = \sub_5ns_5s_5_2_1_U4.din0 ;
assign \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.b  = \sub_5ns_5s_5_2_1_U4.din1 ;
assign \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.ce  = \sub_5ns_5s_5_2_1_U4.ce ;
assign \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.clk  = \sub_5ns_5s_5_2_1_U4.clk ;
assign \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.reset  = \sub_5ns_5s_5_2_1_U4.reset ;
assign \sub_5ns_5s_5_2_1_U4.dout  = \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.s ;
assign \sub_5ns_5s_5_2_1_U4.ce  = 1'h1;
assign \sub_5ns_5s_5_2_1_U4.clk  = ap_clk;
assign \sub_5ns_5s_5_2_1_U4.din0  = 5'h00;
assign \sub_5ns_5s_5_2_1_U4.din1  = { op_5[3], op_5 };
assign grp_fu_305_p2 = \sub_5ns_5s_5_2_1_U4.dout ;
assign \sub_5ns_5s_5_2_1_U4.reset  = ap_rst;
assign \shl_20s_2ns_20_7_1_U6.din1_cast  = \shl_20s_2ns_20_7_1_U6.din1 [1:0];
assign \shl_20s_2ns_20_7_1_U6.din1_mask  = 2'h1;
assign \shl_20s_2ns_20_7_1_U6.ce  = 1'h1;
assign \shl_20s_2ns_20_7_1_U6.clk  = ap_clk;
assign \shl_20s_2ns_20_7_1_U6.din0  = { tmp_reg_1184, tmp_reg_1184, tmp_reg_1184, tmp_reg_1184, or_ln1195_reg_1286, 14'h0000 };
assign \shl_20s_2ns_20_7_1_U6.din1  = { 18'h00000, ret_V_22_reg_1281 };
assign grp_fu_437_p2 = \shl_20s_2ns_20_7_1_U6.dout ;
assign \shl_20s_2ns_20_7_1_U6.reset  = ap_rst;
assign \mul_4s_2s_6_7_1_U1.top_mul_4s_2s_6_7_1_Mul_DSP_0_U.p  = \mul_4s_2s_6_7_1_U1.top_mul_4s_2s_6_7_1_Mul_DSP_0_U.buff4 ;
assign \mul_4s_2s_6_7_1_U1.top_mul_4s_2s_6_7_1_Mul_DSP_0_U.a  = \mul_4s_2s_6_7_1_U1.din0 ;
assign \mul_4s_2s_6_7_1_U1.top_mul_4s_2s_6_7_1_Mul_DSP_0_U.b  = \mul_4s_2s_6_7_1_U1.din1 ;
assign \mul_4s_2s_6_7_1_U1.top_mul_4s_2s_6_7_1_Mul_DSP_0_U.ce  = \mul_4s_2s_6_7_1_U1.ce ;
assign \mul_4s_2s_6_7_1_U1.top_mul_4s_2s_6_7_1_Mul_DSP_0_U.clk  = \mul_4s_2s_6_7_1_U1.clk ;
assign \mul_4s_2s_6_7_1_U1.dout  = \mul_4s_2s_6_7_1_U1.top_mul_4s_2s_6_7_1_Mul_DSP_0_U.p ;
assign \mul_4s_2s_6_7_1_U1.ce  = 1'h1;
assign \mul_4s_2s_6_7_1_U1.clk  = ap_clk;
assign \mul_4s_2s_6_7_1_U1.din0  = op_5;
assign \mul_4s_2s_6_7_1_U1.din1  = op_4;
assign grp_fu_237_p2 = \mul_4s_2s_6_7_1_U1.dout ;
assign \mul_4s_2s_6_7_1_U1.reset  = ap_rst;
assign \add_9ns_9ns_9_2_1_U21.top_add_9ns_9ns_9_2_1_Adder_15_U.ain_s0  = \add_9ns_9ns_9_2_1_U21.top_add_9ns_9ns_9_2_1_Adder_15_U.a ;
assign \add_9ns_9ns_9_2_1_U21.top_add_9ns_9ns_9_2_1_Adder_15_U.bin_s0  = \add_9ns_9ns_9_2_1_U21.top_add_9ns_9ns_9_2_1_Adder_15_U.b ;
assign \add_9ns_9ns_9_2_1_U21.top_add_9ns_9ns_9_2_1_Adder_15_U.s  = { \add_9ns_9ns_9_2_1_U21.top_add_9ns_9ns_9_2_1_Adder_15_U.fas_s2 , \add_9ns_9ns_9_2_1_U21.top_add_9ns_9ns_9_2_1_Adder_15_U.sum_s1  };
assign \add_9ns_9ns_9_2_1_U21.top_add_9ns_9ns_9_2_1_Adder_15_U.u2.a  = \add_9ns_9ns_9_2_1_U21.top_add_9ns_9ns_9_2_1_Adder_15_U.ain_s1 ;
assign \add_9ns_9ns_9_2_1_U21.top_add_9ns_9ns_9_2_1_Adder_15_U.u2.b  = \add_9ns_9ns_9_2_1_U21.top_add_9ns_9ns_9_2_1_Adder_15_U.bin_s1 ;
assign \add_9ns_9ns_9_2_1_U21.top_add_9ns_9ns_9_2_1_Adder_15_U.u2.cin  = \add_9ns_9ns_9_2_1_U21.top_add_9ns_9ns_9_2_1_Adder_15_U.carry_s1 ;
assign \add_9ns_9ns_9_2_1_U21.top_add_9ns_9ns_9_2_1_Adder_15_U.facout_s2  = \add_9ns_9ns_9_2_1_U21.top_add_9ns_9ns_9_2_1_Adder_15_U.u2.cout ;
assign \add_9ns_9ns_9_2_1_U21.top_add_9ns_9ns_9_2_1_Adder_15_U.fas_s2  = \add_9ns_9ns_9_2_1_U21.top_add_9ns_9ns_9_2_1_Adder_15_U.u2.s ;
assign \add_9ns_9ns_9_2_1_U21.top_add_9ns_9ns_9_2_1_Adder_15_U.u1.a  = \add_9ns_9ns_9_2_1_U21.top_add_9ns_9ns_9_2_1_Adder_15_U.a [3:0];
assign \add_9ns_9ns_9_2_1_U21.top_add_9ns_9ns_9_2_1_Adder_15_U.u1.b  = \add_9ns_9ns_9_2_1_U21.top_add_9ns_9ns_9_2_1_Adder_15_U.b [3:0];
assign \add_9ns_9ns_9_2_1_U21.top_add_9ns_9ns_9_2_1_Adder_15_U.u1.cin  = 1'h0;
assign \add_9ns_9ns_9_2_1_U21.top_add_9ns_9ns_9_2_1_Adder_15_U.facout_s1  = \add_9ns_9ns_9_2_1_U21.top_add_9ns_9ns_9_2_1_Adder_15_U.u1.cout ;
assign \add_9ns_9ns_9_2_1_U21.top_add_9ns_9ns_9_2_1_Adder_15_U.fas_s1  = \add_9ns_9ns_9_2_1_U21.top_add_9ns_9ns_9_2_1_Adder_15_U.u1.s ;
assign \add_9ns_9ns_9_2_1_U21.top_add_9ns_9ns_9_2_1_Adder_15_U.a  = \add_9ns_9ns_9_2_1_U21.din0 ;
assign \add_9ns_9ns_9_2_1_U21.top_add_9ns_9ns_9_2_1_Adder_15_U.b  = \add_9ns_9ns_9_2_1_U21.din1 ;
assign \add_9ns_9ns_9_2_1_U21.top_add_9ns_9ns_9_2_1_Adder_15_U.ce  = \add_9ns_9ns_9_2_1_U21.ce ;
assign \add_9ns_9ns_9_2_1_U21.top_add_9ns_9ns_9_2_1_Adder_15_U.clk  = \add_9ns_9ns_9_2_1_U21.clk ;
assign \add_9ns_9ns_9_2_1_U21.top_add_9ns_9ns_9_2_1_Adder_15_U.reset  = \add_9ns_9ns_9_2_1_U21.reset ;
assign \add_9ns_9ns_9_2_1_U21.dout  = \add_9ns_9ns_9_2_1_U21.top_add_9ns_9ns_9_2_1_Adder_15_U.s ;
assign \add_9ns_9ns_9_2_1_U21.ce  = 1'h1;
assign \add_9ns_9ns_9_2_1_U21.clk  = ap_clk;
assign \add_9ns_9ns_9_2_1_U21.din0  = { 1'h0, ret_V_21_reg_1329[2], ret_V_21_reg_1329[2], ret_V_21_reg_1329[2], ret_V_21_reg_1329[2], ret_V_21_reg_1329[2], ret_V_21_reg_1329 };
assign \add_9ns_9ns_9_2_1_U21.din1  = select_ln69_reg_1699;
assign grp_fu_1124_p2 = \add_9ns_9ns_9_2_1_U21.dout ;
assign \add_9ns_9ns_9_2_1_U21.reset  = ap_rst;
assign \add_6ns_6s_6_2_1_U9.top_add_6ns_6s_6_2_1_Adder_6_U.ain_s0  = \add_6ns_6s_6_2_1_U9.top_add_6ns_6s_6_2_1_Adder_6_U.a ;
assign \add_6ns_6s_6_2_1_U9.top_add_6ns_6s_6_2_1_Adder_6_U.bin_s0  = \add_6ns_6s_6_2_1_U9.top_add_6ns_6s_6_2_1_Adder_6_U.b ;
assign \add_6ns_6s_6_2_1_U9.top_add_6ns_6s_6_2_1_Adder_6_U.s  = { \add_6ns_6s_6_2_1_U9.top_add_6ns_6s_6_2_1_Adder_6_U.fas_s2 , \add_6ns_6s_6_2_1_U9.top_add_6ns_6s_6_2_1_Adder_6_U.sum_s1  };
assign \add_6ns_6s_6_2_1_U9.top_add_6ns_6s_6_2_1_Adder_6_U.u2.a  = \add_6ns_6s_6_2_1_U9.top_add_6ns_6s_6_2_1_Adder_6_U.ain_s1 ;
assign \add_6ns_6s_6_2_1_U9.top_add_6ns_6s_6_2_1_Adder_6_U.u2.b  = \add_6ns_6s_6_2_1_U9.top_add_6ns_6s_6_2_1_Adder_6_U.bin_s1 ;
assign \add_6ns_6s_6_2_1_U9.top_add_6ns_6s_6_2_1_Adder_6_U.u2.cin  = \add_6ns_6s_6_2_1_U9.top_add_6ns_6s_6_2_1_Adder_6_U.carry_s1 ;
assign \add_6ns_6s_6_2_1_U9.top_add_6ns_6s_6_2_1_Adder_6_U.facout_s2  = \add_6ns_6s_6_2_1_U9.top_add_6ns_6s_6_2_1_Adder_6_U.u2.cout ;
assign \add_6ns_6s_6_2_1_U9.top_add_6ns_6s_6_2_1_Adder_6_U.fas_s2  = \add_6ns_6s_6_2_1_U9.top_add_6ns_6s_6_2_1_Adder_6_U.u2.s ;
assign \add_6ns_6s_6_2_1_U9.top_add_6ns_6s_6_2_1_Adder_6_U.u1.a  = \add_6ns_6s_6_2_1_U9.top_add_6ns_6s_6_2_1_Adder_6_U.a [2:0];
assign \add_6ns_6s_6_2_1_U9.top_add_6ns_6s_6_2_1_Adder_6_U.u1.b  = \add_6ns_6s_6_2_1_U9.top_add_6ns_6s_6_2_1_Adder_6_U.b [2:0];
assign \add_6ns_6s_6_2_1_U9.top_add_6ns_6s_6_2_1_Adder_6_U.u1.cin  = 1'h0;
assign \add_6ns_6s_6_2_1_U9.top_add_6ns_6s_6_2_1_Adder_6_U.facout_s1  = \add_6ns_6s_6_2_1_U9.top_add_6ns_6s_6_2_1_Adder_6_U.u1.cout ;
assign \add_6ns_6s_6_2_1_U9.top_add_6ns_6s_6_2_1_Adder_6_U.fas_s1  = \add_6ns_6s_6_2_1_U9.top_add_6ns_6s_6_2_1_Adder_6_U.u1.s ;
assign \add_6ns_6s_6_2_1_U9.top_add_6ns_6s_6_2_1_Adder_6_U.a  = \add_6ns_6s_6_2_1_U9.din0 ;
assign \add_6ns_6s_6_2_1_U9.top_add_6ns_6s_6_2_1_Adder_6_U.b  = \add_6ns_6s_6_2_1_U9.din1 ;
assign \add_6ns_6s_6_2_1_U9.top_add_6ns_6s_6_2_1_Adder_6_U.ce  = \add_6ns_6s_6_2_1_U9.ce ;
assign \add_6ns_6s_6_2_1_U9.top_add_6ns_6s_6_2_1_Adder_6_U.clk  = \add_6ns_6s_6_2_1_U9.clk ;
assign \add_6ns_6s_6_2_1_U9.top_add_6ns_6s_6_2_1_Adder_6_U.reset  = \add_6ns_6s_6_2_1_U9.reset ;
assign \add_6ns_6s_6_2_1_U9.dout  = \add_6ns_6s_6_2_1_U9.top_add_6ns_6s_6_2_1_Adder_6_U.s ;
assign \add_6ns_6s_6_2_1_U9.ce  = 1'h1;
assign \add_6ns_6s_6_2_1_U9.clk  = ap_clk;
assign \add_6ns_6s_6_2_1_U9.din0  = { ret_V_23_reg_1384, 3'h0 };
assign \add_6ns_6s_6_2_1_U9.din1  = { op_11_V_reg_1389[3], op_11_V_reg_1389[3], op_11_V_reg_1389 };
assign grp_fu_666_p2 = \add_6ns_6s_6_2_1_U9.dout ;
assign \add_6ns_6s_6_2_1_U9.reset  = ap_rst;
assign \add_4s_4ns_4_2_1_U11.top_add_4s_4ns_4_2_1_Adder_8_U.ain_s0  = \add_4s_4ns_4_2_1_U11.top_add_4s_4ns_4_2_1_Adder_8_U.a ;
assign \add_4s_4ns_4_2_1_U11.top_add_4s_4ns_4_2_1_Adder_8_U.bin_s0  = \add_4s_4ns_4_2_1_U11.top_add_4s_4ns_4_2_1_Adder_8_U.b ;
assign \add_4s_4ns_4_2_1_U11.top_add_4s_4ns_4_2_1_Adder_8_U.s  = { \add_4s_4ns_4_2_1_U11.top_add_4s_4ns_4_2_1_Adder_8_U.fas_s2 , \add_4s_4ns_4_2_1_U11.top_add_4s_4ns_4_2_1_Adder_8_U.sum_s1  };
assign \add_4s_4ns_4_2_1_U11.top_add_4s_4ns_4_2_1_Adder_8_U.u2.a  = \add_4s_4ns_4_2_1_U11.top_add_4s_4ns_4_2_1_Adder_8_U.ain_s1 ;
assign \add_4s_4ns_4_2_1_U11.top_add_4s_4ns_4_2_1_Adder_8_U.u2.b  = \add_4s_4ns_4_2_1_U11.top_add_4s_4ns_4_2_1_Adder_8_U.bin_s1 ;
assign \add_4s_4ns_4_2_1_U11.top_add_4s_4ns_4_2_1_Adder_8_U.u2.cin  = \add_4s_4ns_4_2_1_U11.top_add_4s_4ns_4_2_1_Adder_8_U.carry_s1 ;
assign \add_4s_4ns_4_2_1_U11.top_add_4s_4ns_4_2_1_Adder_8_U.facout_s2  = \add_4s_4ns_4_2_1_U11.top_add_4s_4ns_4_2_1_Adder_8_U.u2.cout ;
assign \add_4s_4ns_4_2_1_U11.top_add_4s_4ns_4_2_1_Adder_8_U.fas_s2  = \add_4s_4ns_4_2_1_U11.top_add_4s_4ns_4_2_1_Adder_8_U.u2.s ;
assign \add_4s_4ns_4_2_1_U11.top_add_4s_4ns_4_2_1_Adder_8_U.u1.a  = \add_4s_4ns_4_2_1_U11.top_add_4s_4ns_4_2_1_Adder_8_U.a [1:0];
assign \add_4s_4ns_4_2_1_U11.top_add_4s_4ns_4_2_1_Adder_8_U.u1.b  = \add_4s_4ns_4_2_1_U11.top_add_4s_4ns_4_2_1_Adder_8_U.b [1:0];
assign \add_4s_4ns_4_2_1_U11.top_add_4s_4ns_4_2_1_Adder_8_U.u1.cin  = 1'h0;
assign \add_4s_4ns_4_2_1_U11.top_add_4s_4ns_4_2_1_Adder_8_U.facout_s1  = \add_4s_4ns_4_2_1_U11.top_add_4s_4ns_4_2_1_Adder_8_U.u1.cout ;
assign \add_4s_4ns_4_2_1_U11.top_add_4s_4ns_4_2_1_Adder_8_U.fas_s1  = \add_4s_4ns_4_2_1_U11.top_add_4s_4ns_4_2_1_Adder_8_U.u1.s ;
assign \add_4s_4ns_4_2_1_U11.top_add_4s_4ns_4_2_1_Adder_8_U.a  = \add_4s_4ns_4_2_1_U11.din0 ;
assign \add_4s_4ns_4_2_1_U11.top_add_4s_4ns_4_2_1_Adder_8_U.b  = \add_4s_4ns_4_2_1_U11.din1 ;
assign \add_4s_4ns_4_2_1_U11.top_add_4s_4ns_4_2_1_Adder_8_U.ce  = \add_4s_4ns_4_2_1_U11.ce ;
assign \add_4s_4ns_4_2_1_U11.top_add_4s_4ns_4_2_1_Adder_8_U.clk  = \add_4s_4ns_4_2_1_U11.clk ;
assign \add_4s_4ns_4_2_1_U11.top_add_4s_4ns_4_2_1_Adder_8_U.reset  = \add_4s_4ns_4_2_1_U11.reset ;
assign \add_4s_4ns_4_2_1_U11.dout  = \add_4s_4ns_4_2_1_U11.top_add_4s_4ns_4_2_1_Adder_8_U.s ;
assign \add_4s_4ns_4_2_1_U11.ce  = 1'h1;
assign \add_4s_4ns_4_2_1_U11.clk  = ap_clk;
assign \add_4s_4ns_4_2_1_U11.din0  = { tmp_3_reg_1475[2], tmp_3_reg_1475 };
assign \add_4s_4ns_4_2_1_U11.din1  = 4'h1;
assign grp_fu_752_p2 = \add_4s_4ns_4_2_1_U11.dout ;
assign \add_4s_4ns_4_2_1_U11.reset  = ap_rst;
assign \add_3s_3ns_3_2_1_U7.top_add_3s_3ns_3_2_1_Adder_4_U.ain_s0  = \add_3s_3ns_3_2_1_U7.top_add_3s_3ns_3_2_1_Adder_4_U.a ;
assign \add_3s_3ns_3_2_1_U7.top_add_3s_3ns_3_2_1_Adder_4_U.bin_s0  = \add_3s_3ns_3_2_1_U7.top_add_3s_3ns_3_2_1_Adder_4_U.b ;
assign \add_3s_3ns_3_2_1_U7.top_add_3s_3ns_3_2_1_Adder_4_U.s  = { \add_3s_3ns_3_2_1_U7.top_add_3s_3ns_3_2_1_Adder_4_U.fas_s2 , \add_3s_3ns_3_2_1_U7.top_add_3s_3ns_3_2_1_Adder_4_U.sum_s1  };
assign \add_3s_3ns_3_2_1_U7.top_add_3s_3ns_3_2_1_Adder_4_U.u2.a  = \add_3s_3ns_3_2_1_U7.top_add_3s_3ns_3_2_1_Adder_4_U.ain_s1 ;
assign \add_3s_3ns_3_2_1_U7.top_add_3s_3ns_3_2_1_Adder_4_U.u2.b  = \add_3s_3ns_3_2_1_U7.top_add_3s_3ns_3_2_1_Adder_4_U.bin_s1 ;
assign \add_3s_3ns_3_2_1_U7.top_add_3s_3ns_3_2_1_Adder_4_U.u2.cin  = \add_3s_3ns_3_2_1_U7.top_add_3s_3ns_3_2_1_Adder_4_U.carry_s1 ;
assign \add_3s_3ns_3_2_1_U7.top_add_3s_3ns_3_2_1_Adder_4_U.facout_s2  = \add_3s_3ns_3_2_1_U7.top_add_3s_3ns_3_2_1_Adder_4_U.u2.cout ;
assign \add_3s_3ns_3_2_1_U7.top_add_3s_3ns_3_2_1_Adder_4_U.fas_s2  = \add_3s_3ns_3_2_1_U7.top_add_3s_3ns_3_2_1_Adder_4_U.u2.s ;
assign \add_3s_3ns_3_2_1_U7.top_add_3s_3ns_3_2_1_Adder_4_U.u1.a  = \add_3s_3ns_3_2_1_U7.top_add_3s_3ns_3_2_1_Adder_4_U.a [0];
assign \add_3s_3ns_3_2_1_U7.top_add_3s_3ns_3_2_1_Adder_4_U.u1.b  = \add_3s_3ns_3_2_1_U7.top_add_3s_3ns_3_2_1_Adder_4_U.b [0];
assign \add_3s_3ns_3_2_1_U7.top_add_3s_3ns_3_2_1_Adder_4_U.u1.cin  = 1'h0;
assign \add_3s_3ns_3_2_1_U7.top_add_3s_3ns_3_2_1_Adder_4_U.facout_s1  = \add_3s_3ns_3_2_1_U7.top_add_3s_3ns_3_2_1_Adder_4_U.u1.cout ;
assign \add_3s_3ns_3_2_1_U7.top_add_3s_3ns_3_2_1_Adder_4_U.fas_s1  = \add_3s_3ns_3_2_1_U7.top_add_3s_3ns_3_2_1_Adder_4_U.u1.s ;
assign \add_3s_3ns_3_2_1_U7.top_add_3s_3ns_3_2_1_Adder_4_U.a  = \add_3s_3ns_3_2_1_U7.din0 ;
assign \add_3s_3ns_3_2_1_U7.top_add_3s_3ns_3_2_1_Adder_4_U.b  = \add_3s_3ns_3_2_1_U7.din1 ;
assign \add_3s_3ns_3_2_1_U7.top_add_3s_3ns_3_2_1_Adder_4_U.ce  = \add_3s_3ns_3_2_1_U7.ce ;
assign \add_3s_3ns_3_2_1_U7.top_add_3s_3ns_3_2_1_Adder_4_U.clk  = \add_3s_3ns_3_2_1_U7.clk ;
assign \add_3s_3ns_3_2_1_U7.top_add_3s_3ns_3_2_1_Adder_4_U.reset  = \add_3s_3ns_3_2_1_U7.reset ;
assign \add_3s_3ns_3_2_1_U7.dout  = \add_3s_3ns_3_2_1_U7.top_add_3s_3ns_3_2_1_Adder_4_U.s ;
assign \add_3s_3ns_3_2_1_U7.ce  = 1'h1;
assign \add_3s_3ns_3_2_1_U7.clk  = ap_clk;
assign \add_3s_3ns_3_2_1_U7.din0  = { op_6[1], op_6 };
assign \add_3s_3ns_3_2_1_U7.din1  = select_ln703_reg_1353;
assign grp_fu_597_p2 = \add_3s_3ns_3_2_1_U7.dout ;
assign \add_3s_3ns_3_2_1_U7.reset  = ap_rst;
assign \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_3_U.ain_s0  = \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_3_U.a ;
assign \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_3_U.bin_s0  = \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_3_U.b ;
assign \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_3_U.s  = { \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_3_U.fas_s2 , \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_3_U.sum_s1  };
assign \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_3_U.u2.a  = \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_3_U.ain_s1 ;
assign \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_3_U.u2.b  = \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_3_U.bin_s1 ;
assign \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_3_U.u2.cin  = \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_3_U.carry_s1 ;
assign \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_3_U.facout_s2  = \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_3_U.u2.cout ;
assign \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_3_U.fas_s2  = \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_3_U.u2.s ;
assign \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_3_U.u1.a  = \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_3_U.a [0];
assign \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_3_U.u1.b  = \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_3_U.b [0];
assign \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_3_U.u1.cin  = 1'h0;
assign \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_3_U.facout_s1  = \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_3_U.u1.cout ;
assign \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_3_U.fas_s1  = \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_3_U.u1.s ;
assign \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_3_U.a  = \add_3ns_3ns_3_2_1_U5.din0 ;
assign \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_3_U.b  = \add_3ns_3ns_3_2_1_U5.din1 ;
assign \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_3_U.ce  = \add_3ns_3ns_3_2_1_U5.ce ;
assign \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_3_U.clk  = \add_3ns_3ns_3_2_1_U5.clk ;
assign \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_3_U.reset  = \add_3ns_3ns_3_2_1_U5.reset ;
assign \add_3ns_3ns_3_2_1_U5.dout  = \add_3ns_3ns_3_2_1_U5.top_add_3ns_3ns_3_2_1_Adder_3_U.s ;
assign \add_3ns_3ns_3_2_1_U5.ce  = 1'h1;
assign \add_3ns_3ns_3_2_1_U5.clk  = ap_clk;
assign \add_3ns_3ns_3_2_1_U5.din0  = ret_V_reg_1227;
assign \add_3ns_3ns_3_2_1_U5.din1  = 3'h1;
assign grp_fu_360_p2 = \add_3ns_3ns_3_2_1_U5.dout ;
assign \add_3ns_3ns_3_2_1_U5.reset  = ap_rst;
assign \add_38s_38s_38_2_1_U16.top_add_38s_38s_38_2_1_Adder_13_U.ain_s0  = \add_38s_38s_38_2_1_U16.top_add_38s_38s_38_2_1_Adder_13_U.a ;
assign \add_38s_38s_38_2_1_U16.top_add_38s_38s_38_2_1_Adder_13_U.bin_s0  = \add_38s_38s_38_2_1_U16.top_add_38s_38s_38_2_1_Adder_13_U.b ;
assign \add_38s_38s_38_2_1_U16.top_add_38s_38s_38_2_1_Adder_13_U.s  = { \add_38s_38s_38_2_1_U16.top_add_38s_38s_38_2_1_Adder_13_U.fas_s2 , \add_38s_38s_38_2_1_U16.top_add_38s_38s_38_2_1_Adder_13_U.sum_s1  };
assign \add_38s_38s_38_2_1_U16.top_add_38s_38s_38_2_1_Adder_13_U.u2.a  = \add_38s_38s_38_2_1_U16.top_add_38s_38s_38_2_1_Adder_13_U.ain_s1 ;
assign \add_38s_38s_38_2_1_U16.top_add_38s_38s_38_2_1_Adder_13_U.u2.b  = \add_38s_38s_38_2_1_U16.top_add_38s_38s_38_2_1_Adder_13_U.bin_s1 ;
assign \add_38s_38s_38_2_1_U16.top_add_38s_38s_38_2_1_Adder_13_U.u2.cin  = \add_38s_38s_38_2_1_U16.top_add_38s_38s_38_2_1_Adder_13_U.carry_s1 ;
assign \add_38s_38s_38_2_1_U16.top_add_38s_38s_38_2_1_Adder_13_U.facout_s2  = \add_38s_38s_38_2_1_U16.top_add_38s_38s_38_2_1_Adder_13_U.u2.cout ;
assign \add_38s_38s_38_2_1_U16.top_add_38s_38s_38_2_1_Adder_13_U.fas_s2  = \add_38s_38s_38_2_1_U16.top_add_38s_38s_38_2_1_Adder_13_U.u2.s ;
assign \add_38s_38s_38_2_1_U16.top_add_38s_38s_38_2_1_Adder_13_U.u1.a  = \add_38s_38s_38_2_1_U16.top_add_38s_38s_38_2_1_Adder_13_U.a [18:0];
assign \add_38s_38s_38_2_1_U16.top_add_38s_38s_38_2_1_Adder_13_U.u1.b  = \add_38s_38s_38_2_1_U16.top_add_38s_38s_38_2_1_Adder_13_U.b [18:0];
assign \add_38s_38s_38_2_1_U16.top_add_38s_38s_38_2_1_Adder_13_U.u1.cin  = 1'h0;
assign \add_38s_38s_38_2_1_U16.top_add_38s_38s_38_2_1_Adder_13_U.facout_s1  = \add_38s_38s_38_2_1_U16.top_add_38s_38s_38_2_1_Adder_13_U.u1.cout ;
assign \add_38s_38s_38_2_1_U16.top_add_38s_38s_38_2_1_Adder_13_U.fas_s1  = \add_38s_38s_38_2_1_U16.top_add_38s_38s_38_2_1_Adder_13_U.u1.s ;
assign \add_38s_38s_38_2_1_U16.top_add_38s_38s_38_2_1_Adder_13_U.a  = \add_38s_38s_38_2_1_U16.din0 ;
assign \add_38s_38s_38_2_1_U16.top_add_38s_38s_38_2_1_Adder_13_U.b  = \add_38s_38s_38_2_1_U16.din1 ;
assign \add_38s_38s_38_2_1_U16.top_add_38s_38s_38_2_1_Adder_13_U.ce  = \add_38s_38s_38_2_1_U16.ce ;
assign \add_38s_38s_38_2_1_U16.top_add_38s_38s_38_2_1_Adder_13_U.clk  = \add_38s_38s_38_2_1_U16.clk ;
assign \add_38s_38s_38_2_1_U16.top_add_38s_38s_38_2_1_Adder_13_U.reset  = \add_38s_38s_38_2_1_U16.reset ;
assign \add_38s_38s_38_2_1_U16.dout  = \add_38s_38s_38_2_1_U16.top_add_38s_38s_38_2_1_Adder_13_U.s ;
assign \add_38s_38s_38_2_1_U16.ce  = 1'h1;
assign \add_38s_38s_38_2_1_U16.clk  = ap_clk;
assign \add_38s_38s_38_2_1_U16.din0  = { op_24_V_reg_1620[31], op_24_V_reg_1620, 5'h00 };
assign \add_38s_38s_38_2_1_U16.din1  = { op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15 };
assign grp_fu_1004_p2 = \add_38s_38s_38_2_1_U16.dout ;
assign \add_38s_38s_38_2_1_U16.reset  = ap_rst;
assign \add_37s_37s_37_2_1_U13.top_add_37s_37s_37_2_1_Adder_10_U.ain_s0  = \add_37s_37s_37_2_1_U13.top_add_37s_37s_37_2_1_Adder_10_U.a ;
assign \add_37s_37s_37_2_1_U13.top_add_37s_37s_37_2_1_Adder_10_U.bin_s0  = \add_37s_37s_37_2_1_U13.top_add_37s_37s_37_2_1_Adder_10_U.b ;
assign \add_37s_37s_37_2_1_U13.top_add_37s_37s_37_2_1_Adder_10_U.s  = { \add_37s_37s_37_2_1_U13.top_add_37s_37s_37_2_1_Adder_10_U.fas_s2 , \add_37s_37s_37_2_1_U13.top_add_37s_37s_37_2_1_Adder_10_U.sum_s1  };
assign \add_37s_37s_37_2_1_U13.top_add_37s_37s_37_2_1_Adder_10_U.u2.a  = \add_37s_37s_37_2_1_U13.top_add_37s_37s_37_2_1_Adder_10_U.ain_s1 ;
assign \add_37s_37s_37_2_1_U13.top_add_37s_37s_37_2_1_Adder_10_U.u2.b  = \add_37s_37s_37_2_1_U13.top_add_37s_37s_37_2_1_Adder_10_U.bin_s1 ;
assign \add_37s_37s_37_2_1_U13.top_add_37s_37s_37_2_1_Adder_10_U.u2.cin  = \add_37s_37s_37_2_1_U13.top_add_37s_37s_37_2_1_Adder_10_U.carry_s1 ;
assign \add_37s_37s_37_2_1_U13.top_add_37s_37s_37_2_1_Adder_10_U.facout_s2  = \add_37s_37s_37_2_1_U13.top_add_37s_37s_37_2_1_Adder_10_U.u2.cout ;
assign \add_37s_37s_37_2_1_U13.top_add_37s_37s_37_2_1_Adder_10_U.fas_s2  = \add_37s_37s_37_2_1_U13.top_add_37s_37s_37_2_1_Adder_10_U.u2.s ;
assign \add_37s_37s_37_2_1_U13.top_add_37s_37s_37_2_1_Adder_10_U.u1.a  = \add_37s_37s_37_2_1_U13.top_add_37s_37s_37_2_1_Adder_10_U.a [17:0];
assign \add_37s_37s_37_2_1_U13.top_add_37s_37s_37_2_1_Adder_10_U.u1.b  = \add_37s_37s_37_2_1_U13.top_add_37s_37s_37_2_1_Adder_10_U.b [17:0];
assign \add_37s_37s_37_2_1_U13.top_add_37s_37s_37_2_1_Adder_10_U.u1.cin  = 1'h0;
assign \add_37s_37s_37_2_1_U13.top_add_37s_37s_37_2_1_Adder_10_U.facout_s1  = \add_37s_37s_37_2_1_U13.top_add_37s_37s_37_2_1_Adder_10_U.u1.cout ;
assign \add_37s_37s_37_2_1_U13.top_add_37s_37s_37_2_1_Adder_10_U.fas_s1  = \add_37s_37s_37_2_1_U13.top_add_37s_37s_37_2_1_Adder_10_U.u1.s ;
assign \add_37s_37s_37_2_1_U13.top_add_37s_37s_37_2_1_Adder_10_U.a  = \add_37s_37s_37_2_1_U13.din0 ;
assign \add_37s_37s_37_2_1_U13.top_add_37s_37s_37_2_1_Adder_10_U.b  = \add_37s_37s_37_2_1_U13.din1 ;
assign \add_37s_37s_37_2_1_U13.top_add_37s_37s_37_2_1_Adder_10_U.ce  = \add_37s_37s_37_2_1_U13.ce ;
assign \add_37s_37s_37_2_1_U13.top_add_37s_37s_37_2_1_Adder_10_U.clk  = \add_37s_37s_37_2_1_U13.clk ;
assign \add_37s_37s_37_2_1_U13.top_add_37s_37s_37_2_1_Adder_10_U.reset  = \add_37s_37s_37_2_1_U13.reset ;
assign \add_37s_37s_37_2_1_U13.dout  = \add_37s_37s_37_2_1_U13.top_add_37s_37s_37_2_1_Adder_10_U.s ;
assign \add_37s_37s_37_2_1_U13.ce  = 1'h1;
assign \add_37s_37s_37_2_1_U13.clk  = ap_clk;
assign \add_37s_37s_37_2_1_U13.din0  = { op_22_V_reg_1568[10], op_22_V_reg_1568[10], op_22_V_reg_1568[10], op_22_V_reg_1568[10], op_22_V_reg_1568[10], op_22_V_reg_1568[10], op_22_V_reg_1568[10], op_22_V_reg_1568[10], op_22_V_reg_1568[10], op_22_V_reg_1568[10], op_22_V_reg_1568[10], op_22_V_reg_1568[10], op_22_V_reg_1568[10], op_22_V_reg_1568[10], op_22_V_reg_1568[10], op_22_V_reg_1568[10], op_22_V_reg_1568[10], op_22_V_reg_1568[10], op_22_V_reg_1568[10], op_22_V_reg_1568[10], op_22_V_reg_1568[10], op_22_V_reg_1568[10], op_22_V_reg_1568, 4'h0 };
assign \add_37s_37s_37_2_1_U13.din1  = { op_13_V_reg_1563[7], op_13_V_reg_1563[7], op_13_V_reg_1563[7], op_13_V_reg_1563[7], op_13_V_reg_1563[7], op_13_V_reg_1563[7], op_13_V_reg_1563[7], op_13_V_reg_1563[7], op_13_V_reg_1563[7], op_13_V_reg_1563[7], op_13_V_reg_1563[7], op_13_V_reg_1563[7], op_13_V_reg_1563[7], op_13_V_reg_1563[7], op_13_V_reg_1563[7], op_13_V_reg_1563[7], op_13_V_reg_1563[7], op_13_V_reg_1563[7], op_13_V_reg_1563[7], op_13_V_reg_1563[7], op_13_V_reg_1563[7], op_13_V_reg_1563[7], op_13_V_reg_1563[7], op_13_V_reg_1563[7], op_13_V_reg_1563[7], op_13_V_reg_1563[7], op_13_V_reg_1563[7], op_13_V_reg_1563[7], op_13_V_reg_1563[7], op_13_V_reg_1563 };
assign grp_fu_935_p2 = \add_37s_37s_37_2_1_U13.dout ;
assign \add_37s_37s_37_2_1_U13.reset  = ap_rst;
assign \add_36s_36s_36_2_1_U19.top_add_36s_36s_36_2_1_Adder_14_U.ain_s0  = \add_36s_36s_36_2_1_U19.top_add_36s_36s_36_2_1_Adder_14_U.a ;
assign \add_36s_36s_36_2_1_U19.top_add_36s_36s_36_2_1_Adder_14_U.bin_s0  = \add_36s_36s_36_2_1_U19.top_add_36s_36s_36_2_1_Adder_14_U.b ;
assign \add_36s_36s_36_2_1_U19.top_add_36s_36s_36_2_1_Adder_14_U.s  = { \add_36s_36s_36_2_1_U19.top_add_36s_36s_36_2_1_Adder_14_U.fas_s2 , \add_36s_36s_36_2_1_U19.top_add_36s_36s_36_2_1_Adder_14_U.sum_s1  };
assign \add_36s_36s_36_2_1_U19.top_add_36s_36s_36_2_1_Adder_14_U.u2.a  = \add_36s_36s_36_2_1_U19.top_add_36s_36s_36_2_1_Adder_14_U.ain_s1 ;
assign \add_36s_36s_36_2_1_U19.top_add_36s_36s_36_2_1_Adder_14_U.u2.b  = \add_36s_36s_36_2_1_U19.top_add_36s_36s_36_2_1_Adder_14_U.bin_s1 ;
assign \add_36s_36s_36_2_1_U19.top_add_36s_36s_36_2_1_Adder_14_U.u2.cin  = \add_36s_36s_36_2_1_U19.top_add_36s_36s_36_2_1_Adder_14_U.carry_s1 ;
assign \add_36s_36s_36_2_1_U19.top_add_36s_36s_36_2_1_Adder_14_U.facout_s2  = \add_36s_36s_36_2_1_U19.top_add_36s_36s_36_2_1_Adder_14_U.u2.cout ;
assign \add_36s_36s_36_2_1_U19.top_add_36s_36s_36_2_1_Adder_14_U.fas_s2  = \add_36s_36s_36_2_1_U19.top_add_36s_36s_36_2_1_Adder_14_U.u2.s ;
assign \add_36s_36s_36_2_1_U19.top_add_36s_36s_36_2_1_Adder_14_U.u1.a  = \add_36s_36s_36_2_1_U19.top_add_36s_36s_36_2_1_Adder_14_U.a [17:0];
assign \add_36s_36s_36_2_1_U19.top_add_36s_36s_36_2_1_Adder_14_U.u1.b  = \add_36s_36s_36_2_1_U19.top_add_36s_36s_36_2_1_Adder_14_U.b [17:0];
assign \add_36s_36s_36_2_1_U19.top_add_36s_36s_36_2_1_Adder_14_U.u1.cin  = 1'h0;
assign \add_36s_36s_36_2_1_U19.top_add_36s_36s_36_2_1_Adder_14_U.facout_s1  = \add_36s_36s_36_2_1_U19.top_add_36s_36s_36_2_1_Adder_14_U.u1.cout ;
assign \add_36s_36s_36_2_1_U19.top_add_36s_36s_36_2_1_Adder_14_U.fas_s1  = \add_36s_36s_36_2_1_U19.top_add_36s_36s_36_2_1_Adder_14_U.u1.s ;
assign \add_36s_36s_36_2_1_U19.top_add_36s_36s_36_2_1_Adder_14_U.a  = \add_36s_36s_36_2_1_U19.din0 ;
assign \add_36s_36s_36_2_1_U19.top_add_36s_36s_36_2_1_Adder_14_U.b  = \add_36s_36s_36_2_1_U19.din1 ;
assign \add_36s_36s_36_2_1_U19.top_add_36s_36s_36_2_1_Adder_14_U.ce  = \add_36s_36s_36_2_1_U19.ce ;
assign \add_36s_36s_36_2_1_U19.top_add_36s_36s_36_2_1_Adder_14_U.clk  = \add_36s_36s_36_2_1_U19.clk ;
assign \add_36s_36s_36_2_1_U19.top_add_36s_36s_36_2_1_Adder_14_U.reset  = \add_36s_36s_36_2_1_U19.reset ;
assign \add_36s_36s_36_2_1_U19.dout  = \add_36s_36s_36_2_1_U19.top_add_36s_36s_36_2_1_Adder_14_U.s ;
assign \add_36s_36s_36_2_1_U19.ce  = 1'h1;
assign \add_36s_36s_36_2_1_U19.clk  = ap_clk;
assign \add_36s_36s_36_2_1_U19.din0  = { op_26_V_reg_1667[31], op_26_V_reg_1667, 3'h0 };
assign \add_36s_36s_36_2_1_U19.din1  = { op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17 };
assign grp_fu_1078_p2 = \add_36s_36s_36_2_1_U19.dout ;
assign \add_36s_36s_36_2_1_U19.reset  = ap_rst;
assign \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_16_U.ain_s0  = \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_16_U.a ;
assign \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_16_U.bin_s0  = \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_16_U.b ;
assign \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_16_U.s  = { \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_16_U.fas_s2 , \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_16_U.sum_s1  };
assign \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_16_U.u2.a  = \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_16_U.ain_s1 ;
assign \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_16_U.u2.b  = \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_16_U.bin_s1 ;
assign \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_16_U.u2.cin  = \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_16_U.carry_s1 ;
assign \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_16_U.facout_s2  = \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_16_U.u2.cout ;
assign \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_16_U.fas_s2  = \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_16_U.u2.s ;
assign \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_16_U.u1.a  = \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_16_U.a [15:0];
assign \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_16_U.u1.b  = \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_16_U.b [15:0];
assign \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_16_U.u1.cin  = 1'h0;
assign \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_16_U.facout_s1  = \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_16_U.u1.cout ;
assign \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_16_U.fas_s1  = \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_16_U.u1.s ;
assign \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_16_U.a  = \add_32s_32ns_32_2_1_U22.din0 ;
assign \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_16_U.b  = \add_32s_32ns_32_2_1_U22.din1 ;
assign \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_16_U.ce  = \add_32s_32ns_32_2_1_U22.ce ;
assign \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_16_U.clk  = \add_32s_32ns_32_2_1_U22.clk ;
assign \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_16_U.reset  = \add_32s_32ns_32_2_1_U22.reset ;
assign \add_32s_32ns_32_2_1_U22.dout  = \add_32s_32ns_32_2_1_U22.top_add_32s_32ns_32_2_1_Adder_16_U.s ;
assign \add_32s_32ns_32_2_1_U22.ce  = 1'h1;
assign \add_32s_32ns_32_2_1_U22.clk  = ap_clk;
assign \add_32s_32ns_32_2_1_U22.din0  = { add_ln69_reg_1719[8], add_ln69_reg_1719[8], add_ln69_reg_1719[8], add_ln69_reg_1719[8], add_ln69_reg_1719[8], add_ln69_reg_1719[8], add_ln69_reg_1719[8], add_ln69_reg_1719[8], add_ln69_reg_1719[8], add_ln69_reg_1719[8], add_ln69_reg_1719[8], add_ln69_reg_1719[8], add_ln69_reg_1719[8], add_ln69_reg_1719[8], add_ln69_reg_1719[8], add_ln69_reg_1719[8], add_ln69_reg_1719[8], add_ln69_reg_1719[8], add_ln69_reg_1719[8], add_ln69_reg_1719[8], add_ln69_reg_1719[8], add_ln69_reg_1719[8], add_ln69_reg_1719[8], add_ln69_reg_1719 };
assign \add_32s_32ns_32_2_1_U22.din1  = ret_V_33_reg_1714;
assign grp_fu_1151_p2 = \add_32s_32ns_32_2_1_U22.dout ;
assign \add_32s_32ns_32_2_1_U22.reset  = ap_rst;
assign \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_12_U.ain_s0  = \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_12_U.a ;
assign \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_12_U.bin_s0  = \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_12_U.b ;
assign \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_12_U.s  = { \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_12_U.fas_s2 , \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_12_U.sum_s1  };
assign \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_12_U.u2.a  = \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_12_U.ain_s1 ;
assign \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_12_U.u2.b  = \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_12_U.bin_s1 ;
assign \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_12_U.u2.cin  = \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_12_U.carry_s1 ;
assign \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_12_U.facout_s2  = \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_12_U.u2.cout ;
assign \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_12_U.fas_s2  = \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_12_U.u2.s ;
assign \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_12_U.u1.a  = \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_12_U.a [15:0];
assign \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_12_U.u1.b  = \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_12_U.b [15:0];
assign \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_12_U.u1.cin  = 1'h0;
assign \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_12_U.facout_s1  = \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_12_U.u1.cout ;
assign \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_12_U.fas_s1  = \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_12_U.u1.s ;
assign \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_12_U.a  = \add_32ns_32s_32_2_1_U15.din0 ;
assign \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_12_U.b  = \add_32ns_32s_32_2_1_U15.din1 ;
assign \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_12_U.ce  = \add_32ns_32s_32_2_1_U15.ce ;
assign \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_12_U.clk  = \add_32ns_32s_32_2_1_U15.clk ;
assign \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_12_U.reset  = \add_32ns_32s_32_2_1_U15.reset ;
assign \add_32ns_32s_32_2_1_U15.dout  = \add_32ns_32s_32_2_1_U15.top_add_32ns_32s_32_2_1_Adder_12_U.s ;
assign \add_32ns_32s_32_2_1_U15.ce  = 1'h1;
assign \add_32ns_32s_32_2_1_U15.clk  = ap_clk;
assign \add_32ns_32s_32_2_1_U15.din0  = ret_V_29_reg_1610;
assign \add_32ns_32s_32_2_1_U15.din1  = { op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14 };
assign grp_fu_984_p2 = \add_32ns_32s_32_2_1_U15.dout ;
assign \add_32ns_32s_32_2_1_U15.reset  = ap_rst;
assign \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.ain_s0  = \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.a ;
assign \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.bin_s0  = \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.b ;
assign \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.s  = { \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.fas_s2 , \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.sum_s1  };
assign \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.a  = \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.ain_s1 ;
assign \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.b  = \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.bin_s1 ;
assign \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.cin  = \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.carry_s1 ;
assign \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.facout_s2  = \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.cout ;
assign \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.fas_s2  = \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.s ;
assign \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.a  = \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.a [15:0];
assign \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.b  = \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.b [15:0];
assign \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.cin  = 1'h0;
assign \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.facout_s1  = \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.cout ;
assign \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.fas_s1  = \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.s ;
assign \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.a  = \add_32ns_32ns_32_2_1_U20.din0 ;
assign \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.b  = \add_32ns_32ns_32_2_1_U20.din1 ;
assign \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.ce  = \add_32ns_32ns_32_2_1_U20.ce ;
assign \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.clk  = \add_32ns_32ns_32_2_1_U20.clk ;
assign \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.reset  = \add_32ns_32ns_32_2_1_U20.reset ;
assign \add_32ns_32ns_32_2_1_U20.dout  = \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.s ;
assign \add_32ns_32ns_32_2_1_U20.ce  = 1'h1;
assign \add_32ns_32ns_32_2_1_U20.clk  = ap_clk;
assign \add_32ns_32ns_32_2_1_U20.din0  = ret_V_33_cast_reg_1692;
assign \add_32ns_32ns_32_2_1_U20.din1  = 32'd1;
assign grp_fu_1104_p2 = \add_32ns_32ns_32_2_1_U20.dout ;
assign \add_32ns_32ns_32_2_1_U20.reset  = ap_rst;
assign \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_11_U.ain_s0  = \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_11_U.a ;
assign \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_11_U.bin_s0  = \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_11_U.b ;
assign \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_11_U.s  = { \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_11_U.fas_s2 , \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_11_U.sum_s1  };
assign \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.a  = \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_11_U.ain_s1 ;
assign \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.b  = \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_11_U.bin_s1 ;
assign \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.cin  = \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_11_U.carry_s1 ;
assign \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_11_U.facout_s2  = \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.cout ;
assign \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_11_U.fas_s2  = \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.s ;
assign \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.a  = \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_11_U.a [15:0];
assign \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.b  = \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_11_U.b [15:0];
assign \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.cin  = 1'h0;
assign \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_11_U.facout_s1  = \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.cout ;
assign \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_11_U.fas_s1  = \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.s ;
assign \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_11_U.a  = \add_32ns_32ns_32_2_1_U18.din0 ;
assign \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_11_U.b  = \add_32ns_32ns_32_2_1_U18.din1 ;
assign \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_11_U.ce  = \add_32ns_32ns_32_2_1_U18.ce ;
assign \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_11_U.clk  = \add_32ns_32ns_32_2_1_U18.clk ;
assign \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_11_U.reset  = \add_32ns_32ns_32_2_1_U18.reset ;
assign \add_32ns_32ns_32_2_1_U18.dout  = \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_11_U.s ;
assign \add_32ns_32ns_32_2_1_U18.ce  = 1'h1;
assign \add_32ns_32ns_32_2_1_U18.clk  = ap_clk;
assign \add_32ns_32ns_32_2_1_U18.din0  = ret_V_31_reg_1657;
assign \add_32ns_32ns_32_2_1_U18.din1  = { 30'h00000000, op_16 };
assign grp_fu_1058_p2 = \add_32ns_32ns_32_2_1_U18.dout ;
assign \add_32ns_32ns_32_2_1_U18.reset  = ap_rst;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.ain_s0  = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.a ;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.bin_s0  = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.b ;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.s  = { \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.fas_s2 , \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.sum_s1  };
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.a  = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.ain_s1 ;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.b  = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.bin_s1 ;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.cin  = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.carry_s1 ;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.facout_s2  = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.cout ;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.fas_s2  = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.s ;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.a  = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.a [15:0];
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.b  = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.b [15:0];
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.cin  = 1'h0;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.facout_s1  = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.cout ;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.fas_s1  = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.s ;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.a  = \add_32ns_32ns_32_2_1_U17.din0 ;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.b  = \add_32ns_32ns_32_2_1_U17.din1 ;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.ce  = \add_32ns_32ns_32_2_1_U17.ce ;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.clk  = \add_32ns_32ns_32_2_1_U17.clk ;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.reset  = \add_32ns_32ns_32_2_1_U17.reset ;
assign \add_32ns_32ns_32_2_1_U17.dout  = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.s ;
assign \add_32ns_32ns_32_2_1_U17.ce  = 1'h1;
assign \add_32ns_32ns_32_2_1_U17.clk  = ap_clk;
assign \add_32ns_32ns_32_2_1_U17.din0  = ret_V_31_cast_reg_1645;
assign \add_32ns_32ns_32_2_1_U17.din1  = 32'd1;
assign grp_fu_1030_p2 = \add_32ns_32ns_32_2_1_U17.dout ;
assign \add_32ns_32ns_32_2_1_U17.reset  = ap_rst;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.ain_s0  = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.a ;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.bin_s0  = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.b ;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.s  = { \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.fas_s2 , \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.sum_s1  };
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.a  = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.ain_s1 ;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.b  = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.bin_s1 ;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.cin  = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.carry_s1 ;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.facout_s2  = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.cout ;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.fas_s2  = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.s ;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.a  = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.a [15:0];
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.b  = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.b [15:0];
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.cin  = 1'h0;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.facout_s1  = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.cout ;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.fas_s1  = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.s ;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.a  = \add_32ns_32ns_32_2_1_U14.din0 ;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.b  = \add_32ns_32ns_32_2_1_U14.din1 ;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.ce  = \add_32ns_32ns_32_2_1_U14.ce ;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.clk  = \add_32ns_32ns_32_2_1_U14.clk ;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.reset  = \add_32ns_32ns_32_2_1_U14.reset ;
assign \add_32ns_32ns_32_2_1_U14.dout  = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.s ;
assign \add_32ns_32ns_32_2_1_U14.ce  = 1'h1;
assign \add_32ns_32ns_32_2_1_U14.clk  = ap_clk;
assign \add_32ns_32ns_32_2_1_U14.din0  = ret_V_29_cast_reg_1598;
assign \add_32ns_32ns_32_2_1_U14.din1  = 32'd1;
assign grp_fu_956_p2 = \add_32ns_32ns_32_2_1_U14.dout ;
assign \add_32ns_32ns_32_2_1_U14.reset  = ap_rst;
assign \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.ain_s0  = \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.a ;
assign \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.bin_s0  = \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.b ;
assign \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.s  = { \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.fas_s2 , \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.sum_s1  };
assign \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.a  = \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.ain_s1 ;
assign \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.b  = \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.bin_s1 ;
assign \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.cin  = \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.carry_s1 ;
assign \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.facout_s2  = \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.cout ;
assign \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.fas_s2  = \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.s ;
assign \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.a  = \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.a [0];
assign \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.b  = \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.b [0];
assign \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.cin  = 1'h0;
assign \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.facout_s1  = \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.cout ;
assign \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.fas_s1  = \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.s ;
assign \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.a  = \add_2ns_2ns_2_2_1_U3.din0 ;
assign \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.b  = \add_2ns_2ns_2_2_1_U3.din1 ;
assign \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.ce  = \add_2ns_2ns_2_2_1_U3.ce ;
assign \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.clk  = \add_2ns_2ns_2_2_1_U3.clk ;
assign \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.reset  = \add_2ns_2ns_2_2_1_U3.reset ;
assign \add_2ns_2ns_2_2_1_U3.dout  = \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.s ;
assign \add_2ns_2ns_2_2_1_U3.ce  = 1'h1;
assign \add_2ns_2ns_2_2_1_U3.clk  = ap_clk;
assign \add_2ns_2ns_2_2_1_U3.din0  = ret_V_3_cast_reg_1194;
assign \add_2ns_2ns_2_2_1_U3.din1  = 2'h1;
assign grp_fu_300_p2 = \add_2ns_2ns_2_2_1_U3.dout ;
assign \add_2ns_2ns_2_2_1_U3.reset  = ap_rst;
assign \add_12ns_12s_12_2_1_U8.top_add_12ns_12s_12_2_1_Adder_5_U.ain_s0  = \add_12ns_12s_12_2_1_U8.top_add_12ns_12s_12_2_1_Adder_5_U.a ;
assign \add_12ns_12s_12_2_1_U8.top_add_12ns_12s_12_2_1_Adder_5_U.bin_s0  = \add_12ns_12s_12_2_1_U8.top_add_12ns_12s_12_2_1_Adder_5_U.b ;
assign \add_12ns_12s_12_2_1_U8.top_add_12ns_12s_12_2_1_Adder_5_U.s  = { \add_12ns_12s_12_2_1_U8.top_add_12ns_12s_12_2_1_Adder_5_U.fas_s2 , \add_12ns_12s_12_2_1_U8.top_add_12ns_12s_12_2_1_Adder_5_U.sum_s1  };
assign \add_12ns_12s_12_2_1_U8.top_add_12ns_12s_12_2_1_Adder_5_U.u2.a  = \add_12ns_12s_12_2_1_U8.top_add_12ns_12s_12_2_1_Adder_5_U.ain_s1 ;
assign \add_12ns_12s_12_2_1_U8.top_add_12ns_12s_12_2_1_Adder_5_U.u2.b  = \add_12ns_12s_12_2_1_U8.top_add_12ns_12s_12_2_1_Adder_5_U.bin_s1 ;
assign \add_12ns_12s_12_2_1_U8.top_add_12ns_12s_12_2_1_Adder_5_U.u2.cin  = \add_12ns_12s_12_2_1_U8.top_add_12ns_12s_12_2_1_Adder_5_U.carry_s1 ;
assign \add_12ns_12s_12_2_1_U8.top_add_12ns_12s_12_2_1_Adder_5_U.facout_s2  = \add_12ns_12s_12_2_1_U8.top_add_12ns_12s_12_2_1_Adder_5_U.u2.cout ;
assign \add_12ns_12s_12_2_1_U8.top_add_12ns_12s_12_2_1_Adder_5_U.fas_s2  = \add_12ns_12s_12_2_1_U8.top_add_12ns_12s_12_2_1_Adder_5_U.u2.s ;
assign \add_12ns_12s_12_2_1_U8.top_add_12ns_12s_12_2_1_Adder_5_U.u1.a  = \add_12ns_12s_12_2_1_U8.top_add_12ns_12s_12_2_1_Adder_5_U.a [5:0];
assign \add_12ns_12s_12_2_1_U8.top_add_12ns_12s_12_2_1_Adder_5_U.u1.b  = \add_12ns_12s_12_2_1_U8.top_add_12ns_12s_12_2_1_Adder_5_U.b [5:0];
assign \add_12ns_12s_12_2_1_U8.top_add_12ns_12s_12_2_1_Adder_5_U.u1.cin  = 1'h0;
assign \add_12ns_12s_12_2_1_U8.top_add_12ns_12s_12_2_1_Adder_5_U.facout_s1  = \add_12ns_12s_12_2_1_U8.top_add_12ns_12s_12_2_1_Adder_5_U.u1.cout ;
assign \add_12ns_12s_12_2_1_U8.top_add_12ns_12s_12_2_1_Adder_5_U.fas_s1  = \add_12ns_12s_12_2_1_U8.top_add_12ns_12s_12_2_1_Adder_5_U.u1.s ;
assign \add_12ns_12s_12_2_1_U8.top_add_12ns_12s_12_2_1_Adder_5_U.a  = \add_12ns_12s_12_2_1_U8.din0 ;
assign \add_12ns_12s_12_2_1_U8.top_add_12ns_12s_12_2_1_Adder_5_U.b  = \add_12ns_12s_12_2_1_U8.din1 ;
assign \add_12ns_12s_12_2_1_U8.top_add_12ns_12s_12_2_1_Adder_5_U.ce  = \add_12ns_12s_12_2_1_U8.ce ;
assign \add_12ns_12s_12_2_1_U8.top_add_12ns_12s_12_2_1_Adder_5_U.clk  = \add_12ns_12s_12_2_1_U8.clk ;
assign \add_12ns_12s_12_2_1_U8.top_add_12ns_12s_12_2_1_Adder_5_U.reset  = \add_12ns_12s_12_2_1_U8.reset ;
assign \add_12ns_12s_12_2_1_U8.dout  = \add_12ns_12s_12_2_1_U8.top_add_12ns_12s_12_2_1_Adder_5_U.s ;
assign \add_12ns_12s_12_2_1_U8.ce  = 1'h1;
assign \add_12ns_12s_12_2_1_U8.clk  = ap_clk;
assign \add_12ns_12s_12_2_1_U8.din0  = { 2'h0, ret_V_21_reg_1329[2], ret_V_21_reg_1329[2], ret_V_21_reg_1329[2], ret_V_21_reg_1329[2], ret_V_21_reg_1329[2], ret_V_21_reg_1329, 2'h0 };
assign \add_12ns_12s_12_2_1_U8.din1  = { op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5 };
assign grp_fu_650_p2 = \add_12ns_12s_12_2_1_U8.dout ;
assign \add_12ns_12s_12_2_1_U8.reset  = ap_rst;
assign \add_11s_11s_11_2_1_U12.top_add_11s_11s_11_2_1_Adder_9_U.ain_s0  = \add_11s_11s_11_2_1_U12.top_add_11s_11s_11_2_1_Adder_9_U.a ;
assign \add_11s_11s_11_2_1_U12.top_add_11s_11s_11_2_1_Adder_9_U.bin_s0  = \add_11s_11s_11_2_1_U12.top_add_11s_11s_11_2_1_Adder_9_U.b ;
assign \add_11s_11s_11_2_1_U12.top_add_11s_11s_11_2_1_Adder_9_U.s  = { \add_11s_11s_11_2_1_U12.top_add_11s_11s_11_2_1_Adder_9_U.fas_s2 , \add_11s_11s_11_2_1_U12.top_add_11s_11s_11_2_1_Adder_9_U.sum_s1  };
assign \add_11s_11s_11_2_1_U12.top_add_11s_11s_11_2_1_Adder_9_U.u2.a  = \add_11s_11s_11_2_1_U12.top_add_11s_11s_11_2_1_Adder_9_U.ain_s1 ;
assign \add_11s_11s_11_2_1_U12.top_add_11s_11s_11_2_1_Adder_9_U.u2.b  = \add_11s_11s_11_2_1_U12.top_add_11s_11s_11_2_1_Adder_9_U.bin_s1 ;
assign \add_11s_11s_11_2_1_U12.top_add_11s_11s_11_2_1_Adder_9_U.u2.cin  = \add_11s_11s_11_2_1_U12.top_add_11s_11s_11_2_1_Adder_9_U.carry_s1 ;
assign \add_11s_11s_11_2_1_U12.top_add_11s_11s_11_2_1_Adder_9_U.facout_s2  = \add_11s_11s_11_2_1_U12.top_add_11s_11s_11_2_1_Adder_9_U.u2.cout ;
assign \add_11s_11s_11_2_1_U12.top_add_11s_11s_11_2_1_Adder_9_U.fas_s2  = \add_11s_11s_11_2_1_U12.top_add_11s_11s_11_2_1_Adder_9_U.u2.s ;
assign \add_11s_11s_11_2_1_U12.top_add_11s_11s_11_2_1_Adder_9_U.u1.a  = \add_11s_11s_11_2_1_U12.top_add_11s_11s_11_2_1_Adder_9_U.a [4:0];
assign \add_11s_11s_11_2_1_U12.top_add_11s_11s_11_2_1_Adder_9_U.u1.b  = \add_11s_11s_11_2_1_U12.top_add_11s_11s_11_2_1_Adder_9_U.b [4:0];
assign \add_11s_11s_11_2_1_U12.top_add_11s_11s_11_2_1_Adder_9_U.u1.cin  = 1'h0;
assign \add_11s_11s_11_2_1_U12.top_add_11s_11s_11_2_1_Adder_9_U.facout_s1  = \add_11s_11s_11_2_1_U12.top_add_11s_11s_11_2_1_Adder_9_U.u1.cout ;
assign \add_11s_11s_11_2_1_U12.top_add_11s_11s_11_2_1_Adder_9_U.fas_s1  = \add_11s_11s_11_2_1_U12.top_add_11s_11s_11_2_1_Adder_9_U.u1.s ;
assign \add_11s_11s_11_2_1_U12.top_add_11s_11s_11_2_1_Adder_9_U.a  = \add_11s_11s_11_2_1_U12.din0 ;
assign \add_11s_11s_11_2_1_U12.top_add_11s_11s_11_2_1_Adder_9_U.b  = \add_11s_11s_11_2_1_U12.din1 ;
assign \add_11s_11s_11_2_1_U12.top_add_11s_11s_11_2_1_Adder_9_U.ce  = \add_11s_11s_11_2_1_U12.ce ;
assign \add_11s_11s_11_2_1_U12.top_add_11s_11s_11_2_1_Adder_9_U.clk  = \add_11s_11s_11_2_1_U12.clk ;
assign \add_11s_11s_11_2_1_U12.top_add_11s_11s_11_2_1_Adder_9_U.reset  = \add_11s_11s_11_2_1_U12.reset ;
assign \add_11s_11s_11_2_1_U12.dout  = \add_11s_11s_11_2_1_U12.top_add_11s_11s_11_2_1_Adder_9_U.s ;
assign \add_11s_11s_11_2_1_U12.ce  = 1'h1;
assign \add_11s_11s_11_2_1_U12.clk  = ap_clk;
assign \add_11s_11s_11_2_1_U12.din0  = { ret_V_27_reg_1543[3], ret_V_27_reg_1543[3], ret_V_27_reg_1543[3], ret_V_27_reg_1543[3], ret_V_27_reg_1543[3], ret_V_27_reg_1543[3], ret_V_27_reg_1543[3], ret_V_27_reg_1543 };
assign \add_11s_11s_11_2_1_U12.din1  = { ret_V_10_reg_1528[9], ret_V_10_reg_1528 };
assign grp_fu_906_p2 = \add_11s_11s_11_2_1_U12.dout ;
assign \add_11s_11s_11_2_1_U12.reset  = ap_rst;
assign \add_10ns_10ns_10_2_1_U10.top_add_10ns_10ns_10_2_1_Adder_7_U.ain_s0  = \add_10ns_10ns_10_2_1_U10.top_add_10ns_10ns_10_2_1_Adder_7_U.a ;
assign \add_10ns_10ns_10_2_1_U10.top_add_10ns_10ns_10_2_1_Adder_7_U.bin_s0  = \add_10ns_10ns_10_2_1_U10.top_add_10ns_10ns_10_2_1_Adder_7_U.b ;
assign \add_10ns_10ns_10_2_1_U10.top_add_10ns_10ns_10_2_1_Adder_7_U.s  = { \add_10ns_10ns_10_2_1_U10.top_add_10ns_10ns_10_2_1_Adder_7_U.fas_s2 , \add_10ns_10ns_10_2_1_U10.top_add_10ns_10ns_10_2_1_Adder_7_U.sum_s1  };
assign \add_10ns_10ns_10_2_1_U10.top_add_10ns_10ns_10_2_1_Adder_7_U.u2.a  = \add_10ns_10ns_10_2_1_U10.top_add_10ns_10ns_10_2_1_Adder_7_U.ain_s1 ;
assign \add_10ns_10ns_10_2_1_U10.top_add_10ns_10ns_10_2_1_Adder_7_U.u2.b  = \add_10ns_10ns_10_2_1_U10.top_add_10ns_10ns_10_2_1_Adder_7_U.bin_s1 ;
assign \add_10ns_10ns_10_2_1_U10.top_add_10ns_10ns_10_2_1_Adder_7_U.u2.cin  = \add_10ns_10ns_10_2_1_U10.top_add_10ns_10ns_10_2_1_Adder_7_U.carry_s1 ;
assign \add_10ns_10ns_10_2_1_U10.top_add_10ns_10ns_10_2_1_Adder_7_U.facout_s2  = \add_10ns_10ns_10_2_1_U10.top_add_10ns_10ns_10_2_1_Adder_7_U.u2.cout ;
assign \add_10ns_10ns_10_2_1_U10.top_add_10ns_10ns_10_2_1_Adder_7_U.fas_s2  = \add_10ns_10ns_10_2_1_U10.top_add_10ns_10ns_10_2_1_Adder_7_U.u2.s ;
assign \add_10ns_10ns_10_2_1_U10.top_add_10ns_10ns_10_2_1_Adder_7_U.u1.a  = \add_10ns_10ns_10_2_1_U10.top_add_10ns_10ns_10_2_1_Adder_7_U.a [4:0];
assign \add_10ns_10ns_10_2_1_U10.top_add_10ns_10ns_10_2_1_Adder_7_U.u1.b  = \add_10ns_10ns_10_2_1_U10.top_add_10ns_10ns_10_2_1_Adder_7_U.b [4:0];
assign \add_10ns_10ns_10_2_1_U10.top_add_10ns_10ns_10_2_1_Adder_7_U.u1.cin  = 1'h0;
assign \add_10ns_10ns_10_2_1_U10.top_add_10ns_10ns_10_2_1_Adder_7_U.facout_s1  = \add_10ns_10ns_10_2_1_U10.top_add_10ns_10ns_10_2_1_Adder_7_U.u1.cout ;
assign \add_10ns_10ns_10_2_1_U10.top_add_10ns_10ns_10_2_1_Adder_7_U.fas_s1  = \add_10ns_10ns_10_2_1_U10.top_add_10ns_10ns_10_2_1_Adder_7_U.u1.s ;
assign \add_10ns_10ns_10_2_1_U10.top_add_10ns_10ns_10_2_1_Adder_7_U.a  = \add_10ns_10ns_10_2_1_U10.din0 ;
assign \add_10ns_10ns_10_2_1_U10.top_add_10ns_10ns_10_2_1_Adder_7_U.b  = \add_10ns_10ns_10_2_1_U10.din1 ;
assign \add_10ns_10ns_10_2_1_U10.top_add_10ns_10ns_10_2_1_Adder_7_U.ce  = \add_10ns_10ns_10_2_1_U10.ce ;
assign \add_10ns_10ns_10_2_1_U10.top_add_10ns_10ns_10_2_1_Adder_7_U.clk  = \add_10ns_10ns_10_2_1_U10.clk ;
assign \add_10ns_10ns_10_2_1_U10.top_add_10ns_10ns_10_2_1_Adder_7_U.reset  = \add_10ns_10ns_10_2_1_U10.reset ;
assign \add_10ns_10ns_10_2_1_U10.dout  = \add_10ns_10ns_10_2_1_U10.top_add_10ns_10ns_10_2_1_Adder_7_U.s ;
assign \add_10ns_10ns_10_2_1_U10.ce  = 1'h1;
assign \add_10ns_10ns_10_2_1_U10.clk  = ap_clk;
assign \add_10ns_10ns_10_2_1_U10.din0  = ret_V_8_reg_1429;
assign \add_10ns_10ns_10_2_1_U10.din1  = 10'h001;
assign grp_fu_731_p2 = \add_10ns_10ns_10_2_1_U10.dout ;
assign \add_10ns_10ns_10_2_1_U10.reset  = ap_rst;
endmodule


// Machine B:
// Processed by function `add_clk_enable_signal` in `verilog_tricks.py`.
// Processed by function `remove_reset_signal` in `verilog_tricks.py`.
module top_B (
  ap_clk,
  ap_start,
  ap_done,
  ap_idle,
  ap_ready,
  op_0,
  op_4,
  op_5,
  op_6,
  op_10,
  op_14,
  op_15,
  op_16,
  op_17,
  op_18,
  op_29,
  op_29_ap_vld,
clk_enable
);
input clk_enable;


input ap_clk;
wire ap_rst;
assign ap_rst = op_29_ap_vld;
input ap_start;
input op_0;
input op_10;
input [3:0] op_14;
input [7:0] op_15;
input [1:0] op_16;
input [7:0] op_17;
input op_18;
input [1:0] op_4;
input [3:0] op_5;
input [1:0] op_6;
output ap_done;
output ap_idle;
output ap_ready;
output [31:0] op_29;
output op_29_ap_vld;


reg [31:0] add_ln691_1_reg_1376;
reg and_ln786_reg_1281;
reg [7:0] ap_CS_fsm = 8'h01;
reg icmp_ln851_2_reg_1255;
reg icmp_ln851_3_reg_1340;
reg icmp_ln851_4_reg_1371;
reg icmp_ln851_5_reg_1393;
reg icmp_ln851_6_reg_1415;
reg [3:0] op_11_V_reg_1301;
reg [7:0] op_13_V_reg_1345;
reg [10:0] op_22_V_reg_1350;
reg [31:0] op_26_V_reg_1398;
reg or_ln785_reg_1271;
reg p_Result_16_reg_1260;
reg p_Result_19_reg_1311;
reg p_Result_20_reg_1327;
reg [3:0] p_Val2_5_reg_1265;
reg [7:0] p_Val2_8_reg_1319;
reg [19:0] r_V_1_reg_1306;
reg [9:0] ret_V_10_reg_1296;
reg [2:0] ret_V_21_reg_1244;
reg [1:0] ret_V_22_reg_1250;
reg [2:0] ret_V_23_reg_1291;
reg [36:0] ret_V_28_reg_1360;
reg [31:0] ret_V_29_cast_reg_1365;
reg [37:0] ret_V_30_reg_1381;
reg [31:0] ret_V_31_cast_reg_1386;
reg [35:0] ret_V_32_reg_1403;
reg [31:0] ret_V_33_cast_reg_1408;
reg sel_tmp11_reg_1286;
reg [3:0] select_ln340_reg_1276;
reg tmp_12_reg_1333;
reg [3:0] trunc_ln851_4_reg_1355;
wire [31:0] _000_;
wire _001_;
wire [7:0] _002_;
wire _003_;
wire _004_;
wire _005_;
wire _006_;
wire _007_;
wire [3:0] _008_;
wire [7:0] _009_;
wire [10:0] _010_;
wire [31:0] _011_;
wire _012_;
wire _013_;
wire _014_;
wire _015_;
wire [2:0] _016_;
wire [7:0] _017_;
wire [19:0] _018_;
wire [9:0] _019_;
wire [2:0] _020_;
wire [1:0] _021_;
wire [2:0] _022_;
wire [36:0] _023_;
wire [31:0] _024_;
wire [37:0] _025_;
wire [31:0] _026_;
wire [35:0] _027_;
wire [31:0] _028_;
wire _029_;
wire [3:0] _030_;
wire _031_;
wire [3:0] _032_;
wire [1:0] _033_;
wire _034_;
wire _035_;
wire _036_;
wire _037_;
wire _038_;
wire _039_;
wire _040_;
wire _041_;
wire _042_;
wire _043_;
wire _044_;
wire _045_;
wire _046_;
wire _047_;
wire _048_;
wire _049_;
wire _050_;
wire _051_;
wire _052_;
wire _053_;
wire [31:0] add_ln691_1_fu_1023_p2;
wire [31:0] add_ln691_2_fu_1107_p2;
wire [31:0] add_ln691_3_fu_1183_p2;
wire [3:0] add_ln691_fu_950_p2;
wire [8:0] add_ln69_fu_1216_p2;
wire and_ln340_1_fu_551_p2;
wire and_ln340_2_fu_844_p2;
wire and_ln340_3_fu_881_p2;
wire and_ln340_fu_525_p2;
wire and_ln785_1_fu_557_p2;
wire and_ln785_3_fu_868_p2;
wire and_ln785_4_fu_887_p2;
wire and_ln785_fu_706_p2;
wire and_ln786_1_fu_791_p2;
wire and_ln786_fu_545_p2;
wire ap_CS_fsm_state1;
wire ap_CS_fsm_state2;
wire ap_CS_fsm_state3;
wire ap_CS_fsm_state4;
wire ap_CS_fsm_state5;
wire ap_CS_fsm_state6;
wire ap_CS_fsm_state7;
wire ap_CS_fsm_state8;
wire [7:0] ap_NS_fsm;
wire ap_clk;
wire ap_done;
wire ap_idle;
wire ap_ready;
wire ap_rst;
wire ap_start;
wire icmp_ln768_fu_427_p2;
wire icmp_ln786_fu_457_p2;
wire icmp_ln851_1_fu_337_p2;
wire icmp_ln851_2_fu_369_p2;
wire icmp_ln851_3_fu_770_p2;
wire icmp_ln851_4_fu_1018_p2;
wire icmp_ln851_5_fu_1094_p2;
wire icmp_ln851_6_fu_1170_p2;
wire icmp_ln851_fu_273_p2;
wire [1:0] lhs_V_fu_662_p3;
wire [1:0] lhs_fu_229_p1;
wire [2:0] lhs_fu_229_p3;
wire [3:0] \mul_4s_2s_6_1_1_U1.din0 ;
wire [1:0] \mul_4s_2s_6_1_1_U1.din1 ;
wire [5:0] \mul_4s_2s_6_1_1_U1.dout ;
wire [3:0] \mul_4s_2s_6_1_1_U1.top_mul_4s_2s_6_1_1_Multiplier_0_U.a ;
wire [1:0] \mul_4s_2s_6_1_1_U1.top_mul_4s_2s_6_1_1_Multiplier_0_U.b ;
wire [5:0] \mul_4s_2s_6_1_1_U1.top_mul_4s_2s_6_1_1_Multiplier_0_U.p ;
wire op_0;
wire op_10;
wire [3:0] op_11_V_fu_717_p3;
wire [7:0] op_13_V_fu_905_p3;
wire [3:0] op_14;
wire [7:0] op_15;
wire [1:0] op_16;
wire [7:0] op_17;
wire op_18;
wire [10:0] op_22_V_fu_978_p2;
wire [31:0] op_24_V_fu_1052_p2;
wire [31:0] op_26_V_fu_1129_p2;
wire [31:0] op_29;
wire op_29_ap_vld;
wire [1:0] op_4;
wire [3:0] op_5;
wire [1:0] op_6;
wire [16:0] op_7_V_fu_682_p4;
wire [1:0] or_ln1195_fu_670_p1;
wire [1:0] or_ln1195_fu_670_p2;
wire or_ln340_1_fu_801_p2;
wire or_ln340_fu_469_p2;
wire or_ln785_1_fu_776_p2;
wire or_ln785_2_fu_701_p2;
wire or_ln785_3_fu_563_p2;
wire or_ln785_4_fu_863_p2;
wire or_ln785_5_fu_893_p2;
wire or_ln785_fu_433_p2;
wire or_ln786_fu_463_p2;
wire overflow_1_fu_785_p2;
wire overflow_fu_445_p2;
wire [7:0] p_Result_11_fu_829_p4;
wire p_Result_12_fu_942_p3;
wire p_Result_13_fu_1029_p3;
wire p_Result_14_fu_1100_p3;
wire p_Result_15_fu_1176_p3;
wire p_Result_16_fu_381_p3;
wire p_Result_17_fu_401_p3;
wire p_Result_18_fu_409_p3;
wire p_Result_1_fu_325_p3;
wire p_Result_3_fu_633_p3;
wire [3:0] p_Result_7_fu_509_p4;
wire [1:0] p_Result_s_18_fu_417_p4;
wire p_Result_s_fu_261_p3;
wire [3:0] p_Val2_5_fu_393_p3;
wire [2:0] p_Val2_6_fu_503_p2;
wire [6:0] p_Val2_9_fu_824_p2;
wire [19:0] r_V_1_fu_726_p2;
wire [5:0] r_V_fu_309_p2;
wire [9:0] ret_V_10_fu_654_p3;
wire [4:0] ret_V_20_fu_245_p2;
wire [2:0] ret_V_21_fu_293_p3;
wire [1:0] ret_V_22_fu_357_p3;
wire [2:0] ret_V_23_fu_587_p2;
wire [11:0] ret_V_24_fu_617_p2;
wire [4:0] ret_V_25_fu_375_p2;
wire [5:0] ret_V_26_fu_922_p2;
wire [3:0] ret_V_27_fu_963_p3;
wire [36:0] ret_V_28_fu_1002_p2;
wire [31:0] ret_V_29_cast_fu_1008_p4;
wire [31:0] ret_V_29_fu_1041_p3;
wire [2:0] ret_V_2_fu_279_p2;
wire [37:0] ret_V_30_fu_1074_p2;
wire [31:0] ret_V_31_fu_1118_p3;
wire [35:0] ret_V_32_fu_1150_p2;
wire [31:0] ret_V_33_fu_1194_p3;
wire [1:0] ret_V_3_cast_fu_315_p4;
wire [1:0] ret_V_4_fu_343_p2;
wire [9:0] ret_V_8_fu_623_p4;
wire [9:0] ret_V_9_fu_641_p2;
wire [2:0] ret_V_fu_251_p4;
wire [4:0] rhs_1_fu_602_p3;
wire [5:0] rhs_2_fu_915_p3;
wire [36:0] rhs_5_fu_1062_p3;
wire [34:0] rhs_7_fu_1139_p3;
wire sel_tmp11_fu_569_p2;
wire sel_tmp24_fu_899_p2;
wire [7:0] select_ln340_1_fu_850_p3;
wire [3:0] select_ln340_fu_531_p3;
wire [8:0] select_ln69_fu_1201_p3;
wire [2:0] select_ln703_fu_579_p3;
wire [7:0] select_ln785_1_fu_874_p3;
wire [3:0] select_ln785_fu_711_p3;
wire [1:0] select_ln850_1_fu_349_p3;
wire [9:0] select_ln850_2_fu_647_p3;
wire [3:0] select_ln850_3_fu_956_p3;
wire [31:0] select_ln850_4_fu_1036_p3;
wire [31:0] select_ln850_5_fu_1112_p3;
wire [31:0] select_ln850_6_fu_1188_p3;
wire [2:0] select_ln850_fu_285_p3;
wire [5:0] sext_ln1192_1_fu_912_p1;
wire [36:0] sext_ln1192_2_fu_998_p1;
wire [37:0] sext_ln1192_3_fu_1070_p1;
wire [35:0] sext_ln1192_4_fu_1146_p1;
wire [9:0] sext_ln1192_fu_609_p1;
wire [4:0] sext_ln1193_1_fu_237_p1;
wire [3:0] sext_ln1193_fu_241_p0;
wire [4:0] sext_ln1193_fu_241_p1;
wire [19:0] sext_ln15_fu_692_p1;
wire [31:0] sext_ln69_1_fu_1048_p1;
wire [7:0] sext_ln69_2_fu_1209_p1;
wire [31:0] sext_ln69_3_fu_1222_p1;
wire [10:0] sext_ln69_fu_975_p1;
wire [3:0] sext_ln703_1_fu_599_p0;
wire [11:0] sext_ln703_1_fu_599_p1;
wire [36:0] sext_ln703_2_fu_988_p1;
wire [7:0] sext_ln703_3_fu_1058_p0;
wire [37:0] sext_ln703_3_fu_1058_p1;
wire [7:0] sext_ln703_4_fu_1135_p0;
wire [35:0] sext_ln703_4_fu_1135_p1;
wire [2:0] sext_ln703_fu_575_p1;
wire [10:0] sext_ln831_fu_971_p1;
wire [3:0] sext_ln850_fu_938_p1;
wire tmp_13_fu_806_p3;
wire [14:0] tmp_16_fu_991_p3;
wire [2:0] tmp_3_fu_928_p4;
wire tmp_7_fu_475_p3;
wire tmp_8_fu_483_p3;
wire [1:0] tmp_fu_675_p1;
wire tmp_fu_675_p3;
wire [2:0] trunc_ln731_fu_389_p1;
wire [2:0] trunc_ln851_1_fu_333_p1;
wire [3:0] trunc_ln851_2_fu_365_p0;
wire [1:0] trunc_ln851_2_fu_365_p1;
wire [2:0] trunc_ln851_3_fu_766_p1;
wire [3:0] trunc_ln851_4_fu_984_p1;
wire [7:0] trunc_ln851_5_fu_1090_p0;
wire [4:0] trunc_ln851_5_fu_1090_p1;
wire [7:0] trunc_ln851_6_fu_1166_p0;
wire [2:0] trunc_ln851_6_fu_1166_p1;
wire [1:0] trunc_ln851_fu_269_p1;
wire xor_ln1499_fu_593_p2;
wire xor_ln340_1_fu_838_p2;
wire xor_ln340_fu_519_p2;
wire xor_ln365_1_fu_497_p2;
wire xor_ln365_2_fu_813_p2;
wire xor_ln365_3_fu_818_p2;
wire xor_ln365_fu_491_p2;
wire xor_ln785_1_fu_780_p2;
wire xor_ln785_2_fu_696_p2;
wire xor_ln785_3_fu_857_p2;
wire xor_ln785_fu_439_p2;
wire xor_ln786_1_fu_539_p2;
wire xor_ln786_2_fu_795_p2;
wire xor_ln786_fu_451_p2;
wire [11:0] zext_ln1192_fu_613_p1;
wire [19:0] zext_ln1393_fu_723_p1;
wire [8:0] zext_ln69_1_fu_1212_p1;
wire [31:0] zext_ln69_fu_1125_p1;


assign add_ln691_1_fu_1023_p2 = { ret_V_28_fu_1002_p2[36], ret_V_28_fu_1002_p2[36], ret_V_28_fu_1002_p2[36], ret_V_28_fu_1002_p2[36], ret_V_28_fu_1002_p2[36], ret_V_28_fu_1002_p2[36], ret_V_28_fu_1002_p2[36], ret_V_28_fu_1002_p2[36], ret_V_28_fu_1002_p2[36], ret_V_28_fu_1002_p2[36], ret_V_28_fu_1002_p2[36], ret_V_28_fu_1002_p2[36], ret_V_28_fu_1002_p2[36], ret_V_28_fu_1002_p2[36], ret_V_28_fu_1002_p2[36], ret_V_28_fu_1002_p2[36], ret_V_28_fu_1002_p2[36], ret_V_28_fu_1002_p2[36], ret_V_28_fu_1002_p2[36], ret_V_28_fu_1002_p2[36], ret_V_28_fu_1002_p2[36], ret_V_28_fu_1002_p2[14:4] } + 1'h1;
assign add_ln691_2_fu_1107_p2 = ret_V_31_cast_reg_1386 + 1'h1;
assign add_ln691_3_fu_1183_p2 = ret_V_33_cast_reg_1408 + 1'h1;
assign add_ln691_fu_950_p2 = $signed(ret_V_26_fu_922_p2[5:3]) + $signed(2'h1);
assign add_ln69_fu_1216_p2 = { ret_V_21_reg_1244[2], ret_V_21_reg_1244[2], ret_V_21_reg_1244[2], ret_V_21_reg_1244[2], ret_V_21_reg_1244[2], ret_V_21_reg_1244 } + select_ln69_fu_1201_p3;
assign op_22_V_fu_978_p2 = $signed(ret_V_27_fu_963_p3) + $signed(ret_V_10_reg_1296);
assign op_24_V_fu_1052_p2 = $signed(ret_V_29_fu_1041_p3) + $signed(op_14);
assign op_26_V_fu_1129_p2 = ret_V_31_fu_1118_p3 + op_16;
assign op_29 = $signed(add_ln69_fu_1216_p2) + $signed(ret_V_33_fu_1194_p3);
assign ret_V_23_fu_587_p2 = $signed(op_6) + $signed(select_ln703_fu_579_p3);
assign ret_V_24_fu_617_p2 = $signed({ 1'h0, ret_V_21_reg_1244[2], ret_V_21_reg_1244[2], ret_V_21_reg_1244[2], ret_V_21_reg_1244[2], ret_V_21_reg_1244[2], ret_V_21_reg_1244, 2'h0 }) + $signed(op_5);
assign ret_V_26_fu_922_p2 = $signed({ ret_V_23_reg_1291, 3'h0 }) + $signed(op_11_V_reg_1301);
assign { ret_V_28_fu_1002_p2[36], ret_V_28_fu_1002_p2[14:0] } = $signed({ op_22_V_reg_1350, 4'h0 }) + $signed(op_13_V_reg_1345);
assign ret_V_2_fu_279_p2 = ret_V_20_fu_245_p2[4:2] + 1'h1;
assign ret_V_30_fu_1074_p2 = $signed({ op_24_V_fu_1052_p2, 5'h00 }) + $signed(op_15);
assign ret_V_32_fu_1150_p2 = $signed({ op_26_V_reg_1398, 3'h0 }) + $signed(op_17);
assign ret_V_4_fu_343_p2 = r_V_fu_309_p2[4:3] + 1'h1;
assign ret_V_9_fu_641_p2 = ret_V_24_fu_617_p2[11:2] + 1'h1;
assign _034_ = ap_CS_fsm[0] & _036_;
assign _035_ = ap_CS_fsm[0] & ap_start;
assign and_ln340_1_fu_551_p2 = or_ln786_fu_463_p2 & or_ln340_fu_469_p2;
assign and_ln340_2_fu_844_p2 = xor_ln786_2_fu_795_p2 & xor_ln340_1_fu_838_p2;
assign and_ln340_3_fu_881_p2 = xor_ln786_2_fu_795_p2 & or_ln340_1_fu_801_p2;
assign and_ln340_fu_525_p2 = xor_ln340_fu_519_p2 & or_ln786_fu_463_p2;
assign and_ln785_1_fu_557_p2 = xor_ln785_fu_439_p2 & and_ln786_fu_545_p2;
assign and_ln785_3_fu_868_p2 = or_ln785_4_fu_863_p2 & and_ln786_1_fu_791_p2;
assign and_ln785_4_fu_887_p2 = xor_ln785_1_fu_780_p2 & and_ln786_1_fu_791_p2;
assign and_ln785_fu_706_p2 = or_ln785_2_fu_701_p2 & and_ln786_reg_1281;
assign and_ln786_1_fu_791_p2 = tmp_12_reg_1333 & p_Result_20_reg_1327;
assign and_ln786_fu_545_p2 = xor_ln786_1_fu_539_p2 & ret_V_25_fu_375_p2[2];
assign overflow_1_fu_785_p2 = xor_ln785_1_fu_780_p2 & or_ln785_1_fu_776_p2;
assign overflow_fu_445_p2 = xor_ln785_fu_439_p2 & or_ln785_fu_433_p2;
assign sel_tmp11_fu_569_p2 = xor_ln365_1_fu_497_p2 & or_ln785_3_fu_563_p2;
assign sel_tmp24_fu_899_p2 = xor_ln365_3_fu_818_p2 & or_ln785_5_fu_893_p2;
assign xor_ln785_fu_439_p2 = ~ ret_V_25_fu_375_p2[4];
assign xor_ln786_fu_451_p2 = ~ ret_V_25_fu_375_p2[2];
assign xor_ln785_1_fu_780_p2 = ~ p_Result_19_reg_1311;
assign xor_ln340_1_fu_838_p2 = ~ or_ln340_1_fu_801_p2;
assign xor_ln786_2_fu_795_p2 = ~ and_ln786_1_fu_791_p2;
assign xor_ln340_fu_519_p2 = ~ or_ln340_fu_469_p2;
assign xor_ln786_1_fu_539_p2 = ~ icmp_ln786_fu_457_p2;
assign xor_ln785_3_fu_857_p2 = ~ or_ln785_1_fu_776_p2;
assign xor_ln785_2_fu_696_p2 = ~ or_ln785_reg_1271;
assign xor_ln365_3_fu_818_p2 = ~ xor_ln365_2_fu_813_p2;
assign xor_ln1499_fu_593_p2 = ~ op_0;
assign xor_ln365_1_fu_497_p2 = ~ xor_ln365_fu_491_p2;
assign p_Val2_9_fu_824_p2 = ~ p_Val2_8_reg_1319[6:0];
assign p_Val2_6_fu_503_p2 = ~ { ret_V_25_fu_375_p2[1:0], 1'h0 };
assign _036_ = ~ ap_start;
assign _037_ = ! r_V_fu_309_p2[2:0];
assign _038_ = ! op_5[1:0];
assign _039_ = ! ret_V_20_fu_245_p2[1:0];
assign \mul_4s_2s_6_1_1_U1.top_mul_4s_2s_6_1_1_Multiplier_0_U.p  = $signed(\mul_4s_2s_6_1_1_U1.top_mul_4s_2s_6_1_1_Multiplier_0_U.a ) * $signed(\mul_4s_2s_6_1_1_U1.top_mul_4s_2s_6_1_1_Multiplier_0_U.b );
assign _040_ = | ret_V_25_fu_375_p2[4:3];
assign _041_ = ret_V_25_fu_375_p2[4:3] != 2'h3;
assign _042_ = | op_11_V_fu_717_p3[2:0];
assign _043_ = | trunc_ln851_4_reg_1355;
assign _044_ = | op_15[4:0];
assign _045_ = | op_17[2:0];
assign or_ln1195_fu_670_p2 = op_4 | { xor_ln1499_fu_593_p2, 1'h0 };
assign or_ln340_1_fu_801_p2 = p_Result_19_reg_1311 | overflow_1_fu_785_p2;
assign or_ln340_fu_469_p2 = ret_V_25_fu_375_p2[4] | overflow_fu_445_p2;
assign or_ln785_1_fu_776_p2 = tmp_12_reg_1333 | p_Result_20_reg_1327;
assign or_ln785_2_fu_701_p2 = xor_ln785_2_fu_696_p2 | p_Result_16_reg_1260;
assign or_ln785_3_fu_563_p2 = and_ln785_1_fu_557_p2 | and_ln340_1_fu_551_p2;
assign or_ln785_4_fu_863_p2 = xor_ln785_3_fu_857_p2 | p_Result_19_reg_1311;
assign or_ln785_5_fu_893_p2 = and_ln785_4_fu_887_p2 | and_ln340_3_fu_881_p2;
assign or_ln785_fu_433_p2 = ret_V_25_fu_375_p2[2] | icmp_ln768_fu_427_p2;
assign or_ln786_fu_463_p2 = xor_ln786_fu_451_p2 | icmp_ln786_fu_457_p2;
always @(posedge ap_clk)
p_Val2_5_reg_1265[0] <= 1'h0;
always @(posedge ap_clk)
op_26_V_reg_1398 <= _011_;
always @(posedge ap_clk)
op_13_V_reg_1345 <= _009_;
always @(posedge ap_clk)
op_22_V_reg_1350 <= _010_;
always @(posedge ap_clk)
trunc_ln851_4_reg_1355 <= _032_;
always @(posedge ap_clk)
ret_V_32_reg_1403 <= _027_;
always @(posedge ap_clk)
ret_V_33_cast_reg_1408 <= _028_;
always @(posedge ap_clk)
icmp_ln851_6_reg_1415 <= _007_;
always @(posedge ap_clk)
ret_V_30_reg_1381 <= _025_;
always @(posedge ap_clk)
ret_V_31_cast_reg_1386 <= _026_;
always @(posedge ap_clk)
icmp_ln851_5_reg_1393 <= _006_;
always @(posedge ap_clk)
ret_V_23_reg_1291 <= _022_;
always @(posedge ap_clk)
ret_V_10_reg_1296 <= _019_;
always @(posedge ap_clk)
op_11_V_reg_1301 <= _008_;
always @(posedge ap_clk)
r_V_1_reg_1306 <= _018_;
always @(posedge ap_clk)
p_Result_19_reg_1311 <= _014_;
always @(posedge ap_clk)
p_Val2_8_reg_1319 <= _017_;
always @(posedge ap_clk)
p_Result_20_reg_1327 <= _015_;
always @(posedge ap_clk)
tmp_12_reg_1333 <= _031_;
always @(posedge ap_clk)
icmp_ln851_3_reg_1340 <= _004_;
always @(posedge ap_clk)
ret_V_21_reg_1244 <= _020_;
always @(posedge ap_clk)
ret_V_22_reg_1250 <= _021_;
always @(posedge ap_clk)
icmp_ln851_2_reg_1255 <= _003_;
always @(posedge ap_clk)
p_Result_16_reg_1260 <= _013_;
always @(posedge ap_clk)
p_Val2_5_reg_1265[3:1] <= _016_;
always @(posedge ap_clk)
or_ln785_reg_1271 <= _012_;
always @(posedge ap_clk)
select_ln340_reg_1276 <= _030_;
always @(posedge ap_clk)
and_ln786_reg_1281 <= _001_;
always @(posedge ap_clk)
sel_tmp11_reg_1286 <= _029_;
always @(posedge ap_clk)
ret_V_28_reg_1360 <= _023_;
always @(posedge ap_clk)
ret_V_29_cast_reg_1365 <= _024_;
always @(posedge ap_clk)
icmp_ln851_4_reg_1371 <= _005_;
always @(posedge ap_clk)
add_ln691_1_reg_1376 <= _000_;
always @(posedge ap_clk)
ap_CS_fsm <= _002_;
assign _033_ = _035_ ? 2'h2 : 2'h1;
assign _046_ = ap_CS_fsm == 1'h1;
function [7:0] _159_;
input [7:0] a;
input [63:0] b;
input [7:0] s;
case (s)
8'b00000001:
_159_ = b[7:0];
8'b00000010:
_159_ = b[15:8];
8'b00000100:
_159_ = b[23:16];
8'b00001000:
_159_ = b[31:24];
8'b00010000:
_159_ = b[39:32];
8'b00100000:
_159_ = b[47:40];
8'b01000000:
_159_ = b[55:48];
8'b10000000:
_159_ = b[63:56];
8'b00000000:
_159_ = a;
default:
_159_ = 8'bx;
endcase
endfunction
assign ap_NS_fsm = _159_(8'hxx, { 6'h00, _033_, 56'h04081020408001 }, { _046_, _053_, _052_, _051_, _050_, _049_, _048_, _047_ });
assign _047_ = ap_CS_fsm == 8'h80;
assign _048_ = ap_CS_fsm == 7'h40;
assign _049_ = ap_CS_fsm == 6'h20;
assign _050_ = ap_CS_fsm == 5'h10;
assign _051_ = ap_CS_fsm == 4'h8;
assign _052_ = ap_CS_fsm == 3'h4;
assign _053_ = ap_CS_fsm == 2'h2;
assign op_29_ap_vld = ap_CS_fsm[7] ? 1'h1 : 1'h0;
assign ap_idle = _034_ ? 1'h1 : 1'h0;
assign _011_ = ap_CS_fsm[5] ? op_26_V_fu_1129_p2 : op_26_V_reg_1398;
assign _032_ = ap_CS_fsm[2] ? op_13_V_fu_905_p3[3:0] : trunc_ln851_4_reg_1355;
assign _010_ = ap_CS_fsm[2] ? op_22_V_fu_978_p2 : op_22_V_reg_1350;
assign _009_ = ap_CS_fsm[2] ? op_13_V_fu_905_p3 : op_13_V_reg_1345;
assign _007_ = ap_CS_fsm[6] ? icmp_ln851_6_fu_1170_p2 : icmp_ln851_6_reg_1415;
assign _028_ = ap_CS_fsm[6] ? ret_V_32_fu_1150_p2[34:3] : ret_V_33_cast_reg_1408;
assign _027_ = ap_CS_fsm[6] ? ret_V_32_fu_1150_p2 : ret_V_32_reg_1403;
assign _006_ = ap_CS_fsm[4] ? icmp_ln851_5_fu_1094_p2 : icmp_ln851_5_reg_1393;
assign _026_ = ap_CS_fsm[4] ? ret_V_30_fu_1074_p2[36:5] : ret_V_31_cast_reg_1386;
assign _025_ = ap_CS_fsm[4] ? ret_V_30_fu_1074_p2 : ret_V_30_reg_1381;
assign _004_ = ap_CS_fsm[1] ? icmp_ln851_3_fu_770_p2 : icmp_ln851_3_reg_1340;
assign _031_ = ap_CS_fsm[1] ? r_V_1_fu_726_p2[19] : tmp_12_reg_1333;
assign _015_ = ap_CS_fsm[1] ? r_V_1_fu_726_p2[18] : p_Result_20_reg_1327;
assign _017_ = ap_CS_fsm[1] ? r_V_1_fu_726_p2[18:11] : p_Val2_8_reg_1319;
assign _014_ = ap_CS_fsm[1] ? r_V_1_fu_726_p2[19] : p_Result_19_reg_1311;
assign _018_ = ap_CS_fsm[1] ? r_V_1_fu_726_p2 : r_V_1_reg_1306;
assign _008_ = ap_CS_fsm[1] ? op_11_V_fu_717_p3 : op_11_V_reg_1301;
assign _019_ = ap_CS_fsm[1] ? ret_V_10_fu_654_p3 : ret_V_10_reg_1296;
assign _022_ = ap_CS_fsm[1] ? ret_V_23_fu_587_p2 : ret_V_23_reg_1291;
assign _029_ = ap_CS_fsm[0] ? sel_tmp11_fu_569_p2 : sel_tmp11_reg_1286;
assign _001_ = ap_CS_fsm[0] ? and_ln786_fu_545_p2 : and_ln786_reg_1281;
assign _030_ = ap_CS_fsm[0] ? select_ln340_fu_531_p3 : select_ln340_reg_1276;
assign _012_ = ap_CS_fsm[0] ? or_ln785_fu_433_p2 : or_ln785_reg_1271;
assign _016_ = ap_CS_fsm[0] ? ret_V_25_fu_375_p2[2:0] : p_Val2_5_reg_1265[3:1];
assign _013_ = ap_CS_fsm[0] ? ret_V_25_fu_375_p2[4] : p_Result_16_reg_1260;
assign _003_ = ap_CS_fsm[0] ? icmp_ln851_2_fu_369_p2 : icmp_ln851_2_reg_1255;
assign _021_ = ap_CS_fsm[0] ? ret_V_22_fu_357_p3 : ret_V_22_reg_1250;
assign _020_ = ap_CS_fsm[0] ? ret_V_21_fu_293_p3 : ret_V_21_reg_1244;
assign _000_ = ap_CS_fsm[3] ? add_ln691_1_fu_1023_p2 : add_ln691_1_reg_1376;
assign _005_ = ap_CS_fsm[3] ? icmp_ln851_4_fu_1018_p2 : icmp_ln851_4_reg_1371;
assign _024_ = ap_CS_fsm[3] ? { ret_V_28_fu_1002_p2[36], ret_V_28_fu_1002_p2[36], ret_V_28_fu_1002_p2[36], ret_V_28_fu_1002_p2[36], ret_V_28_fu_1002_p2[36], ret_V_28_fu_1002_p2[36], ret_V_28_fu_1002_p2[36], ret_V_28_fu_1002_p2[36], ret_V_28_fu_1002_p2[36], ret_V_28_fu_1002_p2[36], ret_V_28_fu_1002_p2[36], ret_V_28_fu_1002_p2[36], ret_V_28_fu_1002_p2[36], ret_V_28_fu_1002_p2[36], ret_V_28_fu_1002_p2[36], ret_V_28_fu_1002_p2[36], ret_V_28_fu_1002_p2[36], ret_V_28_fu_1002_p2[36], ret_V_28_fu_1002_p2[36], ret_V_28_fu_1002_p2[36], ret_V_28_fu_1002_p2[36], ret_V_28_fu_1002_p2[14:4] } : ret_V_29_cast_reg_1365;
assign _023_ = ap_CS_fsm[3] ? { ret_V_28_fu_1002_p2[36], ret_V_28_fu_1002_p2[36], ret_V_28_fu_1002_p2[36], ret_V_28_fu_1002_p2[36], ret_V_28_fu_1002_p2[36], ret_V_28_fu_1002_p2[36], ret_V_28_fu_1002_p2[36], ret_V_28_fu_1002_p2[36], ret_V_28_fu_1002_p2[36], ret_V_28_fu_1002_p2[36], ret_V_28_fu_1002_p2[36], ret_V_28_fu_1002_p2[36], ret_V_28_fu_1002_p2[36], ret_V_28_fu_1002_p2[36], ret_V_28_fu_1002_p2[36], ret_V_28_fu_1002_p2[36], ret_V_28_fu_1002_p2[36], ret_V_28_fu_1002_p2[36], ret_V_28_fu_1002_p2[36], ret_V_28_fu_1002_p2[36], ret_V_28_fu_1002_p2[36], ret_V_28_fu_1002_p2[36], ret_V_28_fu_1002_p2[14:0] } : ret_V_28_reg_1360;
assign _002_ = ap_rst ? 8'h01 : ap_NS_fsm;
assign r_V_1_fu_726_p2 = $signed({ op_4[1], or_ln1195_fu_670_p2, 14'h0000 }) << ret_V_22_reg_1250;
assign ret_V_20_fu_245_p2 = $signed({ op_4, 1'h0 }) - $signed(op_5);
assign ret_V_25_fu_375_p2 = $signed(1'h0) - $signed(op_5);
assign icmp_ln768_fu_427_p2 = _040_ ? 1'h1 : 1'h0;
assign icmp_ln786_fu_457_p2 = _041_ ? 1'h1 : 1'h0;
assign icmp_ln851_1_fu_337_p2 = _037_ ? 1'h1 : 1'h0;
assign icmp_ln851_2_fu_369_p2 = _038_ ? 1'h1 : 1'h0;
assign icmp_ln851_3_fu_770_p2 = _042_ ? 1'h1 : 1'h0;
assign icmp_ln851_4_fu_1018_p2 = _043_ ? 1'h1 : 1'h0;
assign icmp_ln851_5_fu_1094_p2 = _044_ ? 1'h1 : 1'h0;
assign icmp_ln851_6_fu_1170_p2 = _045_ ? 1'h1 : 1'h0;
assign icmp_ln851_fu_273_p2 = _039_ ? 1'h1 : 1'h0;
assign op_11_V_fu_717_p3 = sel_tmp11_reg_1286 ? p_Val2_5_reg_1265 : select_ln785_fu_711_p3;
assign op_13_V_fu_905_p3 = sel_tmp24_fu_899_p2 ? p_Val2_8_reg_1319 : select_ln785_1_fu_874_p3;
assign ret_V_10_fu_654_p3 = ret_V_24_fu_617_p2[11] ? select_ln850_2_fu_647_p3 : { 1'h0, ret_V_24_fu_617_p2[10:2] };
assign ret_V_21_fu_293_p3 = ret_V_20_fu_245_p2[4] ? select_ln850_fu_285_p3 : { 1'h0, ret_V_20_fu_245_p2[3:2] };
assign ret_V_22_fu_357_p3 = r_V_fu_309_p2[5] ? select_ln850_1_fu_349_p3 : r_V_fu_309_p2[4:3];
assign ret_V_27_fu_963_p3 = ret_V_26_fu_922_p2[5] ? select_ln850_3_fu_956_p3 : { 2'h0, ret_V_26_fu_922_p2[4:3] };
assign ret_V_29_fu_1041_p3 = ret_V_28_reg_1360[36] ? select_ln850_4_fu_1036_p3 : ret_V_29_cast_reg_1365;
assign ret_V_31_fu_1118_p3 = ret_V_30_reg_1381[37] ? select_ln850_5_fu_1112_p3 : ret_V_31_cast_reg_1386;
assign ret_V_33_fu_1194_p3 = ret_V_32_reg_1403[35] ? select_ln850_6_fu_1188_p3 : ret_V_33_cast_reg_1408;
assign select_ln340_1_fu_850_p3 = and_ln340_2_fu_844_p2 ? p_Val2_8_reg_1319 : { p_Result_19_reg_1311, p_Val2_9_fu_824_p2 };
assign select_ln340_fu_531_p3 = and_ln340_fu_525_p2 ? { ret_V_25_fu_375_p2[2:0], 1'h0 } : { ret_V_25_fu_375_p2[3], p_Val2_6_fu_503_p2 };
assign select_ln69_fu_1201_p3 = op_18 ? 9'h1ff : 9'h000;
assign select_ln703_fu_579_p3 = op_10 ? 3'h7 : 3'h0;
assign select_ln785_1_fu_874_p3 = and_ln785_3_fu_868_p2 ? p_Val2_8_reg_1319 : select_ln340_1_fu_850_p3;
assign select_ln785_fu_711_p3 = and_ln785_fu_706_p2 ? p_Val2_5_reg_1265 : select_ln340_reg_1276;
assign select_ln850_1_fu_349_p3 = icmp_ln851_1_fu_337_p2 ? r_V_fu_309_p2[4:3] : ret_V_4_fu_343_p2;
assign select_ln850_2_fu_647_p3 = icmp_ln851_2_reg_1255 ? { 1'h1, ret_V_24_fu_617_p2[10:2] } : ret_V_9_fu_641_p2;
assign select_ln850_3_fu_956_p3 = icmp_ln851_3_reg_1340 ? add_ln691_fu_950_p2 : { 2'h3, ret_V_26_fu_922_p2[4:3] };
assign select_ln850_4_fu_1036_p3 = icmp_ln851_4_reg_1371 ? add_ln691_1_reg_1376 : ret_V_29_cast_reg_1365;
assign select_ln850_5_fu_1112_p3 = icmp_ln851_5_reg_1393 ? add_ln691_2_fu_1107_p2 : ret_V_31_cast_reg_1386;
assign select_ln850_6_fu_1188_p3 = icmp_ln851_6_reg_1415 ? add_ln691_3_fu_1183_p2 : ret_V_33_cast_reg_1408;
assign select_ln850_fu_285_p3 = icmp_ln851_fu_273_p2 ? { 1'h1, ret_V_20_fu_245_p2[3:2] } : ret_V_2_fu_279_p2;
assign xor_ln365_2_fu_813_p2 = r_V_1_reg_1306[18] ^ tmp_12_reg_1333;
assign xor_ln365_fu_491_p2 = ret_V_25_fu_375_p2[2] ^ ret_V_25_fu_375_p2[3];
assign ap_CS_fsm_state1 = ap_CS_fsm[0];
assign ap_CS_fsm_state2 = ap_CS_fsm[1];
assign ap_CS_fsm_state3 = ap_CS_fsm[2];
assign ap_CS_fsm_state4 = ap_CS_fsm[3];
assign ap_CS_fsm_state5 = ap_CS_fsm[4];
assign ap_CS_fsm_state6 = ap_CS_fsm[5];
assign ap_CS_fsm_state7 = ap_CS_fsm[6];
assign ap_CS_fsm_state8 = ap_CS_fsm[7];
assign ap_done = op_29_ap_vld;
assign ap_ready = op_29_ap_vld;
assign lhs_V_fu_662_p3 = { xor_ln1499_fu_593_p2, 1'h0 };
assign lhs_fu_229_p1 = op_4;
assign lhs_fu_229_p3 = { op_4, 1'h0 };
assign op_7_V_fu_682_p4 = { op_4[1], or_ln1195_fu_670_p2, 14'h0000 };
assign or_ln1195_fu_670_p1 = op_4;
assign p_Result_11_fu_829_p4 = { p_Result_19_reg_1311, p_Val2_9_fu_824_p2 };
assign p_Result_12_fu_942_p3 = ret_V_26_fu_922_p2[5];
assign p_Result_13_fu_1029_p3 = ret_V_28_reg_1360[36];
assign p_Result_14_fu_1100_p3 = ret_V_30_reg_1381[37];
assign p_Result_15_fu_1176_p3 = ret_V_32_reg_1403[35];
assign p_Result_16_fu_381_p3 = ret_V_25_fu_375_p2[4];
assign p_Result_17_fu_401_p3 = ret_V_25_fu_375_p2[2];
assign p_Result_18_fu_409_p3 = ret_V_25_fu_375_p2[3];
assign p_Result_1_fu_325_p3 = r_V_fu_309_p2[5];
assign p_Result_3_fu_633_p3 = ret_V_24_fu_617_p2[11];
assign p_Result_7_fu_509_p4 = { ret_V_25_fu_375_p2[3], p_Val2_6_fu_503_p2 };
assign p_Result_s_18_fu_417_p4 = ret_V_25_fu_375_p2[4:3];
assign p_Result_s_fu_261_p3 = ret_V_20_fu_245_p2[4];
assign p_Val2_5_fu_393_p3 = { ret_V_25_fu_375_p2[2:0], 1'h0 };
assign ret_V_28_fu_1002_p2[35:15] = { ret_V_28_fu_1002_p2[36], ret_V_28_fu_1002_p2[36], ret_V_28_fu_1002_p2[36], ret_V_28_fu_1002_p2[36], ret_V_28_fu_1002_p2[36], ret_V_28_fu_1002_p2[36], ret_V_28_fu_1002_p2[36], ret_V_28_fu_1002_p2[36], ret_V_28_fu_1002_p2[36], ret_V_28_fu_1002_p2[36], ret_V_28_fu_1002_p2[36], ret_V_28_fu_1002_p2[36], ret_V_28_fu_1002_p2[36], ret_V_28_fu_1002_p2[36], ret_V_28_fu_1002_p2[36], ret_V_28_fu_1002_p2[36], ret_V_28_fu_1002_p2[36], ret_V_28_fu_1002_p2[36], ret_V_28_fu_1002_p2[36], ret_V_28_fu_1002_p2[36], ret_V_28_fu_1002_p2[36] };
assign ret_V_29_cast_fu_1008_p4 = { ret_V_28_fu_1002_p2[36], ret_V_28_fu_1002_p2[36], ret_V_28_fu_1002_p2[36], ret_V_28_fu_1002_p2[36], ret_V_28_fu_1002_p2[36], ret_V_28_fu_1002_p2[36], ret_V_28_fu_1002_p2[36], ret_V_28_fu_1002_p2[36], ret_V_28_fu_1002_p2[36], ret_V_28_fu_1002_p2[36], ret_V_28_fu_1002_p2[36], ret_V_28_fu_1002_p2[36], ret_V_28_fu_1002_p2[36], ret_V_28_fu_1002_p2[36], ret_V_28_fu_1002_p2[36], ret_V_28_fu_1002_p2[36], ret_V_28_fu_1002_p2[36], ret_V_28_fu_1002_p2[36], ret_V_28_fu_1002_p2[36], ret_V_28_fu_1002_p2[36], ret_V_28_fu_1002_p2[36], ret_V_28_fu_1002_p2[14:4] };
assign ret_V_3_cast_fu_315_p4 = r_V_fu_309_p2[4:3];
assign ret_V_8_fu_623_p4 = ret_V_24_fu_617_p2[11:2];
assign ret_V_fu_251_p4 = ret_V_20_fu_245_p2[4:2];
assign rhs_1_fu_602_p3 = { ret_V_21_reg_1244, 2'h0 };
assign rhs_2_fu_915_p3 = { ret_V_23_reg_1291, 3'h0 };
assign rhs_5_fu_1062_p3 = { op_24_V_fu_1052_p2, 5'h00 };
assign rhs_7_fu_1139_p3 = { op_26_V_reg_1398, 3'h0 };
assign sext_ln1192_1_fu_912_p1 = { op_11_V_reg_1301[3], op_11_V_reg_1301[3], op_11_V_reg_1301 };
assign sext_ln1192_2_fu_998_p1 = { op_22_V_reg_1350[10], op_22_V_reg_1350[10], op_22_V_reg_1350[10], op_22_V_reg_1350[10], op_22_V_reg_1350[10], op_22_V_reg_1350[10], op_22_V_reg_1350[10], op_22_V_reg_1350[10], op_22_V_reg_1350[10], op_22_V_reg_1350[10], op_22_V_reg_1350[10], op_22_V_reg_1350[10], op_22_V_reg_1350[10], op_22_V_reg_1350[10], op_22_V_reg_1350[10], op_22_V_reg_1350[10], op_22_V_reg_1350[10], op_22_V_reg_1350[10], op_22_V_reg_1350[10], op_22_V_reg_1350[10], op_22_V_reg_1350[10], op_22_V_reg_1350[10], op_22_V_reg_1350, 4'h0 };
assign sext_ln1192_3_fu_1070_p1 = { op_24_V_fu_1052_p2[31], op_24_V_fu_1052_p2, 5'h00 };
assign sext_ln1192_4_fu_1146_p1 = { op_26_V_reg_1398[31], op_26_V_reg_1398, 3'h0 };
assign sext_ln1192_fu_609_p1 = { ret_V_21_reg_1244[2], ret_V_21_reg_1244[2], ret_V_21_reg_1244[2], ret_V_21_reg_1244[2], ret_V_21_reg_1244[2], ret_V_21_reg_1244, 2'h0 };
assign sext_ln1193_1_fu_237_p1 = { op_4[1], op_4[1], op_4, 1'h0 };
assign sext_ln1193_fu_241_p0 = op_5;
assign sext_ln1193_fu_241_p1 = { op_5[3], op_5 };
assign sext_ln15_fu_692_p1 = { op_4[1], op_4[1], op_4[1], op_4[1], or_ln1195_fu_670_p2, 14'h0000 };
assign sext_ln69_1_fu_1048_p1 = { op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14 };
assign sext_ln69_2_fu_1209_p1 = { ret_V_21_reg_1244[2], ret_V_21_reg_1244[2], ret_V_21_reg_1244[2], ret_V_21_reg_1244[2], ret_V_21_reg_1244[2], ret_V_21_reg_1244 };
assign sext_ln69_3_fu_1222_p1 = { add_ln69_fu_1216_p2[8], add_ln69_fu_1216_p2[8], add_ln69_fu_1216_p2[8], add_ln69_fu_1216_p2[8], add_ln69_fu_1216_p2[8], add_ln69_fu_1216_p2[8], add_ln69_fu_1216_p2[8], add_ln69_fu_1216_p2[8], add_ln69_fu_1216_p2[8], add_ln69_fu_1216_p2[8], add_ln69_fu_1216_p2[8], add_ln69_fu_1216_p2[8], add_ln69_fu_1216_p2[8], add_ln69_fu_1216_p2[8], add_ln69_fu_1216_p2[8], add_ln69_fu_1216_p2[8], add_ln69_fu_1216_p2[8], add_ln69_fu_1216_p2[8], add_ln69_fu_1216_p2[8], add_ln69_fu_1216_p2[8], add_ln69_fu_1216_p2[8], add_ln69_fu_1216_p2[8], add_ln69_fu_1216_p2[8], add_ln69_fu_1216_p2 };
assign sext_ln69_fu_975_p1 = { ret_V_10_reg_1296[9], ret_V_10_reg_1296 };
assign sext_ln703_1_fu_599_p0 = op_5;
assign sext_ln703_1_fu_599_p1 = { op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5 };
assign sext_ln703_2_fu_988_p1 = { op_13_V_reg_1345[7], op_13_V_reg_1345[7], op_13_V_reg_1345[7], op_13_V_reg_1345[7], op_13_V_reg_1345[7], op_13_V_reg_1345[7], op_13_V_reg_1345[7], op_13_V_reg_1345[7], op_13_V_reg_1345[7], op_13_V_reg_1345[7], op_13_V_reg_1345[7], op_13_V_reg_1345[7], op_13_V_reg_1345[7], op_13_V_reg_1345[7], op_13_V_reg_1345[7], op_13_V_reg_1345[7], op_13_V_reg_1345[7], op_13_V_reg_1345[7], op_13_V_reg_1345[7], op_13_V_reg_1345[7], op_13_V_reg_1345[7], op_13_V_reg_1345[7], op_13_V_reg_1345[7], op_13_V_reg_1345[7], op_13_V_reg_1345[7], op_13_V_reg_1345[7], op_13_V_reg_1345[7], op_13_V_reg_1345[7], op_13_V_reg_1345[7], op_13_V_reg_1345 };
assign sext_ln703_3_fu_1058_p0 = op_15;
assign sext_ln703_3_fu_1058_p1 = { op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15 };
assign sext_ln703_4_fu_1135_p0 = op_17;
assign sext_ln703_4_fu_1135_p1 = { op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17 };
assign sext_ln703_fu_575_p1 = { op_6[1], op_6 };
assign sext_ln831_fu_971_p1 = { ret_V_27_fu_963_p3[3], ret_V_27_fu_963_p3[3], ret_V_27_fu_963_p3[3], ret_V_27_fu_963_p3[3], ret_V_27_fu_963_p3[3], ret_V_27_fu_963_p3[3], ret_V_27_fu_963_p3[3], ret_V_27_fu_963_p3 };
assign sext_ln850_fu_938_p1 = { ret_V_26_fu_922_p2[5], ret_V_26_fu_922_p2[5:3] };
assign tmp_13_fu_806_p3 = r_V_1_reg_1306[18];
assign tmp_16_fu_991_p3 = { op_22_V_reg_1350, 4'h0 };
assign tmp_3_fu_928_p4 = ret_V_26_fu_922_p2[5:3];
assign tmp_7_fu_475_p3 = ret_V_25_fu_375_p2[3];
assign tmp_8_fu_483_p3 = ret_V_25_fu_375_p2[2];
assign tmp_fu_675_p1 = op_4;
assign tmp_fu_675_p3 = op_4[1];
assign trunc_ln731_fu_389_p1 = ret_V_25_fu_375_p2[2:0];
assign trunc_ln851_1_fu_333_p1 = r_V_fu_309_p2[2:0];
assign trunc_ln851_2_fu_365_p0 = op_5;
assign trunc_ln851_2_fu_365_p1 = op_5[1:0];
assign trunc_ln851_3_fu_766_p1 = op_11_V_fu_717_p3[2:0];
assign trunc_ln851_4_fu_984_p1 = op_13_V_fu_905_p3[3:0];
assign trunc_ln851_5_fu_1090_p0 = op_15;
assign trunc_ln851_5_fu_1090_p1 = op_15[4:0];
assign trunc_ln851_6_fu_1166_p0 = op_17;
assign trunc_ln851_6_fu_1166_p1 = op_17[2:0];
assign trunc_ln851_fu_269_p1 = ret_V_20_fu_245_p2[1:0];
assign zext_ln1192_fu_613_p1 = { 2'h0, ret_V_21_reg_1244[2], ret_V_21_reg_1244[2], ret_V_21_reg_1244[2], ret_V_21_reg_1244[2], ret_V_21_reg_1244[2], ret_V_21_reg_1244, 2'h0 };
assign zext_ln1393_fu_723_p1 = { 18'h00000, ret_V_22_reg_1250 };
assign zext_ln69_1_fu_1212_p1 = { 1'h0, ret_V_21_reg_1244[2], ret_V_21_reg_1244[2], ret_V_21_reg_1244[2], ret_V_21_reg_1244[2], ret_V_21_reg_1244[2], ret_V_21_reg_1244 };
assign zext_ln69_fu_1125_p1 = { 30'h00000000, op_16 };
assign \mul_4s_2s_6_1_1_U1.top_mul_4s_2s_6_1_1_Multiplier_0_U.a  = \mul_4s_2s_6_1_1_U1.din0 ;
assign \mul_4s_2s_6_1_1_U1.top_mul_4s_2s_6_1_1_Multiplier_0_U.b  = \mul_4s_2s_6_1_1_U1.din1 ;
assign \mul_4s_2s_6_1_1_U1.dout  = \mul_4s_2s_6_1_1_U1.top_mul_4s_2s_6_1_1_Multiplier_0_U.p ;
assign \mul_4s_2s_6_1_1_U1.din0  = op_5;
assign \mul_4s_2s_6_1_1_U1.din1  = op_4;
assign r_V_fu_309_p2 = \mul_4s_2s_6_1_1_U1.dout ;
endmodule


// Product machine:
module top_A_times_top_B (ap_start, op_0, op_10, op_14, op_15, op_16, op_17, op_18, op_4, op_5, op_6, ap_clk, unsafe_signal);
input ap_start;
input op_0;
input op_10;
input [3:0] op_14;
input [7:0] op_15;
input [1:0] op_16;
input [7:0] op_17;
input op_18;
input [1:0] op_4;
input [3:0] op_5;
input [1:0] op_6;
input ap_clk;
output unsafe_signal;
reg _setup;
initial _setup = 1'b0;
always @ (posedge ap_clk) _setup <= 1'b1;
reg ap_start_internal;
always @ (posedge ap_clk) if (!_setup) ap_start_internal <= ap_start;
reg op_0_internal;
always @ (posedge ap_clk) if (!_setup) op_0_internal <= op_0;
reg op_10_internal;
always @ (posedge ap_clk) if (!_setup) op_10_internal <= op_10;
reg [3:0] op_14_internal;
always @ (posedge ap_clk) if (!_setup) op_14_internal <= op_14;
reg [7:0] op_15_internal;
always @ (posedge ap_clk) if (!_setup) op_15_internal <= op_15;
reg [1:0] op_16_internal;
always @ (posedge ap_clk) if (!_setup) op_16_internal <= op_16;
reg [7:0] op_17_internal;
always @ (posedge ap_clk) if (!_setup) op_17_internal <= op_17;
reg op_18_internal;
always @ (posedge ap_clk) if (!_setup) op_18_internal <= op_18;
reg [1:0] op_4_internal;
always @ (posedge ap_clk) if (!_setup) op_4_internal <= op_4;
reg [3:0] op_5_internal;
always @ (posedge ap_clk) if (!_setup) op_5_internal <= op_5;
reg [1:0] op_6_internal;
always @ (posedge ap_clk) if (!_setup) op_6_internal <= op_6;
wire ap_done_A;
wire ap_done_B;
wire ap_done_eq;
assign ap_done_eq = ap_done_A == ap_done_B;
wire ap_idle_A;
wire ap_idle_B;
wire ap_idle_eq;
assign ap_idle_eq = ap_idle_A == ap_idle_B;
wire ap_ready_A;
wire ap_ready_B;
wire ap_ready_eq;
assign ap_ready_eq = ap_ready_A == ap_ready_B;
wire [31:0] op_29_A;
wire [31:0] op_29_B;
wire op_29_eq;
assign op_29_eq = op_29_A == op_29_B;
wire op_29_ap_vld_A;
wire op_29_ap_vld_B;
wire clk_enable_A;
wire clk_enable_B;
assign clk_enable_A = _setup & (~op_29_ap_vld_A | op_29_ap_vld_B);
assign clk_enable_B = _setup;
wire divergent;
assign divergent = ~(ap_done_eq & ap_idle_eq & ap_ready_eq & op_29_eq);
assign unsafe_signal = op_29_ap_vld_A & op_29_ap_vld_B & divergent;
top_A instance_A (
    .ap_clk(ap_clk),
    .clk_enable(clk_enable_A),
    .ap_start(ap_start_internal),
    .op_0(op_0_internal),
    .op_10(op_10_internal),
    .op_14(op_14_internal),
    .op_15(op_15_internal),
    .op_16(op_16_internal),
    .op_17(op_17_internal),
    .op_18(op_18_internal),
    .op_4(op_4_internal),
    .op_5(op_5_internal),
    .op_6(op_6_internal),
    .ap_done(ap_done_A),
    .ap_idle(ap_idle_A),
    .ap_ready(ap_ready_A),
    .op_29(op_29_A),
    .op_29_ap_vld(op_29_ap_vld_A)
);
top_B instance_B (
    .ap_clk(ap_clk),
    .clk_enable(clk_enable_B),
    .ap_start(ap_start_internal),
    .op_0(op_0_internal),
    .op_10(op_10_internal),
    .op_14(op_14_internal),
    .op_15(op_15_internal),
    .op_16(op_16_internal),
    .op_17(op_17_internal),
    .op_18(op_18_internal),
    .op_4(op_4_internal),
    .op_5(op_5_internal),
    .op_6(op_6_internal),
    .ap_done(ap_done_B),
    .ap_idle(ap_idle_B),
    .ap_ready(ap_ready_B),
    .op_29(op_29_B),
    .op_29_ap_vld(op_29_ap_vld_B)
);
endmodule
