// Processed by function `construct_kairos` in `verilog_tricks.py`.
// Machine A:
// Processed by function `add_clk_enable_signal` in `verilog_tricks.py`.
// Processed by function `remove_reset_signal` in `verilog_tricks.py`.
module top_A (
  ap_clk,
  ap_start,
  ap_done,
  ap_idle,
  ap_ready,
  op_0,
  op_1,
  op_2,
  op_6,
  op_10,
  op_12,
  op_13,
  op_15,
  op_16,
  op_18,
  op_19,
  op_31,
  op_31_ap_vld,
clk_enable
);
input clk_enable;


input ap_clk;
wire ap_rst;
assign ap_rst = op_31_ap_vld;
input ap_start;
input [7:0] op_0;
input [3:0] op_1;
input [1:0] op_10;
input [3:0] op_12;
input [1:0] op_13;
input [31:0] op_15;
input [31:0] op_16;
input [3:0] op_18;
input [31:0] op_19;
input op_2;
input op_6;
output ap_done;
output ap_idle;
output ap_ready;
output [31:0] op_31;
output op_31_ap_vld;


reg [31:0] add_ln691_3_reg_987;
reg [31:0] add_ln69_reg_931;
reg [7:0] ap_CS_fsm = 8'h01;
reg icmp_ln851_1_reg_951;
reg icmp_ln851_3_reg_982;
reg [31:0] op_27_V_reg_966;
reg op_3_V_reg_912;
reg r_1_reg_925;
reg [3:0] r_reg_920;
reg [13:0] ret_V_16_reg_941;
reg [31:0] ret_V_19_reg_961;
reg [31:0] ret_V_20_cast_reg_976;
reg [42:0] ret_V_21_reg_971;
reg [4:0] ret_V_4_reg_936;
reg [31:0] tmp_5_reg_956;
reg [6:0] tmp_reg_946;
wire [31:0] _000_;
wire [31:0] _001_;
wire [7:0] _002_;
wire _003_;
wire _004_;
wire [31:0] _005_;
wire _006_;
wire _007_;
wire [3:0] _008_;
wire [13:0] _009_;
wire [31:0] _010_;
wire [31:0] _011_;
wire [42:0] _012_;
wire [4:0] _013_;
wire [31:0] _014_;
wire [6:0] _015_;
wire [1:0] _016_;
wire _017_;
wire _018_;
wire _019_;
wire _020_;
wire _021_;
wire _022_;
wire _023_;
wire _024_;
wire _025_;
wire _026_;
wire _027_;
wire _028_;
wire _029_;
wire _030_;
wire _031_;
wire _032_;
wire _033_;
wire _034_;
wire _035_;
wire [31:0] add_ln691_2_fu_748_p2;
wire [31:0] add_ln691_3_fu_825_p2;
wire [7:0] add_ln691_fu_636_p2;
wire [31:0] add_ln69_fu_390_p2;
wire and_ln340_fu_303_p2;
wire and_ln785_1_fu_333_p2;
wire and_ln785_fu_327_p2;
wire ap_CS_fsm_state1;
wire ap_CS_fsm_state2;
wire ap_CS_fsm_state3;
wire ap_CS_fsm_state4;
wire ap_CS_fsm_state5;
wire ap_CS_fsm_state6;
wire ap_CS_fsm_state7;
wire ap_CS_fsm_state8;
wire [7:0] ap_NS_fsm;
wire ap_clk;
wire ap_done;
wire ap_idle;
wire ap_ready;
wire ap_rst;
wire ap_start;
wire icmp_ln768_1_fu_486_p2;
wire icmp_ln768_fu_249_p2;
wire icmp_ln786_1_fu_509_p2;
wire icmp_ln786_fu_279_p2;
wire icmp_ln851_1_fu_613_p2;
wire icmp_ln851_2_fu_742_p2;
wire icmp_ln851_3_fu_819_p2;
wire icmp_ln851_fu_436_p2;
wire newsignbit_fu_235_p1;
wire [7:0] op_0;
wire [3:0] op_1;
wire [1:0] op_10;
wire [5:0] op_11_V_fu_619_p3;
wire [3:0] op_12;
wire [1:0] op_13;
wire [31:0] op_15;
wire [31:0] op_16;
wire [2:0] op_17_V_fu_838_p1;
wire [3:0] op_18;
wire [31:0] op_19;
wire op_2;
wire [7:0] op_22_V_fu_661_p2;
wire [31:0] op_27_V_fu_779_p2;
wire [31:0] op_29_V_fu_879_p4;
wire [31:0] op_31;
wire op_31_ap_vld;
wire op_3_V_fu_345_p2;
wire op_6;
wire [7:0] op_9_V_fu_540_p3;
wire or_ln340_fu_291_p2;
wire or_ln384_fu_534_p2;
wire or_ln785_1_fu_492_p2;
wire or_ln785_2_fu_321_p2;
wire or_ln785_3_fu_339_p2;
wire or_ln785_fu_255_p2;
wire or_ln786_1_fu_515_p2;
wire or_ln786_fu_285_p2;
wire overflow_1_fu_498_p2;
wire overflow_fu_267_p2;
wire [3:0] p_Result_1_fu_476_p4;
wire p_Result_5_fu_629_p3;
wire p_Result_6_fu_730_p3;
wire p_Result_7_fu_842_p3;
wire p_Result_8_fu_227_p3;
wire p_Result_9_fu_470_p2;
wire p_Result_s_18_fu_424_p3;
wire [2:0] p_Result_s_fu_239_p4;
wire [32:0] p_Val2_11_fu_873_p2;
wire [7:0] p_Val2_3_fu_462_p3;
wire [32:0] p_Val2_6_fu_683_p2;
wire r_1_fu_367_p2;
wire [3:0] r_fu_356_p3;
wire [1:0] ret_2_fu_372_p3;
wire [8:0] ret_V_14_fu_408_p2;
wire [4:0] ret_V_15_fu_451_p3;
wire [13:0] ret_V_16_fu_593_p2;
wire [31:0] ret_V_17_cast_fu_720_p4;
wire [7:0] ret_V_17_fu_649_p3;
wire [35:0] ret_V_18_fu_714_p2;
wire [31:0] ret_V_19_fu_762_p3;
wire [31:0] ret_V_20_cast_fu_805_p4;
wire [31:0] ret_V_20_fu_774_p2;
wire [42:0] ret_V_21_fu_799_p2;
wire [31:0] ret_V_22_fu_893_p2;
wire [5:0] ret_V_2_fu_442_p2;
wire [4:0] ret_V_4_fu_555_p2;
wire [5:0] ret_V_fu_414_p4;
wire [1:0] ret_fu_380_p2;
wire [12:0] rhs_1_fu_581_p3;
wire [32:0] rhs_2_fu_679_p1;
wire [34:0] rhs_3_fu_703_p3;
wire [41:0] rhs_6_fu_788_p3;
wire [32:0] rhs_7_fu_865_p3;
wire select_ln1192_fu_400_p0;
wire [8:0] select_ln1192_fu_400_p3;
wire [4:0] select_ln1193_fu_548_p3;
wire [31:0] select_ln353_fu_858_p3;
wire [7:0] select_ln384_fu_526_p3;
wire [7:0] select_ln850_1_fu_642_p3;
wire [31:0] select_ln850_2_fu_754_p3;
wire [5:0] select_ln850_3_fu_573_p3;
wire [31:0] select_ln850_4_fu_853_p3;
wire [5:0] select_ln850_fu_565_p3;
wire [13:0] sext_ln1192_1_fu_589_p1;
wire [32:0] sext_ln1192_2_fu_667_p1;
wire [35:0] sext_ln1192_3_fu_710_p1;
wire [31:0] sext_ln1192_4_fu_770_p1;
wire [42:0] sext_ln1192_5_fu_795_p1;
wire [31:0] sext_ln1192_6_fu_889_p1;
wire [13:0] sext_ln1192_fu_561_p1;
wire [3:0] sext_ln703_1_fu_699_p0;
wire [35:0] sext_ln703_1_fu_699_p1;
wire [31:0] sext_ln703_2_fu_784_p0;
wire [42:0] sext_ln703_2_fu_784_p1;
wire [8:0] sext_ln703_fu_396_p1;
wire [7:0] sext_ln850_fu_626_p1;
wire [3:0] shl_ln1497_fu_351_p2;
wire [1:0] tmp_4_fu_831_p3;
wire [8:0] tmp_6_fu_671_p3;
wire [1:0] trunc_ln1497_fu_363_p1;
wire trunc_ln728_fu_458_p1;
wire [6:0] trunc_ln851_1_fu_609_p1;
wire [3:0] trunc_ln851_2_fu_738_p0;
wire [2:0] trunc_ln851_2_fu_738_p1;
wire [31:0] trunc_ln851_3_fu_815_p0;
wire [9:0] trunc_ln851_3_fu_815_p1;
wire [2:0] trunc_ln851_fu_432_p1;
wire underflow_1_fu_521_p2;
wire xor_ln340_fu_297_p2;
wire xor_ln785_1_fu_315_p2;
wire xor_ln785_fu_261_p2;
wire xor_ln786_1_fu_503_p2;
wire xor_ln786_2_fu_309_p2;
wire xor_ln786_fu_273_p2;
wire [32:0] zext_ln1192_fu_849_p1;
wire [31:0] zext_ln69_1_fu_386_p1;
wire [7:0] zext_ln69_fu_657_p1;
wire [4:0] zext_ln703_fu_448_p1;


assign add_ln691_2_fu_748_p2 = ret_V_18_fu_714_p2[34:3] + 1'h1;
assign add_ln691_3_fu_825_p2 = ret_V_21_fu_799_p2[41:10] + 1'h1;
assign add_ln691_fu_636_p2 = $signed(tmp_reg_946) + $signed(2'h1);
assign add_ln69_fu_390_p2 = ret_fu_380_p2 + op_15;
assign op_22_V_fu_661_p2 = ret_V_17_fu_649_p3 + op_10;
assign op_27_V_fu_779_p2 = add_ln69_reg_931 + ret_V_20_fu_774_p2;
assign op_31 = ret_V_22_fu_893_p2 + op_19;
assign p_Val2_11_fu_873_p2 = { select_ln353_fu_858_p3, 1'h0 } + { r_1_reg_925, r_1_reg_925, 1'h0 };
assign { p_Val2_6_fu_683_p2[32], p_Val2_6_fu_683_p2[8:0] } = $signed({ op_22_V_fu_661_p2, 1'h0 }) + $signed({ ret_V_4_reg_936, 1'h0 });
assign ret_V_14_fu_408_p2 = $signed(select_ln1192_fu_400_p3) + $signed(op_0);
assign ret_V_16_fu_593_p2 = $signed({ select_ln850_3_fu_573_p3, 7'h00 }) + $signed(op_9_V_fu_540_p3);
assign ret_V_18_fu_714_p2 = $signed({ tmp_5_reg_956, 3'h0 }) + $signed(op_12);
assign ret_V_20_fu_774_p2 = $signed(ret_V_19_reg_961) + $signed(op_13);
assign ret_V_21_fu_799_p2 = $signed({ op_27_V_reg_966, 10'h000 }) + $signed(op_16);
assign ret_V_22_fu_893_p2 = $signed(p_Val2_11_fu_873_p2[32:1]) + $signed(op_18);
assign ret_V_2_fu_442_p2 = ret_V_14_fu_408_p2[8:3] + 1'h1;
assign _017_ = ap_CS_fsm[0] & _019_;
assign _018_ = ap_CS_fsm[0] & ap_start;
assign and_ln340_fu_303_p2 = xor_ln340_fu_297_p2 & or_ln786_fu_285_p2;
assign and_ln785_1_fu_333_p2 = op_1[0] & and_ln785_fu_327_p2;
assign and_ln785_fu_327_p2 = xor_ln786_2_fu_309_p2 & or_ln785_2_fu_321_p2;
assign op_3_V_fu_345_p2 = or_ln785_3_fu_339_p2 & op_1[0];
assign overflow_1_fu_498_p2 = r_1_reg_925 & or_ln785_1_fu_492_p2;
assign overflow_fu_267_p2 = xor_ln785_fu_261_p2 & or_ln785_fu_255_p2;
assign ret_fu_380_p2 = r_fu_356_p3[1:0] & ret_2_fu_372_p3;
assign underflow_1_fu_521_p2 = or_ln786_1_fu_515_p2 & op_3_V_reg_912;
assign r_1_fu_367_p2 = ~ op_3_V_reg_912;
assign xor_ln786_fu_273_p2 = ~ op_1[0];
assign xor_ln785_fu_261_p2 = ~ op_1[3];
assign xor_ln340_fu_297_p2 = ~ or_ln340_fu_291_p2;
assign xor_ln785_1_fu_315_p2 = ~ or_ln785_fu_255_p2;
assign xor_ln786_2_fu_309_p2 = ~ icmp_ln786_fu_279_p2;
assign xor_ln786_1_fu_503_p2 = ~ p_Result_9_fu_470_p2;
assign _019_ = ~ ap_start;
assign _020_ = ! ret_V_14_fu_408_p2[2:0];
assign _021_ = | ret_V_15_fu_451_p3[4:1];
assign _022_ = | op_1[3:1];
assign _023_ = ret_V_15_fu_451_p3[4:1] != 4'hf;
assign _024_ = op_1[3:1] != 3'h7;
assign _025_ = | op_9_V_fu_540_p3[6:0];
assign _026_ = | op_12[2:0];
assign _027_ = | op_16[9:0];
assign or_ln340_fu_291_p2 = op_1[3] | overflow_fu_267_p2;
assign or_ln384_fu_534_p2 = underflow_1_fu_521_p2 | overflow_1_fu_498_p2;
assign or_ln785_1_fu_492_p2 = p_Result_9_fu_470_p2 | icmp_ln768_1_fu_486_p2;
assign or_ln785_2_fu_321_p2 = xor_ln785_1_fu_315_p2 | op_1[3];
assign or_ln785_3_fu_339_p2 = and_ln785_1_fu_333_p2 | and_ln340_fu_303_p2;
assign or_ln785_fu_255_p2 = op_1[0] | icmp_ln768_fu_249_p2;
assign or_ln786_1_fu_515_p2 = xor_ln786_1_fu_503_p2 | icmp_ln786_1_fu_509_p2;
assign or_ln786_fu_285_p2 = xor_ln786_fu_273_p2 | icmp_ln786_fu_279_p2;
always @(posedge ap_clk)
tmp_5_reg_956 <= _014_;
always @(posedge ap_clk)
ret_V_19_reg_961 <= _010_;
always @(posedge ap_clk)
op_3_V_reg_912 <= _006_;
always @(posedge ap_clk)
op_27_V_reg_966 <= _005_;
always @(posedge ap_clk)
ret_V_4_reg_936 <= _013_;
always @(posedge ap_clk)
ret_V_16_reg_941 <= _009_;
always @(posedge ap_clk)
tmp_reg_946 <= _015_;
always @(posedge ap_clk)
icmp_ln851_1_reg_951 <= _003_;
always @(posedge ap_clk)
r_reg_920 <= _008_;
always @(posedge ap_clk)
r_1_reg_925 <= _007_;
always @(posedge ap_clk)
add_ln69_reg_931 <= _001_;
always @(posedge ap_clk)
ret_V_21_reg_971 <= _012_;
always @(posedge ap_clk)
ret_V_20_cast_reg_976 <= _011_;
always @(posedge ap_clk)
icmp_ln851_3_reg_982 <= _004_;
always @(posedge ap_clk)
add_ln691_3_reg_987 <= _000_;
always @(posedge ap_clk)
ap_CS_fsm <= _002_;
assign _016_ = _018_ ? 2'h2 : 2'h1;
assign _028_ = ap_CS_fsm == 1'h1;
function [7:0] _104_;
input [7:0] a;
input [63:0] b;
input [7:0] s;
case (s)
8'b00000001:
_104_ = b[7:0];
8'b00000010:
_104_ = b[15:8];
8'b00000100:
_104_ = b[23:16];
8'b00001000:
_104_ = b[31:24];
8'b00010000:
_104_ = b[39:32];
8'b00100000:
_104_ = b[47:40];
8'b01000000:
_104_ = b[55:48];
8'b10000000:
_104_ = b[63:56];
8'b00000000:
_104_ = a;
default:
_104_ = 8'bx;
endcase
endfunction
assign ap_NS_fsm = _104_(8'hxx, { 6'h00, _016_, 56'h04081020408001 }, { _028_, _035_, _034_, _033_, _032_, _031_, _030_, _029_ });
assign _029_ = ap_CS_fsm == 8'h80;
assign _030_ = ap_CS_fsm == 7'h40;
assign _031_ = ap_CS_fsm == 6'h20;
assign _032_ = ap_CS_fsm == 5'h10;
assign _033_ = ap_CS_fsm == 4'h8;
assign _034_ = ap_CS_fsm == 3'h4;
assign _035_ = ap_CS_fsm == 2'h2;
assign op_31_ap_vld = ap_CS_fsm[7] ? 1'h1 : 1'h0;
assign ap_idle = _017_ ? 1'h1 : 1'h0;
assign _014_ = ap_CS_fsm[3] ? { p_Val2_6_fu_683_p2[32], p_Val2_6_fu_683_p2[32], p_Val2_6_fu_683_p2[32], p_Val2_6_fu_683_p2[32], p_Val2_6_fu_683_p2[32], p_Val2_6_fu_683_p2[32], p_Val2_6_fu_683_p2[32], p_Val2_6_fu_683_p2[32], p_Val2_6_fu_683_p2[32], p_Val2_6_fu_683_p2[32], p_Val2_6_fu_683_p2[32], p_Val2_6_fu_683_p2[32], p_Val2_6_fu_683_p2[32], p_Val2_6_fu_683_p2[32], p_Val2_6_fu_683_p2[32], p_Val2_6_fu_683_p2[32], p_Val2_6_fu_683_p2[32], p_Val2_6_fu_683_p2[32], p_Val2_6_fu_683_p2[32], p_Val2_6_fu_683_p2[32], p_Val2_6_fu_683_p2[32], p_Val2_6_fu_683_p2[32], p_Val2_6_fu_683_p2[32], p_Val2_6_fu_683_p2[32], p_Val2_6_fu_683_p2[8:1] } : tmp_5_reg_956;
assign _010_ = ap_CS_fsm[4] ? ret_V_19_fu_762_p3 : ret_V_19_reg_961;
assign _006_ = ap_CS_fsm[0] ? op_3_V_fu_345_p2 : op_3_V_reg_912;
assign _005_ = ap_CS_fsm[5] ? op_27_V_fu_779_p2 : op_27_V_reg_966;
assign _003_ = ap_CS_fsm[2] ? icmp_ln851_1_fu_613_p2 : icmp_ln851_1_reg_951;
assign _015_ = ap_CS_fsm[2] ? ret_V_16_fu_593_p2[13:7] : tmp_reg_946;
assign _009_ = ap_CS_fsm[2] ? ret_V_16_fu_593_p2 : ret_V_16_reg_941;
assign _013_ = ap_CS_fsm[2] ? ret_V_4_fu_555_p2 : ret_V_4_reg_936;
assign _001_ = ap_CS_fsm[1] ? add_ln69_fu_390_p2 : add_ln69_reg_931;
assign _007_ = ap_CS_fsm[1] ? r_1_fu_367_p2 : r_1_reg_925;
assign _008_ = ap_CS_fsm[1] ? r_fu_356_p3 : r_reg_920;
assign _000_ = ap_CS_fsm[6] ? add_ln691_3_fu_825_p2 : add_ln691_3_reg_987;
assign _004_ = ap_CS_fsm[6] ? icmp_ln851_3_fu_819_p2 : icmp_ln851_3_reg_982;
assign _011_ = ap_CS_fsm[6] ? ret_V_21_fu_799_p2[41:10] : ret_V_20_cast_reg_976;
assign _012_ = ap_CS_fsm[6] ? ret_V_21_fu_799_p2 : ret_V_21_reg_971;
assign _002_ = ap_rst ? 8'h01 : ap_NS_fsm;
assign ret_V_4_fu_555_p2 = select_ln1193_fu_548_p3 - r_reg_920;
assign icmp_ln768_1_fu_486_p2 = _021_ ? 1'h1 : 1'h0;
assign icmp_ln768_fu_249_p2 = _022_ ? 1'h1 : 1'h0;
assign icmp_ln786_1_fu_509_p2 = _023_ ? 1'h1 : 1'h0;
assign icmp_ln786_fu_279_p2 = _024_ ? 1'h1 : 1'h0;
assign icmp_ln851_1_fu_613_p2 = _025_ ? 1'h1 : 1'h0;
assign icmp_ln851_2_fu_742_p2 = _026_ ? 1'h1 : 1'h0;
assign icmp_ln851_3_fu_819_p2 = _027_ ? 1'h1 : 1'h0;
assign icmp_ln851_fu_436_p2 = _020_ ? 1'h1 : 1'h0;
assign op_9_V_fu_540_p3 = or_ln384_fu_534_p2 ? select_ln384_fu_526_p3 : { ret_V_15_fu_451_p3[0], 7'h00 };
assign p_Result_9_fu_470_p2 = ret_V_15_fu_451_p3[0] ? 1'h1 : 1'h0;
assign r_fu_356_p3 = op_2 ? { op_1[2:0], 1'h0 } : op_1;
assign ret_2_fu_372_p3 = op_3_V_reg_912 ? 2'h0 : 2'h3;
assign ret_V_15_fu_451_p3 = op_3_V_reg_912 ? 5'h1f : { 1'h0, r_reg_920 };
assign ret_V_17_fu_649_p3 = ret_V_16_reg_941[13] ? select_ln850_1_fu_642_p3 : { tmp_reg_946[6], tmp_reg_946 };
assign ret_V_19_fu_762_p3 = ret_V_18_fu_714_p2[35] ? select_ln850_2_fu_754_p3 : ret_V_18_fu_714_p2[34:3];
assign select_ln1192_fu_400_p3 = op_6 ? 9'h1f8 : 9'h000;
assign select_ln1193_fu_548_p3 = op_3_V_reg_912 ? 5'h1f : 5'h00;
assign select_ln353_fu_858_p3 = ret_V_21_reg_971[42] ? select_ln850_4_fu_853_p3 : ret_V_20_cast_reg_976;
assign select_ln384_fu_526_p3 = overflow_1_fu_498_p2 ? 8'h7f : 8'h80;
assign select_ln850_1_fu_642_p3 = icmp_ln851_1_reg_951 ? add_ln691_fu_636_p2 : { tmp_reg_946[6], tmp_reg_946 };
assign select_ln850_2_fu_754_p3 = icmp_ln851_2_fu_742_p2 ? add_ln691_2_fu_748_p2 : ret_V_18_fu_714_p2[34:3];
assign select_ln850_3_fu_573_p3 = ret_V_14_fu_408_p2[8] ? select_ln850_fu_565_p3 : { 1'h0, ret_V_14_fu_408_p2[7:3] };
assign select_ln850_4_fu_853_p3 = icmp_ln851_3_reg_982 ? add_ln691_3_reg_987 : ret_V_20_cast_reg_976;
assign select_ln850_fu_565_p3 = icmp_ln851_fu_436_p2 ? { 1'h1, ret_V_14_fu_408_p2[7:3] } : ret_V_2_fu_442_p2;
assign ap_CS_fsm_state1 = ap_CS_fsm[0];
assign ap_CS_fsm_state2 = ap_CS_fsm[1];
assign ap_CS_fsm_state3 = ap_CS_fsm[2];
assign ap_CS_fsm_state4 = ap_CS_fsm[3];
assign ap_CS_fsm_state5 = ap_CS_fsm[4];
assign ap_CS_fsm_state6 = ap_CS_fsm[5];
assign ap_CS_fsm_state7 = ap_CS_fsm[6];
assign ap_CS_fsm_state8 = ap_CS_fsm[7];
assign ap_done = op_31_ap_vld;
assign ap_ready = op_31_ap_vld;
assign newsignbit_fu_235_p1 = op_1[0];
assign op_11_V_fu_619_p3 = { ret_V_4_reg_936, 1'h0 };
assign op_17_V_fu_838_p1 = { r_1_reg_925, r_1_reg_925, 1'h0 };
assign op_29_V_fu_879_p4 = p_Val2_11_fu_873_p2[32:1];
assign p_Result_1_fu_476_p4 = ret_V_15_fu_451_p3[4:1];
assign p_Result_5_fu_629_p3 = ret_V_16_reg_941[13];
assign p_Result_6_fu_730_p3 = ret_V_18_fu_714_p2[35];
assign p_Result_7_fu_842_p3 = ret_V_21_reg_971[42];
assign p_Result_8_fu_227_p3 = op_1[3];
assign p_Result_s_18_fu_424_p3 = ret_V_14_fu_408_p2[8];
assign p_Result_s_fu_239_p4 = op_1[3:1];
assign p_Val2_3_fu_462_p3 = { ret_V_15_fu_451_p3[0], 7'h00 };
assign p_Val2_6_fu_683_p2[31:9] = { p_Val2_6_fu_683_p2[32], p_Val2_6_fu_683_p2[32], p_Val2_6_fu_683_p2[32], p_Val2_6_fu_683_p2[32], p_Val2_6_fu_683_p2[32], p_Val2_6_fu_683_p2[32], p_Val2_6_fu_683_p2[32], p_Val2_6_fu_683_p2[32], p_Val2_6_fu_683_p2[32], p_Val2_6_fu_683_p2[32], p_Val2_6_fu_683_p2[32], p_Val2_6_fu_683_p2[32], p_Val2_6_fu_683_p2[32], p_Val2_6_fu_683_p2[32], p_Val2_6_fu_683_p2[32], p_Val2_6_fu_683_p2[32], p_Val2_6_fu_683_p2[32], p_Val2_6_fu_683_p2[32], p_Val2_6_fu_683_p2[32], p_Val2_6_fu_683_p2[32], p_Val2_6_fu_683_p2[32], p_Val2_6_fu_683_p2[32], p_Val2_6_fu_683_p2[32] };
assign ret_V_17_cast_fu_720_p4 = ret_V_18_fu_714_p2[34:3];
assign ret_V_20_cast_fu_805_p4 = ret_V_21_fu_799_p2[41:10];
assign ret_V_fu_414_p4 = ret_V_14_fu_408_p2[8:3];
assign rhs_1_fu_581_p3 = { select_ln850_3_fu_573_p3, 7'h00 };
assign rhs_2_fu_679_p1 = { op_22_V_fu_661_p2[7], op_22_V_fu_661_p2[7], op_22_V_fu_661_p2[7], op_22_V_fu_661_p2[7], op_22_V_fu_661_p2[7], op_22_V_fu_661_p2[7], op_22_V_fu_661_p2[7], op_22_V_fu_661_p2[7], op_22_V_fu_661_p2[7], op_22_V_fu_661_p2[7], op_22_V_fu_661_p2[7], op_22_V_fu_661_p2[7], op_22_V_fu_661_p2[7], op_22_V_fu_661_p2[7], op_22_V_fu_661_p2[7], op_22_V_fu_661_p2[7], op_22_V_fu_661_p2[7], op_22_V_fu_661_p2[7], op_22_V_fu_661_p2[7], op_22_V_fu_661_p2[7], op_22_V_fu_661_p2[7], op_22_V_fu_661_p2[7], op_22_V_fu_661_p2[7], op_22_V_fu_661_p2[7], op_22_V_fu_661_p2, 1'h0 };
assign rhs_3_fu_703_p3 = { tmp_5_reg_956, 3'h0 };
assign rhs_6_fu_788_p3 = { op_27_V_reg_966, 10'h000 };
assign rhs_7_fu_865_p3 = { select_ln353_fu_858_p3, 1'h0 };
assign select_ln1192_fu_400_p0 = op_6;
assign sext_ln1192_1_fu_589_p1 = { select_ln850_3_fu_573_p3[5], select_ln850_3_fu_573_p3, 7'h00 };
assign sext_ln1192_2_fu_667_p1 = { ret_V_4_reg_936[4], ret_V_4_reg_936[4], ret_V_4_reg_936[4], ret_V_4_reg_936[4], ret_V_4_reg_936[4], ret_V_4_reg_936[4], ret_V_4_reg_936[4], ret_V_4_reg_936[4], ret_V_4_reg_936[4], ret_V_4_reg_936[4], ret_V_4_reg_936[4], ret_V_4_reg_936[4], ret_V_4_reg_936[4], ret_V_4_reg_936[4], ret_V_4_reg_936[4], ret_V_4_reg_936[4], ret_V_4_reg_936[4], ret_V_4_reg_936[4], ret_V_4_reg_936[4], ret_V_4_reg_936[4], ret_V_4_reg_936[4], ret_V_4_reg_936[4], ret_V_4_reg_936[4], ret_V_4_reg_936[4], ret_V_4_reg_936[4], ret_V_4_reg_936[4], ret_V_4_reg_936[4], ret_V_4_reg_936, 1'h0 };
assign sext_ln1192_3_fu_710_p1 = { tmp_5_reg_956[31], tmp_5_reg_956, 3'h0 };
assign sext_ln1192_4_fu_770_p1 = { op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13 };
assign sext_ln1192_5_fu_795_p1 = { op_27_V_reg_966[31], op_27_V_reg_966, 10'h000 };
assign sext_ln1192_6_fu_889_p1 = { op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18 };
assign sext_ln1192_fu_561_p1 = { op_9_V_fu_540_p3[7], op_9_V_fu_540_p3[7], op_9_V_fu_540_p3[7], op_9_V_fu_540_p3[7], op_9_V_fu_540_p3[7], op_9_V_fu_540_p3[7], op_9_V_fu_540_p3 };
assign sext_ln703_1_fu_699_p0 = op_12;
assign sext_ln703_1_fu_699_p1 = { op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12 };
assign sext_ln703_2_fu_784_p0 = op_16;
assign sext_ln703_2_fu_784_p1 = { op_16[31], op_16[31], op_16[31], op_16[31], op_16[31], op_16[31], op_16[31], op_16[31], op_16[31], op_16[31], op_16[31], op_16 };
assign sext_ln703_fu_396_p1 = { op_0[7], op_0 };
assign sext_ln850_fu_626_p1 = { tmp_reg_946[6], tmp_reg_946 };
assign shl_ln1497_fu_351_p2 = { op_1[2:0], 1'h0 };
assign tmp_4_fu_831_p3 = { r_1_reg_925, 1'h0 };
assign tmp_6_fu_671_p3 = { op_22_V_fu_661_p2, 1'h0 };
assign trunc_ln1497_fu_363_p1 = r_fu_356_p3[1:0];
assign trunc_ln728_fu_458_p1 = ret_V_15_fu_451_p3[0];
assign trunc_ln851_1_fu_609_p1 = op_9_V_fu_540_p3[6:0];
assign trunc_ln851_2_fu_738_p0 = op_12;
assign trunc_ln851_2_fu_738_p1 = op_12[2:0];
assign trunc_ln851_3_fu_815_p0 = op_16;
assign trunc_ln851_3_fu_815_p1 = op_16[9:0];
assign trunc_ln851_fu_432_p1 = ret_V_14_fu_408_p2[2:0];
assign zext_ln1192_fu_849_p1 = { 30'h00000000, r_1_reg_925, r_1_reg_925, 1'h0 };
assign zext_ln69_1_fu_386_p1 = { 30'h00000000, ret_fu_380_p2 };
assign zext_ln69_fu_657_p1 = { 6'h00, op_10 };
assign zext_ln703_fu_448_p1 = { 1'h0, r_reg_920 };
endmodule


// Machine B:
// Processed by function `add_clk_enable_signal` in `verilog_tricks.py`.
// Processed by function `remove_reset_signal` in `verilog_tricks.py`.
module top_B (
  ap_clk,
  ap_start,
  ap_done,
  ap_idle,
  ap_ready,
  op_0,
  op_1,
  op_2,
  op_6,
  op_10,
  op_12,
  op_13,
  op_15,
  op_16,
  op_18,
  op_19,
  op_31,
  op_31_ap_vld,
clk_enable
);
input clk_enable;


input ap_clk;
wire ap_rst;
assign ap_rst = op_31_ap_vld;
input ap_start;
input [7:0] op_0;
input [3:0] op_1;
input [1:0] op_10;
input [3:0] op_12;
input [1:0] op_13;
input [31:0] op_15;
input [31:0] op_16;
input [3:0] op_18;
input [31:0] op_19;
input op_2;
input op_6;
output ap_done;
output ap_idle;
output ap_ready;
output [31:0] op_31;
output op_31_ap_vld;


reg [6:0] \add_14s_14s_14_2_1_U4.top_add_14s_14s_14_2_1_Adder_3_U.ain_s1 ;
reg [6:0] \add_14s_14s_14_2_1_U4.top_add_14s_14s_14_2_1_Adder_3_U.bin_s1 ;
reg \add_14s_14s_14_2_1_U4.top_add_14s_14s_14_2_1_Adder_3_U.carry_s1 ;
reg [6:0] \add_14s_14s_14_2_1_U4.top_add_14s_14s_14_2_1_Adder_3_U.sum_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.ain_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.bin_s1 ;
reg \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.carry_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.sum_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_8_U.ain_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_8_U.bin_s1 ;
reg \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_8_U.carry_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_8_U.sum_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_8_U.ain_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_8_U.bin_s1 ;
reg \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_8_U.carry_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_8_U.sum_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.ain_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.bin_s1 ;
reg \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.carry_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.sum_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_8_U.ain_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_8_U.bin_s1 ;
reg \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_8_U.carry_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_8_U.sum_s1 ;
reg [15:0] \add_32ns_32s_32_2_1_U10.top_add_32ns_32s_32_2_1_Adder_9_U.ain_s1 ;
reg [15:0] \add_32ns_32s_32_2_1_U10.top_add_32ns_32s_32_2_1_Adder_9_U.bin_s1 ;
reg \add_32ns_32s_32_2_1_U10.top_add_32ns_32s_32_2_1_Adder_9_U.carry_s1 ;
reg [15:0] \add_32ns_32s_32_2_1_U10.top_add_32ns_32s_32_2_1_Adder_9_U.sum_s1 ;
reg [15:0] \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.ain_s1 ;
reg [15:0] \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.bin_s1 ;
reg \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.carry_s1 ;
reg [15:0] \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.sum_s1 ;
reg [16:0] \add_33ns_33ns_33_2_1_U15.top_add_33ns_33ns_33_2_1_Adder_11_U.ain_s1 ;
reg [16:0] \add_33ns_33ns_33_2_1_U15.top_add_33ns_33ns_33_2_1_Adder_11_U.bin_s1 ;
reg \add_33ns_33ns_33_2_1_U15.top_add_33ns_33ns_33_2_1_Adder_11_U.carry_s1 ;
reg [15:0] \add_33ns_33ns_33_2_1_U15.top_add_33ns_33ns_33_2_1_Adder_11_U.sum_s1 ;
reg [16:0] \add_33s_33s_33_2_1_U7.top_add_33s_33s_33_2_1_Adder_6_U.ain_s1 ;
reg [16:0] \add_33s_33s_33_2_1_U7.top_add_33s_33s_33_2_1_Adder_6_U.bin_s1 ;
reg \add_33s_33s_33_2_1_U7.top_add_33s_33s_33_2_1_Adder_6_U.carry_s1 ;
reg [15:0] \add_33s_33s_33_2_1_U7.top_add_33s_33s_33_2_1_Adder_6_U.sum_s1 ;
reg [17:0] \add_36s_36s_36_2_1_U8.top_add_36s_36s_36_2_1_Adder_7_U.ain_s1 ;
reg [17:0] \add_36s_36s_36_2_1_U8.top_add_36s_36s_36_2_1_Adder_7_U.bin_s1 ;
reg \add_36s_36s_36_2_1_U8.top_add_36s_36s_36_2_1_Adder_7_U.carry_s1 ;
reg [17:0] \add_36s_36s_36_2_1_U8.top_add_36s_36s_36_2_1_Adder_7_U.sum_s1 ;
reg [21:0] \add_43s_43s_43_2_1_U13.top_add_43s_43s_43_2_1_Adder_10_U.ain_s1 ;
reg [21:0] \add_43s_43s_43_2_1_U13.top_add_43s_43s_43_2_1_Adder_10_U.bin_s1 ;
reg \add_43s_43s_43_2_1_U13.top_add_43s_43s_43_2_1_Adder_10_U.carry_s1 ;
reg [20:0] \add_43s_43s_43_2_1_U13.top_add_43s_43s_43_2_1_Adder_10_U.sum_s1 ;
reg [2:0] \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.ain_s1 ;
reg [2:0] \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.bin_s1 ;
reg \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.carry_s1 ;
reg [2:0] \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.sum_s1 ;
reg [3:0] \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.ain_s1 ;
reg [3:0] \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.bin_s1 ;
reg \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.carry_s1 ;
reg [3:0] \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.sum_s1 ;
reg [3:0] \add_8s_8ns_8_2_1_U5.top_add_8s_8ns_8_2_1_Adder_4_U.ain_s1 ;
reg [3:0] \add_8s_8ns_8_2_1_U5.top_add_8s_8ns_8_2_1_Adder_4_U.bin_s1 ;
reg \add_8s_8ns_8_2_1_U5.top_add_8s_8ns_8_2_1_Adder_4_U.carry_s1 ;
reg [3:0] \add_8s_8ns_8_2_1_U5.top_add_8s_8ns_8_2_1_Adder_4_U.sum_s1 ;
reg [4:0] \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.ain_s1 ;
reg [4:0] \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.bin_s1 ;
reg \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.carry_s1 ;
reg [3:0] \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.sum_s1 ;
reg [31:0] add_ln691_2_reg_1115;
reg [31:0] add_ln691_3_reg_1182;
reg [7:0] add_ln691_reg_1053;
reg [31:0] add_ln69_reg_1145;
reg and_ln340_reg_891;
reg [36:0] ap_CS_fsm = 37'h0000000001;
reg icmp_ln768_1_reg_970;
reg icmp_ln768_reg_868;
reg icmp_ln786_1_reg_975;
reg icmp_ln786_reg_873;
reg icmp_ln851_1_reg_1026;
reg icmp_ln851_2_reg_1098;
reg icmp_ln851_3_reg_1165;
reg icmp_ln851_reg_954;
reg newsignbit_reg_860;
reg [7:0] op_22_V_reg_1068;
reg [31:0] op_27_V_reg_1150;
reg [31:0] op_29_V_reg_1202;
reg op_3_V_reg_901;
reg [7:0] op_9_V_reg_996;
reg or_ln785_reg_885;
reg overflow_1_reg_990;
reg [3:0] p_Result_1_reg_948;
reg p_Result_8_reg_853;
reg p_Result_9_reg_964;
reg [7:0] p_Val2_3_reg_959;
reg r_1_reg_931;
reg [3:0] r_reg_879;
reg [8:0] ret_V_14_reg_914;
reg [13:0] ret_V_16_reg_1036;
reg [31:0] ret_V_17_cast_reg_1108;
reg [7:0] ret_V_17_reg_1058;
reg [35:0] ret_V_18_reg_1103;
reg [31:0] ret_V_19_reg_1120;
reg [31:0] ret_V_20_cast_reg_1175;
reg [31:0] ret_V_20_reg_1140;
reg [42:0] ret_V_21_reg_1170;
reg [31:0] ret_V_22_reg_1212;
reg [5:0] ret_V_2_reg_985;
reg [4:0] ret_V_4_reg_1031;
reg [5:0] ret_V_reg_919;
reg [1:0] ret_reg_980;
reg [8:0] select_ln1192_reg_896;
reg [4:0] select_ln1193_reg_1001;
reg [31:0] select_ln353_reg_1187;
reg [5:0] select_ln850_3_reg_1006;
reg [7:0] sext_ln850_reg_1046;
reg [2:0] \sub_5ns_5ns_5_2_1_U3.top_sub_5ns_5ns_5_2_1_Adder_2_U.ain_s1 ;
reg [2:0] \sub_5ns_5ns_5_2_1_U3.top_sub_5ns_5ns_5_2_1_Adder_2_U.bin_s1 ;
reg \sub_5ns_5ns_5_2_1_U3.top_sub_5ns_5ns_5_2_1_Adder_2_U.carry_s1 ;
reg [1:0] \sub_5ns_5ns_5_2_1_U3.top_sub_5ns_5ns_5_2_1_Adder_2_U.sum_s1 ;
reg [31:0] tmp_5_reg_1083;
reg [6:0] tmp_reg_1041;
reg trunc_ln728_reg_943;
reg [6:0] trunc_ln851_1_reg_1011;
reg [2:0] trunc_ln851_reg_926;
reg [4:0] zext_ln703_reg_938;
wire [31:0] _000_;
wire [31:0] _001_;
wire [7:0] _002_;
wire [31:0] _003_;
wire _004_;
wire [36:0] _005_;
wire _006_;
wire _007_;
wire _008_;
wire _009_;
wire _010_;
wire _011_;
wire _012_;
wire _013_;
wire _014_;
wire [7:0] _015_;
wire [31:0] _016_;
wire [31:0] _017_;
wire _018_;
wire [7:0] _019_;
wire _020_;
wire _021_;
wire [3:0] _022_;
wire _023_;
wire _024_;
wire _025_;
wire _026_;
wire [3:0] _027_;
wire [8:0] _028_;
wire [13:0] _029_;
wire [31:0] _030_;
wire [7:0] _031_;
wire [35:0] _032_;
wire [31:0] _033_;
wire [31:0] _034_;
wire [31:0] _035_;
wire [42:0] _036_;
wire [31:0] _037_;
wire [5:0] _038_;
wire [4:0] _039_;
wire [5:0] _040_;
wire [1:0] _041_;
wire [5:0] _042_;
wire [4:0] _043_;
wire [31:0] _044_;
wire [5:0] _045_;
wire [7:0] _046_;
wire [31:0] _047_;
wire [6:0] _048_;
wire _049_;
wire [6:0] _050_;
wire [2:0] _051_;
wire [3:0] _052_;
wire [1:0] _053_;
wire _054_;
wire _055_;
wire _056_;
wire _057_;
wire _058_;
wire _059_;
wire _060_;
wire [6:0] _061_;
wire [6:0] _062_;
wire _063_;
wire [6:0] _064_;
wire [7:0] _065_;
wire [7:0] _066_;
wire [15:0] _067_;
wire [15:0] _068_;
wire _069_;
wire [15:0] _070_;
wire [16:0] _071_;
wire [16:0] _072_;
wire [15:0] _073_;
wire [15:0] _074_;
wire _075_;
wire [15:0] _076_;
wire [16:0] _077_;
wire [16:0] _078_;
wire [15:0] _079_;
wire [15:0] _080_;
wire _081_;
wire [15:0] _082_;
wire [16:0] _083_;
wire [16:0] _084_;
wire [15:0] _085_;
wire [15:0] _086_;
wire _087_;
wire [15:0] _088_;
wire [16:0] _089_;
wire [16:0] _090_;
wire [15:0] _091_;
wire [15:0] _092_;
wire _093_;
wire [15:0] _094_;
wire [16:0] _095_;
wire [16:0] _096_;
wire [15:0] _097_;
wire [15:0] _098_;
wire _099_;
wire [15:0] _100_;
wire [16:0] _101_;
wire [16:0] _102_;
wire [15:0] _103_;
wire [15:0] _104_;
wire _105_;
wire [15:0] _106_;
wire [16:0] _107_;
wire [16:0] _108_;
wire [16:0] _109_;
wire [16:0] _110_;
wire _111_;
wire [15:0] _112_;
wire [16:0] _113_;
wire [17:0] _114_;
wire [16:0] _115_;
wire [16:0] _116_;
wire _117_;
wire [15:0] _118_;
wire [16:0] _119_;
wire [17:0] _120_;
wire [17:0] _121_;
wire [17:0] _122_;
wire _123_;
wire [17:0] _124_;
wire [18:0] _125_;
wire [18:0] _126_;
wire [21:0] _127_;
wire [21:0] _128_;
wire _129_;
wire [20:0] _130_;
wire [21:0] _131_;
wire [22:0] _132_;
wire [2:0] _133_;
wire [2:0] _134_;
wire _135_;
wire [2:0] _136_;
wire [3:0] _137_;
wire [3:0] _138_;
wire [3:0] _139_;
wire [3:0] _140_;
wire _141_;
wire [3:0] _142_;
wire [4:0] _143_;
wire [4:0] _144_;
wire [3:0] _145_;
wire [3:0] _146_;
wire _147_;
wire [3:0] _148_;
wire [4:0] _149_;
wire [4:0] _150_;
wire [4:0] _151_;
wire [4:0] _152_;
wire _153_;
wire [3:0] _154_;
wire [4:0] _155_;
wire [5:0] _156_;
wire [2:0] _157_;
wire [2:0] _158_;
wire _159_;
wire [1:0] _160_;
wire [2:0] _161_;
wire [3:0] _162_;
wire _163_;
wire _164_;
wire _165_;
wire _166_;
wire _167_;
wire _168_;
wire _169_;
wire _170_;
wire _171_;
wire _172_;
wire _173_;
wire _174_;
wire _175_;
wire _176_;
wire _177_;
wire _178_;
wire _179_;
wire _180_;
wire _181_;
wire _182_;
wire _183_;
wire _184_;
wire _185_;
wire _186_;
wire _187_;
wire _188_;
wire _189_;
wire _190_;
wire _191_;
wire _192_;
wire _193_;
wire _194_;
wire _195_;
wire _196_;
wire _197_;
wire _198_;
wire _199_;
wire _200_;
wire _201_;
wire _202_;
wire _203_;
wire _204_;
wire _205_;
wire _206_;
wire \add_14s_14s_14_2_1_U4.ce ;
wire \add_14s_14s_14_2_1_U4.clk ;
wire [13:0] \add_14s_14s_14_2_1_U4.din0 ;
wire [13:0] \add_14s_14s_14_2_1_U4.din1 ;
wire [13:0] \add_14s_14s_14_2_1_U4.dout ;
wire \add_14s_14s_14_2_1_U4.reset ;
wire [13:0] \add_14s_14s_14_2_1_U4.top_add_14s_14s_14_2_1_Adder_3_U.a ;
wire [13:0] \add_14s_14s_14_2_1_U4.top_add_14s_14s_14_2_1_Adder_3_U.ain_s0 ;
wire [13:0] \add_14s_14s_14_2_1_U4.top_add_14s_14s_14_2_1_Adder_3_U.b ;
wire [13:0] \add_14s_14s_14_2_1_U4.top_add_14s_14s_14_2_1_Adder_3_U.bin_s0 ;
wire \add_14s_14s_14_2_1_U4.top_add_14s_14s_14_2_1_Adder_3_U.ce ;
wire \add_14s_14s_14_2_1_U4.top_add_14s_14s_14_2_1_Adder_3_U.clk ;
wire \add_14s_14s_14_2_1_U4.top_add_14s_14s_14_2_1_Adder_3_U.facout_s1 ;
wire \add_14s_14s_14_2_1_U4.top_add_14s_14s_14_2_1_Adder_3_U.facout_s2 ;
wire [6:0] \add_14s_14s_14_2_1_U4.top_add_14s_14s_14_2_1_Adder_3_U.fas_s1 ;
wire [6:0] \add_14s_14s_14_2_1_U4.top_add_14s_14s_14_2_1_Adder_3_U.fas_s2 ;
wire \add_14s_14s_14_2_1_U4.top_add_14s_14s_14_2_1_Adder_3_U.reset ;
wire [13:0] \add_14s_14s_14_2_1_U4.top_add_14s_14s_14_2_1_Adder_3_U.s ;
wire [6:0] \add_14s_14s_14_2_1_U4.top_add_14s_14s_14_2_1_Adder_3_U.u1.a ;
wire [6:0] \add_14s_14s_14_2_1_U4.top_add_14s_14s_14_2_1_Adder_3_U.u1.b ;
wire \add_14s_14s_14_2_1_U4.top_add_14s_14s_14_2_1_Adder_3_U.u1.cin ;
wire \add_14s_14s_14_2_1_U4.top_add_14s_14s_14_2_1_Adder_3_U.u1.cout ;
wire [6:0] \add_14s_14s_14_2_1_U4.top_add_14s_14s_14_2_1_Adder_3_U.u1.s ;
wire [6:0] \add_14s_14s_14_2_1_U4.top_add_14s_14s_14_2_1_Adder_3_U.u2.a ;
wire [6:0] \add_14s_14s_14_2_1_U4.top_add_14s_14s_14_2_1_Adder_3_U.u2.b ;
wire \add_14s_14s_14_2_1_U4.top_add_14s_14s_14_2_1_Adder_3_U.u2.cin ;
wire \add_14s_14s_14_2_1_U4.top_add_14s_14s_14_2_1_Adder_3_U.u2.cout ;
wire [6:0] \add_14s_14s_14_2_1_U4.top_add_14s_14s_14_2_1_Adder_3_U.u2.s ;
wire \add_32ns_32ns_32_2_1_U11.ce ;
wire \add_32ns_32ns_32_2_1_U11.clk ;
wire [31:0] \add_32ns_32ns_32_2_1_U11.din0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U11.din1 ;
wire [31:0] \add_32ns_32ns_32_2_1_U11.dout ;
wire \add_32ns_32ns_32_2_1_U11.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.a ;
wire [31:0] \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.ain_s0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.b ;
wire [31:0] \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.bin_s0 ;
wire \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.ce ;
wire \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.clk ;
wire \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.facout_s1 ;
wire \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.facout_s2 ;
wire [15:0] \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.fas_s1 ;
wire [15:0] \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.fas_s2 ;
wire \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.u1.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.u1.b ;
wire \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.u1.cin ;
wire \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.u1.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.u1.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.u2.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.u2.b ;
wire \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.u2.cin ;
wire \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.u2.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.u2.s ;
wire \add_32ns_32ns_32_2_1_U12.ce ;
wire \add_32ns_32ns_32_2_1_U12.clk ;
wire [31:0] \add_32ns_32ns_32_2_1_U12.din0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U12.din1 ;
wire [31:0] \add_32ns_32ns_32_2_1_U12.dout ;
wire \add_32ns_32ns_32_2_1_U12.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_8_U.a ;
wire [31:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_8_U.ain_s0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_8_U.b ;
wire [31:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_8_U.bin_s0 ;
wire \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_8_U.ce ;
wire \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_8_U.clk ;
wire \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_8_U.facout_s1 ;
wire \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_8_U.facout_s2 ;
wire [15:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_8_U.fas_s1 ;
wire [15:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_8_U.fas_s2 ;
wire \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_8_U.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_8_U.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_8_U.u1.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_8_U.u1.b ;
wire \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_8_U.u1.cin ;
wire \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_8_U.u1.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_8_U.u1.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_8_U.u2.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_8_U.u2.b ;
wire \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_8_U.u2.cin ;
wire \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_8_U.u2.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_8_U.u2.s ;
wire \add_32ns_32ns_32_2_1_U14.ce ;
wire \add_32ns_32ns_32_2_1_U14.clk ;
wire [31:0] \add_32ns_32ns_32_2_1_U14.din0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U14.din1 ;
wire [31:0] \add_32ns_32ns_32_2_1_U14.dout ;
wire \add_32ns_32ns_32_2_1_U14.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_8_U.a ;
wire [31:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_8_U.ain_s0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_8_U.b ;
wire [31:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_8_U.bin_s0 ;
wire \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_8_U.ce ;
wire \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_8_U.clk ;
wire \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_8_U.facout_s1 ;
wire \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_8_U.facout_s2 ;
wire [15:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_8_U.fas_s1 ;
wire [15:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_8_U.fas_s2 ;
wire \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_8_U.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_8_U.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_8_U.u1.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_8_U.u1.b ;
wire \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_8_U.u1.cin ;
wire \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_8_U.u1.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_8_U.u1.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_8_U.u2.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_8_U.u2.b ;
wire \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_8_U.u2.cin ;
wire \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_8_U.u2.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_8_U.u2.s ;
wire \add_32ns_32ns_32_2_1_U17.ce ;
wire \add_32ns_32ns_32_2_1_U17.clk ;
wire [31:0] \add_32ns_32ns_32_2_1_U17.din0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U17.din1 ;
wire [31:0] \add_32ns_32ns_32_2_1_U17.dout ;
wire \add_32ns_32ns_32_2_1_U17.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.a ;
wire [31:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.ain_s0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.b ;
wire [31:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.bin_s0 ;
wire \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.ce ;
wire \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.clk ;
wire \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.facout_s1 ;
wire \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.facout_s2 ;
wire [15:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.fas_s1 ;
wire [15:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.fas_s2 ;
wire \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.u1.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.u1.b ;
wire \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.u1.cin ;
wire \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.u1.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.u1.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.u2.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.u2.b ;
wire \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.u2.cin ;
wire \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.u2.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.u2.s ;
wire \add_32ns_32ns_32_2_1_U9.ce ;
wire \add_32ns_32ns_32_2_1_U9.clk ;
wire [31:0] \add_32ns_32ns_32_2_1_U9.din0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U9.din1 ;
wire [31:0] \add_32ns_32ns_32_2_1_U9.dout ;
wire \add_32ns_32ns_32_2_1_U9.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_8_U.a ;
wire [31:0] \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_8_U.ain_s0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_8_U.b ;
wire [31:0] \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_8_U.bin_s0 ;
wire \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_8_U.ce ;
wire \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_8_U.clk ;
wire \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_8_U.facout_s1 ;
wire \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_8_U.facout_s2 ;
wire [15:0] \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_8_U.fas_s1 ;
wire [15:0] \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_8_U.fas_s2 ;
wire \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_8_U.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_8_U.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_8_U.u1.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_8_U.u1.b ;
wire \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_8_U.u1.cin ;
wire \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_8_U.u1.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_8_U.u1.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_8_U.u2.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_8_U.u2.b ;
wire \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_8_U.u2.cin ;
wire \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_8_U.u2.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_8_U.u2.s ;
wire \add_32ns_32s_32_2_1_U10.ce ;
wire \add_32ns_32s_32_2_1_U10.clk ;
wire [31:0] \add_32ns_32s_32_2_1_U10.din0 ;
wire [31:0] \add_32ns_32s_32_2_1_U10.din1 ;
wire [31:0] \add_32ns_32s_32_2_1_U10.dout ;
wire \add_32ns_32s_32_2_1_U10.reset ;
wire [31:0] \add_32ns_32s_32_2_1_U10.top_add_32ns_32s_32_2_1_Adder_9_U.a ;
wire [31:0] \add_32ns_32s_32_2_1_U10.top_add_32ns_32s_32_2_1_Adder_9_U.ain_s0 ;
wire [31:0] \add_32ns_32s_32_2_1_U10.top_add_32ns_32s_32_2_1_Adder_9_U.b ;
wire [31:0] \add_32ns_32s_32_2_1_U10.top_add_32ns_32s_32_2_1_Adder_9_U.bin_s0 ;
wire \add_32ns_32s_32_2_1_U10.top_add_32ns_32s_32_2_1_Adder_9_U.ce ;
wire \add_32ns_32s_32_2_1_U10.top_add_32ns_32s_32_2_1_Adder_9_U.clk ;
wire \add_32ns_32s_32_2_1_U10.top_add_32ns_32s_32_2_1_Adder_9_U.facout_s1 ;
wire \add_32ns_32s_32_2_1_U10.top_add_32ns_32s_32_2_1_Adder_9_U.facout_s2 ;
wire [15:0] \add_32ns_32s_32_2_1_U10.top_add_32ns_32s_32_2_1_Adder_9_U.fas_s1 ;
wire [15:0] \add_32ns_32s_32_2_1_U10.top_add_32ns_32s_32_2_1_Adder_9_U.fas_s2 ;
wire \add_32ns_32s_32_2_1_U10.top_add_32ns_32s_32_2_1_Adder_9_U.reset ;
wire [31:0] \add_32ns_32s_32_2_1_U10.top_add_32ns_32s_32_2_1_Adder_9_U.s ;
wire [15:0] \add_32ns_32s_32_2_1_U10.top_add_32ns_32s_32_2_1_Adder_9_U.u1.a ;
wire [15:0] \add_32ns_32s_32_2_1_U10.top_add_32ns_32s_32_2_1_Adder_9_U.u1.b ;
wire \add_32ns_32s_32_2_1_U10.top_add_32ns_32s_32_2_1_Adder_9_U.u1.cin ;
wire \add_32ns_32s_32_2_1_U10.top_add_32ns_32s_32_2_1_Adder_9_U.u1.cout ;
wire [15:0] \add_32ns_32s_32_2_1_U10.top_add_32ns_32s_32_2_1_Adder_9_U.u1.s ;
wire [15:0] \add_32ns_32s_32_2_1_U10.top_add_32ns_32s_32_2_1_Adder_9_U.u2.a ;
wire [15:0] \add_32ns_32s_32_2_1_U10.top_add_32ns_32s_32_2_1_Adder_9_U.u2.b ;
wire \add_32ns_32s_32_2_1_U10.top_add_32ns_32s_32_2_1_Adder_9_U.u2.cin ;
wire \add_32ns_32s_32_2_1_U10.top_add_32ns_32s_32_2_1_Adder_9_U.u2.cout ;
wire [15:0] \add_32ns_32s_32_2_1_U10.top_add_32ns_32s_32_2_1_Adder_9_U.u2.s ;
wire \add_32ns_32s_32_2_1_U16.ce ;
wire \add_32ns_32s_32_2_1_U16.clk ;
wire [31:0] \add_32ns_32s_32_2_1_U16.din0 ;
wire [31:0] \add_32ns_32s_32_2_1_U16.din1 ;
wire [31:0] \add_32ns_32s_32_2_1_U16.dout ;
wire \add_32ns_32s_32_2_1_U16.reset ;
wire [31:0] \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.a ;
wire [31:0] \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.ain_s0 ;
wire [31:0] \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.b ;
wire [31:0] \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.bin_s0 ;
wire \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.ce ;
wire \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.clk ;
wire \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.facout_s1 ;
wire \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.facout_s2 ;
wire [15:0] \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.fas_s1 ;
wire [15:0] \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.fas_s2 ;
wire \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.reset ;
wire [31:0] \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.s ;
wire [15:0] \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.u1.a ;
wire [15:0] \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.u1.b ;
wire \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.u1.cin ;
wire \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.u1.cout ;
wire [15:0] \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.u1.s ;
wire [15:0] \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.u2.a ;
wire [15:0] \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.u2.b ;
wire \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.u2.cin ;
wire \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.u2.cout ;
wire [15:0] \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.u2.s ;
wire \add_33ns_33ns_33_2_1_U15.ce ;
wire \add_33ns_33ns_33_2_1_U15.clk ;
wire [32:0] \add_33ns_33ns_33_2_1_U15.din0 ;
wire [32:0] \add_33ns_33ns_33_2_1_U15.din1 ;
wire [32:0] \add_33ns_33ns_33_2_1_U15.dout ;
wire \add_33ns_33ns_33_2_1_U15.reset ;
wire [32:0] \add_33ns_33ns_33_2_1_U15.top_add_33ns_33ns_33_2_1_Adder_11_U.a ;
wire [32:0] \add_33ns_33ns_33_2_1_U15.top_add_33ns_33ns_33_2_1_Adder_11_U.ain_s0 ;
wire [32:0] \add_33ns_33ns_33_2_1_U15.top_add_33ns_33ns_33_2_1_Adder_11_U.b ;
wire [32:0] \add_33ns_33ns_33_2_1_U15.top_add_33ns_33ns_33_2_1_Adder_11_U.bin_s0 ;
wire \add_33ns_33ns_33_2_1_U15.top_add_33ns_33ns_33_2_1_Adder_11_U.ce ;
wire \add_33ns_33ns_33_2_1_U15.top_add_33ns_33ns_33_2_1_Adder_11_U.clk ;
wire \add_33ns_33ns_33_2_1_U15.top_add_33ns_33ns_33_2_1_Adder_11_U.facout_s1 ;
wire \add_33ns_33ns_33_2_1_U15.top_add_33ns_33ns_33_2_1_Adder_11_U.facout_s2 ;
wire [15:0] \add_33ns_33ns_33_2_1_U15.top_add_33ns_33ns_33_2_1_Adder_11_U.fas_s1 ;
wire [16:0] \add_33ns_33ns_33_2_1_U15.top_add_33ns_33ns_33_2_1_Adder_11_U.fas_s2 ;
wire \add_33ns_33ns_33_2_1_U15.top_add_33ns_33ns_33_2_1_Adder_11_U.reset ;
wire [32:0] \add_33ns_33ns_33_2_1_U15.top_add_33ns_33ns_33_2_1_Adder_11_U.s ;
wire [15:0] \add_33ns_33ns_33_2_1_U15.top_add_33ns_33ns_33_2_1_Adder_11_U.u1.a ;
wire [15:0] \add_33ns_33ns_33_2_1_U15.top_add_33ns_33ns_33_2_1_Adder_11_U.u1.b ;
wire \add_33ns_33ns_33_2_1_U15.top_add_33ns_33ns_33_2_1_Adder_11_U.u1.cin ;
wire \add_33ns_33ns_33_2_1_U15.top_add_33ns_33ns_33_2_1_Adder_11_U.u1.cout ;
wire [15:0] \add_33ns_33ns_33_2_1_U15.top_add_33ns_33ns_33_2_1_Adder_11_U.u1.s ;
wire [16:0] \add_33ns_33ns_33_2_1_U15.top_add_33ns_33ns_33_2_1_Adder_11_U.u2.a ;
wire [16:0] \add_33ns_33ns_33_2_1_U15.top_add_33ns_33ns_33_2_1_Adder_11_U.u2.b ;
wire \add_33ns_33ns_33_2_1_U15.top_add_33ns_33ns_33_2_1_Adder_11_U.u2.cin ;
wire \add_33ns_33ns_33_2_1_U15.top_add_33ns_33ns_33_2_1_Adder_11_U.u2.cout ;
wire [16:0] \add_33ns_33ns_33_2_1_U15.top_add_33ns_33ns_33_2_1_Adder_11_U.u2.s ;
wire \add_33s_33s_33_2_1_U7.ce ;
wire \add_33s_33s_33_2_1_U7.clk ;
wire [32:0] \add_33s_33s_33_2_1_U7.din0 ;
wire [32:0] \add_33s_33s_33_2_1_U7.din1 ;
wire [32:0] \add_33s_33s_33_2_1_U7.dout ;
wire \add_33s_33s_33_2_1_U7.reset ;
wire [32:0] \add_33s_33s_33_2_1_U7.top_add_33s_33s_33_2_1_Adder_6_U.a ;
wire [32:0] \add_33s_33s_33_2_1_U7.top_add_33s_33s_33_2_1_Adder_6_U.ain_s0 ;
wire [32:0] \add_33s_33s_33_2_1_U7.top_add_33s_33s_33_2_1_Adder_6_U.b ;
wire [32:0] \add_33s_33s_33_2_1_U7.top_add_33s_33s_33_2_1_Adder_6_U.bin_s0 ;
wire \add_33s_33s_33_2_1_U7.top_add_33s_33s_33_2_1_Adder_6_U.ce ;
wire \add_33s_33s_33_2_1_U7.top_add_33s_33s_33_2_1_Adder_6_U.clk ;
wire \add_33s_33s_33_2_1_U7.top_add_33s_33s_33_2_1_Adder_6_U.facout_s1 ;
wire \add_33s_33s_33_2_1_U7.top_add_33s_33s_33_2_1_Adder_6_U.facout_s2 ;
wire [15:0] \add_33s_33s_33_2_1_U7.top_add_33s_33s_33_2_1_Adder_6_U.fas_s1 ;
wire [16:0] \add_33s_33s_33_2_1_U7.top_add_33s_33s_33_2_1_Adder_6_U.fas_s2 ;
wire \add_33s_33s_33_2_1_U7.top_add_33s_33s_33_2_1_Adder_6_U.reset ;
wire [32:0] \add_33s_33s_33_2_1_U7.top_add_33s_33s_33_2_1_Adder_6_U.s ;
wire [15:0] \add_33s_33s_33_2_1_U7.top_add_33s_33s_33_2_1_Adder_6_U.u1.a ;
wire [15:0] \add_33s_33s_33_2_1_U7.top_add_33s_33s_33_2_1_Adder_6_U.u1.b ;
wire \add_33s_33s_33_2_1_U7.top_add_33s_33s_33_2_1_Adder_6_U.u1.cin ;
wire \add_33s_33s_33_2_1_U7.top_add_33s_33s_33_2_1_Adder_6_U.u1.cout ;
wire [15:0] \add_33s_33s_33_2_1_U7.top_add_33s_33s_33_2_1_Adder_6_U.u1.s ;
wire [16:0] \add_33s_33s_33_2_1_U7.top_add_33s_33s_33_2_1_Adder_6_U.u2.a ;
wire [16:0] \add_33s_33s_33_2_1_U7.top_add_33s_33s_33_2_1_Adder_6_U.u2.b ;
wire \add_33s_33s_33_2_1_U7.top_add_33s_33s_33_2_1_Adder_6_U.u2.cin ;
wire \add_33s_33s_33_2_1_U7.top_add_33s_33s_33_2_1_Adder_6_U.u2.cout ;
wire [16:0] \add_33s_33s_33_2_1_U7.top_add_33s_33s_33_2_1_Adder_6_U.u2.s ;
wire \add_36s_36s_36_2_1_U8.ce ;
wire \add_36s_36s_36_2_1_U8.clk ;
wire [35:0] \add_36s_36s_36_2_1_U8.din0 ;
wire [35:0] \add_36s_36s_36_2_1_U8.din1 ;
wire [35:0] \add_36s_36s_36_2_1_U8.dout ;
wire \add_36s_36s_36_2_1_U8.reset ;
wire [35:0] \add_36s_36s_36_2_1_U8.top_add_36s_36s_36_2_1_Adder_7_U.a ;
wire [35:0] \add_36s_36s_36_2_1_U8.top_add_36s_36s_36_2_1_Adder_7_U.ain_s0 ;
wire [35:0] \add_36s_36s_36_2_1_U8.top_add_36s_36s_36_2_1_Adder_7_U.b ;
wire [35:0] \add_36s_36s_36_2_1_U8.top_add_36s_36s_36_2_1_Adder_7_U.bin_s0 ;
wire \add_36s_36s_36_2_1_U8.top_add_36s_36s_36_2_1_Adder_7_U.ce ;
wire \add_36s_36s_36_2_1_U8.top_add_36s_36s_36_2_1_Adder_7_U.clk ;
wire \add_36s_36s_36_2_1_U8.top_add_36s_36s_36_2_1_Adder_7_U.facout_s1 ;
wire \add_36s_36s_36_2_1_U8.top_add_36s_36s_36_2_1_Adder_7_U.facout_s2 ;
wire [17:0] \add_36s_36s_36_2_1_U8.top_add_36s_36s_36_2_1_Adder_7_U.fas_s1 ;
wire [17:0] \add_36s_36s_36_2_1_U8.top_add_36s_36s_36_2_1_Adder_7_U.fas_s2 ;
wire \add_36s_36s_36_2_1_U8.top_add_36s_36s_36_2_1_Adder_7_U.reset ;
wire [35:0] \add_36s_36s_36_2_1_U8.top_add_36s_36s_36_2_1_Adder_7_U.s ;
wire [17:0] \add_36s_36s_36_2_1_U8.top_add_36s_36s_36_2_1_Adder_7_U.u1.a ;
wire [17:0] \add_36s_36s_36_2_1_U8.top_add_36s_36s_36_2_1_Adder_7_U.u1.b ;
wire \add_36s_36s_36_2_1_U8.top_add_36s_36s_36_2_1_Adder_7_U.u1.cin ;
wire \add_36s_36s_36_2_1_U8.top_add_36s_36s_36_2_1_Adder_7_U.u1.cout ;
wire [17:0] \add_36s_36s_36_2_1_U8.top_add_36s_36s_36_2_1_Adder_7_U.u1.s ;
wire [17:0] \add_36s_36s_36_2_1_U8.top_add_36s_36s_36_2_1_Adder_7_U.u2.a ;
wire [17:0] \add_36s_36s_36_2_1_U8.top_add_36s_36s_36_2_1_Adder_7_U.u2.b ;
wire \add_36s_36s_36_2_1_U8.top_add_36s_36s_36_2_1_Adder_7_U.u2.cin ;
wire \add_36s_36s_36_2_1_U8.top_add_36s_36s_36_2_1_Adder_7_U.u2.cout ;
wire [17:0] \add_36s_36s_36_2_1_U8.top_add_36s_36s_36_2_1_Adder_7_U.u2.s ;
wire \add_43s_43s_43_2_1_U13.ce ;
wire \add_43s_43s_43_2_1_U13.clk ;
wire [42:0] \add_43s_43s_43_2_1_U13.din0 ;
wire [42:0] \add_43s_43s_43_2_1_U13.din1 ;
wire [42:0] \add_43s_43s_43_2_1_U13.dout ;
wire \add_43s_43s_43_2_1_U13.reset ;
wire [42:0] \add_43s_43s_43_2_1_U13.top_add_43s_43s_43_2_1_Adder_10_U.a ;
wire [42:0] \add_43s_43s_43_2_1_U13.top_add_43s_43s_43_2_1_Adder_10_U.ain_s0 ;
wire [42:0] \add_43s_43s_43_2_1_U13.top_add_43s_43s_43_2_1_Adder_10_U.b ;
wire [42:0] \add_43s_43s_43_2_1_U13.top_add_43s_43s_43_2_1_Adder_10_U.bin_s0 ;
wire \add_43s_43s_43_2_1_U13.top_add_43s_43s_43_2_1_Adder_10_U.ce ;
wire \add_43s_43s_43_2_1_U13.top_add_43s_43s_43_2_1_Adder_10_U.clk ;
wire \add_43s_43s_43_2_1_U13.top_add_43s_43s_43_2_1_Adder_10_U.facout_s1 ;
wire \add_43s_43s_43_2_1_U13.top_add_43s_43s_43_2_1_Adder_10_U.facout_s2 ;
wire [20:0] \add_43s_43s_43_2_1_U13.top_add_43s_43s_43_2_1_Adder_10_U.fas_s1 ;
wire [21:0] \add_43s_43s_43_2_1_U13.top_add_43s_43s_43_2_1_Adder_10_U.fas_s2 ;
wire \add_43s_43s_43_2_1_U13.top_add_43s_43s_43_2_1_Adder_10_U.reset ;
wire [42:0] \add_43s_43s_43_2_1_U13.top_add_43s_43s_43_2_1_Adder_10_U.s ;
wire [20:0] \add_43s_43s_43_2_1_U13.top_add_43s_43s_43_2_1_Adder_10_U.u1.a ;
wire [20:0] \add_43s_43s_43_2_1_U13.top_add_43s_43s_43_2_1_Adder_10_U.u1.b ;
wire \add_43s_43s_43_2_1_U13.top_add_43s_43s_43_2_1_Adder_10_U.u1.cin ;
wire \add_43s_43s_43_2_1_U13.top_add_43s_43s_43_2_1_Adder_10_U.u1.cout ;
wire [20:0] \add_43s_43s_43_2_1_U13.top_add_43s_43s_43_2_1_Adder_10_U.u1.s ;
wire [21:0] \add_43s_43s_43_2_1_U13.top_add_43s_43s_43_2_1_Adder_10_U.u2.a ;
wire [21:0] \add_43s_43s_43_2_1_U13.top_add_43s_43s_43_2_1_Adder_10_U.u2.b ;
wire \add_43s_43s_43_2_1_U13.top_add_43s_43s_43_2_1_Adder_10_U.u2.cin ;
wire \add_43s_43s_43_2_1_U13.top_add_43s_43s_43_2_1_Adder_10_U.u2.cout ;
wire [21:0] \add_43s_43s_43_2_1_U13.top_add_43s_43s_43_2_1_Adder_10_U.u2.s ;
wire \add_6ns_6ns_6_2_1_U2.ce ;
wire \add_6ns_6ns_6_2_1_U2.clk ;
wire [5:0] \add_6ns_6ns_6_2_1_U2.din0 ;
wire [5:0] \add_6ns_6ns_6_2_1_U2.din1 ;
wire [5:0] \add_6ns_6ns_6_2_1_U2.dout ;
wire \add_6ns_6ns_6_2_1_U2.reset ;
wire [5:0] \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.a ;
wire [5:0] \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.ain_s0 ;
wire [5:0] \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.b ;
wire [5:0] \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.bin_s0 ;
wire \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.ce ;
wire \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.clk ;
wire \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.facout_s1 ;
wire \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.facout_s2 ;
wire [2:0] \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.fas_s1 ;
wire [2:0] \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.fas_s2 ;
wire \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.reset ;
wire [5:0] \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.s ;
wire [2:0] \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.u1.a ;
wire [2:0] \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.u1.b ;
wire \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.u1.cin ;
wire \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.u1.cout ;
wire [2:0] \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.u1.s ;
wire [2:0] \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.u2.a ;
wire [2:0] \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.u2.b ;
wire \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.u2.cin ;
wire \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.u2.cout ;
wire [2:0] \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.u2.s ;
wire \add_8ns_8ns_8_2_1_U6.ce ;
wire \add_8ns_8ns_8_2_1_U6.clk ;
wire [7:0] \add_8ns_8ns_8_2_1_U6.din0 ;
wire [7:0] \add_8ns_8ns_8_2_1_U6.din1 ;
wire [7:0] \add_8ns_8ns_8_2_1_U6.dout ;
wire \add_8ns_8ns_8_2_1_U6.reset ;
wire [7:0] \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.a ;
wire [7:0] \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.ain_s0 ;
wire [7:0] \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.b ;
wire [7:0] \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.bin_s0 ;
wire \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.ce ;
wire \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.clk ;
wire \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.facout_s1 ;
wire \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.facout_s2 ;
wire [3:0] \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.fas_s1 ;
wire [3:0] \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.fas_s2 ;
wire \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.reset ;
wire [7:0] \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.s ;
wire [3:0] \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.u1.a ;
wire [3:0] \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.u1.b ;
wire \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.u1.cin ;
wire \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.u1.cout ;
wire [3:0] \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.u1.s ;
wire [3:0] \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.u2.a ;
wire [3:0] \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.u2.b ;
wire \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.u2.cin ;
wire \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.u2.cout ;
wire [3:0] \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.u2.s ;
wire \add_8s_8ns_8_2_1_U5.ce ;
wire \add_8s_8ns_8_2_1_U5.clk ;
wire [7:0] \add_8s_8ns_8_2_1_U5.din0 ;
wire [7:0] \add_8s_8ns_8_2_1_U5.din1 ;
wire [7:0] \add_8s_8ns_8_2_1_U5.dout ;
wire \add_8s_8ns_8_2_1_U5.reset ;
wire [7:0] \add_8s_8ns_8_2_1_U5.top_add_8s_8ns_8_2_1_Adder_4_U.a ;
wire [7:0] \add_8s_8ns_8_2_1_U5.top_add_8s_8ns_8_2_1_Adder_4_U.ain_s0 ;
wire [7:0] \add_8s_8ns_8_2_1_U5.top_add_8s_8ns_8_2_1_Adder_4_U.b ;
wire [7:0] \add_8s_8ns_8_2_1_U5.top_add_8s_8ns_8_2_1_Adder_4_U.bin_s0 ;
wire \add_8s_8ns_8_2_1_U5.top_add_8s_8ns_8_2_1_Adder_4_U.ce ;
wire \add_8s_8ns_8_2_1_U5.top_add_8s_8ns_8_2_1_Adder_4_U.clk ;
wire \add_8s_8ns_8_2_1_U5.top_add_8s_8ns_8_2_1_Adder_4_U.facout_s1 ;
wire \add_8s_8ns_8_2_1_U5.top_add_8s_8ns_8_2_1_Adder_4_U.facout_s2 ;
wire [3:0] \add_8s_8ns_8_2_1_U5.top_add_8s_8ns_8_2_1_Adder_4_U.fas_s1 ;
wire [3:0] \add_8s_8ns_8_2_1_U5.top_add_8s_8ns_8_2_1_Adder_4_U.fas_s2 ;
wire \add_8s_8ns_8_2_1_U5.top_add_8s_8ns_8_2_1_Adder_4_U.reset ;
wire [7:0] \add_8s_8ns_8_2_1_U5.top_add_8s_8ns_8_2_1_Adder_4_U.s ;
wire [3:0] \add_8s_8ns_8_2_1_U5.top_add_8s_8ns_8_2_1_Adder_4_U.u1.a ;
wire [3:0] \add_8s_8ns_8_2_1_U5.top_add_8s_8ns_8_2_1_Adder_4_U.u1.b ;
wire \add_8s_8ns_8_2_1_U5.top_add_8s_8ns_8_2_1_Adder_4_U.u1.cin ;
wire \add_8s_8ns_8_2_1_U5.top_add_8s_8ns_8_2_1_Adder_4_U.u1.cout ;
wire [3:0] \add_8s_8ns_8_2_1_U5.top_add_8s_8ns_8_2_1_Adder_4_U.u1.s ;
wire [3:0] \add_8s_8ns_8_2_1_U5.top_add_8s_8ns_8_2_1_Adder_4_U.u2.a ;
wire [3:0] \add_8s_8ns_8_2_1_U5.top_add_8s_8ns_8_2_1_Adder_4_U.u2.b ;
wire \add_8s_8ns_8_2_1_U5.top_add_8s_8ns_8_2_1_Adder_4_U.u2.cin ;
wire \add_8s_8ns_8_2_1_U5.top_add_8s_8ns_8_2_1_Adder_4_U.u2.cout ;
wire [3:0] \add_8s_8ns_8_2_1_U5.top_add_8s_8ns_8_2_1_Adder_4_U.u2.s ;
wire \add_9ns_9s_9_2_1_U1.ce ;
wire \add_9ns_9s_9_2_1_U1.clk ;
wire [8:0] \add_9ns_9s_9_2_1_U1.din0 ;
wire [8:0] \add_9ns_9s_9_2_1_U1.din1 ;
wire [8:0] \add_9ns_9s_9_2_1_U1.dout ;
wire \add_9ns_9s_9_2_1_U1.reset ;
wire [8:0] \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.a ;
wire [8:0] \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.ain_s0 ;
wire [8:0] \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.b ;
wire [8:0] \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.bin_s0 ;
wire \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.ce ;
wire \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.clk ;
wire \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.facout_s1 ;
wire \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.facout_s2 ;
wire [3:0] \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.fas_s1 ;
wire [4:0] \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.fas_s2 ;
wire \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.reset ;
wire [8:0] \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.s ;
wire [3:0] \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.u1.a ;
wire [3:0] \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.u1.b ;
wire \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.u1.cin ;
wire \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.u1.cout ;
wire [3:0] \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.u1.s ;
wire [4:0] \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.u2.a ;
wire [4:0] \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.u2.b ;
wire \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.u2.cin ;
wire \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.u2.cout ;
wire [4:0] \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.u2.s ;
wire and_ln340_fu_310_p2;
wire and_ln785_1_fu_345_p2;
wire and_ln785_fu_339_p2;
wire ap_CS_fsm_state1;
wire ap_CS_fsm_state10;
wire ap_CS_fsm_state11;
wire ap_CS_fsm_state12;
wire ap_CS_fsm_state13;
wire ap_CS_fsm_state14;
wire ap_CS_fsm_state15;
wire ap_CS_fsm_state16;
wire ap_CS_fsm_state17;
wire ap_CS_fsm_state18;
wire ap_CS_fsm_state19;
wire ap_CS_fsm_state2;
wire ap_CS_fsm_state20;
wire ap_CS_fsm_state21;
wire ap_CS_fsm_state22;
wire ap_CS_fsm_state23;
wire ap_CS_fsm_state24;
wire ap_CS_fsm_state25;
wire ap_CS_fsm_state26;
wire ap_CS_fsm_state27;
wire ap_CS_fsm_state28;
wire ap_CS_fsm_state29;
wire ap_CS_fsm_state3;
wire ap_CS_fsm_state30;
wire ap_CS_fsm_state31;
wire ap_CS_fsm_state32;
wire ap_CS_fsm_state33;
wire ap_CS_fsm_state34;
wire ap_CS_fsm_state35;
wire ap_CS_fsm_state36;
wire ap_CS_fsm_state37;
wire ap_CS_fsm_state4;
wire ap_CS_fsm_state5;
wire ap_CS_fsm_state6;
wire ap_CS_fsm_state7;
wire ap_CS_fsm_state8;
wire ap_CS_fsm_state9;
wire [36:0] ap_NS_fsm;
wire ap_clk;
wire ap_done;
wire ap_idle;
wire ap_ready;
wire ap_rst;
wire ap_start;
wire [8:0] grp_fu_364_p1;
wire [8:0] grp_fu_364_p2;
wire [5:0] grp_fu_420_p2;
wire [4:0] grp_fu_534_p2;
wire [13:0] grp_fu_552_p0;
wire [13:0] grp_fu_552_p1;
wire [13:0] grp_fu_552_p2;
wire [7:0] grp_fu_576_p0;
wire [7:0] grp_fu_576_p2;
wire [7:0] grp_fu_605_p1;
wire [7:0] grp_fu_605_p2;
wire [32:0] grp_fu_632_p0;
wire [32:0] grp_fu_632_p1;
wire [32:0] grp_fu_632_p2;
wire [35:0] grp_fu_663_p0;
wire [35:0] grp_fu_663_p1;
wire [35:0] grp_fu_663_p2;
wire [31:0] grp_fu_689_p2;
wire [31:0] grp_fu_717_p1;
wire [31:0] grp_fu_717_p2;
wire [31:0] grp_fu_725_p0;
wire [31:0] grp_fu_725_p2;
wire [31:0] grp_fu_731_p2;
wire [42:0] grp_fu_750_p0;
wire [42:0] grp_fu_750_p1;
wire [42:0] grp_fu_750_p2;
wire [31:0] grp_fu_776_p2;
wire [32:0] grp_fu_822_p0;
wire [32:0] grp_fu_822_p1;
wire [32:0] grp_fu_822_p2;
wire [31:0] grp_fu_842_p1;
wire [31:0] grp_fu_842_p2;
wire [31:0] grp_fu_847_p2;
wire icmp_ln768_1_fu_445_p2;
wire icmp_ln768_fu_249_p2;
wire icmp_ln786_1_fu_450_p2;
wire icmp_ln786_fu_255_p2;
wire icmp_ln851_1_fu_558_p2;
wire icmp_ln851_2_fu_673_p2;
wire icmp_ln851_3_fu_760_p2;
wire icmp_ln851_fu_415_p2;
wire newsignbit_fu_235_p1;
wire [7:0] op_0;
wire [3:0] op_1;
wire [1:0] op_10;
wire [5:0] op_11_V_fu_610_p3;
wire [3:0] op_12;
wire [1:0] op_13;
wire [31:0] op_15;
wire [31:0] op_16;
wire [2:0] op_17_V_fu_807_p1;
wire [3:0] op_18;
wire [31:0] op_19;
wire op_2;
wire [31:0] op_31;
wire op_31_ap_vld;
wire op_3_V_fu_355_p2;
wire op_6;
wire [7:0] op_9_V_fu_504_p3;
wire or_ln340_fu_299_p2;
wire or_ln384_fu_499_p2;
wire or_ln785_1_fu_461_p2;
wire or_ln785_2_fu_334_p2;
wire or_ln785_3_fu_350_p2;
wire or_ln785_fu_275_p2;
wire or_ln786_1_fu_482_p2;
wire or_ln786_fu_294_p2;
wire overflow_1_fu_465_p2;
wire overflow_fu_284_p2;
wire p_Result_5_fu_582_p3;
wire p_Result_6_fu_694_p3;
wire p_Result_7_fu_781_p3;
wire p_Result_9_fu_439_p2;
wire p_Result_s_18_fu_470_p3;
wire [2:0] p_Result_s_fu_239_p4;
wire [7:0] p_Val2_3_fu_432_p3;
wire r_1_fu_383_p2;
wire [3:0] r_fu_267_p3;
wire [1:0] ret_2_fu_425_p3;
wire [4:0] ret_V_15_fu_391_p3;
wire [7:0] ret_V_17_fu_594_p3;
wire [31:0] ret_V_19_fu_706_p3;
wire [1:0] ret_fu_455_p2;
wire [12:0] rhs_1_fu_541_p3;
wire [34:0] rhs_3_fu_652_p3;
wire [41:0] rhs_6_fu_739_p3;
wire select_ln1192_fu_316_p0;
wire [8:0] select_ln1192_fu_316_p3;
wire [4:0] select_ln1193_fu_511_p3;
wire [31:0] select_ln353_fu_793_p3;
wire [7:0] select_ln384_fu_492_p3;
wire [7:0] select_ln850_1_fu_589_p3;
wire [31:0] select_ln850_2_fu_701_p3;
wire [5:0] select_ln850_3_fu_523_p3;
wire [31:0] select_ln850_4_fu_788_p3;
wire [5:0] select_ln850_fu_518_p3;
wire [3:0] sext_ln703_1_fu_648_p0;
wire [31:0] sext_ln703_2_fu_735_p0;
wire [7:0] sext_ln850_fu_573_p1;
wire [3:0] shl_ln1497_fu_261_p2;
wire \sub_5ns_5ns_5_2_1_U3.ce ;
wire \sub_5ns_5ns_5_2_1_U3.clk ;
wire [4:0] \sub_5ns_5ns_5_2_1_U3.din0 ;
wire [4:0] \sub_5ns_5ns_5_2_1_U3.din1 ;
wire [4:0] \sub_5ns_5ns_5_2_1_U3.dout ;
wire \sub_5ns_5ns_5_2_1_U3.reset ;
wire [4:0] \sub_5ns_5ns_5_2_1_U3.top_sub_5ns_5ns_5_2_1_Adder_2_U.a ;
wire [4:0] \sub_5ns_5ns_5_2_1_U3.top_sub_5ns_5ns_5_2_1_Adder_2_U.ain_s0 ;
wire [4:0] \sub_5ns_5ns_5_2_1_U3.top_sub_5ns_5ns_5_2_1_Adder_2_U.b ;
wire [4:0] \sub_5ns_5ns_5_2_1_U3.top_sub_5ns_5ns_5_2_1_Adder_2_U.bin_s0 ;
wire \sub_5ns_5ns_5_2_1_U3.top_sub_5ns_5ns_5_2_1_Adder_2_U.ce ;
wire \sub_5ns_5ns_5_2_1_U3.top_sub_5ns_5ns_5_2_1_Adder_2_U.clk ;
wire \sub_5ns_5ns_5_2_1_U3.top_sub_5ns_5ns_5_2_1_Adder_2_U.facout_s1 ;
wire \sub_5ns_5ns_5_2_1_U3.top_sub_5ns_5ns_5_2_1_Adder_2_U.facout_s2 ;
wire [1:0] \sub_5ns_5ns_5_2_1_U3.top_sub_5ns_5ns_5_2_1_Adder_2_U.fas_s1 ;
wire [2:0] \sub_5ns_5ns_5_2_1_U3.top_sub_5ns_5ns_5_2_1_Adder_2_U.fas_s2 ;
wire \sub_5ns_5ns_5_2_1_U3.top_sub_5ns_5ns_5_2_1_Adder_2_U.reset ;
wire [4:0] \sub_5ns_5ns_5_2_1_U3.top_sub_5ns_5ns_5_2_1_Adder_2_U.s ;
wire [1:0] \sub_5ns_5ns_5_2_1_U3.top_sub_5ns_5ns_5_2_1_Adder_2_U.u1.a ;
wire [1:0] \sub_5ns_5ns_5_2_1_U3.top_sub_5ns_5ns_5_2_1_Adder_2_U.u1.b ;
wire \sub_5ns_5ns_5_2_1_U3.top_sub_5ns_5ns_5_2_1_Adder_2_U.u1.cin ;
wire \sub_5ns_5ns_5_2_1_U3.top_sub_5ns_5ns_5_2_1_Adder_2_U.u1.cout ;
wire [1:0] \sub_5ns_5ns_5_2_1_U3.top_sub_5ns_5ns_5_2_1_Adder_2_U.u1.s ;
wire [2:0] \sub_5ns_5ns_5_2_1_U3.top_sub_5ns_5ns_5_2_1_Adder_2_U.u2.a ;
wire [2:0] \sub_5ns_5ns_5_2_1_U3.top_sub_5ns_5ns_5_2_1_Adder_2_U.u2.b ;
wire \sub_5ns_5ns_5_2_1_U3.top_sub_5ns_5ns_5_2_1_Adder_2_U.u2.cin ;
wire \sub_5ns_5ns_5_2_1_U3.top_sub_5ns_5ns_5_2_1_Adder_2_U.u2.cout ;
wire [2:0] \sub_5ns_5ns_5_2_1_U3.top_sub_5ns_5ns_5_2_1_Adder_2_U.u2.s ;
wire [1:0] tmp_4_fu_800_p3;
wire [8:0] tmp_6_fu_621_p3;
wire [1:0] trunc_ln1497_fu_412_p1;
wire trunc_ln728_fu_398_p1;
wire [6:0] trunc_ln851_1_fu_530_p1;
wire [3:0] trunc_ln851_2_fu_669_p0;
wire [2:0] trunc_ln851_2_fu_669_p1;
wire [31:0] trunc_ln851_3_fu_756_p0;
wire [9:0] trunc_ln851_3_fu_756_p1;
wire [2:0] trunc_ln851_fu_379_p1;
wire underflow_1_fu_487_p2;
wire xor_ln340_fu_304_p2;
wire xor_ln785_1_fu_329_p2;
wire xor_ln785_fu_279_p2;
wire xor_ln786_1_fu_477_p2;
wire xor_ln786_2_fu_324_p2;
wire xor_ln786_fu_289_p2;
wire [4:0] zext_ln703_fu_388_p1;


assign _054_ = icmp_ln851_2_reg_1098 & ap_CS_fsm[20];
assign _055_ = icmp_ln851_3_reg_1165 & ap_CS_fsm[29];
assign _056_ = ap_CS_fsm[11] & icmp_ln851_1_reg_1026;
assign _057_ = _059_ & ap_CS_fsm[0];
assign _058_ = ap_start & ap_CS_fsm[0];
assign and_ln340_fu_310_p2 = xor_ln340_fu_304_p2 & or_ln786_fu_294_p2;
assign and_ln785_1_fu_345_p2 = newsignbit_reg_860 & and_ln785_fu_339_p2;
assign and_ln785_fu_339_p2 = xor_ln786_2_fu_324_p2 & or_ln785_2_fu_334_p2;
assign op_3_V_fu_355_p2 = or_ln785_3_fu_350_p2 & newsignbit_reg_860;
assign overflow_1_fu_465_p2 = r_1_reg_931 & or_ln785_1_fu_461_p2;
assign overflow_fu_284_p2 = xor_ln785_fu_279_p2 & or_ln785_reg_885;
assign ret_fu_455_p2 = r_reg_879[1:0] & ret_2_fu_425_p3;
assign underflow_1_fu_487_p2 = or_ln786_1_fu_482_p2 & op_3_V_reg_901;
assign xor_ln786_fu_289_p2 = ~ newsignbit_reg_860;
assign xor_ln785_fu_279_p2 = ~ p_Result_8_reg_853;
assign xor_ln340_fu_304_p2 = ~ or_ln340_fu_299_p2;
assign xor_ln785_1_fu_329_p2 = ~ or_ln785_reg_885;
assign xor_ln786_2_fu_324_p2 = ~ icmp_ln786_reg_873;
assign xor_ln786_1_fu_477_p2 = ~ p_Result_9_reg_964;
assign r_1_fu_383_p2 = ~ op_3_V_reg_901;
assign _059_ = ~ ap_start;
assign _060_ = ! trunc_ln851_reg_926;
always @(posedge \add_14s_14s_14_2_1_U4.top_add_14s_14s_14_2_1_Adder_3_U.clk )
\add_14s_14s_14_2_1_U4.top_add_14s_14s_14_2_1_Adder_3_U.bin_s1  <= _062_;
always @(posedge \add_14s_14s_14_2_1_U4.top_add_14s_14s_14_2_1_Adder_3_U.clk )
\add_14s_14s_14_2_1_U4.top_add_14s_14s_14_2_1_Adder_3_U.ain_s1  <= _061_;
always @(posedge \add_14s_14s_14_2_1_U4.top_add_14s_14s_14_2_1_Adder_3_U.clk )
\add_14s_14s_14_2_1_U4.top_add_14s_14s_14_2_1_Adder_3_U.sum_s1  <= _064_;
always @(posedge \add_14s_14s_14_2_1_U4.top_add_14s_14s_14_2_1_Adder_3_U.clk )
\add_14s_14s_14_2_1_U4.top_add_14s_14s_14_2_1_Adder_3_U.carry_s1  <= _063_;
assign _062_ = \add_14s_14s_14_2_1_U4.top_add_14s_14s_14_2_1_Adder_3_U.ce  ? \add_14s_14s_14_2_1_U4.top_add_14s_14s_14_2_1_Adder_3_U.b [13:7] : \add_14s_14s_14_2_1_U4.top_add_14s_14s_14_2_1_Adder_3_U.bin_s1 ;
assign _061_ = \add_14s_14s_14_2_1_U4.top_add_14s_14s_14_2_1_Adder_3_U.ce  ? \add_14s_14s_14_2_1_U4.top_add_14s_14s_14_2_1_Adder_3_U.a [13:7] : \add_14s_14s_14_2_1_U4.top_add_14s_14s_14_2_1_Adder_3_U.ain_s1 ;
assign _063_ = \add_14s_14s_14_2_1_U4.top_add_14s_14s_14_2_1_Adder_3_U.ce  ? \add_14s_14s_14_2_1_U4.top_add_14s_14s_14_2_1_Adder_3_U.facout_s1  : \add_14s_14s_14_2_1_U4.top_add_14s_14s_14_2_1_Adder_3_U.carry_s1 ;
assign _064_ = \add_14s_14s_14_2_1_U4.top_add_14s_14s_14_2_1_Adder_3_U.ce  ? \add_14s_14s_14_2_1_U4.top_add_14s_14s_14_2_1_Adder_3_U.fas_s1  : \add_14s_14s_14_2_1_U4.top_add_14s_14s_14_2_1_Adder_3_U.sum_s1 ;
assign _065_ = \add_14s_14s_14_2_1_U4.top_add_14s_14s_14_2_1_Adder_3_U.u1.a  + \add_14s_14s_14_2_1_U4.top_add_14s_14s_14_2_1_Adder_3_U.u1.b ;
assign { \add_14s_14s_14_2_1_U4.top_add_14s_14s_14_2_1_Adder_3_U.u1.cout , \add_14s_14s_14_2_1_U4.top_add_14s_14s_14_2_1_Adder_3_U.u1.s  } = _065_ + \add_14s_14s_14_2_1_U4.top_add_14s_14s_14_2_1_Adder_3_U.u1.cin ;
assign _066_ = \add_14s_14s_14_2_1_U4.top_add_14s_14s_14_2_1_Adder_3_U.u2.a  + \add_14s_14s_14_2_1_U4.top_add_14s_14s_14_2_1_Adder_3_U.u2.b ;
assign { \add_14s_14s_14_2_1_U4.top_add_14s_14s_14_2_1_Adder_3_U.u2.cout , \add_14s_14s_14_2_1_U4.top_add_14s_14s_14_2_1_Adder_3_U.u2.s  } = _066_ + \add_14s_14s_14_2_1_U4.top_add_14s_14s_14_2_1_Adder_3_U.u2.cin ;
always @(posedge \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.clk )
\add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.bin_s1  <= _068_;
always @(posedge \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.clk )
\add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.ain_s1  <= _067_;
always @(posedge \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.clk )
\add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.sum_s1  <= _070_;
always @(posedge \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.clk )
\add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.carry_s1  <= _069_;
assign _068_ = \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.ce  ? \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.b [31:16] : \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.bin_s1 ;
assign _067_ = \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.ce  ? \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.a [31:16] : \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.ain_s1 ;
assign _069_ = \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.ce  ? \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.facout_s1  : \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.carry_s1 ;
assign _070_ = \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.ce  ? \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.fas_s1  : \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.sum_s1 ;
assign _071_ = \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.u1.a  + \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.u1.b ;
assign { \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.u1.cout , \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.u1.s  } = _071_ + \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.u1.cin ;
assign _072_ = \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.u2.a  + \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.u2.b ;
assign { \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.u2.cout , \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.u2.s  } = _072_ + \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.u2.cin ;
always @(posedge \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_8_U.clk )
\add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_8_U.bin_s1  <= _074_;
always @(posedge \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_8_U.clk )
\add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_8_U.ain_s1  <= _073_;
always @(posedge \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_8_U.clk )
\add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_8_U.sum_s1  <= _076_;
always @(posedge \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_8_U.clk )
\add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_8_U.carry_s1  <= _075_;
assign _074_ = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_8_U.ce  ? \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_8_U.b [31:16] : \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_8_U.bin_s1 ;
assign _073_ = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_8_U.ce  ? \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_8_U.a [31:16] : \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_8_U.ain_s1 ;
assign _075_ = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_8_U.ce  ? \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_8_U.facout_s1  : \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_8_U.carry_s1 ;
assign _076_ = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_8_U.ce  ? \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_8_U.fas_s1  : \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_8_U.sum_s1 ;
assign _077_ = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_8_U.u1.a  + \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_8_U.u1.b ;
assign { \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_8_U.u1.cout , \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_8_U.u1.s  } = _077_ + \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_8_U.u1.cin ;
assign _078_ = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_8_U.u2.a  + \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_8_U.u2.b ;
assign { \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_8_U.u2.cout , \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_8_U.u2.s  } = _078_ + \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_8_U.u2.cin ;
always @(posedge \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_8_U.clk )
\add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_8_U.bin_s1  <= _080_;
always @(posedge \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_8_U.clk )
\add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_8_U.ain_s1  <= _079_;
always @(posedge \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_8_U.clk )
\add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_8_U.sum_s1  <= _082_;
always @(posedge \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_8_U.clk )
\add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_8_U.carry_s1  <= _081_;
assign _080_ = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_8_U.ce  ? \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_8_U.b [31:16] : \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_8_U.bin_s1 ;
assign _079_ = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_8_U.ce  ? \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_8_U.a [31:16] : \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_8_U.ain_s1 ;
assign _081_ = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_8_U.ce  ? \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_8_U.facout_s1  : \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_8_U.carry_s1 ;
assign _082_ = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_8_U.ce  ? \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_8_U.fas_s1  : \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_8_U.sum_s1 ;
assign _083_ = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_8_U.u1.a  + \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_8_U.u1.b ;
assign { \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_8_U.u1.cout , \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_8_U.u1.s  } = _083_ + \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_8_U.u1.cin ;
assign _084_ = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_8_U.u2.a  + \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_8_U.u2.b ;
assign { \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_8_U.u2.cout , \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_8_U.u2.s  } = _084_ + \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_8_U.u2.cin ;
always @(posedge \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.clk )
\add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.bin_s1  <= _086_;
always @(posedge \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.clk )
\add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.ain_s1  <= _085_;
always @(posedge \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.clk )
\add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.sum_s1  <= _088_;
always @(posedge \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.clk )
\add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.carry_s1  <= _087_;
assign _086_ = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.ce  ? \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.b [31:16] : \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.bin_s1 ;
assign _085_ = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.ce  ? \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.a [31:16] : \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.ain_s1 ;
assign _087_ = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.ce  ? \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.facout_s1  : \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.carry_s1 ;
assign _088_ = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.ce  ? \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.fas_s1  : \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.sum_s1 ;
assign _089_ = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.u1.a  + \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.u1.b ;
assign { \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.u1.cout , \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.u1.s  } = _089_ + \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.u1.cin ;
assign _090_ = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.u2.a  + \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.u2.b ;
assign { \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.u2.cout , \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.u2.s  } = _090_ + \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.u2.cin ;
always @(posedge \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_8_U.clk )
\add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_8_U.bin_s1  <= _092_;
always @(posedge \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_8_U.clk )
\add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_8_U.ain_s1  <= _091_;
always @(posedge \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_8_U.clk )
\add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_8_U.sum_s1  <= _094_;
always @(posedge \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_8_U.clk )
\add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_8_U.carry_s1  <= _093_;
assign _092_ = \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_8_U.ce  ? \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_8_U.b [31:16] : \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_8_U.bin_s1 ;
assign _091_ = \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_8_U.ce  ? \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_8_U.a [31:16] : \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_8_U.ain_s1 ;
assign _093_ = \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_8_U.ce  ? \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_8_U.facout_s1  : \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_8_U.carry_s1 ;
assign _094_ = \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_8_U.ce  ? \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_8_U.fas_s1  : \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_8_U.sum_s1 ;
assign _095_ = \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_8_U.u1.a  + \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_8_U.u1.b ;
assign { \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_8_U.u1.cout , \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_8_U.u1.s  } = _095_ + \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_8_U.u1.cin ;
assign _096_ = \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_8_U.u2.a  + \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_8_U.u2.b ;
assign { \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_8_U.u2.cout , \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_8_U.u2.s  } = _096_ + \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_8_U.u2.cin ;
always @(posedge \add_32ns_32s_32_2_1_U10.top_add_32ns_32s_32_2_1_Adder_9_U.clk )
\add_32ns_32s_32_2_1_U10.top_add_32ns_32s_32_2_1_Adder_9_U.bin_s1  <= _098_;
always @(posedge \add_32ns_32s_32_2_1_U10.top_add_32ns_32s_32_2_1_Adder_9_U.clk )
\add_32ns_32s_32_2_1_U10.top_add_32ns_32s_32_2_1_Adder_9_U.ain_s1  <= _097_;
always @(posedge \add_32ns_32s_32_2_1_U10.top_add_32ns_32s_32_2_1_Adder_9_U.clk )
\add_32ns_32s_32_2_1_U10.top_add_32ns_32s_32_2_1_Adder_9_U.sum_s1  <= _100_;
always @(posedge \add_32ns_32s_32_2_1_U10.top_add_32ns_32s_32_2_1_Adder_9_U.clk )
\add_32ns_32s_32_2_1_U10.top_add_32ns_32s_32_2_1_Adder_9_U.carry_s1  <= _099_;
assign _098_ = \add_32ns_32s_32_2_1_U10.top_add_32ns_32s_32_2_1_Adder_9_U.ce  ? \add_32ns_32s_32_2_1_U10.top_add_32ns_32s_32_2_1_Adder_9_U.b [31:16] : \add_32ns_32s_32_2_1_U10.top_add_32ns_32s_32_2_1_Adder_9_U.bin_s1 ;
assign _097_ = \add_32ns_32s_32_2_1_U10.top_add_32ns_32s_32_2_1_Adder_9_U.ce  ? \add_32ns_32s_32_2_1_U10.top_add_32ns_32s_32_2_1_Adder_9_U.a [31:16] : \add_32ns_32s_32_2_1_U10.top_add_32ns_32s_32_2_1_Adder_9_U.ain_s1 ;
assign _099_ = \add_32ns_32s_32_2_1_U10.top_add_32ns_32s_32_2_1_Adder_9_U.ce  ? \add_32ns_32s_32_2_1_U10.top_add_32ns_32s_32_2_1_Adder_9_U.facout_s1  : \add_32ns_32s_32_2_1_U10.top_add_32ns_32s_32_2_1_Adder_9_U.carry_s1 ;
assign _100_ = \add_32ns_32s_32_2_1_U10.top_add_32ns_32s_32_2_1_Adder_9_U.ce  ? \add_32ns_32s_32_2_1_U10.top_add_32ns_32s_32_2_1_Adder_9_U.fas_s1  : \add_32ns_32s_32_2_1_U10.top_add_32ns_32s_32_2_1_Adder_9_U.sum_s1 ;
assign _101_ = \add_32ns_32s_32_2_1_U10.top_add_32ns_32s_32_2_1_Adder_9_U.u1.a  + \add_32ns_32s_32_2_1_U10.top_add_32ns_32s_32_2_1_Adder_9_U.u1.b ;
assign { \add_32ns_32s_32_2_1_U10.top_add_32ns_32s_32_2_1_Adder_9_U.u1.cout , \add_32ns_32s_32_2_1_U10.top_add_32ns_32s_32_2_1_Adder_9_U.u1.s  } = _101_ + \add_32ns_32s_32_2_1_U10.top_add_32ns_32s_32_2_1_Adder_9_U.u1.cin ;
assign _102_ = \add_32ns_32s_32_2_1_U10.top_add_32ns_32s_32_2_1_Adder_9_U.u2.a  + \add_32ns_32s_32_2_1_U10.top_add_32ns_32s_32_2_1_Adder_9_U.u2.b ;
assign { \add_32ns_32s_32_2_1_U10.top_add_32ns_32s_32_2_1_Adder_9_U.u2.cout , \add_32ns_32s_32_2_1_U10.top_add_32ns_32s_32_2_1_Adder_9_U.u2.s  } = _102_ + \add_32ns_32s_32_2_1_U10.top_add_32ns_32s_32_2_1_Adder_9_U.u2.cin ;
always @(posedge \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.clk )
\add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.bin_s1  <= _104_;
always @(posedge \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.clk )
\add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.ain_s1  <= _103_;
always @(posedge \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.clk )
\add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.sum_s1  <= _106_;
always @(posedge \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.clk )
\add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.carry_s1  <= _105_;
assign _104_ = \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.ce  ? \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.b [31:16] : \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.bin_s1 ;
assign _103_ = \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.ce  ? \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.a [31:16] : \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.ain_s1 ;
assign _105_ = \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.ce  ? \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.facout_s1  : \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.carry_s1 ;
assign _106_ = \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.ce  ? \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.fas_s1  : \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.sum_s1 ;
assign _107_ = \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.u1.a  + \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.u1.b ;
assign { \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.u1.cout , \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.u1.s  } = _107_ + \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.u1.cin ;
assign _108_ = \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.u2.a  + \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.u2.b ;
assign { \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.u2.cout , \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.u2.s  } = _108_ + \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.u2.cin ;
always @(posedge \add_33ns_33ns_33_2_1_U15.top_add_33ns_33ns_33_2_1_Adder_11_U.clk )
\add_33ns_33ns_33_2_1_U15.top_add_33ns_33ns_33_2_1_Adder_11_U.bin_s1  <= _110_;
always @(posedge \add_33ns_33ns_33_2_1_U15.top_add_33ns_33ns_33_2_1_Adder_11_U.clk )
\add_33ns_33ns_33_2_1_U15.top_add_33ns_33ns_33_2_1_Adder_11_U.ain_s1  <= _109_;
always @(posedge \add_33ns_33ns_33_2_1_U15.top_add_33ns_33ns_33_2_1_Adder_11_U.clk )
\add_33ns_33ns_33_2_1_U15.top_add_33ns_33ns_33_2_1_Adder_11_U.sum_s1  <= _112_;
always @(posedge \add_33ns_33ns_33_2_1_U15.top_add_33ns_33ns_33_2_1_Adder_11_U.clk )
\add_33ns_33ns_33_2_1_U15.top_add_33ns_33ns_33_2_1_Adder_11_U.carry_s1  <= _111_;
assign _110_ = \add_33ns_33ns_33_2_1_U15.top_add_33ns_33ns_33_2_1_Adder_11_U.ce  ? \add_33ns_33ns_33_2_1_U15.top_add_33ns_33ns_33_2_1_Adder_11_U.b [32:16] : \add_33ns_33ns_33_2_1_U15.top_add_33ns_33ns_33_2_1_Adder_11_U.bin_s1 ;
assign _109_ = \add_33ns_33ns_33_2_1_U15.top_add_33ns_33ns_33_2_1_Adder_11_U.ce  ? \add_33ns_33ns_33_2_1_U15.top_add_33ns_33ns_33_2_1_Adder_11_U.a [32:16] : \add_33ns_33ns_33_2_1_U15.top_add_33ns_33ns_33_2_1_Adder_11_U.ain_s1 ;
assign _111_ = \add_33ns_33ns_33_2_1_U15.top_add_33ns_33ns_33_2_1_Adder_11_U.ce  ? \add_33ns_33ns_33_2_1_U15.top_add_33ns_33ns_33_2_1_Adder_11_U.facout_s1  : \add_33ns_33ns_33_2_1_U15.top_add_33ns_33ns_33_2_1_Adder_11_U.carry_s1 ;
assign _112_ = \add_33ns_33ns_33_2_1_U15.top_add_33ns_33ns_33_2_1_Adder_11_U.ce  ? \add_33ns_33ns_33_2_1_U15.top_add_33ns_33ns_33_2_1_Adder_11_U.fas_s1  : \add_33ns_33ns_33_2_1_U15.top_add_33ns_33ns_33_2_1_Adder_11_U.sum_s1 ;
assign _113_ = \add_33ns_33ns_33_2_1_U15.top_add_33ns_33ns_33_2_1_Adder_11_U.u1.a  + \add_33ns_33ns_33_2_1_U15.top_add_33ns_33ns_33_2_1_Adder_11_U.u1.b ;
assign { \add_33ns_33ns_33_2_1_U15.top_add_33ns_33ns_33_2_1_Adder_11_U.u1.cout , \add_33ns_33ns_33_2_1_U15.top_add_33ns_33ns_33_2_1_Adder_11_U.u1.s  } = _113_ + \add_33ns_33ns_33_2_1_U15.top_add_33ns_33ns_33_2_1_Adder_11_U.u1.cin ;
assign _114_ = \add_33ns_33ns_33_2_1_U15.top_add_33ns_33ns_33_2_1_Adder_11_U.u2.a  + \add_33ns_33ns_33_2_1_U15.top_add_33ns_33ns_33_2_1_Adder_11_U.u2.b ;
assign { \add_33ns_33ns_33_2_1_U15.top_add_33ns_33ns_33_2_1_Adder_11_U.u2.cout , \add_33ns_33ns_33_2_1_U15.top_add_33ns_33ns_33_2_1_Adder_11_U.u2.s  } = _114_ + \add_33ns_33ns_33_2_1_U15.top_add_33ns_33ns_33_2_1_Adder_11_U.u2.cin ;
always @(posedge \add_33s_33s_33_2_1_U7.top_add_33s_33s_33_2_1_Adder_6_U.clk )
\add_33s_33s_33_2_1_U7.top_add_33s_33s_33_2_1_Adder_6_U.bin_s1  <= _116_;
always @(posedge \add_33s_33s_33_2_1_U7.top_add_33s_33s_33_2_1_Adder_6_U.clk )
\add_33s_33s_33_2_1_U7.top_add_33s_33s_33_2_1_Adder_6_U.ain_s1  <= _115_;
always @(posedge \add_33s_33s_33_2_1_U7.top_add_33s_33s_33_2_1_Adder_6_U.clk )
\add_33s_33s_33_2_1_U7.top_add_33s_33s_33_2_1_Adder_6_U.sum_s1  <= _118_;
always @(posedge \add_33s_33s_33_2_1_U7.top_add_33s_33s_33_2_1_Adder_6_U.clk )
\add_33s_33s_33_2_1_U7.top_add_33s_33s_33_2_1_Adder_6_U.carry_s1  <= _117_;
assign _116_ = \add_33s_33s_33_2_1_U7.top_add_33s_33s_33_2_1_Adder_6_U.ce  ? \add_33s_33s_33_2_1_U7.top_add_33s_33s_33_2_1_Adder_6_U.b [32:16] : \add_33s_33s_33_2_1_U7.top_add_33s_33s_33_2_1_Adder_6_U.bin_s1 ;
assign _115_ = \add_33s_33s_33_2_1_U7.top_add_33s_33s_33_2_1_Adder_6_U.ce  ? \add_33s_33s_33_2_1_U7.top_add_33s_33s_33_2_1_Adder_6_U.a [32:16] : \add_33s_33s_33_2_1_U7.top_add_33s_33s_33_2_1_Adder_6_U.ain_s1 ;
assign _117_ = \add_33s_33s_33_2_1_U7.top_add_33s_33s_33_2_1_Adder_6_U.ce  ? \add_33s_33s_33_2_1_U7.top_add_33s_33s_33_2_1_Adder_6_U.facout_s1  : \add_33s_33s_33_2_1_U7.top_add_33s_33s_33_2_1_Adder_6_U.carry_s1 ;
assign _118_ = \add_33s_33s_33_2_1_U7.top_add_33s_33s_33_2_1_Adder_6_U.ce  ? \add_33s_33s_33_2_1_U7.top_add_33s_33s_33_2_1_Adder_6_U.fas_s1  : \add_33s_33s_33_2_1_U7.top_add_33s_33s_33_2_1_Adder_6_U.sum_s1 ;
assign _119_ = \add_33s_33s_33_2_1_U7.top_add_33s_33s_33_2_1_Adder_6_U.u1.a  + \add_33s_33s_33_2_1_U7.top_add_33s_33s_33_2_1_Adder_6_U.u1.b ;
assign { \add_33s_33s_33_2_1_U7.top_add_33s_33s_33_2_1_Adder_6_U.u1.cout , \add_33s_33s_33_2_1_U7.top_add_33s_33s_33_2_1_Adder_6_U.u1.s  } = _119_ + \add_33s_33s_33_2_1_U7.top_add_33s_33s_33_2_1_Adder_6_U.u1.cin ;
assign _120_ = \add_33s_33s_33_2_1_U7.top_add_33s_33s_33_2_1_Adder_6_U.u2.a  + \add_33s_33s_33_2_1_U7.top_add_33s_33s_33_2_1_Adder_6_U.u2.b ;
assign { \add_33s_33s_33_2_1_U7.top_add_33s_33s_33_2_1_Adder_6_U.u2.cout , \add_33s_33s_33_2_1_U7.top_add_33s_33s_33_2_1_Adder_6_U.u2.s  } = _120_ + \add_33s_33s_33_2_1_U7.top_add_33s_33s_33_2_1_Adder_6_U.u2.cin ;
always @(posedge \add_36s_36s_36_2_1_U8.top_add_36s_36s_36_2_1_Adder_7_U.clk )
\add_36s_36s_36_2_1_U8.top_add_36s_36s_36_2_1_Adder_7_U.bin_s1  <= _122_;
always @(posedge \add_36s_36s_36_2_1_U8.top_add_36s_36s_36_2_1_Adder_7_U.clk )
\add_36s_36s_36_2_1_U8.top_add_36s_36s_36_2_1_Adder_7_U.ain_s1  <= _121_;
always @(posedge \add_36s_36s_36_2_1_U8.top_add_36s_36s_36_2_1_Adder_7_U.clk )
\add_36s_36s_36_2_1_U8.top_add_36s_36s_36_2_1_Adder_7_U.sum_s1  <= _124_;
always @(posedge \add_36s_36s_36_2_1_U8.top_add_36s_36s_36_2_1_Adder_7_U.clk )
\add_36s_36s_36_2_1_U8.top_add_36s_36s_36_2_1_Adder_7_U.carry_s1  <= _123_;
assign _122_ = \add_36s_36s_36_2_1_U8.top_add_36s_36s_36_2_1_Adder_7_U.ce  ? \add_36s_36s_36_2_1_U8.top_add_36s_36s_36_2_1_Adder_7_U.b [35:18] : \add_36s_36s_36_2_1_U8.top_add_36s_36s_36_2_1_Adder_7_U.bin_s1 ;
assign _121_ = \add_36s_36s_36_2_1_U8.top_add_36s_36s_36_2_1_Adder_7_U.ce  ? \add_36s_36s_36_2_1_U8.top_add_36s_36s_36_2_1_Adder_7_U.a [35:18] : \add_36s_36s_36_2_1_U8.top_add_36s_36s_36_2_1_Adder_7_U.ain_s1 ;
assign _123_ = \add_36s_36s_36_2_1_U8.top_add_36s_36s_36_2_1_Adder_7_U.ce  ? \add_36s_36s_36_2_1_U8.top_add_36s_36s_36_2_1_Adder_7_U.facout_s1  : \add_36s_36s_36_2_1_U8.top_add_36s_36s_36_2_1_Adder_7_U.carry_s1 ;
assign _124_ = \add_36s_36s_36_2_1_U8.top_add_36s_36s_36_2_1_Adder_7_U.ce  ? \add_36s_36s_36_2_1_U8.top_add_36s_36s_36_2_1_Adder_7_U.fas_s1  : \add_36s_36s_36_2_1_U8.top_add_36s_36s_36_2_1_Adder_7_U.sum_s1 ;
assign _125_ = \add_36s_36s_36_2_1_U8.top_add_36s_36s_36_2_1_Adder_7_U.u1.a  + \add_36s_36s_36_2_1_U8.top_add_36s_36s_36_2_1_Adder_7_U.u1.b ;
assign { \add_36s_36s_36_2_1_U8.top_add_36s_36s_36_2_1_Adder_7_U.u1.cout , \add_36s_36s_36_2_1_U8.top_add_36s_36s_36_2_1_Adder_7_U.u1.s  } = _125_ + \add_36s_36s_36_2_1_U8.top_add_36s_36s_36_2_1_Adder_7_U.u1.cin ;
assign _126_ = \add_36s_36s_36_2_1_U8.top_add_36s_36s_36_2_1_Adder_7_U.u2.a  + \add_36s_36s_36_2_1_U8.top_add_36s_36s_36_2_1_Adder_7_U.u2.b ;
assign { \add_36s_36s_36_2_1_U8.top_add_36s_36s_36_2_1_Adder_7_U.u2.cout , \add_36s_36s_36_2_1_U8.top_add_36s_36s_36_2_1_Adder_7_U.u2.s  } = _126_ + \add_36s_36s_36_2_1_U8.top_add_36s_36s_36_2_1_Adder_7_U.u2.cin ;
always @(posedge \add_43s_43s_43_2_1_U13.top_add_43s_43s_43_2_1_Adder_10_U.clk )
\add_43s_43s_43_2_1_U13.top_add_43s_43s_43_2_1_Adder_10_U.bin_s1  <= _128_;
always @(posedge \add_43s_43s_43_2_1_U13.top_add_43s_43s_43_2_1_Adder_10_U.clk )
\add_43s_43s_43_2_1_U13.top_add_43s_43s_43_2_1_Adder_10_U.ain_s1  <= _127_;
always @(posedge \add_43s_43s_43_2_1_U13.top_add_43s_43s_43_2_1_Adder_10_U.clk )
\add_43s_43s_43_2_1_U13.top_add_43s_43s_43_2_1_Adder_10_U.sum_s1  <= _130_;
always @(posedge \add_43s_43s_43_2_1_U13.top_add_43s_43s_43_2_1_Adder_10_U.clk )
\add_43s_43s_43_2_1_U13.top_add_43s_43s_43_2_1_Adder_10_U.carry_s1  <= _129_;
assign _128_ = \add_43s_43s_43_2_1_U13.top_add_43s_43s_43_2_1_Adder_10_U.ce  ? \add_43s_43s_43_2_1_U13.top_add_43s_43s_43_2_1_Adder_10_U.b [42:21] : \add_43s_43s_43_2_1_U13.top_add_43s_43s_43_2_1_Adder_10_U.bin_s1 ;
assign _127_ = \add_43s_43s_43_2_1_U13.top_add_43s_43s_43_2_1_Adder_10_U.ce  ? \add_43s_43s_43_2_1_U13.top_add_43s_43s_43_2_1_Adder_10_U.a [42:21] : \add_43s_43s_43_2_1_U13.top_add_43s_43s_43_2_1_Adder_10_U.ain_s1 ;
assign _129_ = \add_43s_43s_43_2_1_U13.top_add_43s_43s_43_2_1_Adder_10_U.ce  ? \add_43s_43s_43_2_1_U13.top_add_43s_43s_43_2_1_Adder_10_U.facout_s1  : \add_43s_43s_43_2_1_U13.top_add_43s_43s_43_2_1_Adder_10_U.carry_s1 ;
assign _130_ = \add_43s_43s_43_2_1_U13.top_add_43s_43s_43_2_1_Adder_10_U.ce  ? \add_43s_43s_43_2_1_U13.top_add_43s_43s_43_2_1_Adder_10_U.fas_s1  : \add_43s_43s_43_2_1_U13.top_add_43s_43s_43_2_1_Adder_10_U.sum_s1 ;
assign _131_ = \add_43s_43s_43_2_1_U13.top_add_43s_43s_43_2_1_Adder_10_U.u1.a  + \add_43s_43s_43_2_1_U13.top_add_43s_43s_43_2_1_Adder_10_U.u1.b ;
assign { \add_43s_43s_43_2_1_U13.top_add_43s_43s_43_2_1_Adder_10_U.u1.cout , \add_43s_43s_43_2_1_U13.top_add_43s_43s_43_2_1_Adder_10_U.u1.s  } = _131_ + \add_43s_43s_43_2_1_U13.top_add_43s_43s_43_2_1_Adder_10_U.u1.cin ;
assign _132_ = \add_43s_43s_43_2_1_U13.top_add_43s_43s_43_2_1_Adder_10_U.u2.a  + \add_43s_43s_43_2_1_U13.top_add_43s_43s_43_2_1_Adder_10_U.u2.b ;
assign { \add_43s_43s_43_2_1_U13.top_add_43s_43s_43_2_1_Adder_10_U.u2.cout , \add_43s_43s_43_2_1_U13.top_add_43s_43s_43_2_1_Adder_10_U.u2.s  } = _132_ + \add_43s_43s_43_2_1_U13.top_add_43s_43s_43_2_1_Adder_10_U.u2.cin ;
always @(posedge \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.clk )
\add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.bin_s1  <= _134_;
always @(posedge \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.clk )
\add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.ain_s1  <= _133_;
always @(posedge \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.clk )
\add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.sum_s1  <= _136_;
always @(posedge \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.clk )
\add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.carry_s1  <= _135_;
assign _134_ = \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.ce  ? \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.b [5:3] : \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.bin_s1 ;
assign _133_ = \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.ce  ? \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.a [5:3] : \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.ain_s1 ;
assign _135_ = \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.ce  ? \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.facout_s1  : \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.carry_s1 ;
assign _136_ = \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.ce  ? \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.fas_s1  : \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.sum_s1 ;
assign _137_ = \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.u1.a  + \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.u1.b ;
assign { \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.u1.cout , \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.u1.s  } = _137_ + \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.u1.cin ;
assign _138_ = \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.u2.a  + \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.u2.b ;
assign { \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.u2.cout , \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.u2.s  } = _138_ + \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.u2.cin ;
always @(posedge \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.clk )
\add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.bin_s1  <= _140_;
always @(posedge \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.clk )
\add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.ain_s1  <= _139_;
always @(posedge \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.clk )
\add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.sum_s1  <= _142_;
always @(posedge \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.clk )
\add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.carry_s1  <= _141_;
assign _140_ = \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.ce  ? \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.b [7:4] : \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.bin_s1 ;
assign _139_ = \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.ce  ? \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.a [7:4] : \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.ain_s1 ;
assign _141_ = \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.ce  ? \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.facout_s1  : \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.carry_s1 ;
assign _142_ = \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.ce  ? \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.fas_s1  : \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.sum_s1 ;
assign _143_ = \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.u1.a  + \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.u1.b ;
assign { \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.u1.cout , \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.u1.s  } = _143_ + \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.u1.cin ;
assign _144_ = \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.u2.a  + \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.u2.b ;
assign { \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.u2.cout , \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.u2.s  } = _144_ + \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.u2.cin ;
always @(posedge \add_8s_8ns_8_2_1_U5.top_add_8s_8ns_8_2_1_Adder_4_U.clk )
\add_8s_8ns_8_2_1_U5.top_add_8s_8ns_8_2_1_Adder_4_U.bin_s1  <= _146_;
always @(posedge \add_8s_8ns_8_2_1_U5.top_add_8s_8ns_8_2_1_Adder_4_U.clk )
\add_8s_8ns_8_2_1_U5.top_add_8s_8ns_8_2_1_Adder_4_U.ain_s1  <= _145_;
always @(posedge \add_8s_8ns_8_2_1_U5.top_add_8s_8ns_8_2_1_Adder_4_U.clk )
\add_8s_8ns_8_2_1_U5.top_add_8s_8ns_8_2_1_Adder_4_U.sum_s1  <= _148_;
always @(posedge \add_8s_8ns_8_2_1_U5.top_add_8s_8ns_8_2_1_Adder_4_U.clk )
\add_8s_8ns_8_2_1_U5.top_add_8s_8ns_8_2_1_Adder_4_U.carry_s1  <= _147_;
assign _146_ = \add_8s_8ns_8_2_1_U5.top_add_8s_8ns_8_2_1_Adder_4_U.ce  ? \add_8s_8ns_8_2_1_U5.top_add_8s_8ns_8_2_1_Adder_4_U.b [7:4] : \add_8s_8ns_8_2_1_U5.top_add_8s_8ns_8_2_1_Adder_4_U.bin_s1 ;
assign _145_ = \add_8s_8ns_8_2_1_U5.top_add_8s_8ns_8_2_1_Adder_4_U.ce  ? \add_8s_8ns_8_2_1_U5.top_add_8s_8ns_8_2_1_Adder_4_U.a [7:4] : \add_8s_8ns_8_2_1_U5.top_add_8s_8ns_8_2_1_Adder_4_U.ain_s1 ;
assign _147_ = \add_8s_8ns_8_2_1_U5.top_add_8s_8ns_8_2_1_Adder_4_U.ce  ? \add_8s_8ns_8_2_1_U5.top_add_8s_8ns_8_2_1_Adder_4_U.facout_s1  : \add_8s_8ns_8_2_1_U5.top_add_8s_8ns_8_2_1_Adder_4_U.carry_s1 ;
assign _148_ = \add_8s_8ns_8_2_1_U5.top_add_8s_8ns_8_2_1_Adder_4_U.ce  ? \add_8s_8ns_8_2_1_U5.top_add_8s_8ns_8_2_1_Adder_4_U.fas_s1  : \add_8s_8ns_8_2_1_U5.top_add_8s_8ns_8_2_1_Adder_4_U.sum_s1 ;
assign _149_ = \add_8s_8ns_8_2_1_U5.top_add_8s_8ns_8_2_1_Adder_4_U.u1.a  + \add_8s_8ns_8_2_1_U5.top_add_8s_8ns_8_2_1_Adder_4_U.u1.b ;
assign { \add_8s_8ns_8_2_1_U5.top_add_8s_8ns_8_2_1_Adder_4_U.u1.cout , \add_8s_8ns_8_2_1_U5.top_add_8s_8ns_8_2_1_Adder_4_U.u1.s  } = _149_ + \add_8s_8ns_8_2_1_U5.top_add_8s_8ns_8_2_1_Adder_4_U.u1.cin ;
assign _150_ = \add_8s_8ns_8_2_1_U5.top_add_8s_8ns_8_2_1_Adder_4_U.u2.a  + \add_8s_8ns_8_2_1_U5.top_add_8s_8ns_8_2_1_Adder_4_U.u2.b ;
assign { \add_8s_8ns_8_2_1_U5.top_add_8s_8ns_8_2_1_Adder_4_U.u2.cout , \add_8s_8ns_8_2_1_U5.top_add_8s_8ns_8_2_1_Adder_4_U.u2.s  } = _150_ + \add_8s_8ns_8_2_1_U5.top_add_8s_8ns_8_2_1_Adder_4_U.u2.cin ;
always @(posedge \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.clk )
\add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.bin_s1  <= _152_;
always @(posedge \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.clk )
\add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.ain_s1  <= _151_;
always @(posedge \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.clk )
\add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.sum_s1  <= _154_;
always @(posedge \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.clk )
\add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.carry_s1  <= _153_;
assign _152_ = \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.ce  ? \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.b [8:4] : \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.bin_s1 ;
assign _151_ = \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.ce  ? \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.a [8:4] : \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.ain_s1 ;
assign _153_ = \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.ce  ? \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.facout_s1  : \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.carry_s1 ;
assign _154_ = \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.ce  ? \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.fas_s1  : \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.sum_s1 ;
assign _155_ = \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.u1.a  + \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.u1.b ;
assign { \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.u1.cout , \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.u1.s  } = _155_ + \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.u1.cin ;
assign _156_ = \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.u2.a  + \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.u2.b ;
assign { \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.u2.cout , \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.u2.s  } = _156_ + \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.u2.cin ;
assign \sub_5ns_5ns_5_2_1_U3.top_sub_5ns_5ns_5_2_1_Adder_2_U.bin_s0  = ~ \sub_5ns_5ns_5_2_1_U3.top_sub_5ns_5ns_5_2_1_Adder_2_U.b ;
always @(posedge \sub_5ns_5ns_5_2_1_U3.top_sub_5ns_5ns_5_2_1_Adder_2_U.clk )
\sub_5ns_5ns_5_2_1_U3.top_sub_5ns_5ns_5_2_1_Adder_2_U.bin_s1  <= _158_;
always @(posedge \sub_5ns_5ns_5_2_1_U3.top_sub_5ns_5ns_5_2_1_Adder_2_U.clk )
\sub_5ns_5ns_5_2_1_U3.top_sub_5ns_5ns_5_2_1_Adder_2_U.ain_s1  <= _157_;
always @(posedge \sub_5ns_5ns_5_2_1_U3.top_sub_5ns_5ns_5_2_1_Adder_2_U.clk )
\sub_5ns_5ns_5_2_1_U3.top_sub_5ns_5ns_5_2_1_Adder_2_U.sum_s1  <= _160_;
always @(posedge \sub_5ns_5ns_5_2_1_U3.top_sub_5ns_5ns_5_2_1_Adder_2_U.clk )
\sub_5ns_5ns_5_2_1_U3.top_sub_5ns_5ns_5_2_1_Adder_2_U.carry_s1  <= _159_;
assign _158_ = \sub_5ns_5ns_5_2_1_U3.top_sub_5ns_5ns_5_2_1_Adder_2_U.ce  ? \sub_5ns_5ns_5_2_1_U3.top_sub_5ns_5ns_5_2_1_Adder_2_U.bin_s0 [4:2] : \sub_5ns_5ns_5_2_1_U3.top_sub_5ns_5ns_5_2_1_Adder_2_U.bin_s1 ;
assign _157_ = \sub_5ns_5ns_5_2_1_U3.top_sub_5ns_5ns_5_2_1_Adder_2_U.ce  ? \sub_5ns_5ns_5_2_1_U3.top_sub_5ns_5ns_5_2_1_Adder_2_U.a [4:2] : \sub_5ns_5ns_5_2_1_U3.top_sub_5ns_5ns_5_2_1_Adder_2_U.ain_s1 ;
assign _159_ = \sub_5ns_5ns_5_2_1_U3.top_sub_5ns_5ns_5_2_1_Adder_2_U.ce  ? \sub_5ns_5ns_5_2_1_U3.top_sub_5ns_5ns_5_2_1_Adder_2_U.facout_s1  : \sub_5ns_5ns_5_2_1_U3.top_sub_5ns_5ns_5_2_1_Adder_2_U.carry_s1 ;
assign _160_ = \sub_5ns_5ns_5_2_1_U3.top_sub_5ns_5ns_5_2_1_Adder_2_U.ce  ? \sub_5ns_5ns_5_2_1_U3.top_sub_5ns_5ns_5_2_1_Adder_2_U.fas_s1  : \sub_5ns_5ns_5_2_1_U3.top_sub_5ns_5ns_5_2_1_Adder_2_U.sum_s1 ;
assign _161_ = \sub_5ns_5ns_5_2_1_U3.top_sub_5ns_5ns_5_2_1_Adder_2_U.u1.a  + \sub_5ns_5ns_5_2_1_U3.top_sub_5ns_5ns_5_2_1_Adder_2_U.u1.b ;
assign { \sub_5ns_5ns_5_2_1_U3.top_sub_5ns_5ns_5_2_1_Adder_2_U.u1.cout , \sub_5ns_5ns_5_2_1_U3.top_sub_5ns_5ns_5_2_1_Adder_2_U.u1.s  } = _161_ + \sub_5ns_5ns_5_2_1_U3.top_sub_5ns_5ns_5_2_1_Adder_2_U.u1.cin ;
assign _162_ = \sub_5ns_5ns_5_2_1_U3.top_sub_5ns_5ns_5_2_1_Adder_2_U.u2.a  + \sub_5ns_5ns_5_2_1_U3.top_sub_5ns_5ns_5_2_1_Adder_2_U.u2.b ;
assign { \sub_5ns_5ns_5_2_1_U3.top_sub_5ns_5ns_5_2_1_Adder_2_U.u2.cout , \sub_5ns_5ns_5_2_1_U3.top_sub_5ns_5ns_5_2_1_Adder_2_U.u2.s  } = _162_ + \sub_5ns_5ns_5_2_1_U3.top_sub_5ns_5ns_5_2_1_Adder_2_U.u2.cin ;
assign _163_ = | p_Result_1_reg_948;
assign _164_ = | op_1[3:1];
assign _165_ = p_Result_1_reg_948 != 4'hf;
assign _166_ = op_1[3:1] != 3'h7;
assign _167_ = | trunc_ln851_1_reg_1011;
assign _168_ = | op_12[2:0];
assign _169_ = | op_16[9:0];
assign or_ln340_fu_299_p2 = p_Result_8_reg_853 | overflow_fu_284_p2;
assign or_ln384_fu_499_p2 = underflow_1_fu_487_p2 | overflow_1_reg_990;
assign or_ln785_1_fu_461_p2 = p_Result_9_reg_964 | icmp_ln768_1_reg_970;
assign or_ln785_2_fu_334_p2 = xor_ln785_1_fu_329_p2 | p_Result_8_reg_853;
assign or_ln785_3_fu_350_p2 = and_ln785_1_fu_345_p2 | and_ln340_reg_891;
assign or_ln785_fu_275_p2 = newsignbit_reg_860 | icmp_ln768_reg_868;
assign or_ln786_1_fu_482_p2 = xor_ln786_1_fu_477_p2 | icmp_ln786_1_reg_975;
assign or_ln786_fu_294_p2 = xor_ln786_fu_289_p2 | icmp_ln786_reg_873;
always @(posedge ap_clk)
select_ln1192_reg_896[2:0] <= 3'h0;
always @(posedge ap_clk)
zext_ln703_reg_938[4] <= 1'h0;
always @(posedge ap_clk)
p_Val2_3_reg_959[6:0] <= 7'h00;
always @(posedge ap_clk)
tmp_5_reg_1083 <= _047_;
always @(posedge ap_clk)
sext_ln850_reg_1046 <= _046_;
always @(posedge ap_clk)
select_ln353_reg_1187 <= _044_;
always @(posedge ap_clk)
ret_V_22_reg_1212 <= _037_;
always @(posedge ap_clk)
ret_V_21_reg_1170 <= _036_;
always @(posedge ap_clk)
ret_V_20_cast_reg_1175 <= _034_;
always @(posedge ap_clk)
ret_V_19_reg_1120 <= _033_;
always @(posedge ap_clk)
ret_V_17_reg_1058 <= _031_;
always @(posedge ap_clk)
ret_V_18_reg_1103 <= _032_;
always @(posedge ap_clk)
ret_V_17_cast_reg_1108 <= _030_;
always @(posedge ap_clk)
ret_V_4_reg_1031 <= _039_;
always @(posedge ap_clk)
ret_V_16_reg_1036 <= _029_;
always @(posedge ap_clk)
tmp_reg_1041 <= _048_;
always @(posedge ap_clk)
ret_V_14_reg_914 <= _028_;
always @(posedge ap_clk)
ret_V_reg_919 <= _040_;
always @(posedge ap_clk)
trunc_ln851_reg_926 <= _051_;
always @(posedge ap_clk)
r_1_reg_931 <= _026_;
always @(posedge ap_clk)
zext_ln703_reg_938[3:0] <= _052_;
always @(posedge ap_clk)
trunc_ln728_reg_943 <= _049_;
always @(posedge ap_clk)
p_Result_1_reg_948 <= _022_;
always @(posedge ap_clk)
ret_V_2_reg_985 <= _038_;
always @(posedge ap_clk)
overflow_1_reg_990 <= _021_;
always @(posedge ap_clk)
or_ln785_reg_885 <= _020_;
always @(posedge ap_clk)
op_9_V_reg_996 <= _019_;
always @(posedge ap_clk)
select_ln1193_reg_1001 <= _043_;
always @(posedge ap_clk)
select_ln850_3_reg_1006 <= _045_;
always @(posedge ap_clk)
trunc_ln851_1_reg_1011 <= _050_;
always @(posedge ap_clk)
op_3_V_reg_901 <= _018_;
always @(posedge ap_clk)
op_29_V_reg_1202 <= _017_;
always @(posedge ap_clk)
op_27_V_reg_1150 <= _016_;
always @(posedge ap_clk)
op_22_V_reg_1068 <= _015_;
always @(posedge ap_clk)
icmp_ln851_3_reg_1165 <= _012_;
always @(posedge ap_clk)
icmp_ln851_2_reg_1098 <= _011_;
always @(posedge ap_clk)
icmp_ln851_1_reg_1026 <= _010_;
always @(posedge ap_clk)
p_Result_8_reg_853 <= _023_;
always @(posedge ap_clk)
newsignbit_reg_860 <= _014_;
always @(posedge ap_clk)
icmp_ln768_reg_868 <= _007_;
always @(posedge ap_clk)
icmp_ln786_reg_873 <= _009_;
always @(posedge ap_clk)
r_reg_879 <= _027_;
always @(posedge ap_clk)
icmp_ln851_reg_954 <= _013_;
always @(posedge ap_clk)
p_Val2_3_reg_959[7] <= _025_;
always @(posedge ap_clk)
p_Result_9_reg_964 <= _024_;
always @(posedge ap_clk)
icmp_ln768_1_reg_970 <= _006_;
always @(posedge ap_clk)
icmp_ln786_1_reg_975 <= _008_;
always @(posedge ap_clk)
ret_reg_980 <= _041_;
always @(posedge ap_clk)
and_ln340_reg_891 <= _004_;
always @(posedge ap_clk)
select_ln1192_reg_896[8:3] <= _042_;
always @(posedge ap_clk)
ret_V_20_reg_1140 <= _035_;
always @(posedge ap_clk)
add_ln69_reg_1145 <= _003_;
always @(posedge ap_clk)
add_ln691_reg_1053 <= _002_;
always @(posedge ap_clk)
add_ln691_3_reg_1182 <= _001_;
always @(posedge ap_clk)
add_ln691_2_reg_1115 <= _000_;
always @(posedge ap_clk)
ap_CS_fsm <= _005_;
assign _053_ = _058_ ? 2'h2 : 2'h1;
assign _170_ = ap_CS_fsm == 1'h1;
function [36:0] _507_;
input [36:0] a;
input [1368:0] b;
input [36:0] s;
case (s)
37'b0000000000000000000000000000000000001:
_507_ = b[36:0];
37'b0000000000000000000000000000000000010:
_507_ = b[73:37];
37'b0000000000000000000000000000000000100:
_507_ = b[110:74];
37'b0000000000000000000000000000000001000:
_507_ = b[147:111];
37'b0000000000000000000000000000000010000:
_507_ = b[184:148];
37'b0000000000000000000000000000000100000:
_507_ = b[221:185];
37'b0000000000000000000000000000001000000:
_507_ = b[258:222];
37'b0000000000000000000000000000010000000:
_507_ = b[295:259];
37'b0000000000000000000000000000100000000:
_507_ = b[332:296];
37'b0000000000000000000000000001000000000:
_507_ = b[369:333];
37'b0000000000000000000000000010000000000:
_507_ = b[406:370];
37'b0000000000000000000000000100000000000:
_507_ = b[443:407];
37'b0000000000000000000000001000000000000:
_507_ = b[480:444];
37'b0000000000000000000000010000000000000:
_507_ = b[517:481];
37'b0000000000000000000000100000000000000:
_507_ = b[554:518];
37'b0000000000000000000001000000000000000:
_507_ = b[591:555];
37'b0000000000000000000010000000000000000:
_507_ = b[628:592];
37'b0000000000000000000100000000000000000:
_507_ = b[665:629];
37'b0000000000000000001000000000000000000:
_507_ = b[702:666];
37'b0000000000000000010000000000000000000:
_507_ = b[739:703];
37'b0000000000000000100000000000000000000:
_507_ = b[776:740];
37'b0000000000000001000000000000000000000:
_507_ = b[813:777];
37'b0000000000000010000000000000000000000:
_507_ = b[850:814];
37'b0000000000000100000000000000000000000:
_507_ = b[887:851];
37'b0000000000001000000000000000000000000:
_507_ = b[924:888];
37'b0000000000010000000000000000000000000:
_507_ = b[961:925];
37'b0000000000100000000000000000000000000:
_507_ = b[998:962];
37'b0000000001000000000000000000000000000:
_507_ = b[1035:999];
37'b0000000010000000000000000000000000000:
_507_ = b[1072:1036];
37'b0000000100000000000000000000000000000:
_507_ = b[1109:1073];
37'b0000001000000000000000000000000000000:
_507_ = b[1146:1110];
37'b0000010000000000000000000000000000000:
_507_ = b[1183:1147];
37'b0000100000000000000000000000000000000:
_507_ = b[1220:1184];
37'b0001000000000000000000000000000000000:
_507_ = b[1257:1221];
37'b0010000000000000000000000000000000000:
_507_ = b[1294:1258];
37'b0100000000000000000000000000000000000:
_507_ = b[1331:1295];
37'b1000000000000000000000000000000000000:
_507_ = b[1368:1332];
37'b0000000000000000000000000000000000000:
_507_ = a;
default:
_507_ = 37'bx;
endcase
endfunction
assign ap_NS_fsm = _507_(37'hxxxxxxxxxx, { 35'h000000000, _053_, 1332'h000000002000000002000000002000000002000000002000000002000000002000000002000000002000000002000000002000000002000000002000000002000000002000000002000000002000000002000000002000000002000000002000000002000000002000000002000000002000000002000000002000000002000000002000000002000000002000000002000000002000000002000000002000000000000000001 }, { _170_, _206_, _205_, _204_, _203_, _202_, _201_, _200_, _199_, _198_, _197_, _196_, _195_, _194_, _193_, _192_, _191_, _190_, _189_, _188_, _187_, _186_, _185_, _184_, _183_, _182_, _181_, _180_, _179_, _178_, _177_, _176_, _175_, _174_, _173_, _172_, _171_ });
assign _171_ = ap_CS_fsm == 37'h1000000000;
assign _172_ = ap_CS_fsm == 36'h800000000;
assign _173_ = ap_CS_fsm == 35'h400000000;
assign _174_ = ap_CS_fsm == 34'h200000000;
assign _175_ = ap_CS_fsm == 33'h100000000;
assign _176_ = ap_CS_fsm == 32'd2147483648;
assign _177_ = ap_CS_fsm == 31'h40000000;
assign _178_ = ap_CS_fsm == 30'h20000000;
assign _179_ = ap_CS_fsm == 29'h10000000;
assign _180_ = ap_CS_fsm == 28'h8000000;
assign _181_ = ap_CS_fsm == 27'h4000000;
assign _182_ = ap_CS_fsm == 26'h2000000;
assign _183_ = ap_CS_fsm == 25'h1000000;
assign _184_ = ap_CS_fsm == 24'h800000;
assign _185_ = ap_CS_fsm == 23'h400000;
assign _186_ = ap_CS_fsm == 22'h200000;
assign _187_ = ap_CS_fsm == 21'h100000;
assign _188_ = ap_CS_fsm == 20'h80000;
assign _189_ = ap_CS_fsm == 19'h40000;
assign _190_ = ap_CS_fsm == 18'h20000;
assign _191_ = ap_CS_fsm == 17'h10000;
assign _192_ = ap_CS_fsm == 16'h8000;
assign _193_ = ap_CS_fsm == 15'h4000;
assign _194_ = ap_CS_fsm == 14'h2000;
assign _195_ = ap_CS_fsm == 13'h1000;
assign _196_ = ap_CS_fsm == 12'h800;
assign _197_ = ap_CS_fsm == 11'h400;
assign _198_ = ap_CS_fsm == 10'h200;
assign _199_ = ap_CS_fsm == 9'h100;
assign _200_ = ap_CS_fsm == 8'h80;
assign _201_ = ap_CS_fsm == 7'h40;
assign _202_ = ap_CS_fsm == 6'h20;
assign _203_ = ap_CS_fsm == 5'h10;
assign _204_ = ap_CS_fsm == 4'h8;
assign _205_ = ap_CS_fsm == 3'h4;
assign _206_ = ap_CS_fsm == 2'h2;
assign op_31_ap_vld = ap_CS_fsm[36] ? 1'h1 : 1'h0;
assign ap_idle = _057_ ? 1'h1 : 1'h0;
assign _047_ = ap_CS_fsm[16] ? grp_fu_632_p2[32:1] : tmp_5_reg_1083;
assign _046_ = ap_CS_fsm[10] ? { tmp_reg_1041[6], tmp_reg_1041 } : sext_ln850_reg_1046;
assign _044_ = ap_CS_fsm[30] ? select_ln353_fu_793_p3 : select_ln353_reg_1187;
assign _037_ = ap_CS_fsm[34] ? grp_fu_842_p2 : ret_V_22_reg_1212;
assign _034_ = ap_CS_fsm[27] ? grp_fu_750_p2[41:10] : ret_V_20_cast_reg_1175;
assign _036_ = ap_CS_fsm[27] ? grp_fu_750_p2 : ret_V_21_reg_1170;
assign _033_ = ap_CS_fsm[21] ? ret_V_19_fu_706_p3 : ret_V_19_reg_1120;
assign _031_ = ap_CS_fsm[12] ? ret_V_17_fu_594_p3 : ret_V_17_reg_1058;
assign _030_ = ap_CS_fsm[18] ? grp_fu_663_p2[34:3] : ret_V_17_cast_reg_1108;
assign _032_ = ap_CS_fsm[18] ? grp_fu_663_p2 : ret_V_18_reg_1103;
assign _048_ = ap_CS_fsm[9] ? grp_fu_552_p2[13:7] : tmp_reg_1041;
assign _029_ = ap_CS_fsm[9] ? grp_fu_552_p2 : ret_V_16_reg_1036;
assign _039_ = ap_CS_fsm[9] ? grp_fu_534_p2 : ret_V_4_reg_1031;
assign _022_ = ap_CS_fsm[4] ? ret_V_15_fu_391_p3[4:1] : p_Result_1_reg_948;
assign _049_ = ap_CS_fsm[4] ? ret_V_15_fu_391_p3[0] : trunc_ln728_reg_943;
assign _052_ = ap_CS_fsm[4] ? r_reg_879 : zext_ln703_reg_938[3:0];
assign _026_ = ap_CS_fsm[4] ? r_1_fu_383_p2 : r_1_reg_931;
assign _051_ = ap_CS_fsm[4] ? grp_fu_364_p2[2:0] : trunc_ln851_reg_926;
assign _040_ = ap_CS_fsm[4] ? grp_fu_364_p2[8:3] : ret_V_reg_919;
assign _028_ = ap_CS_fsm[4] ? grp_fu_364_p2 : ret_V_14_reg_914;
assign _021_ = ap_CS_fsm[6] ? overflow_1_fu_465_p2 : overflow_1_reg_990;
assign _038_ = ap_CS_fsm[6] ? grp_fu_420_p2 : ret_V_2_reg_985;
assign _020_ = ap_CS_fsm[1] ? or_ln785_fu_275_p2 : or_ln785_reg_885;
assign _050_ = ap_CS_fsm[7] ? op_9_V_fu_504_p3[6:0] : trunc_ln851_1_reg_1011;
assign _045_ = ap_CS_fsm[7] ? select_ln850_3_fu_523_p3 : select_ln850_3_reg_1006;
assign _043_ = ap_CS_fsm[7] ? select_ln1193_fu_511_p3 : select_ln1193_reg_1001;
assign _019_ = ap_CS_fsm[7] ? op_9_V_fu_504_p3 : op_9_V_reg_996;
assign _018_ = ap_CS_fsm[3] ? op_3_V_fu_355_p2 : op_3_V_reg_901;
assign _017_ = ap_CS_fsm[32] ? grp_fu_822_p2[32:1] : op_29_V_reg_1202;
assign _016_ = ap_CS_fsm[25] ? grp_fu_731_p2 : op_27_V_reg_1150;
assign _015_ = ap_CS_fsm[14] ? grp_fu_605_p2 : op_22_V_reg_1068;
assign _012_ = ap_CS_fsm[26] ? icmp_ln851_3_fu_760_p2 : icmp_ln851_3_reg_1165;
assign _011_ = ap_CS_fsm[17] ? icmp_ln851_2_fu_673_p2 : icmp_ln851_2_reg_1098;
assign _010_ = ap_CS_fsm[8] ? icmp_ln851_1_fu_558_p2 : icmp_ln851_1_reg_1026;
assign _027_ = ap_CS_fsm[0] ? r_fu_267_p3 : r_reg_879;
assign _009_ = ap_CS_fsm[0] ? icmp_ln786_fu_255_p2 : icmp_ln786_reg_873;
assign _007_ = ap_CS_fsm[0] ? icmp_ln768_fu_249_p2 : icmp_ln768_reg_868;
assign _014_ = ap_CS_fsm[0] ? op_1[0] : newsignbit_reg_860;
assign _023_ = ap_CS_fsm[0] ? op_1[3] : p_Result_8_reg_853;
assign _041_ = ap_CS_fsm[5] ? ret_fu_455_p2 : ret_reg_980;
assign _008_ = ap_CS_fsm[5] ? icmp_ln786_1_fu_450_p2 : icmp_ln786_1_reg_975;
assign _006_ = ap_CS_fsm[5] ? icmp_ln768_1_fu_445_p2 : icmp_ln768_1_reg_970;
assign _024_ = ap_CS_fsm[5] ? p_Result_9_fu_439_p2 : p_Result_9_reg_964;
assign _025_ = ap_CS_fsm[5] ? trunc_ln728_reg_943 : p_Val2_3_reg_959[7];
assign _013_ = ap_CS_fsm[5] ? icmp_ln851_fu_415_p2 : icmp_ln851_reg_954;
assign _042_ = ap_CS_fsm[2] ? select_ln1192_fu_316_p3[8:3] : select_ln1192_reg_896[8:3];
assign _004_ = ap_CS_fsm[2] ? and_ln340_fu_310_p2 : and_ln340_reg_891;
assign _003_ = ap_CS_fsm[23] ? grp_fu_725_p2 : add_ln69_reg_1145;
assign _035_ = ap_CS_fsm[23] ? grp_fu_717_p2 : ret_V_20_reg_1140;
assign _002_ = _056_ ? grp_fu_576_p2 : add_ln691_reg_1053;
assign _001_ = _055_ ? grp_fu_776_p2 : add_ln691_3_reg_1182;
assign _000_ = _054_ ? grp_fu_689_p2 : add_ln691_2_reg_1115;
assign _005_ = ap_rst ? 37'h0000000001 : ap_NS_fsm;
assign icmp_ln768_1_fu_445_p2 = _163_ ? 1'h1 : 1'h0;
assign icmp_ln768_fu_249_p2 = _164_ ? 1'h1 : 1'h0;
assign icmp_ln786_1_fu_450_p2 = _165_ ? 1'h1 : 1'h0;
assign icmp_ln786_fu_255_p2 = _166_ ? 1'h1 : 1'h0;
assign icmp_ln851_1_fu_558_p2 = _167_ ? 1'h1 : 1'h0;
assign icmp_ln851_2_fu_673_p2 = _168_ ? 1'h1 : 1'h0;
assign icmp_ln851_3_fu_760_p2 = _169_ ? 1'h1 : 1'h0;
assign icmp_ln851_fu_415_p2 = _060_ ? 1'h1 : 1'h0;
assign op_9_V_fu_504_p3 = or_ln384_fu_499_p2 ? select_ln384_fu_492_p3 : p_Val2_3_reg_959;
assign p_Result_9_fu_439_p2 = trunc_ln728_reg_943 ? 1'h1 : 1'h0;
assign r_fu_267_p3 = op_2 ? { op_1[2:0], 1'h0 } : op_1;
assign ret_2_fu_425_p3 = r_1_reg_931 ? 2'h3 : 2'h0;
assign ret_V_15_fu_391_p3 = op_3_V_reg_901 ? 5'h1f : { 1'h0, r_reg_879 };
assign ret_V_17_fu_594_p3 = ret_V_16_reg_1036[13] ? select_ln850_1_fu_589_p3 : sext_ln850_reg_1046;
assign ret_V_19_fu_706_p3 = ret_V_18_reg_1103[35] ? select_ln850_2_fu_701_p3 : ret_V_17_cast_reg_1108;
assign select_ln1192_fu_316_p3 = op_6 ? 9'h1f8 : 9'h000;
assign select_ln1193_fu_511_p3 = op_3_V_reg_901 ? 5'h1f : 5'h00;
assign select_ln353_fu_793_p3 = ret_V_21_reg_1170[42] ? select_ln850_4_fu_788_p3 : ret_V_20_cast_reg_1175;
assign select_ln384_fu_492_p3 = overflow_1_reg_990 ? 8'h7f : 8'h80;
assign select_ln850_1_fu_589_p3 = icmp_ln851_1_reg_1026 ? add_ln691_reg_1053 : sext_ln850_reg_1046;
assign select_ln850_2_fu_701_p3 = icmp_ln851_2_reg_1098 ? add_ln691_2_reg_1115 : ret_V_17_cast_reg_1108;
assign select_ln850_3_fu_523_p3 = ret_V_14_reg_914[8] ? select_ln850_fu_518_p3 : ret_V_reg_919;
assign select_ln850_4_fu_788_p3 = icmp_ln851_3_reg_1165 ? add_ln691_3_reg_1182 : ret_V_20_cast_reg_1175;
assign select_ln850_fu_518_p3 = icmp_ln851_reg_954 ? ret_V_reg_919 : ret_V_2_reg_985;
assign ap_CS_fsm_state1 = ap_CS_fsm[0];
assign ap_CS_fsm_state10 = ap_CS_fsm[9];
assign ap_CS_fsm_state11 = ap_CS_fsm[10];
assign ap_CS_fsm_state12 = ap_CS_fsm[11];
assign ap_CS_fsm_state13 = ap_CS_fsm[12];
assign ap_CS_fsm_state14 = ap_CS_fsm[13];
assign ap_CS_fsm_state15 = ap_CS_fsm[14];
assign ap_CS_fsm_state16 = ap_CS_fsm[15];
assign ap_CS_fsm_state17 = ap_CS_fsm[16];
assign ap_CS_fsm_state18 = ap_CS_fsm[17];
assign ap_CS_fsm_state19 = ap_CS_fsm[18];
assign ap_CS_fsm_state2 = ap_CS_fsm[1];
assign ap_CS_fsm_state20 = ap_CS_fsm[19];
assign ap_CS_fsm_state21 = ap_CS_fsm[20];
assign ap_CS_fsm_state22 = ap_CS_fsm[21];
assign ap_CS_fsm_state23 = ap_CS_fsm[22];
assign ap_CS_fsm_state24 = ap_CS_fsm[23];
assign ap_CS_fsm_state25 = ap_CS_fsm[24];
assign ap_CS_fsm_state26 = ap_CS_fsm[25];
assign ap_CS_fsm_state27 = ap_CS_fsm[26];
assign ap_CS_fsm_state28 = ap_CS_fsm[27];
assign ap_CS_fsm_state29 = ap_CS_fsm[28];
assign ap_CS_fsm_state3 = ap_CS_fsm[2];
assign ap_CS_fsm_state30 = ap_CS_fsm[29];
assign ap_CS_fsm_state31 = ap_CS_fsm[30];
assign ap_CS_fsm_state32 = ap_CS_fsm[31];
assign ap_CS_fsm_state33 = ap_CS_fsm[32];
assign ap_CS_fsm_state34 = ap_CS_fsm[33];
assign ap_CS_fsm_state35 = ap_CS_fsm[34];
assign ap_CS_fsm_state36 = ap_CS_fsm[35];
assign ap_CS_fsm_state37 = ap_CS_fsm[36];
assign ap_CS_fsm_state4 = ap_CS_fsm[3];
assign ap_CS_fsm_state5 = ap_CS_fsm[4];
assign ap_CS_fsm_state6 = ap_CS_fsm[5];
assign ap_CS_fsm_state7 = ap_CS_fsm[6];
assign ap_CS_fsm_state8 = ap_CS_fsm[7];
assign ap_CS_fsm_state9 = ap_CS_fsm[8];
assign ap_done = op_31_ap_vld;
assign ap_ready = op_31_ap_vld;
assign grp_fu_364_p1 = { op_0[7], op_0 };
assign grp_fu_552_p0 = { select_ln850_3_reg_1006[5], select_ln850_3_reg_1006, 7'h00 };
assign grp_fu_552_p1 = { op_9_V_reg_996[7], op_9_V_reg_996[7], op_9_V_reg_996[7], op_9_V_reg_996[7], op_9_V_reg_996[7], op_9_V_reg_996[7], op_9_V_reg_996 };
assign grp_fu_576_p0 = { tmp_reg_1041[6], tmp_reg_1041 };
assign grp_fu_605_p1 = { 6'h00, op_10 };
assign grp_fu_632_p0 = { op_22_V_reg_1068[7], op_22_V_reg_1068[7], op_22_V_reg_1068[7], op_22_V_reg_1068[7], op_22_V_reg_1068[7], op_22_V_reg_1068[7], op_22_V_reg_1068[7], op_22_V_reg_1068[7], op_22_V_reg_1068[7], op_22_V_reg_1068[7], op_22_V_reg_1068[7], op_22_V_reg_1068[7], op_22_V_reg_1068[7], op_22_V_reg_1068[7], op_22_V_reg_1068[7], op_22_V_reg_1068[7], op_22_V_reg_1068[7], op_22_V_reg_1068[7], op_22_V_reg_1068[7], op_22_V_reg_1068[7], op_22_V_reg_1068[7], op_22_V_reg_1068[7], op_22_V_reg_1068[7], op_22_V_reg_1068[7], op_22_V_reg_1068, 1'h0 };
assign grp_fu_632_p1 = { ret_V_4_reg_1031[4], ret_V_4_reg_1031[4], ret_V_4_reg_1031[4], ret_V_4_reg_1031[4], ret_V_4_reg_1031[4], ret_V_4_reg_1031[4], ret_V_4_reg_1031[4], ret_V_4_reg_1031[4], ret_V_4_reg_1031[4], ret_V_4_reg_1031[4], ret_V_4_reg_1031[4], ret_V_4_reg_1031[4], ret_V_4_reg_1031[4], ret_V_4_reg_1031[4], ret_V_4_reg_1031[4], ret_V_4_reg_1031[4], ret_V_4_reg_1031[4], ret_V_4_reg_1031[4], ret_V_4_reg_1031[4], ret_V_4_reg_1031[4], ret_V_4_reg_1031[4], ret_V_4_reg_1031[4], ret_V_4_reg_1031[4], ret_V_4_reg_1031[4], ret_V_4_reg_1031[4], ret_V_4_reg_1031[4], ret_V_4_reg_1031[4], ret_V_4_reg_1031, 1'h0 };
assign grp_fu_663_p0 = { tmp_5_reg_1083[31], tmp_5_reg_1083, 3'h0 };
assign grp_fu_663_p1 = { op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12 };
assign grp_fu_717_p1 = { op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13 };
assign grp_fu_725_p0 = { 30'h00000000, ret_reg_980 };
assign grp_fu_750_p0 = { op_27_V_reg_1150[31], op_27_V_reg_1150, 10'h000 };
assign grp_fu_750_p1 = { op_16[31], op_16[31], op_16[31], op_16[31], op_16[31], op_16[31], op_16[31], op_16[31], op_16[31], op_16[31], op_16[31], op_16 };
assign grp_fu_822_p0 = { select_ln353_reg_1187, 1'h0 };
assign grp_fu_822_p1 = { 30'h00000000, r_1_reg_931, r_1_reg_931, 1'h0 };
assign grp_fu_842_p1 = { op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18 };
assign newsignbit_fu_235_p1 = op_1[0];
assign op_11_V_fu_610_p3 = { ret_V_4_reg_1031, 1'h0 };
assign op_17_V_fu_807_p1 = { r_1_reg_931, r_1_reg_931, 1'h0 };
assign op_31 = grp_fu_847_p2;
assign p_Result_5_fu_582_p3 = ret_V_16_reg_1036[13];
assign p_Result_6_fu_694_p3 = ret_V_18_reg_1103[35];
assign p_Result_7_fu_781_p3 = ret_V_21_reg_1170[42];
assign p_Result_s_18_fu_470_p3 = ret_V_14_reg_914[8];
assign p_Result_s_fu_239_p4 = op_1[3:1];
assign p_Val2_3_fu_432_p3 = { trunc_ln728_reg_943, 7'h00 };
assign rhs_1_fu_541_p3 = { select_ln850_3_reg_1006, 7'h00 };
assign rhs_3_fu_652_p3 = { tmp_5_reg_1083, 3'h0 };
assign rhs_6_fu_739_p3 = { op_27_V_reg_1150, 10'h000 };
assign select_ln1192_fu_316_p0 = op_6;
assign sext_ln703_1_fu_648_p0 = op_12;
assign sext_ln703_2_fu_735_p0 = op_16;
assign sext_ln850_fu_573_p1 = { tmp_reg_1041[6], tmp_reg_1041 };
assign shl_ln1497_fu_261_p2 = { op_1[2:0], 1'h0 };
assign tmp_4_fu_800_p3 = { r_1_reg_931, 1'h0 };
assign tmp_6_fu_621_p3 = { op_22_V_reg_1068, 1'h0 };
assign trunc_ln1497_fu_412_p1 = r_reg_879[1:0];
assign trunc_ln728_fu_398_p1 = ret_V_15_fu_391_p3[0];
assign trunc_ln851_1_fu_530_p1 = op_9_V_fu_504_p3[6:0];
assign trunc_ln851_2_fu_669_p0 = op_12;
assign trunc_ln851_2_fu_669_p1 = op_12[2:0];
assign trunc_ln851_3_fu_756_p0 = op_16;
assign trunc_ln851_3_fu_756_p1 = op_16[9:0];
assign trunc_ln851_fu_379_p1 = grp_fu_364_p2[2:0];
assign zext_ln703_fu_388_p1 = { 1'h0, r_reg_879 };
assign \sub_5ns_5ns_5_2_1_U3.top_sub_5ns_5ns_5_2_1_Adder_2_U.ain_s0  = \sub_5ns_5ns_5_2_1_U3.top_sub_5ns_5ns_5_2_1_Adder_2_U.a ;
assign \sub_5ns_5ns_5_2_1_U3.top_sub_5ns_5ns_5_2_1_Adder_2_U.s  = { \sub_5ns_5ns_5_2_1_U3.top_sub_5ns_5ns_5_2_1_Adder_2_U.fas_s2 , \sub_5ns_5ns_5_2_1_U3.top_sub_5ns_5ns_5_2_1_Adder_2_U.sum_s1  };
assign \sub_5ns_5ns_5_2_1_U3.top_sub_5ns_5ns_5_2_1_Adder_2_U.u2.a  = \sub_5ns_5ns_5_2_1_U3.top_sub_5ns_5ns_5_2_1_Adder_2_U.ain_s1 ;
assign \sub_5ns_5ns_5_2_1_U3.top_sub_5ns_5ns_5_2_1_Adder_2_U.u2.b  = \sub_5ns_5ns_5_2_1_U3.top_sub_5ns_5ns_5_2_1_Adder_2_U.bin_s1 ;
assign \sub_5ns_5ns_5_2_1_U3.top_sub_5ns_5ns_5_2_1_Adder_2_U.u2.cin  = \sub_5ns_5ns_5_2_1_U3.top_sub_5ns_5ns_5_2_1_Adder_2_U.carry_s1 ;
assign \sub_5ns_5ns_5_2_1_U3.top_sub_5ns_5ns_5_2_1_Adder_2_U.facout_s2  = \sub_5ns_5ns_5_2_1_U3.top_sub_5ns_5ns_5_2_1_Adder_2_U.u2.cout ;
assign \sub_5ns_5ns_5_2_1_U3.top_sub_5ns_5ns_5_2_1_Adder_2_U.fas_s2  = \sub_5ns_5ns_5_2_1_U3.top_sub_5ns_5ns_5_2_1_Adder_2_U.u2.s ;
assign \sub_5ns_5ns_5_2_1_U3.top_sub_5ns_5ns_5_2_1_Adder_2_U.u1.a  = \sub_5ns_5ns_5_2_1_U3.top_sub_5ns_5ns_5_2_1_Adder_2_U.a [1:0];
assign \sub_5ns_5ns_5_2_1_U3.top_sub_5ns_5ns_5_2_1_Adder_2_U.u1.b  = \sub_5ns_5ns_5_2_1_U3.top_sub_5ns_5ns_5_2_1_Adder_2_U.bin_s0 [1:0];
assign \sub_5ns_5ns_5_2_1_U3.top_sub_5ns_5ns_5_2_1_Adder_2_U.u1.cin  = 1'h1;
assign \sub_5ns_5ns_5_2_1_U3.top_sub_5ns_5ns_5_2_1_Adder_2_U.facout_s1  = \sub_5ns_5ns_5_2_1_U3.top_sub_5ns_5ns_5_2_1_Adder_2_U.u1.cout ;
assign \sub_5ns_5ns_5_2_1_U3.top_sub_5ns_5ns_5_2_1_Adder_2_U.fas_s1  = \sub_5ns_5ns_5_2_1_U3.top_sub_5ns_5ns_5_2_1_Adder_2_U.u1.s ;
assign \sub_5ns_5ns_5_2_1_U3.top_sub_5ns_5ns_5_2_1_Adder_2_U.a  = \sub_5ns_5ns_5_2_1_U3.din0 ;
assign \sub_5ns_5ns_5_2_1_U3.top_sub_5ns_5ns_5_2_1_Adder_2_U.b  = \sub_5ns_5ns_5_2_1_U3.din1 ;
assign \sub_5ns_5ns_5_2_1_U3.top_sub_5ns_5ns_5_2_1_Adder_2_U.ce  = \sub_5ns_5ns_5_2_1_U3.ce ;
assign \sub_5ns_5ns_5_2_1_U3.top_sub_5ns_5ns_5_2_1_Adder_2_U.clk  = \sub_5ns_5ns_5_2_1_U3.clk ;
assign \sub_5ns_5ns_5_2_1_U3.top_sub_5ns_5ns_5_2_1_Adder_2_U.reset  = \sub_5ns_5ns_5_2_1_U3.reset ;
assign \sub_5ns_5ns_5_2_1_U3.dout  = \sub_5ns_5ns_5_2_1_U3.top_sub_5ns_5ns_5_2_1_Adder_2_U.s ;
assign \sub_5ns_5ns_5_2_1_U3.ce  = 1'h1;
assign \sub_5ns_5ns_5_2_1_U3.clk  = ap_clk;
assign \sub_5ns_5ns_5_2_1_U3.din0  = select_ln1193_reg_1001;
assign \sub_5ns_5ns_5_2_1_U3.din1  = zext_ln703_reg_938;
assign grp_fu_534_p2 = \sub_5ns_5ns_5_2_1_U3.dout ;
assign \sub_5ns_5ns_5_2_1_U3.reset  = ap_rst;
assign \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.ain_s0  = \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.a ;
assign \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.bin_s0  = \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.b ;
assign \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.s  = { \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.fas_s2 , \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.sum_s1  };
assign \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.u2.a  = \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.ain_s1 ;
assign \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.u2.b  = \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.bin_s1 ;
assign \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.u2.cin  = \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.carry_s1 ;
assign \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.facout_s2  = \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.u2.cout ;
assign \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.fas_s2  = \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.u2.s ;
assign \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.u1.a  = \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.a [3:0];
assign \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.u1.b  = \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.b [3:0];
assign \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.u1.cin  = 1'h0;
assign \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.facout_s1  = \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.u1.cout ;
assign \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.fas_s1  = \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.u1.s ;
assign \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.a  = \add_9ns_9s_9_2_1_U1.din0 ;
assign \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.b  = \add_9ns_9s_9_2_1_U1.din1 ;
assign \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.ce  = \add_9ns_9s_9_2_1_U1.ce ;
assign \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.clk  = \add_9ns_9s_9_2_1_U1.clk ;
assign \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.reset  = \add_9ns_9s_9_2_1_U1.reset ;
assign \add_9ns_9s_9_2_1_U1.dout  = \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.s ;
assign \add_9ns_9s_9_2_1_U1.ce  = 1'h1;
assign \add_9ns_9s_9_2_1_U1.clk  = ap_clk;
assign \add_9ns_9s_9_2_1_U1.din0  = select_ln1192_reg_896;
assign \add_9ns_9s_9_2_1_U1.din1  = { op_0[7], op_0 };
assign grp_fu_364_p2 = \add_9ns_9s_9_2_1_U1.dout ;
assign \add_9ns_9s_9_2_1_U1.reset  = ap_rst;
assign \add_8s_8ns_8_2_1_U5.top_add_8s_8ns_8_2_1_Adder_4_U.ain_s0  = \add_8s_8ns_8_2_1_U5.top_add_8s_8ns_8_2_1_Adder_4_U.a ;
assign \add_8s_8ns_8_2_1_U5.top_add_8s_8ns_8_2_1_Adder_4_U.bin_s0  = \add_8s_8ns_8_2_1_U5.top_add_8s_8ns_8_2_1_Adder_4_U.b ;
assign \add_8s_8ns_8_2_1_U5.top_add_8s_8ns_8_2_1_Adder_4_U.s  = { \add_8s_8ns_8_2_1_U5.top_add_8s_8ns_8_2_1_Adder_4_U.fas_s2 , \add_8s_8ns_8_2_1_U5.top_add_8s_8ns_8_2_1_Adder_4_U.sum_s1  };
assign \add_8s_8ns_8_2_1_U5.top_add_8s_8ns_8_2_1_Adder_4_U.u2.a  = \add_8s_8ns_8_2_1_U5.top_add_8s_8ns_8_2_1_Adder_4_U.ain_s1 ;
assign \add_8s_8ns_8_2_1_U5.top_add_8s_8ns_8_2_1_Adder_4_U.u2.b  = \add_8s_8ns_8_2_1_U5.top_add_8s_8ns_8_2_1_Adder_4_U.bin_s1 ;
assign \add_8s_8ns_8_2_1_U5.top_add_8s_8ns_8_2_1_Adder_4_U.u2.cin  = \add_8s_8ns_8_2_1_U5.top_add_8s_8ns_8_2_1_Adder_4_U.carry_s1 ;
assign \add_8s_8ns_8_2_1_U5.top_add_8s_8ns_8_2_1_Adder_4_U.facout_s2  = \add_8s_8ns_8_2_1_U5.top_add_8s_8ns_8_2_1_Adder_4_U.u2.cout ;
assign \add_8s_8ns_8_2_1_U5.top_add_8s_8ns_8_2_1_Adder_4_U.fas_s2  = \add_8s_8ns_8_2_1_U5.top_add_8s_8ns_8_2_1_Adder_4_U.u2.s ;
assign \add_8s_8ns_8_2_1_U5.top_add_8s_8ns_8_2_1_Adder_4_U.u1.a  = \add_8s_8ns_8_2_1_U5.top_add_8s_8ns_8_2_1_Adder_4_U.a [3:0];
assign \add_8s_8ns_8_2_1_U5.top_add_8s_8ns_8_2_1_Adder_4_U.u1.b  = \add_8s_8ns_8_2_1_U5.top_add_8s_8ns_8_2_1_Adder_4_U.b [3:0];
assign \add_8s_8ns_8_2_1_U5.top_add_8s_8ns_8_2_1_Adder_4_U.u1.cin  = 1'h0;
assign \add_8s_8ns_8_2_1_U5.top_add_8s_8ns_8_2_1_Adder_4_U.facout_s1  = \add_8s_8ns_8_2_1_U5.top_add_8s_8ns_8_2_1_Adder_4_U.u1.cout ;
assign \add_8s_8ns_8_2_1_U5.top_add_8s_8ns_8_2_1_Adder_4_U.fas_s1  = \add_8s_8ns_8_2_1_U5.top_add_8s_8ns_8_2_1_Adder_4_U.u1.s ;
assign \add_8s_8ns_8_2_1_U5.top_add_8s_8ns_8_2_1_Adder_4_U.a  = \add_8s_8ns_8_2_1_U5.din0 ;
assign \add_8s_8ns_8_2_1_U5.top_add_8s_8ns_8_2_1_Adder_4_U.b  = \add_8s_8ns_8_2_1_U5.din1 ;
assign \add_8s_8ns_8_2_1_U5.top_add_8s_8ns_8_2_1_Adder_4_U.ce  = \add_8s_8ns_8_2_1_U5.ce ;
assign \add_8s_8ns_8_2_1_U5.top_add_8s_8ns_8_2_1_Adder_4_U.clk  = \add_8s_8ns_8_2_1_U5.clk ;
assign \add_8s_8ns_8_2_1_U5.top_add_8s_8ns_8_2_1_Adder_4_U.reset  = \add_8s_8ns_8_2_1_U5.reset ;
assign \add_8s_8ns_8_2_1_U5.dout  = \add_8s_8ns_8_2_1_U5.top_add_8s_8ns_8_2_1_Adder_4_U.s ;
assign \add_8s_8ns_8_2_1_U5.ce  = 1'h1;
assign \add_8s_8ns_8_2_1_U5.clk  = ap_clk;
assign \add_8s_8ns_8_2_1_U5.din0  = { tmp_reg_1041[6], tmp_reg_1041 };
assign \add_8s_8ns_8_2_1_U5.din1  = 8'h01;
assign grp_fu_576_p2 = \add_8s_8ns_8_2_1_U5.dout ;
assign \add_8s_8ns_8_2_1_U5.reset  = ap_rst;
assign \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.ain_s0  = \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.a ;
assign \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.bin_s0  = \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.b ;
assign \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.s  = { \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.fas_s2 , \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.sum_s1  };
assign \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.u2.a  = \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.ain_s1 ;
assign \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.u2.b  = \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.bin_s1 ;
assign \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.u2.cin  = \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.carry_s1 ;
assign \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.facout_s2  = \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.u2.cout ;
assign \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.fas_s2  = \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.u2.s ;
assign \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.u1.a  = \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.a [3:0];
assign \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.u1.b  = \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.b [3:0];
assign \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.u1.cin  = 1'h0;
assign \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.facout_s1  = \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.u1.cout ;
assign \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.fas_s1  = \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.u1.s ;
assign \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.a  = \add_8ns_8ns_8_2_1_U6.din0 ;
assign \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.b  = \add_8ns_8ns_8_2_1_U6.din1 ;
assign \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.ce  = \add_8ns_8ns_8_2_1_U6.ce ;
assign \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.clk  = \add_8ns_8ns_8_2_1_U6.clk ;
assign \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.reset  = \add_8ns_8ns_8_2_1_U6.reset ;
assign \add_8ns_8ns_8_2_1_U6.dout  = \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.s ;
assign \add_8ns_8ns_8_2_1_U6.ce  = 1'h1;
assign \add_8ns_8ns_8_2_1_U6.clk  = ap_clk;
assign \add_8ns_8ns_8_2_1_U6.din0  = ret_V_17_reg_1058;
assign \add_8ns_8ns_8_2_1_U6.din1  = { 6'h00, op_10 };
assign grp_fu_605_p2 = \add_8ns_8ns_8_2_1_U6.dout ;
assign \add_8ns_8ns_8_2_1_U6.reset  = ap_rst;
assign \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.ain_s0  = \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.a ;
assign \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.bin_s0  = \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.b ;
assign \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.s  = { \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.fas_s2 , \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.sum_s1  };
assign \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.u2.a  = \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.ain_s1 ;
assign \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.u2.b  = \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.bin_s1 ;
assign \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.u2.cin  = \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.carry_s1 ;
assign \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.facout_s2  = \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.u2.cout ;
assign \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.fas_s2  = \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.u2.s ;
assign \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.u1.a  = \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.a [2:0];
assign \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.u1.b  = \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.b [2:0];
assign \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.u1.cin  = 1'h0;
assign \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.facout_s1  = \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.u1.cout ;
assign \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.fas_s1  = \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.u1.s ;
assign \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.a  = \add_6ns_6ns_6_2_1_U2.din0 ;
assign \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.b  = \add_6ns_6ns_6_2_1_U2.din1 ;
assign \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.ce  = \add_6ns_6ns_6_2_1_U2.ce ;
assign \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.clk  = \add_6ns_6ns_6_2_1_U2.clk ;
assign \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.reset  = \add_6ns_6ns_6_2_1_U2.reset ;
assign \add_6ns_6ns_6_2_1_U2.dout  = \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.s ;
assign \add_6ns_6ns_6_2_1_U2.ce  = 1'h1;
assign \add_6ns_6ns_6_2_1_U2.clk  = ap_clk;
assign \add_6ns_6ns_6_2_1_U2.din0  = ret_V_reg_919;
assign \add_6ns_6ns_6_2_1_U2.din1  = 6'h01;
assign grp_fu_420_p2 = \add_6ns_6ns_6_2_1_U2.dout ;
assign \add_6ns_6ns_6_2_1_U2.reset  = ap_rst;
assign \add_43s_43s_43_2_1_U13.top_add_43s_43s_43_2_1_Adder_10_U.ain_s0  = \add_43s_43s_43_2_1_U13.top_add_43s_43s_43_2_1_Adder_10_U.a ;
assign \add_43s_43s_43_2_1_U13.top_add_43s_43s_43_2_1_Adder_10_U.bin_s0  = \add_43s_43s_43_2_1_U13.top_add_43s_43s_43_2_1_Adder_10_U.b ;
assign \add_43s_43s_43_2_1_U13.top_add_43s_43s_43_2_1_Adder_10_U.s  = { \add_43s_43s_43_2_1_U13.top_add_43s_43s_43_2_1_Adder_10_U.fas_s2 , \add_43s_43s_43_2_1_U13.top_add_43s_43s_43_2_1_Adder_10_U.sum_s1  };
assign \add_43s_43s_43_2_1_U13.top_add_43s_43s_43_2_1_Adder_10_U.u2.a  = \add_43s_43s_43_2_1_U13.top_add_43s_43s_43_2_1_Adder_10_U.ain_s1 ;
assign \add_43s_43s_43_2_1_U13.top_add_43s_43s_43_2_1_Adder_10_U.u2.b  = \add_43s_43s_43_2_1_U13.top_add_43s_43s_43_2_1_Adder_10_U.bin_s1 ;
assign \add_43s_43s_43_2_1_U13.top_add_43s_43s_43_2_1_Adder_10_U.u2.cin  = \add_43s_43s_43_2_1_U13.top_add_43s_43s_43_2_1_Adder_10_U.carry_s1 ;
assign \add_43s_43s_43_2_1_U13.top_add_43s_43s_43_2_1_Adder_10_U.facout_s2  = \add_43s_43s_43_2_1_U13.top_add_43s_43s_43_2_1_Adder_10_U.u2.cout ;
assign \add_43s_43s_43_2_1_U13.top_add_43s_43s_43_2_1_Adder_10_U.fas_s2  = \add_43s_43s_43_2_1_U13.top_add_43s_43s_43_2_1_Adder_10_U.u2.s ;
assign \add_43s_43s_43_2_1_U13.top_add_43s_43s_43_2_1_Adder_10_U.u1.a  = \add_43s_43s_43_2_1_U13.top_add_43s_43s_43_2_1_Adder_10_U.a [20:0];
assign \add_43s_43s_43_2_1_U13.top_add_43s_43s_43_2_1_Adder_10_U.u1.b  = \add_43s_43s_43_2_1_U13.top_add_43s_43s_43_2_1_Adder_10_U.b [20:0];
assign \add_43s_43s_43_2_1_U13.top_add_43s_43s_43_2_1_Adder_10_U.u1.cin  = 1'h0;
assign \add_43s_43s_43_2_1_U13.top_add_43s_43s_43_2_1_Adder_10_U.facout_s1  = \add_43s_43s_43_2_1_U13.top_add_43s_43s_43_2_1_Adder_10_U.u1.cout ;
assign \add_43s_43s_43_2_1_U13.top_add_43s_43s_43_2_1_Adder_10_U.fas_s1  = \add_43s_43s_43_2_1_U13.top_add_43s_43s_43_2_1_Adder_10_U.u1.s ;
assign \add_43s_43s_43_2_1_U13.top_add_43s_43s_43_2_1_Adder_10_U.a  = \add_43s_43s_43_2_1_U13.din0 ;
assign \add_43s_43s_43_2_1_U13.top_add_43s_43s_43_2_1_Adder_10_U.b  = \add_43s_43s_43_2_1_U13.din1 ;
assign \add_43s_43s_43_2_1_U13.top_add_43s_43s_43_2_1_Adder_10_U.ce  = \add_43s_43s_43_2_1_U13.ce ;
assign \add_43s_43s_43_2_1_U13.top_add_43s_43s_43_2_1_Adder_10_U.clk  = \add_43s_43s_43_2_1_U13.clk ;
assign \add_43s_43s_43_2_1_U13.top_add_43s_43s_43_2_1_Adder_10_U.reset  = \add_43s_43s_43_2_1_U13.reset ;
assign \add_43s_43s_43_2_1_U13.dout  = \add_43s_43s_43_2_1_U13.top_add_43s_43s_43_2_1_Adder_10_U.s ;
assign \add_43s_43s_43_2_1_U13.ce  = 1'h1;
assign \add_43s_43s_43_2_1_U13.clk  = ap_clk;
assign \add_43s_43s_43_2_1_U13.din0  = { op_27_V_reg_1150[31], op_27_V_reg_1150, 10'h000 };
assign \add_43s_43s_43_2_1_U13.din1  = { op_16[31], op_16[31], op_16[31], op_16[31], op_16[31], op_16[31], op_16[31], op_16[31], op_16[31], op_16[31], op_16[31], op_16 };
assign grp_fu_750_p2 = \add_43s_43s_43_2_1_U13.dout ;
assign \add_43s_43s_43_2_1_U13.reset  = ap_rst;
assign \add_36s_36s_36_2_1_U8.top_add_36s_36s_36_2_1_Adder_7_U.ain_s0  = \add_36s_36s_36_2_1_U8.top_add_36s_36s_36_2_1_Adder_7_U.a ;
assign \add_36s_36s_36_2_1_U8.top_add_36s_36s_36_2_1_Adder_7_U.bin_s0  = \add_36s_36s_36_2_1_U8.top_add_36s_36s_36_2_1_Adder_7_U.b ;
assign \add_36s_36s_36_2_1_U8.top_add_36s_36s_36_2_1_Adder_7_U.s  = { \add_36s_36s_36_2_1_U8.top_add_36s_36s_36_2_1_Adder_7_U.fas_s2 , \add_36s_36s_36_2_1_U8.top_add_36s_36s_36_2_1_Adder_7_U.sum_s1  };
assign \add_36s_36s_36_2_1_U8.top_add_36s_36s_36_2_1_Adder_7_U.u2.a  = \add_36s_36s_36_2_1_U8.top_add_36s_36s_36_2_1_Adder_7_U.ain_s1 ;
assign \add_36s_36s_36_2_1_U8.top_add_36s_36s_36_2_1_Adder_7_U.u2.b  = \add_36s_36s_36_2_1_U8.top_add_36s_36s_36_2_1_Adder_7_U.bin_s1 ;
assign \add_36s_36s_36_2_1_U8.top_add_36s_36s_36_2_1_Adder_7_U.u2.cin  = \add_36s_36s_36_2_1_U8.top_add_36s_36s_36_2_1_Adder_7_U.carry_s1 ;
assign \add_36s_36s_36_2_1_U8.top_add_36s_36s_36_2_1_Adder_7_U.facout_s2  = \add_36s_36s_36_2_1_U8.top_add_36s_36s_36_2_1_Adder_7_U.u2.cout ;
assign \add_36s_36s_36_2_1_U8.top_add_36s_36s_36_2_1_Adder_7_U.fas_s2  = \add_36s_36s_36_2_1_U8.top_add_36s_36s_36_2_1_Adder_7_U.u2.s ;
assign \add_36s_36s_36_2_1_U8.top_add_36s_36s_36_2_1_Adder_7_U.u1.a  = \add_36s_36s_36_2_1_U8.top_add_36s_36s_36_2_1_Adder_7_U.a [17:0];
assign \add_36s_36s_36_2_1_U8.top_add_36s_36s_36_2_1_Adder_7_U.u1.b  = \add_36s_36s_36_2_1_U8.top_add_36s_36s_36_2_1_Adder_7_U.b [17:0];
assign \add_36s_36s_36_2_1_U8.top_add_36s_36s_36_2_1_Adder_7_U.u1.cin  = 1'h0;
assign \add_36s_36s_36_2_1_U8.top_add_36s_36s_36_2_1_Adder_7_U.facout_s1  = \add_36s_36s_36_2_1_U8.top_add_36s_36s_36_2_1_Adder_7_U.u1.cout ;
assign \add_36s_36s_36_2_1_U8.top_add_36s_36s_36_2_1_Adder_7_U.fas_s1  = \add_36s_36s_36_2_1_U8.top_add_36s_36s_36_2_1_Adder_7_U.u1.s ;
assign \add_36s_36s_36_2_1_U8.top_add_36s_36s_36_2_1_Adder_7_U.a  = \add_36s_36s_36_2_1_U8.din0 ;
assign \add_36s_36s_36_2_1_U8.top_add_36s_36s_36_2_1_Adder_7_U.b  = \add_36s_36s_36_2_1_U8.din1 ;
assign \add_36s_36s_36_2_1_U8.top_add_36s_36s_36_2_1_Adder_7_U.ce  = \add_36s_36s_36_2_1_U8.ce ;
assign \add_36s_36s_36_2_1_U8.top_add_36s_36s_36_2_1_Adder_7_U.clk  = \add_36s_36s_36_2_1_U8.clk ;
assign \add_36s_36s_36_2_1_U8.top_add_36s_36s_36_2_1_Adder_7_U.reset  = \add_36s_36s_36_2_1_U8.reset ;
assign \add_36s_36s_36_2_1_U8.dout  = \add_36s_36s_36_2_1_U8.top_add_36s_36s_36_2_1_Adder_7_U.s ;
assign \add_36s_36s_36_2_1_U8.ce  = 1'h1;
assign \add_36s_36s_36_2_1_U8.clk  = ap_clk;
assign \add_36s_36s_36_2_1_U8.din0  = { tmp_5_reg_1083[31], tmp_5_reg_1083, 3'h0 };
assign \add_36s_36s_36_2_1_U8.din1  = { op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12 };
assign grp_fu_663_p2 = \add_36s_36s_36_2_1_U8.dout ;
assign \add_36s_36s_36_2_1_U8.reset  = ap_rst;
assign \add_33s_33s_33_2_1_U7.top_add_33s_33s_33_2_1_Adder_6_U.ain_s0  = \add_33s_33s_33_2_1_U7.top_add_33s_33s_33_2_1_Adder_6_U.a ;
assign \add_33s_33s_33_2_1_U7.top_add_33s_33s_33_2_1_Adder_6_U.bin_s0  = \add_33s_33s_33_2_1_U7.top_add_33s_33s_33_2_1_Adder_6_U.b ;
assign \add_33s_33s_33_2_1_U7.top_add_33s_33s_33_2_1_Adder_6_U.s  = { \add_33s_33s_33_2_1_U7.top_add_33s_33s_33_2_1_Adder_6_U.fas_s2 , \add_33s_33s_33_2_1_U7.top_add_33s_33s_33_2_1_Adder_6_U.sum_s1  };
assign \add_33s_33s_33_2_1_U7.top_add_33s_33s_33_2_1_Adder_6_U.u2.a  = \add_33s_33s_33_2_1_U7.top_add_33s_33s_33_2_1_Adder_6_U.ain_s1 ;
assign \add_33s_33s_33_2_1_U7.top_add_33s_33s_33_2_1_Adder_6_U.u2.b  = \add_33s_33s_33_2_1_U7.top_add_33s_33s_33_2_1_Adder_6_U.bin_s1 ;
assign \add_33s_33s_33_2_1_U7.top_add_33s_33s_33_2_1_Adder_6_U.u2.cin  = \add_33s_33s_33_2_1_U7.top_add_33s_33s_33_2_1_Adder_6_U.carry_s1 ;
assign \add_33s_33s_33_2_1_U7.top_add_33s_33s_33_2_1_Adder_6_U.facout_s2  = \add_33s_33s_33_2_1_U7.top_add_33s_33s_33_2_1_Adder_6_U.u2.cout ;
assign \add_33s_33s_33_2_1_U7.top_add_33s_33s_33_2_1_Adder_6_U.fas_s2  = \add_33s_33s_33_2_1_U7.top_add_33s_33s_33_2_1_Adder_6_U.u2.s ;
assign \add_33s_33s_33_2_1_U7.top_add_33s_33s_33_2_1_Adder_6_U.u1.a  = \add_33s_33s_33_2_1_U7.top_add_33s_33s_33_2_1_Adder_6_U.a [15:0];
assign \add_33s_33s_33_2_1_U7.top_add_33s_33s_33_2_1_Adder_6_U.u1.b  = \add_33s_33s_33_2_1_U7.top_add_33s_33s_33_2_1_Adder_6_U.b [15:0];
assign \add_33s_33s_33_2_1_U7.top_add_33s_33s_33_2_1_Adder_6_U.u1.cin  = 1'h0;
assign \add_33s_33s_33_2_1_U7.top_add_33s_33s_33_2_1_Adder_6_U.facout_s1  = \add_33s_33s_33_2_1_U7.top_add_33s_33s_33_2_1_Adder_6_U.u1.cout ;
assign \add_33s_33s_33_2_1_U7.top_add_33s_33s_33_2_1_Adder_6_U.fas_s1  = \add_33s_33s_33_2_1_U7.top_add_33s_33s_33_2_1_Adder_6_U.u1.s ;
assign \add_33s_33s_33_2_1_U7.top_add_33s_33s_33_2_1_Adder_6_U.a  = \add_33s_33s_33_2_1_U7.din0 ;
assign \add_33s_33s_33_2_1_U7.top_add_33s_33s_33_2_1_Adder_6_U.b  = \add_33s_33s_33_2_1_U7.din1 ;
assign \add_33s_33s_33_2_1_U7.top_add_33s_33s_33_2_1_Adder_6_U.ce  = \add_33s_33s_33_2_1_U7.ce ;
assign \add_33s_33s_33_2_1_U7.top_add_33s_33s_33_2_1_Adder_6_U.clk  = \add_33s_33s_33_2_1_U7.clk ;
assign \add_33s_33s_33_2_1_U7.top_add_33s_33s_33_2_1_Adder_6_U.reset  = \add_33s_33s_33_2_1_U7.reset ;
assign \add_33s_33s_33_2_1_U7.dout  = \add_33s_33s_33_2_1_U7.top_add_33s_33s_33_2_1_Adder_6_U.s ;
assign \add_33s_33s_33_2_1_U7.ce  = 1'h1;
assign \add_33s_33s_33_2_1_U7.clk  = ap_clk;
assign \add_33s_33s_33_2_1_U7.din0  = { op_22_V_reg_1068[7], op_22_V_reg_1068[7], op_22_V_reg_1068[7], op_22_V_reg_1068[7], op_22_V_reg_1068[7], op_22_V_reg_1068[7], op_22_V_reg_1068[7], op_22_V_reg_1068[7], op_22_V_reg_1068[7], op_22_V_reg_1068[7], op_22_V_reg_1068[7], op_22_V_reg_1068[7], op_22_V_reg_1068[7], op_22_V_reg_1068[7], op_22_V_reg_1068[7], op_22_V_reg_1068[7], op_22_V_reg_1068[7], op_22_V_reg_1068[7], op_22_V_reg_1068[7], op_22_V_reg_1068[7], op_22_V_reg_1068[7], op_22_V_reg_1068[7], op_22_V_reg_1068[7], op_22_V_reg_1068[7], op_22_V_reg_1068, 1'h0 };
assign \add_33s_33s_33_2_1_U7.din1  = { ret_V_4_reg_1031[4], ret_V_4_reg_1031[4], ret_V_4_reg_1031[4], ret_V_4_reg_1031[4], ret_V_4_reg_1031[4], ret_V_4_reg_1031[4], ret_V_4_reg_1031[4], ret_V_4_reg_1031[4], ret_V_4_reg_1031[4], ret_V_4_reg_1031[4], ret_V_4_reg_1031[4], ret_V_4_reg_1031[4], ret_V_4_reg_1031[4], ret_V_4_reg_1031[4], ret_V_4_reg_1031[4], ret_V_4_reg_1031[4], ret_V_4_reg_1031[4], ret_V_4_reg_1031[4], ret_V_4_reg_1031[4], ret_V_4_reg_1031[4], ret_V_4_reg_1031[4], ret_V_4_reg_1031[4], ret_V_4_reg_1031[4], ret_V_4_reg_1031[4], ret_V_4_reg_1031[4], ret_V_4_reg_1031[4], ret_V_4_reg_1031[4], ret_V_4_reg_1031, 1'h0 };
assign grp_fu_632_p2 = \add_33s_33s_33_2_1_U7.dout ;
assign \add_33s_33s_33_2_1_U7.reset  = ap_rst;
assign \add_33ns_33ns_33_2_1_U15.top_add_33ns_33ns_33_2_1_Adder_11_U.ain_s0  = \add_33ns_33ns_33_2_1_U15.top_add_33ns_33ns_33_2_1_Adder_11_U.a ;
assign \add_33ns_33ns_33_2_1_U15.top_add_33ns_33ns_33_2_1_Adder_11_U.bin_s0  = \add_33ns_33ns_33_2_1_U15.top_add_33ns_33ns_33_2_1_Adder_11_U.b ;
assign \add_33ns_33ns_33_2_1_U15.top_add_33ns_33ns_33_2_1_Adder_11_U.s  = { \add_33ns_33ns_33_2_1_U15.top_add_33ns_33ns_33_2_1_Adder_11_U.fas_s2 , \add_33ns_33ns_33_2_1_U15.top_add_33ns_33ns_33_2_1_Adder_11_U.sum_s1  };
assign \add_33ns_33ns_33_2_1_U15.top_add_33ns_33ns_33_2_1_Adder_11_U.u2.a  = \add_33ns_33ns_33_2_1_U15.top_add_33ns_33ns_33_2_1_Adder_11_U.ain_s1 ;
assign \add_33ns_33ns_33_2_1_U15.top_add_33ns_33ns_33_2_1_Adder_11_U.u2.b  = \add_33ns_33ns_33_2_1_U15.top_add_33ns_33ns_33_2_1_Adder_11_U.bin_s1 ;
assign \add_33ns_33ns_33_2_1_U15.top_add_33ns_33ns_33_2_1_Adder_11_U.u2.cin  = \add_33ns_33ns_33_2_1_U15.top_add_33ns_33ns_33_2_1_Adder_11_U.carry_s1 ;
assign \add_33ns_33ns_33_2_1_U15.top_add_33ns_33ns_33_2_1_Adder_11_U.facout_s2  = \add_33ns_33ns_33_2_1_U15.top_add_33ns_33ns_33_2_1_Adder_11_U.u2.cout ;
assign \add_33ns_33ns_33_2_1_U15.top_add_33ns_33ns_33_2_1_Adder_11_U.fas_s2  = \add_33ns_33ns_33_2_1_U15.top_add_33ns_33ns_33_2_1_Adder_11_U.u2.s ;
assign \add_33ns_33ns_33_2_1_U15.top_add_33ns_33ns_33_2_1_Adder_11_U.u1.a  = \add_33ns_33ns_33_2_1_U15.top_add_33ns_33ns_33_2_1_Adder_11_U.a [15:0];
assign \add_33ns_33ns_33_2_1_U15.top_add_33ns_33ns_33_2_1_Adder_11_U.u1.b  = \add_33ns_33ns_33_2_1_U15.top_add_33ns_33ns_33_2_1_Adder_11_U.b [15:0];
assign \add_33ns_33ns_33_2_1_U15.top_add_33ns_33ns_33_2_1_Adder_11_U.u1.cin  = 1'h0;
assign \add_33ns_33ns_33_2_1_U15.top_add_33ns_33ns_33_2_1_Adder_11_U.facout_s1  = \add_33ns_33ns_33_2_1_U15.top_add_33ns_33ns_33_2_1_Adder_11_U.u1.cout ;
assign \add_33ns_33ns_33_2_1_U15.top_add_33ns_33ns_33_2_1_Adder_11_U.fas_s1  = \add_33ns_33ns_33_2_1_U15.top_add_33ns_33ns_33_2_1_Adder_11_U.u1.s ;
assign \add_33ns_33ns_33_2_1_U15.top_add_33ns_33ns_33_2_1_Adder_11_U.a  = \add_33ns_33ns_33_2_1_U15.din0 ;
assign \add_33ns_33ns_33_2_1_U15.top_add_33ns_33ns_33_2_1_Adder_11_U.b  = \add_33ns_33ns_33_2_1_U15.din1 ;
assign \add_33ns_33ns_33_2_1_U15.top_add_33ns_33ns_33_2_1_Adder_11_U.ce  = \add_33ns_33ns_33_2_1_U15.ce ;
assign \add_33ns_33ns_33_2_1_U15.top_add_33ns_33ns_33_2_1_Adder_11_U.clk  = \add_33ns_33ns_33_2_1_U15.clk ;
assign \add_33ns_33ns_33_2_1_U15.top_add_33ns_33ns_33_2_1_Adder_11_U.reset  = \add_33ns_33ns_33_2_1_U15.reset ;
assign \add_33ns_33ns_33_2_1_U15.dout  = \add_33ns_33ns_33_2_1_U15.top_add_33ns_33ns_33_2_1_Adder_11_U.s ;
assign \add_33ns_33ns_33_2_1_U15.ce  = 1'h1;
assign \add_33ns_33ns_33_2_1_U15.clk  = ap_clk;
assign \add_33ns_33ns_33_2_1_U15.din0  = { select_ln353_reg_1187, 1'h0 };
assign \add_33ns_33ns_33_2_1_U15.din1  = { 30'h00000000, r_1_reg_931, r_1_reg_931, 1'h0 };
assign grp_fu_822_p2 = \add_33ns_33ns_33_2_1_U15.dout ;
assign \add_33ns_33ns_33_2_1_U15.reset  = ap_rst;
assign \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.ain_s0  = \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.a ;
assign \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.bin_s0  = \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.b ;
assign \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.s  = { \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.fas_s2 , \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.sum_s1  };
assign \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.u2.a  = \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.ain_s1 ;
assign \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.u2.b  = \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.bin_s1 ;
assign \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.u2.cin  = \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.carry_s1 ;
assign \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.facout_s2  = \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.u2.cout ;
assign \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.fas_s2  = \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.u2.s ;
assign \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.u1.a  = \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.a [15:0];
assign \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.u1.b  = \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.b [15:0];
assign \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.u1.cin  = 1'h0;
assign \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.facout_s1  = \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.u1.cout ;
assign \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.fas_s1  = \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.u1.s ;
assign \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.a  = \add_32ns_32s_32_2_1_U16.din0 ;
assign \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.b  = \add_32ns_32s_32_2_1_U16.din1 ;
assign \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.ce  = \add_32ns_32s_32_2_1_U16.ce ;
assign \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.clk  = \add_32ns_32s_32_2_1_U16.clk ;
assign \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.reset  = \add_32ns_32s_32_2_1_U16.reset ;
assign \add_32ns_32s_32_2_1_U16.dout  = \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.s ;
assign \add_32ns_32s_32_2_1_U16.ce  = 1'h1;
assign \add_32ns_32s_32_2_1_U16.clk  = ap_clk;
assign \add_32ns_32s_32_2_1_U16.din0  = op_29_V_reg_1202;
assign \add_32ns_32s_32_2_1_U16.din1  = { op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18 };
assign grp_fu_842_p2 = \add_32ns_32s_32_2_1_U16.dout ;
assign \add_32ns_32s_32_2_1_U16.reset  = ap_rst;
assign \add_32ns_32s_32_2_1_U10.top_add_32ns_32s_32_2_1_Adder_9_U.ain_s0  = \add_32ns_32s_32_2_1_U10.top_add_32ns_32s_32_2_1_Adder_9_U.a ;
assign \add_32ns_32s_32_2_1_U10.top_add_32ns_32s_32_2_1_Adder_9_U.bin_s0  = \add_32ns_32s_32_2_1_U10.top_add_32ns_32s_32_2_1_Adder_9_U.b ;
assign \add_32ns_32s_32_2_1_U10.top_add_32ns_32s_32_2_1_Adder_9_U.s  = { \add_32ns_32s_32_2_1_U10.top_add_32ns_32s_32_2_1_Adder_9_U.fas_s2 , \add_32ns_32s_32_2_1_U10.top_add_32ns_32s_32_2_1_Adder_9_U.sum_s1  };
assign \add_32ns_32s_32_2_1_U10.top_add_32ns_32s_32_2_1_Adder_9_U.u2.a  = \add_32ns_32s_32_2_1_U10.top_add_32ns_32s_32_2_1_Adder_9_U.ain_s1 ;
assign \add_32ns_32s_32_2_1_U10.top_add_32ns_32s_32_2_1_Adder_9_U.u2.b  = \add_32ns_32s_32_2_1_U10.top_add_32ns_32s_32_2_1_Adder_9_U.bin_s1 ;
assign \add_32ns_32s_32_2_1_U10.top_add_32ns_32s_32_2_1_Adder_9_U.u2.cin  = \add_32ns_32s_32_2_1_U10.top_add_32ns_32s_32_2_1_Adder_9_U.carry_s1 ;
assign \add_32ns_32s_32_2_1_U10.top_add_32ns_32s_32_2_1_Adder_9_U.facout_s2  = \add_32ns_32s_32_2_1_U10.top_add_32ns_32s_32_2_1_Adder_9_U.u2.cout ;
assign \add_32ns_32s_32_2_1_U10.top_add_32ns_32s_32_2_1_Adder_9_U.fas_s2  = \add_32ns_32s_32_2_1_U10.top_add_32ns_32s_32_2_1_Adder_9_U.u2.s ;
assign \add_32ns_32s_32_2_1_U10.top_add_32ns_32s_32_2_1_Adder_9_U.u1.a  = \add_32ns_32s_32_2_1_U10.top_add_32ns_32s_32_2_1_Adder_9_U.a [15:0];
assign \add_32ns_32s_32_2_1_U10.top_add_32ns_32s_32_2_1_Adder_9_U.u1.b  = \add_32ns_32s_32_2_1_U10.top_add_32ns_32s_32_2_1_Adder_9_U.b [15:0];
assign \add_32ns_32s_32_2_1_U10.top_add_32ns_32s_32_2_1_Adder_9_U.u1.cin  = 1'h0;
assign \add_32ns_32s_32_2_1_U10.top_add_32ns_32s_32_2_1_Adder_9_U.facout_s1  = \add_32ns_32s_32_2_1_U10.top_add_32ns_32s_32_2_1_Adder_9_U.u1.cout ;
assign \add_32ns_32s_32_2_1_U10.top_add_32ns_32s_32_2_1_Adder_9_U.fas_s1  = \add_32ns_32s_32_2_1_U10.top_add_32ns_32s_32_2_1_Adder_9_U.u1.s ;
assign \add_32ns_32s_32_2_1_U10.top_add_32ns_32s_32_2_1_Adder_9_U.a  = \add_32ns_32s_32_2_1_U10.din0 ;
assign \add_32ns_32s_32_2_1_U10.top_add_32ns_32s_32_2_1_Adder_9_U.b  = \add_32ns_32s_32_2_1_U10.din1 ;
assign \add_32ns_32s_32_2_1_U10.top_add_32ns_32s_32_2_1_Adder_9_U.ce  = \add_32ns_32s_32_2_1_U10.ce ;
assign \add_32ns_32s_32_2_1_U10.top_add_32ns_32s_32_2_1_Adder_9_U.clk  = \add_32ns_32s_32_2_1_U10.clk ;
assign \add_32ns_32s_32_2_1_U10.top_add_32ns_32s_32_2_1_Adder_9_U.reset  = \add_32ns_32s_32_2_1_U10.reset ;
assign \add_32ns_32s_32_2_1_U10.dout  = \add_32ns_32s_32_2_1_U10.top_add_32ns_32s_32_2_1_Adder_9_U.s ;
assign \add_32ns_32s_32_2_1_U10.ce  = 1'h1;
assign \add_32ns_32s_32_2_1_U10.clk  = ap_clk;
assign \add_32ns_32s_32_2_1_U10.din0  = ret_V_19_reg_1120;
assign \add_32ns_32s_32_2_1_U10.din1  = { op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13 };
assign grp_fu_717_p2 = \add_32ns_32s_32_2_1_U10.dout ;
assign \add_32ns_32s_32_2_1_U10.reset  = ap_rst;
assign \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_8_U.ain_s0  = \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_8_U.a ;
assign \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_8_U.bin_s0  = \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_8_U.b ;
assign \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_8_U.s  = { \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_8_U.fas_s2 , \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_8_U.sum_s1  };
assign \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_8_U.u2.a  = \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_8_U.ain_s1 ;
assign \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_8_U.u2.b  = \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_8_U.bin_s1 ;
assign \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_8_U.u2.cin  = \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_8_U.carry_s1 ;
assign \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_8_U.facout_s2  = \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_8_U.u2.cout ;
assign \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_8_U.fas_s2  = \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_8_U.u2.s ;
assign \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_8_U.u1.a  = \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_8_U.a [15:0];
assign \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_8_U.u1.b  = \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_8_U.b [15:0];
assign \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_8_U.u1.cin  = 1'h0;
assign \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_8_U.facout_s1  = \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_8_U.u1.cout ;
assign \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_8_U.fas_s1  = \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_8_U.u1.s ;
assign \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_8_U.a  = \add_32ns_32ns_32_2_1_U9.din0 ;
assign \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_8_U.b  = \add_32ns_32ns_32_2_1_U9.din1 ;
assign \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_8_U.ce  = \add_32ns_32ns_32_2_1_U9.ce ;
assign \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_8_U.clk  = \add_32ns_32ns_32_2_1_U9.clk ;
assign \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_8_U.reset  = \add_32ns_32ns_32_2_1_U9.reset ;
assign \add_32ns_32ns_32_2_1_U9.dout  = \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_8_U.s ;
assign \add_32ns_32ns_32_2_1_U9.ce  = 1'h1;
assign \add_32ns_32ns_32_2_1_U9.clk  = ap_clk;
assign \add_32ns_32ns_32_2_1_U9.din0  = ret_V_17_cast_reg_1108;
assign \add_32ns_32ns_32_2_1_U9.din1  = 32'd1;
assign grp_fu_689_p2 = \add_32ns_32ns_32_2_1_U9.dout ;
assign \add_32ns_32ns_32_2_1_U9.reset  = ap_rst;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.ain_s0  = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.a ;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.bin_s0  = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.b ;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.s  = { \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.fas_s2 , \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.sum_s1  };
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.u2.a  = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.ain_s1 ;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.u2.b  = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.bin_s1 ;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.u2.cin  = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.carry_s1 ;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.facout_s2  = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.u2.cout ;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.fas_s2  = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.u2.s ;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.u1.a  = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.a [15:0];
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.u1.b  = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.b [15:0];
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.u1.cin  = 1'h0;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.facout_s1  = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.u1.cout ;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.fas_s1  = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.u1.s ;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.a  = \add_32ns_32ns_32_2_1_U17.din0 ;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.b  = \add_32ns_32ns_32_2_1_U17.din1 ;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.ce  = \add_32ns_32ns_32_2_1_U17.ce ;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.clk  = \add_32ns_32ns_32_2_1_U17.clk ;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.reset  = \add_32ns_32ns_32_2_1_U17.reset ;
assign \add_32ns_32ns_32_2_1_U17.dout  = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_8_U.s ;
assign \add_32ns_32ns_32_2_1_U17.ce  = 1'h1;
assign \add_32ns_32ns_32_2_1_U17.clk  = ap_clk;
assign \add_32ns_32ns_32_2_1_U17.din0  = ret_V_22_reg_1212;
assign \add_32ns_32ns_32_2_1_U17.din1  = op_19;
assign grp_fu_847_p2 = \add_32ns_32ns_32_2_1_U17.dout ;
assign \add_32ns_32ns_32_2_1_U17.reset  = ap_rst;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_8_U.ain_s0  = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_8_U.a ;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_8_U.bin_s0  = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_8_U.b ;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_8_U.s  = { \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_8_U.fas_s2 , \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_8_U.sum_s1  };
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_8_U.u2.a  = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_8_U.ain_s1 ;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_8_U.u2.b  = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_8_U.bin_s1 ;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_8_U.u2.cin  = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_8_U.carry_s1 ;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_8_U.facout_s2  = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_8_U.u2.cout ;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_8_U.fas_s2  = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_8_U.u2.s ;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_8_U.u1.a  = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_8_U.a [15:0];
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_8_U.u1.b  = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_8_U.b [15:0];
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_8_U.u1.cin  = 1'h0;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_8_U.facout_s1  = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_8_U.u1.cout ;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_8_U.fas_s1  = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_8_U.u1.s ;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_8_U.a  = \add_32ns_32ns_32_2_1_U14.din0 ;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_8_U.b  = \add_32ns_32ns_32_2_1_U14.din1 ;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_8_U.ce  = \add_32ns_32ns_32_2_1_U14.ce ;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_8_U.clk  = \add_32ns_32ns_32_2_1_U14.clk ;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_8_U.reset  = \add_32ns_32ns_32_2_1_U14.reset ;
assign \add_32ns_32ns_32_2_1_U14.dout  = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_8_U.s ;
assign \add_32ns_32ns_32_2_1_U14.ce  = 1'h1;
assign \add_32ns_32ns_32_2_1_U14.clk  = ap_clk;
assign \add_32ns_32ns_32_2_1_U14.din0  = ret_V_20_cast_reg_1175;
assign \add_32ns_32ns_32_2_1_U14.din1  = 32'd1;
assign grp_fu_776_p2 = \add_32ns_32ns_32_2_1_U14.dout ;
assign \add_32ns_32ns_32_2_1_U14.reset  = ap_rst;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_8_U.ain_s0  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_8_U.a ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_8_U.bin_s0  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_8_U.b ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_8_U.s  = { \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_8_U.fas_s2 , \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_8_U.sum_s1  };
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_8_U.u2.a  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_8_U.ain_s1 ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_8_U.u2.b  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_8_U.bin_s1 ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_8_U.u2.cin  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_8_U.carry_s1 ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_8_U.facout_s2  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_8_U.u2.cout ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_8_U.fas_s2  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_8_U.u2.s ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_8_U.u1.a  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_8_U.a [15:0];
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_8_U.u1.b  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_8_U.b [15:0];
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_8_U.u1.cin  = 1'h0;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_8_U.facout_s1  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_8_U.u1.cout ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_8_U.fas_s1  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_8_U.u1.s ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_8_U.a  = \add_32ns_32ns_32_2_1_U12.din0 ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_8_U.b  = \add_32ns_32ns_32_2_1_U12.din1 ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_8_U.ce  = \add_32ns_32ns_32_2_1_U12.ce ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_8_U.clk  = \add_32ns_32ns_32_2_1_U12.clk ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_8_U.reset  = \add_32ns_32ns_32_2_1_U12.reset ;
assign \add_32ns_32ns_32_2_1_U12.dout  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_8_U.s ;
assign \add_32ns_32ns_32_2_1_U12.ce  = 1'h1;
assign \add_32ns_32ns_32_2_1_U12.clk  = ap_clk;
assign \add_32ns_32ns_32_2_1_U12.din0  = add_ln69_reg_1145;
assign \add_32ns_32ns_32_2_1_U12.din1  = ret_V_20_reg_1140;
assign grp_fu_731_p2 = \add_32ns_32ns_32_2_1_U12.dout ;
assign \add_32ns_32ns_32_2_1_U12.reset  = ap_rst;
assign \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.ain_s0  = \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.a ;
assign \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.bin_s0  = \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.b ;
assign \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.s  = { \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.fas_s2 , \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.sum_s1  };
assign \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.u2.a  = \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.ain_s1 ;
assign \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.u2.b  = \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.bin_s1 ;
assign \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.u2.cin  = \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.carry_s1 ;
assign \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.facout_s2  = \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.u2.cout ;
assign \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.fas_s2  = \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.u2.s ;
assign \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.u1.a  = \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.a [15:0];
assign \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.u1.b  = \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.b [15:0];
assign \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.u1.cin  = 1'h0;
assign \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.facout_s1  = \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.u1.cout ;
assign \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.fas_s1  = \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.u1.s ;
assign \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.a  = \add_32ns_32ns_32_2_1_U11.din0 ;
assign \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.b  = \add_32ns_32ns_32_2_1_U11.din1 ;
assign \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.ce  = \add_32ns_32ns_32_2_1_U11.ce ;
assign \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.clk  = \add_32ns_32ns_32_2_1_U11.clk ;
assign \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.reset  = \add_32ns_32ns_32_2_1_U11.reset ;
assign \add_32ns_32ns_32_2_1_U11.dout  = \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_8_U.s ;
assign \add_32ns_32ns_32_2_1_U11.ce  = 1'h1;
assign \add_32ns_32ns_32_2_1_U11.clk  = ap_clk;
assign \add_32ns_32ns_32_2_1_U11.din0  = { 30'h00000000, ret_reg_980 };
assign \add_32ns_32ns_32_2_1_U11.din1  = op_15;
assign grp_fu_725_p2 = \add_32ns_32ns_32_2_1_U11.dout ;
assign \add_32ns_32ns_32_2_1_U11.reset  = ap_rst;
assign \add_14s_14s_14_2_1_U4.top_add_14s_14s_14_2_1_Adder_3_U.ain_s0  = \add_14s_14s_14_2_1_U4.top_add_14s_14s_14_2_1_Adder_3_U.a ;
assign \add_14s_14s_14_2_1_U4.top_add_14s_14s_14_2_1_Adder_3_U.bin_s0  = \add_14s_14s_14_2_1_U4.top_add_14s_14s_14_2_1_Adder_3_U.b ;
assign \add_14s_14s_14_2_1_U4.top_add_14s_14s_14_2_1_Adder_3_U.s  = { \add_14s_14s_14_2_1_U4.top_add_14s_14s_14_2_1_Adder_3_U.fas_s2 , \add_14s_14s_14_2_1_U4.top_add_14s_14s_14_2_1_Adder_3_U.sum_s1  };
assign \add_14s_14s_14_2_1_U4.top_add_14s_14s_14_2_1_Adder_3_U.u2.a  = \add_14s_14s_14_2_1_U4.top_add_14s_14s_14_2_1_Adder_3_U.ain_s1 ;
assign \add_14s_14s_14_2_1_U4.top_add_14s_14s_14_2_1_Adder_3_U.u2.b  = \add_14s_14s_14_2_1_U4.top_add_14s_14s_14_2_1_Adder_3_U.bin_s1 ;
assign \add_14s_14s_14_2_1_U4.top_add_14s_14s_14_2_1_Adder_3_U.u2.cin  = \add_14s_14s_14_2_1_U4.top_add_14s_14s_14_2_1_Adder_3_U.carry_s1 ;
assign \add_14s_14s_14_2_1_U4.top_add_14s_14s_14_2_1_Adder_3_U.facout_s2  = \add_14s_14s_14_2_1_U4.top_add_14s_14s_14_2_1_Adder_3_U.u2.cout ;
assign \add_14s_14s_14_2_1_U4.top_add_14s_14s_14_2_1_Adder_3_U.fas_s2  = \add_14s_14s_14_2_1_U4.top_add_14s_14s_14_2_1_Adder_3_U.u2.s ;
assign \add_14s_14s_14_2_1_U4.top_add_14s_14s_14_2_1_Adder_3_U.u1.a  = \add_14s_14s_14_2_1_U4.top_add_14s_14s_14_2_1_Adder_3_U.a [6:0];
assign \add_14s_14s_14_2_1_U4.top_add_14s_14s_14_2_1_Adder_3_U.u1.b  = \add_14s_14s_14_2_1_U4.top_add_14s_14s_14_2_1_Adder_3_U.b [6:0];
assign \add_14s_14s_14_2_1_U4.top_add_14s_14s_14_2_1_Adder_3_U.u1.cin  = 1'h0;
assign \add_14s_14s_14_2_1_U4.top_add_14s_14s_14_2_1_Adder_3_U.facout_s1  = \add_14s_14s_14_2_1_U4.top_add_14s_14s_14_2_1_Adder_3_U.u1.cout ;
assign \add_14s_14s_14_2_1_U4.top_add_14s_14s_14_2_1_Adder_3_U.fas_s1  = \add_14s_14s_14_2_1_U4.top_add_14s_14s_14_2_1_Adder_3_U.u1.s ;
assign \add_14s_14s_14_2_1_U4.top_add_14s_14s_14_2_1_Adder_3_U.a  = \add_14s_14s_14_2_1_U4.din0 ;
assign \add_14s_14s_14_2_1_U4.top_add_14s_14s_14_2_1_Adder_3_U.b  = \add_14s_14s_14_2_1_U4.din1 ;
assign \add_14s_14s_14_2_1_U4.top_add_14s_14s_14_2_1_Adder_3_U.ce  = \add_14s_14s_14_2_1_U4.ce ;
assign \add_14s_14s_14_2_1_U4.top_add_14s_14s_14_2_1_Adder_3_U.clk  = \add_14s_14s_14_2_1_U4.clk ;
assign \add_14s_14s_14_2_1_U4.top_add_14s_14s_14_2_1_Adder_3_U.reset  = \add_14s_14s_14_2_1_U4.reset ;
assign \add_14s_14s_14_2_1_U4.dout  = \add_14s_14s_14_2_1_U4.top_add_14s_14s_14_2_1_Adder_3_U.s ;
assign \add_14s_14s_14_2_1_U4.ce  = 1'h1;
assign \add_14s_14s_14_2_1_U4.clk  = ap_clk;
assign \add_14s_14s_14_2_1_U4.din0  = { select_ln850_3_reg_1006[5], select_ln850_3_reg_1006, 7'h00 };
assign \add_14s_14s_14_2_1_U4.din1  = { op_9_V_reg_996[7], op_9_V_reg_996[7], op_9_V_reg_996[7], op_9_V_reg_996[7], op_9_V_reg_996[7], op_9_V_reg_996[7], op_9_V_reg_996 };
assign grp_fu_552_p2 = \add_14s_14s_14_2_1_U4.dout ;
assign \add_14s_14s_14_2_1_U4.reset  = ap_rst;
endmodule


// Product machine:
module top_A_times_top_B (ap_start, op_0, op_1, op_10, op_12, op_13, op_15, op_16, op_18, op_19, op_2, op_6, ap_clk, unsafe_signal);
input ap_start;
input [7:0] op_0;
input [3:0] op_1;
input [1:0] op_10;
input [3:0] op_12;
input [1:0] op_13;
input [31:0] op_15;
input [31:0] op_16;
input [3:0] op_18;
input [31:0] op_19;
input op_2;
input op_6;
input ap_clk;
output unsafe_signal;
reg _setup;
initial _setup = 1'b0;
always @ (posedge ap_clk) _setup <= 1'b1;
reg ap_start_internal;
always @ (posedge ap_clk) if (!_setup) ap_start_internal <= ap_start;
reg [7:0] op_0_internal;
always @ (posedge ap_clk) if (!_setup) op_0_internal <= op_0;
reg [3:0] op_1_internal;
always @ (posedge ap_clk) if (!_setup) op_1_internal <= op_1;
reg [1:0] op_10_internal;
always @ (posedge ap_clk) if (!_setup) op_10_internal <= op_10;
reg [3:0] op_12_internal;
always @ (posedge ap_clk) if (!_setup) op_12_internal <= op_12;
reg [1:0] op_13_internal;
always @ (posedge ap_clk) if (!_setup) op_13_internal <= op_13;
reg [31:0] op_15_internal;
always @ (posedge ap_clk) if (!_setup) op_15_internal <= op_15;
reg [31:0] op_16_internal;
always @ (posedge ap_clk) if (!_setup) op_16_internal <= op_16;
reg [3:0] op_18_internal;
always @ (posedge ap_clk) if (!_setup) op_18_internal <= op_18;
reg [31:0] op_19_internal;
always @ (posedge ap_clk) if (!_setup) op_19_internal <= op_19;
reg op_2_internal;
always @ (posedge ap_clk) if (!_setup) op_2_internal <= op_2;
reg op_6_internal;
always @ (posedge ap_clk) if (!_setup) op_6_internal <= op_6;
wire ap_done_A;
wire ap_done_B;
wire ap_done_eq;
assign ap_done_eq = ap_done_A == ap_done_B;
wire ap_idle_A;
wire ap_idle_B;
wire ap_idle_eq;
assign ap_idle_eq = ap_idle_A == ap_idle_B;
wire ap_ready_A;
wire ap_ready_B;
wire ap_ready_eq;
assign ap_ready_eq = ap_ready_A == ap_ready_B;
wire [31:0] op_31_A;
wire [31:0] op_31_B;
wire op_31_eq;
assign op_31_eq = op_31_A == op_31_B;
wire op_31_ap_vld_A;
wire op_31_ap_vld_B;
wire clk_enable_A;
wire clk_enable_B;
assign clk_enable_A = _setup & (~op_31_ap_vld_A | op_31_ap_vld_B);
assign clk_enable_B = _setup;
wire divergent;
assign divergent = ~(ap_done_eq & ap_idle_eq & ap_ready_eq & op_31_eq);
assign unsafe_signal = op_31_ap_vld_A & op_31_ap_vld_B & divergent;
top_A instance_A (
    .ap_clk(ap_clk),
    .clk_enable(clk_enable_A),
    .ap_start(ap_start_internal),
    .op_0(op_0_internal),
    .op_1(op_1_internal),
    .op_10(op_10_internal),
    .op_12(op_12_internal),
    .op_13(op_13_internal),
    .op_15(op_15_internal),
    .op_16(op_16_internal),
    .op_18(op_18_internal),
    .op_19(op_19_internal),
    .op_2(op_2_internal),
    .op_6(op_6_internal),
    .ap_done(ap_done_A),
    .ap_idle(ap_idle_A),
    .ap_ready(ap_ready_A),
    .op_31(op_31_A),
    .op_31_ap_vld(op_31_ap_vld_A)
);
top_B instance_B (
    .ap_clk(ap_clk),
    .clk_enable(clk_enable_B),
    .ap_start(ap_start_internal),
    .op_0(op_0_internal),
    .op_1(op_1_internal),
    .op_10(op_10_internal),
    .op_12(op_12_internal),
    .op_13(op_13_internal),
    .op_15(op_15_internal),
    .op_16(op_16_internal),
    .op_18(op_18_internal),
    .op_19(op_19_internal),
    .op_2(op_2_internal),
    .op_6(op_6_internal),
    .ap_done(ap_done_B),
    .ap_idle(ap_idle_B),
    .ap_ready(ap_ready_B),
    .op_31(op_31_B),
    .op_31_ap_vld(op_31_ap_vld_B)
);
endmodule
