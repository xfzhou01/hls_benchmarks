// Processed by function `construct_kairos` in `verilog_tricks.py`.
// Machine A:
// Processed by function `add_clk_enable_signal` in `verilog_tricks.py`.
// Processed by function `remove_reset_signal` in `verilog_tricks.py`.
module top_A (
  ap_clk,
  ap_start,
  ap_done,
  ap_idle,
  ap_ready,
  op_0,
  op_2,
  op_3,
  op_6,
  op_7,
  op_10,
  op_11,
  op_12,
  op_16,
  op_17,
  op_18,
  op_19,
  op_31,
  op_31_ap_vld,
clk_enable
);
input clk_enable;


input ap_clk;
wire ap_rst;
assign ap_rst = op_31_ap_vld;
input ap_start;
input [15:0] op_0;
input [15:0] op_10;
input op_11;
input op_12;
input [3:0] op_16;
input [1:0] op_17;
input op_18;
input [3:0] op_19;
input op_2;
input [7:0] op_3;
input [1:0] op_6;
input [31:0] op_7;
output ap_done;
output ap_idle;
output ap_ready;
output [31:0] op_31;
output op_31_ap_vld;


reg [4:0] \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.ain_s1 ;
reg [4:0] \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.bin_s1 ;
reg \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.carry_s1 ;
reg [4:0] \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.sum_s1 ;
reg [4:0] \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.ain_s1 ;
reg [4:0] \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.bin_s1 ;
reg \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.carry_s1 ;
reg [4:0] \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.sum_s1 ;
reg [4:0] \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.ain_s1 ;
reg [4:0] \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.bin_s1 ;
reg \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.carry_s1 ;
reg [4:0] \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.sum_s1 ;
reg [8:0] \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.ain_s1 ;
reg [8:0] \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.bin_s1 ;
reg \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.carry_s1 ;
reg [7:0] \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.sum_s1 ;
reg \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.ain_s1 ;
reg \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.bin_s1 ;
reg \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.carry_s1 ;
reg \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.sum_s1 ;
reg \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.ain_s1 ;
reg \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.bin_s1 ;
reg \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.carry_s1 ;
reg \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.sum_s1 ;
reg \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.ain_s1 ;
reg \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.bin_s1 ;
reg \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.carry_s1 ;
reg \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.sum_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.ain_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.bin_s1 ;
reg \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.carry_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.sum_s1 ;
reg [16:0] \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.ain_s1 ;
reg [16:0] \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.bin_s1 ;
reg \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.carry_s1 ;
reg [16:0] \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.sum_s1 ;
reg [2:0] \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.ain_s1 ;
reg [2:0] \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.bin_s1 ;
reg \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.carry_s1 ;
reg [1:0] \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.sum_s1 ;
reg [2:0] \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.ain_s1 ;
reg [2:0] \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.bin_s1 ;
reg \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.carry_s1 ;
reg [1:0] \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.sum_s1 ;
reg [2:0] \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.ain_s1 ;
reg [2:0] \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.bin_s1 ;
reg \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.carry_s1 ;
reg [1:0] \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.sum_s1 ;
reg [2:0] \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.ain_s1 ;
reg [2:0] \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.bin_s1 ;
reg \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.carry_s1 ;
reg [1:0] \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.sum_s1 ;
reg [2:0] \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.ain_s1 ;
reg [2:0] \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.bin_s1 ;
reg \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.carry_s1 ;
reg [2:0] \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.sum_s1 ;
reg [3:0] \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.ain_s1 ;
reg [3:0] \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.bin_s1 ;
reg \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.carry_s1 ;
reg [3:0] \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.sum_s1 ;
reg [4:0] \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.ain_s1 ;
reg [4:0] \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.bin_s1 ;
reg \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.carry_s1 ;
reg [3:0] \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.sum_s1 ;
reg [31:0] add_ln691_1_reg_1261;
reg [7:0] add_ln691_reg_1114;
reg [4:0] add_ln69_1_reg_1184;
reg [9:0] add_ln69_2_reg_1214;
reg [4:0] add_ln69_3_reg_1189;
reg [1:0] add_ln69_4_reg_1144;
reg [1:0] add_ln69_5_reg_1194;
reg [5:0] add_ln69_6_reg_1219;
reg [9:0] add_ln69_reg_1179;
reg [32:0] ap_CS_fsm = 33'h000000001;
reg icmp_ln768_reg_984;
reg icmp_ln786_reg_989;
reg icmp_ln850_1_reg_944;
reg icmp_ln850_2_reg_949;
reg icmp_ln850_3_reg_1032;
reg icmp_ln850_reg_939;
reg icmp_ln851_1_reg_1067;
reg icmp_ln851_reg_874;
reg [3:0] op_14_V_reg_1124;
reg [3:0] op_1_V_reg_1016;
reg [4:0] op_21_V_reg_1052;
reg [9:0] op_30_V_reg_1229;
reg or_ln785_reg_1000;
reg p_Result_7_reg_970;
reg p_Result_8_reg_977;
reg [3:0] p_Val2_s_reg_1006;
reg [7:0] r_reg_995;
reg [8:0] ret_V_17_reg_879;
reg [1:0] ret_V_18_reg_896;
reg [7:0] ret_V_19_reg_907;
reg [31:0] ret_V_21_cast_reg_1254;
reg [7:0] ret_V_21_reg_918;
reg ret_V_22_reg_954;
reg [4:0] ret_V_24_reg_1042;
reg [16:0] ret_V_25_reg_1072;
reg [7:0] ret_V_26_reg_1134;
reg [33:0] ret_V_27_reg_1249;
reg [1:0] ret_V_2_reg_891;
reg [1:0] ret_V_reg_884;
reg [1:0] ret_reg_1129;
reg [4:0] select_ln1192_reg_960;
reg [1:0] select_ln1347_1_reg_1087;
reg [1:0] select_ln1347_reg_1082;
reg [3:0] select_ln340_reg_1011;
reg [1:0] select_ln69_1_reg_1139;
reg [1:0] select_ln69_2_reg_1099;
reg [4:0] select_ln69_reg_1047;
reg [8:0] select_ln703_reg_857;
reg [7:0] sext_ln353_reg_902;
reg [7:0] sext_ln850_reg_1092;
reg [7:0] \shl_32s_8ns_32_7_1_U3.din1_cast_array[0] ;
reg [7:0] \shl_32s_8ns_32_7_1_U3.din1_cast_array[1] ;
reg [7:0] \shl_32s_8ns_32_7_1_U3.din1_cast_array[2] ;
reg [7:0] \shl_32s_8ns_32_7_1_U3.din1_cast_array[3] ;
reg [7:0] \shl_32s_8ns_32_7_1_U3.din1_cast_array[4] ;
reg [7:0] \shl_32s_8ns_32_7_1_U3.din1_cast_array[5] ;
reg [31:0] \shl_32s_8ns_32_7_1_U3.dout_array[0] ;
reg [31:0] \shl_32s_8ns_32_7_1_U3.dout_array[1] ;
reg [31:0] \shl_32s_8ns_32_7_1_U3.dout_array[2] ;
reg [31:0] \shl_32s_8ns_32_7_1_U3.dout_array[3] ;
reg [31:0] \shl_32s_8ns_32_7_1_U3.dout_array[4] ;
reg [31:0] \shl_32s_8ns_32_7_1_U3.dout_array[5] ;
reg [31:0] shl_ln1299_reg_1021;
reg \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.ain_s1 ;
reg \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.bin_s1 ;
reg \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.carry_s1 ;
reg \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.sum_s1 ;
reg [1:0] \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.ain_s1 ;
reg [1:0] \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.bin_s1 ;
reg \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.carry_s1 ;
reg [1:0] \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.sum_s1 ;
reg [6:0] tmp_reg_1077;
reg [2:0] trunc_ln703_reg_965;
reg [6:0] trunc_ln851_1_reg_924;
reg [6:0] trunc_ln851_2_reg_1027;
reg [6:0] trunc_ln851_reg_913;
wire [31:0] _000_;
wire [7:0] _001_;
wire [4:0] _002_;
wire [9:0] _003_;
wire [4:0] _004_;
wire [1:0] _005_;
wire [1:0] _006_;
wire [5:0] _007_;
wire [9:0] _008_;
wire [32:0] _009_;
wire _010_;
wire _011_;
wire _012_;
wire _013_;
wire _014_;
wire _015_;
wire _016_;
wire _017_;
wire [3:0] _018_;
wire [2:0] _019_;
wire [4:0] _020_;
wire [9:0] _021_;
wire _022_;
wire _023_;
wire _024_;
wire [2:0] _025_;
wire [7:0] _026_;
wire [8:0] _027_;
wire [1:0] _028_;
wire [7:0] _029_;
wire [31:0] _030_;
wire _031_;
wire _032_;
wire [4:0] _033_;
wire [16:0] _034_;
wire [7:0] _035_;
wire [33:0] _036_;
wire [1:0] _037_;
wire [1:0] _038_;
wire [1:0] _039_;
wire [1:0] _040_;
wire [1:0] _041_;
wire [1:0] _042_;
wire [2:0] _043_;
wire [1:0] _044_;
wire [1:0] _045_;
wire [4:0] _046_;
wire [1:0] _047_;
wire [7:0] _048_;
wire [7:0] _049_;
wire [31:0] _050_;
wire [6:0] _051_;
wire [2:0] _052_;
wire [6:0] _053_;
wire [6:0] _054_;
wire [1:0] _055_;
wire _056_;
wire _057_;
wire _058_;
wire _059_;
wire _060_;
wire _061_;
wire _062_;
wire [4:0] _063_;
wire [4:0] _064_;
wire _065_;
wire [4:0] _066_;
wire [5:0] _067_;
wire [5:0] _068_;
wire [4:0] _069_;
wire [4:0] _070_;
wire _071_;
wire [4:0] _072_;
wire [5:0] _073_;
wire [5:0] _074_;
wire [4:0] _075_;
wire [4:0] _076_;
wire _077_;
wire [4:0] _078_;
wire [5:0] _079_;
wire [5:0] _080_;
wire [8:0] _081_;
wire [8:0] _082_;
wire _083_;
wire [7:0] _084_;
wire [8:0] _085_;
wire [9:0] _086_;
wire _087_;
wire _088_;
wire _089_;
wire _090_;
wire [1:0] _091_;
wire [1:0] _092_;
wire _093_;
wire _094_;
wire _095_;
wire _096_;
wire [1:0] _097_;
wire [1:0] _098_;
wire _099_;
wire _100_;
wire _101_;
wire _102_;
wire [1:0] _103_;
wire [1:0] _104_;
wire [15:0] _105_;
wire [15:0] _106_;
wire _107_;
wire [15:0] _108_;
wire [16:0] _109_;
wire [16:0] _110_;
wire [16:0] _111_;
wire [16:0] _112_;
wire _113_;
wire [16:0] _114_;
wire [17:0] _115_;
wire [17:0] _116_;
wire [2:0] _117_;
wire [2:0] _118_;
wire _119_;
wire [1:0] _120_;
wire [2:0] _121_;
wire [3:0] _122_;
wire [2:0] _123_;
wire [2:0] _124_;
wire _125_;
wire [1:0] _126_;
wire [2:0] _127_;
wire [3:0] _128_;
wire [2:0] _129_;
wire [2:0] _130_;
wire _131_;
wire [1:0] _132_;
wire [2:0] _133_;
wire [3:0] _134_;
wire [2:0] _135_;
wire [2:0] _136_;
wire _137_;
wire [1:0] _138_;
wire [2:0] _139_;
wire [3:0] _140_;
wire [2:0] _141_;
wire [2:0] _142_;
wire _143_;
wire [2:0] _144_;
wire [3:0] _145_;
wire [3:0] _146_;
wire [3:0] _147_;
wire [3:0] _148_;
wire _149_;
wire [3:0] _150_;
wire [4:0] _151_;
wire [4:0] _152_;
wire [4:0] _153_;
wire [4:0] _154_;
wire _155_;
wire [3:0] _156_;
wire [4:0] _157_;
wire [5:0] _158_;
wire [7:0] _159_;
wire [7:0] _160_;
wire [7:0] _161_;
wire [7:0] _162_;
wire [7:0] _163_;
wire [7:0] _164_;
wire [31:0] _165_;
wire [31:0] _166_;
wire [31:0] _167_;
wire [31:0] _168_;
wire [31:0] _169_;
wire [31:0] _170_;
wire [7:0] _171_;
wire [31:0] _172_;
wire [7:0] _173_;
wire [31:0] _174_;
wire [7:0] _175_;
wire [31:0] _176_;
wire [7:0] _177_;
wire [31:0] _178_;
wire [7:0] _179_;
wire [31:0] _180_;
wire [7:0] _181_;
wire [31:0] _182_;
wire [31:0] _183_;
wire [31:0] _184_;
wire [31:0] _185_;
wire _186_;
wire _187_;
wire _188_;
wire _189_;
wire [1:0] _190_;
wire [1:0] _191_;
wire [1:0] _192_;
wire [1:0] _193_;
wire _194_;
wire [1:0] _195_;
wire [2:0] _196_;
wire [2:0] _197_;
wire _198_;
wire _199_;
wire _200_;
wire _201_;
wire _202_;
wire _203_;
wire _204_;
wire _205_;
wire _206_;
wire _207_;
wire _208_;
wire _209_;
wire _210_;
wire _211_;
wire _212_;
wire _213_;
wire _214_;
wire _215_;
wire _216_;
wire _217_;
wire _218_;
wire _219_;
wire _220_;
wire _221_;
wire _222_;
wire _223_;
wire _224_;
wire _225_;
wire _226_;
wire _227_;
wire _228_;
wire _229_;
wire _230_;
wire _231_;
wire _232_;
wire _233_;
wire _234_;
wire _235_;
wire _236_;
wire _237_;
wire \add_10s_10ns_10_2_1_U11.ce ;
wire \add_10s_10ns_10_2_1_U11.clk ;
wire [9:0] \add_10s_10ns_10_2_1_U11.din0 ;
wire [9:0] \add_10s_10ns_10_2_1_U11.din1 ;
wire [9:0] \add_10s_10ns_10_2_1_U11.dout ;
wire \add_10s_10ns_10_2_1_U11.reset ;
wire [9:0] \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.a ;
wire [9:0] \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.ain_s0 ;
wire [9:0] \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.b ;
wire [9:0] \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.bin_s0 ;
wire \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.ce ;
wire \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.clk ;
wire \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.facout_s1 ;
wire \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.facout_s2 ;
wire [4:0] \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.fas_s1 ;
wire [4:0] \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.fas_s2 ;
wire \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.reset ;
wire [9:0] \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.s ;
wire [4:0] \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.u1.a ;
wire [4:0] \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.u1.b ;
wire \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.u1.cin ;
wire \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.u1.cout ;
wire [4:0] \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.u1.s ;
wire [4:0] \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.u2.a ;
wire [4:0] \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.u2.b ;
wire \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.u2.cin ;
wire \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.u2.cout ;
wire [4:0] \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.u2.s ;
wire \add_10s_10ns_10_2_1_U15.ce ;
wire \add_10s_10ns_10_2_1_U15.clk ;
wire [9:0] \add_10s_10ns_10_2_1_U15.din0 ;
wire [9:0] \add_10s_10ns_10_2_1_U15.din1 ;
wire [9:0] \add_10s_10ns_10_2_1_U15.dout ;
wire \add_10s_10ns_10_2_1_U15.reset ;
wire [9:0] \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.a ;
wire [9:0] \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.ain_s0 ;
wire [9:0] \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.b ;
wire [9:0] \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.bin_s0 ;
wire \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.ce ;
wire \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.clk ;
wire \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.facout_s1 ;
wire \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.facout_s2 ;
wire [4:0] \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.fas_s1 ;
wire [4:0] \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.fas_s2 ;
wire \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.reset ;
wire [9:0] \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.s ;
wire [4:0] \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.u1.a ;
wire [4:0] \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.u1.b ;
wire \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.u1.cin ;
wire \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.u1.cout ;
wire [4:0] \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.u1.s ;
wire [4:0] \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.u2.a ;
wire [4:0] \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.u2.b ;
wire \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.u2.cin ;
wire \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.u2.cout ;
wire [4:0] \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.u2.s ;
wire \add_10s_10ns_10_2_1_U17.ce ;
wire \add_10s_10ns_10_2_1_U17.clk ;
wire [9:0] \add_10s_10ns_10_2_1_U17.din0 ;
wire [9:0] \add_10s_10ns_10_2_1_U17.din1 ;
wire [9:0] \add_10s_10ns_10_2_1_U17.dout ;
wire \add_10s_10ns_10_2_1_U17.reset ;
wire [9:0] \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.a ;
wire [9:0] \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.ain_s0 ;
wire [9:0] \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.b ;
wire [9:0] \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.bin_s0 ;
wire \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.ce ;
wire \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.clk ;
wire \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.facout_s1 ;
wire \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.facout_s2 ;
wire [4:0] \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.fas_s1 ;
wire [4:0] \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.fas_s2 ;
wire \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.reset ;
wire [9:0] \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.s ;
wire [4:0] \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.u1.a ;
wire [4:0] \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.u1.b ;
wire \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.u1.cin ;
wire \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.u1.cout ;
wire [4:0] \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.u1.s ;
wire [4:0] \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.u2.a ;
wire [4:0] \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.u2.b ;
wire \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.u2.cin ;
wire \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.u2.cout ;
wire [4:0] \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.u2.s ;
wire \add_17s_17s_17_2_1_U6.ce ;
wire \add_17s_17s_17_2_1_U6.clk ;
wire [16:0] \add_17s_17s_17_2_1_U6.din0 ;
wire [16:0] \add_17s_17s_17_2_1_U6.din1 ;
wire [16:0] \add_17s_17s_17_2_1_U6.dout ;
wire \add_17s_17s_17_2_1_U6.reset ;
wire [16:0] \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.a ;
wire [16:0] \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.ain_s0 ;
wire [16:0] \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.b ;
wire [16:0] \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.bin_s0 ;
wire \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.ce ;
wire \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.clk ;
wire \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.facout_s1 ;
wire \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.facout_s2 ;
wire [7:0] \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.fas_s1 ;
wire [8:0] \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.fas_s2 ;
wire \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.reset ;
wire [16:0] \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.s ;
wire [7:0] \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.u1.a ;
wire [7:0] \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.u1.b ;
wire \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.u1.cin ;
wire \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.u1.cout ;
wire [7:0] \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.u1.s ;
wire [8:0] \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.u2.a ;
wire [8:0] \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.u2.b ;
wire \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.u2.cin ;
wire \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.u2.cout ;
wire [8:0] \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.u2.s ;
wire \add_2ns_2ns_2_2_1_U10.ce ;
wire \add_2ns_2ns_2_2_1_U10.clk ;
wire [1:0] \add_2ns_2ns_2_2_1_U10.din0 ;
wire [1:0] \add_2ns_2ns_2_2_1_U10.din1 ;
wire [1:0] \add_2ns_2ns_2_2_1_U10.dout ;
wire \add_2ns_2ns_2_2_1_U10.reset ;
wire [1:0] \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.a ;
wire [1:0] \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.ain_s0 ;
wire [1:0] \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.b ;
wire [1:0] \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.bin_s0 ;
wire \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.ce ;
wire \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.clk ;
wire \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.facout_s1 ;
wire \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.facout_s2 ;
wire \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.fas_s1 ;
wire \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.fas_s2 ;
wire \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.reset ;
wire [1:0] \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.s ;
wire \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.a ;
wire \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.b ;
wire \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.cin ;
wire \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.cout ;
wire \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.s ;
wire \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.a ;
wire \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.b ;
wire \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.cin ;
wire \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.cout ;
wire \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.s ;
wire \add_2ns_2ns_2_2_1_U14.ce ;
wire \add_2ns_2ns_2_2_1_U14.clk ;
wire [1:0] \add_2ns_2ns_2_2_1_U14.din0 ;
wire [1:0] \add_2ns_2ns_2_2_1_U14.din1 ;
wire [1:0] \add_2ns_2ns_2_2_1_U14.dout ;
wire \add_2ns_2ns_2_2_1_U14.reset ;
wire [1:0] \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.a ;
wire [1:0] \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.ain_s0 ;
wire [1:0] \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.b ;
wire [1:0] \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.bin_s0 ;
wire \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.ce ;
wire \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.clk ;
wire \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.facout_s1 ;
wire \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.facout_s2 ;
wire \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.fas_s1 ;
wire \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.fas_s2 ;
wire \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.reset ;
wire [1:0] \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.s ;
wire \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.a ;
wire \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.b ;
wire \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.cin ;
wire \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.cout ;
wire \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.s ;
wire \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.a ;
wire \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.b ;
wire \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.cin ;
wire \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.cout ;
wire \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.s ;
wire \add_2ns_2ns_2_2_1_U2.ce ;
wire \add_2ns_2ns_2_2_1_U2.clk ;
wire [1:0] \add_2ns_2ns_2_2_1_U2.din0 ;
wire [1:0] \add_2ns_2ns_2_2_1_U2.din1 ;
wire [1:0] \add_2ns_2ns_2_2_1_U2.dout ;
wire \add_2ns_2ns_2_2_1_U2.reset ;
wire [1:0] \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.a ;
wire [1:0] \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.ain_s0 ;
wire [1:0] \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.b ;
wire [1:0] \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.bin_s0 ;
wire \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.ce ;
wire \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.clk ;
wire \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.facout_s1 ;
wire \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.facout_s2 ;
wire \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.fas_s1 ;
wire \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.fas_s2 ;
wire \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.reset ;
wire [1:0] \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.s ;
wire \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.a ;
wire \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.b ;
wire \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.cin ;
wire \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.cout ;
wire \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.s ;
wire \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.a ;
wire \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.b ;
wire \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.cin ;
wire \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.cout ;
wire \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.s ;
wire \add_32ns_32ns_32_2_1_U19.ce ;
wire \add_32ns_32ns_32_2_1_U19.clk ;
wire [31:0] \add_32ns_32ns_32_2_1_U19.din0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U19.din1 ;
wire [31:0] \add_32ns_32ns_32_2_1_U19.dout ;
wire \add_32ns_32ns_32_2_1_U19.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.a ;
wire [31:0] \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.ain_s0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.b ;
wire [31:0] \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.bin_s0 ;
wire \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.ce ;
wire \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.clk ;
wire \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.facout_s1 ;
wire \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.facout_s2 ;
wire [15:0] \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.fas_s1 ;
wire [15:0] \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.fas_s2 ;
wire \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.u1.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.u1.b ;
wire \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.u1.cin ;
wire \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.u1.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.u1.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.u2.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.u2.b ;
wire \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.u2.cin ;
wire \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.u2.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.u2.s ;
wire \add_34s_34s_34_2_1_U18.ce ;
wire \add_34s_34s_34_2_1_U18.clk ;
wire [33:0] \add_34s_34s_34_2_1_U18.din0 ;
wire [33:0] \add_34s_34s_34_2_1_U18.din1 ;
wire [33:0] \add_34s_34s_34_2_1_U18.dout ;
wire \add_34s_34s_34_2_1_U18.reset ;
wire [33:0] \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.a ;
wire [33:0] \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.ain_s0 ;
wire [33:0] \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.b ;
wire [33:0] \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.bin_s0 ;
wire \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.ce ;
wire \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.clk ;
wire \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.facout_s1 ;
wire \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.facout_s2 ;
wire [16:0] \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.fas_s1 ;
wire [16:0] \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.fas_s2 ;
wire \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.reset ;
wire [33:0] \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.s ;
wire [16:0] \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.u1.a ;
wire [16:0] \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.u1.b ;
wire \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.u1.cin ;
wire \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.u1.cout ;
wire [16:0] \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.u1.s ;
wire [16:0] \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.u2.a ;
wire [16:0] \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.u2.b ;
wire \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.u2.cin ;
wire \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.u2.cout ;
wire [16:0] \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.u2.s ;
wire \add_5ns_5ns_5_2_1_U13.ce ;
wire \add_5ns_5ns_5_2_1_U13.clk ;
wire [4:0] \add_5ns_5ns_5_2_1_U13.din0 ;
wire [4:0] \add_5ns_5ns_5_2_1_U13.din1 ;
wire [4:0] \add_5ns_5ns_5_2_1_U13.dout ;
wire \add_5ns_5ns_5_2_1_U13.reset ;
wire [4:0] \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.a ;
wire [4:0] \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.ain_s0 ;
wire [4:0] \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.b ;
wire [4:0] \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.bin_s0 ;
wire \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.ce ;
wire \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.clk ;
wire \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.facout_s1 ;
wire \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.facout_s2 ;
wire [1:0] \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.fas_s1 ;
wire [2:0] \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.fas_s2 ;
wire \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.reset ;
wire [4:0] \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.s ;
wire [1:0] \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.u1.a ;
wire [1:0] \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.u1.b ;
wire \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.u1.cin ;
wire \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.u1.cout ;
wire [1:0] \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.u1.s ;
wire [2:0] \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.u2.a ;
wire [2:0] \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.u2.b ;
wire \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.u2.cin ;
wire \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.u2.cout ;
wire [2:0] \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.u2.s ;
wire \add_5ns_5ns_5_2_1_U5.ce ;
wire \add_5ns_5ns_5_2_1_U5.clk ;
wire [4:0] \add_5ns_5ns_5_2_1_U5.din0 ;
wire [4:0] \add_5ns_5ns_5_2_1_U5.din1 ;
wire [4:0] \add_5ns_5ns_5_2_1_U5.dout ;
wire \add_5ns_5ns_5_2_1_U5.reset ;
wire [4:0] \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.a ;
wire [4:0] \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.ain_s0 ;
wire [4:0] \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.b ;
wire [4:0] \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.bin_s0 ;
wire \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.ce ;
wire \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.clk ;
wire \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.facout_s1 ;
wire \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.facout_s2 ;
wire [1:0] \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.fas_s1 ;
wire [2:0] \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.fas_s2 ;
wire \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.reset ;
wire [4:0] \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.s ;
wire [1:0] \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.u1.a ;
wire [1:0] \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.u1.b ;
wire \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.u1.cin ;
wire \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.u1.cout ;
wire [1:0] \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.u1.s ;
wire [2:0] \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.u2.a ;
wire [2:0] \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.u2.b ;
wire \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.u2.cin ;
wire \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.u2.cout ;
wire [2:0] \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.u2.s ;
wire \add_5ns_5s_5_2_1_U4.ce ;
wire \add_5ns_5s_5_2_1_U4.clk ;
wire [4:0] \add_5ns_5s_5_2_1_U4.din0 ;
wire [4:0] \add_5ns_5s_5_2_1_U4.din1 ;
wire [4:0] \add_5ns_5s_5_2_1_U4.dout ;
wire \add_5ns_5s_5_2_1_U4.reset ;
wire [4:0] \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.a ;
wire [4:0] \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.ain_s0 ;
wire [4:0] \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.b ;
wire [4:0] \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.bin_s0 ;
wire \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.ce ;
wire \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.clk ;
wire \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.facout_s1 ;
wire \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.facout_s2 ;
wire [1:0] \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.fas_s1 ;
wire [2:0] \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.fas_s2 ;
wire \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.reset ;
wire [4:0] \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.s ;
wire [1:0] \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.u1.a ;
wire [1:0] \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.u1.b ;
wire \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.u1.cin ;
wire \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.u1.cout ;
wire [1:0] \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.u1.s ;
wire [2:0] \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.u2.a ;
wire [2:0] \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.u2.b ;
wire \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.u2.cin ;
wire \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.u2.cout ;
wire [2:0] \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.u2.s ;
wire \add_5s_5s_5_2_1_U12.ce ;
wire \add_5s_5s_5_2_1_U12.clk ;
wire [4:0] \add_5s_5s_5_2_1_U12.din0 ;
wire [4:0] \add_5s_5s_5_2_1_U12.din1 ;
wire [4:0] \add_5s_5s_5_2_1_U12.dout ;
wire \add_5s_5s_5_2_1_U12.reset ;
wire [4:0] \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.a ;
wire [4:0] \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.ain_s0 ;
wire [4:0] \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.b ;
wire [4:0] \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.bin_s0 ;
wire \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.ce ;
wire \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.clk ;
wire \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.facout_s1 ;
wire \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.facout_s2 ;
wire [1:0] \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.fas_s1 ;
wire [2:0] \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.fas_s2 ;
wire \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.reset ;
wire [4:0] \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.s ;
wire [1:0] \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.u1.a ;
wire [1:0] \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.u1.b ;
wire \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.u1.cin ;
wire \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.u1.cout ;
wire [1:0] \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.u1.s ;
wire [2:0] \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.u2.a ;
wire [2:0] \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.u2.b ;
wire \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.u2.cin ;
wire \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.u2.cout ;
wire [2:0] \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.u2.s ;
wire \add_6s_6ns_6_2_1_U16.ce ;
wire \add_6s_6ns_6_2_1_U16.clk ;
wire [5:0] \add_6s_6ns_6_2_1_U16.din0 ;
wire [5:0] \add_6s_6ns_6_2_1_U16.din1 ;
wire [5:0] \add_6s_6ns_6_2_1_U16.dout ;
wire \add_6s_6ns_6_2_1_U16.reset ;
wire [5:0] \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.a ;
wire [5:0] \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.ain_s0 ;
wire [5:0] \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.b ;
wire [5:0] \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.bin_s0 ;
wire \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.ce ;
wire \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.clk ;
wire \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.facout_s1 ;
wire \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.facout_s2 ;
wire [2:0] \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.fas_s1 ;
wire [2:0] \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.fas_s2 ;
wire \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.reset ;
wire [5:0] \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.s ;
wire [2:0] \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.u1.a ;
wire [2:0] \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.u1.b ;
wire \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.u1.cin ;
wire \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.u1.cout ;
wire [2:0] \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.u1.s ;
wire [2:0] \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.u2.a ;
wire [2:0] \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.u2.b ;
wire \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.u2.cin ;
wire \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.u2.cout ;
wire [2:0] \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.u2.s ;
wire \add_8s_8ns_8_2_1_U7.ce ;
wire \add_8s_8ns_8_2_1_U7.clk ;
wire [7:0] \add_8s_8ns_8_2_1_U7.din0 ;
wire [7:0] \add_8s_8ns_8_2_1_U7.din1 ;
wire [7:0] \add_8s_8ns_8_2_1_U7.dout ;
wire \add_8s_8ns_8_2_1_U7.reset ;
wire [7:0] \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.a ;
wire [7:0] \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.ain_s0 ;
wire [7:0] \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.b ;
wire [7:0] \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.bin_s0 ;
wire \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.ce ;
wire \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.clk ;
wire \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.facout_s1 ;
wire \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.facout_s2 ;
wire [3:0] \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.fas_s1 ;
wire [3:0] \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.fas_s2 ;
wire \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.reset ;
wire [7:0] \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.s ;
wire [3:0] \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.u1.a ;
wire [3:0] \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.u1.b ;
wire \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.u1.cin ;
wire \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.u1.cout ;
wire [3:0] \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.u1.s ;
wire [3:0] \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.u2.a ;
wire [3:0] \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.u2.b ;
wire \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.u2.cin ;
wire \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.u2.cout ;
wire [3:0] \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.u2.s ;
wire \add_9ns_9s_9_2_1_U1.ce ;
wire \add_9ns_9s_9_2_1_U1.clk ;
wire [8:0] \add_9ns_9s_9_2_1_U1.din0 ;
wire [8:0] \add_9ns_9s_9_2_1_U1.din1 ;
wire [8:0] \add_9ns_9s_9_2_1_U1.dout ;
wire \add_9ns_9s_9_2_1_U1.reset ;
wire [8:0] \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.a ;
wire [8:0] \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.ain_s0 ;
wire [8:0] \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.b ;
wire [8:0] \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.bin_s0 ;
wire \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.ce ;
wire \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.clk ;
wire \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.facout_s1 ;
wire \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.facout_s2 ;
wire [3:0] \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.fas_s1 ;
wire [4:0] \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.fas_s2 ;
wire \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.reset ;
wire [8:0] \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.s ;
wire [3:0] \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.u1.a ;
wire [3:0] \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.u1.b ;
wire \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.u1.cin ;
wire \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.u1.cout ;
wire [3:0] \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.u1.s ;
wire [4:0] \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.u2.a ;
wire [4:0] \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.u2.b ;
wire \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.u2.cin ;
wire \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.u2.cout ;
wire [4:0] \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.u2.s ;
wire and_ln340_fu_491_p2;
wire and_ln785_1_fu_526_p2;
wire and_ln785_fu_520_p2;
wire and_ln850_1_fu_368_p2;
wire and_ln850_2_fu_568_p2;
wire and_ln850_fu_350_p2;
wire ap_CS_fsm_state1;
wire ap_CS_fsm_state10;
wire ap_CS_fsm_state11;
wire ap_CS_fsm_state12;
wire ap_CS_fsm_state13;
wire ap_CS_fsm_state14;
wire ap_CS_fsm_state15;
wire ap_CS_fsm_state16;
wire ap_CS_fsm_state17;
wire ap_CS_fsm_state18;
wire ap_CS_fsm_state19;
wire ap_CS_fsm_state2;
wire ap_CS_fsm_state20;
wire ap_CS_fsm_state21;
wire ap_CS_fsm_state22;
wire ap_CS_fsm_state23;
wire ap_CS_fsm_state24;
wire ap_CS_fsm_state25;
wire ap_CS_fsm_state26;
wire ap_CS_fsm_state27;
wire ap_CS_fsm_state28;
wire ap_CS_fsm_state29;
wire ap_CS_fsm_state3;
wire ap_CS_fsm_state30;
wire ap_CS_fsm_state31;
wire ap_CS_fsm_state32;
wire ap_CS_fsm_state33;
wire ap_CS_fsm_state4;
wire ap_CS_fsm_state5;
wire ap_CS_fsm_state6;
wire ap_CS_fsm_state7;
wire ap_CS_fsm_state8;
wire ap_CS_fsm_state9;
wire [32:0] ap_NS_fsm;
wire ap_clk;
wire ap_done;
wire ap_idle;
wire ap_ready;
wire ap_rst;
wire ap_start;
wire [8:0] grp_fu_235_p1;
wire [8:0] grp_fu_235_p2;
wire [1:0] grp_fu_256_p2;
wire [31:0] grp_fu_315_p0;
wire [31:0] grp_fu_315_p1;
wire [31:0] grp_fu_315_p2;
wire [4:0] grp_fu_549_p1;
wire [4:0] grp_fu_549_p2;
wire [4:0] grp_fu_587_p2;
wire [16:0] grp_fu_606_p0;
wire [16:0] grp_fu_606_p1;
wire [16:0] grp_fu_606_p2;
wire [7:0] grp_fu_649_p0;
wire [7:0] grp_fu_649_p2;
wire [3:0] grp_fu_671_p0;
wire [3:0] grp_fu_671_p1;
wire [3:0] grp_fu_671_p2;
wire [1:0] grp_fu_677_p2;
wire [1:0] grp_fu_685_p1;
wire [1:0] grp_fu_685_p2;
wire [9:0] grp_fu_741_p0;
wire [9:0] grp_fu_741_p1;
wire [9:0] grp_fu_741_p2;
wire [4:0] grp_fu_747_p0;
wire [4:0] grp_fu_747_p1;
wire [4:0] grp_fu_747_p2;
wire [4:0] grp_fu_753_p0;
wire [4:0] grp_fu_753_p1;
wire [4:0] grp_fu_753_p2;
wire [1:0] grp_fu_759_p2;
wire [9:0] grp_fu_766_p0;
wire [9:0] grp_fu_766_p2;
wire [5:0] grp_fu_777_p0;
wire [5:0] grp_fu_777_p1;
wire [5:0] grp_fu_777_p2;
wire [9:0] grp_fu_786_p0;
wire [9:0] grp_fu_786_p2;
wire [33:0] grp_fu_806_p0;
wire [33:0] grp_fu_806_p1;
wire [33:0] grp_fu_806_p2;
wire [31:0] grp_fu_822_p2;
wire icmp_ln768_fu_416_p2;
wire icmp_ln786_fu_422_p2;
wire icmp_ln850_1_fu_326_p2;
wire icmp_ln850_2_fu_331_p2;
wire icmp_ln850_3_fu_541_p2;
wire icmp_ln850_fu_321_p2;
wire icmp_ln851_1_fu_616_p2;
wire icmp_ln851_fu_240_p2;
wire [7:0] lhs_fu_283_p3;
wire [15:0] op_0;
wire [15:0] op_10;
wire op_11;
wire op_12;
wire [3:0] op_16;
wire [1:0] op_17;
wire op_18;
wire [3:0] op_19;
wire [3:0] op_1_V_fu_531_p3;
wire op_2;
wire [7:0] op_3;
wire [31:0] op_31;
wire op_31_ap_vld;
wire [1:0] op_6;
wire [31:0] op_7;
wire or_ln340_fu_480_p2;
wire or_ln785_1_fu_515_p2;
wire or_ln785_fu_449_p2;
wire or_ln786_fu_475_p2;
wire overflow_fu_465_p2;
wire p_Result_1_fu_343_p3;
wire p_Result_2_fu_561_p3;
wire p_Result_5_fu_690_p3;
wire p_Result_6_fu_827_p3;
wire p_Result_s_12_fu_261_p3;
wire [12:0] p_Result_s_fu_406_p4;
wire [3:0] p_Val2_s_fu_453_p3;
wire [7:0] r_fu_443_p3;
wire ret_V_10_fu_554_p3;
wire [1:0] ret_V_18_fu_273_p3;
wire [7:0] ret_V_19_fu_290_p1;
wire [7:0] ret_V_19_fu_290_p2;
wire ret_V_20_fu_355_p2;
wire [7:0] ret_V_21_fu_299_p1;
wire [7:0] ret_V_21_fu_299_p2;
wire ret_V_22_fu_372_p2;
wire ret_V_23_fu_573_p2;
wire [7:0] ret_V_26_fu_702_p3;
wire ret_V_5_fu_336_p3;
wire ret_V_8_fu_361_p3;
wire [14:0] rhs_2_fu_595_p3;
wire [1:0] select_ln1192_fu_378_p3;
wire [1:0] select_ln1347_1_fu_639_p3;
wire [1:0] select_ln1347_fu_632_p3;
wire [3:0] select_ln340_fu_497_p3;
wire [1:0] select_ln69_1_fu_709_p3;
wire [1:0] select_ln69_2_fu_655_p3;
wire [4:0] select_ln69_fu_579_p3;
wire [8:0] select_ln703_fu_219_p3;
wire [7:0] select_ln850_1_fu_697_p3;
wire [31:0] select_ln850_2_fu_837_p3;
wire [6:0] select_ln850_4_fu_435_p3;
wire [1:0] select_ln850_fu_268_p3;
wire [15:0] sext_ln1192_fu_591_p0;
wire [7:0] sext_ln1299_fu_312_p0;
wire [7:0] sext_ln353_fu_280_p1;
wire [3:0] sext_ln69_1_fu_720_p1;
wire [3:0] sext_ln703_2_fu_791_p0;
wire [7:0] sext_ln703_fu_227_p0;
wire [7:0] sext_ln850_fu_646_p1;
wire \shl_32s_8ns_32_7_1_U3.ce ;
wire \shl_32s_8ns_32_7_1_U3.clk ;
wire [31:0] \shl_32s_8ns_32_7_1_U3.din0 ;
wire [31:0] \shl_32s_8ns_32_7_1_U3.din1 ;
wire [7:0] \shl_32s_8ns_32_7_1_U3.din1_cast ;
wire [7:0] \shl_32s_8ns_32_7_1_U3.din1_mask ;
wire [31:0] \shl_32s_8ns_32_7_1_U3.dout ;
wire \shl_32s_8ns_32_7_1_U3.reset ;
wire \sub_2ns_2ns_2_2_1_U9.ce ;
wire \sub_2ns_2ns_2_2_1_U9.clk ;
wire [1:0] \sub_2ns_2ns_2_2_1_U9.din0 ;
wire [1:0] \sub_2ns_2ns_2_2_1_U9.din1 ;
wire [1:0] \sub_2ns_2ns_2_2_1_U9.dout ;
wire \sub_2ns_2ns_2_2_1_U9.reset ;
wire [1:0] \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.a ;
wire [1:0] \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.ain_s0 ;
wire [1:0] \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.b ;
wire [1:0] \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.bin_s0 ;
wire \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.ce ;
wire \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.clk ;
wire \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.facout_s1 ;
wire \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.facout_s2 ;
wire \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.fas_s1 ;
wire \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.fas_s2 ;
wire \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.reset ;
wire [1:0] \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.s ;
wire \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.u1.a ;
wire \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.u1.b ;
wire \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.u1.cin ;
wire \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.u1.cout ;
wire \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.u1.s ;
wire \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.u2.a ;
wire \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.u2.b ;
wire \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.u2.cin ;
wire \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.u2.cout ;
wire \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.u2.s ;
wire \sub_4s_4ns_4_2_1_U8.ce ;
wire \sub_4s_4ns_4_2_1_U8.clk ;
wire [3:0] \sub_4s_4ns_4_2_1_U8.din0 ;
wire [3:0] \sub_4s_4ns_4_2_1_U8.din1 ;
wire [3:0] \sub_4s_4ns_4_2_1_U8.dout ;
wire \sub_4s_4ns_4_2_1_U8.reset ;
wire [3:0] \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.a ;
wire [3:0] \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.ain_s0 ;
wire [3:0] \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.b ;
wire [3:0] \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.bin_s0 ;
wire \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.ce ;
wire \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.clk ;
wire \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.facout_s1 ;
wire \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.facout_s2 ;
wire [1:0] \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.fas_s1 ;
wire [1:0] \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.fas_s2 ;
wire \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.reset ;
wire [3:0] \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.s ;
wire [1:0] \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.u1.a ;
wire [1:0] \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.u1.b ;
wire \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.u1.cin ;
wire \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.u1.cout ;
wire [1:0] \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.u1.s ;
wire [1:0] \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.u2.a ;
wire [1:0] \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.u2.b ;
wire \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.u2.cin ;
wire \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.u2.cout ;
wire [1:0] \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.u2.s ;
wire [10:0] tmp_11_fu_795_p3;
wire tmp_9_fu_428_p3;
wire [7:0] trunc_ln1192_fu_231_p0;
wire [6:0] trunc_ln1192_fu_231_p1;
wire [2:0] trunc_ln703_fu_386_p1;
wire [6:0] trunc_ln851_1_fu_304_p1;
wire [6:0] trunc_ln851_2_fu_537_p1;
wire [15:0] trunc_ln851_3_fu_612_p0;
wire [9:0] trunc_ln851_3_fu_612_p1;
wire [3:0] trunc_ln851_4_fu_834_p0;
wire trunc_ln851_4_fu_834_p1;
wire [6:0] trunc_ln851_fu_295_p1;
wire xor_ln340_fu_485_p2;
wire xor_ln785_1_fu_510_p2;
wire xor_ln785_fu_460_p2;
wire xor_ln786_1_fu_505_p2;
wire xor_ln786_fu_470_p2;


assign _056_ = icmp_ln851_1_reg_1067 & ap_CS_fsm[20];
assign _057_ = _060_ & ap_CS_fsm[4];
assign _058_ = _061_ & ap_CS_fsm[0];
assign _059_ = ap_start & ap_CS_fsm[0];
assign and_ln340_fu_491_p2 = xor_ln340_fu_485_p2 & or_ln786_fu_475_p2;
assign and_ln785_1_fu_526_p2 = p_Result_8_reg_977 & and_ln785_fu_520_p2;
assign and_ln785_fu_520_p2 = xor_ln786_1_fu_505_p2 & or_ln785_1_fu_515_p2;
assign and_ln850_1_fu_368_p2 = icmp_ln850_2_reg_949 & icmp_ln850_1_reg_944;
assign and_ln850_2_fu_568_p2 = shl_ln1299_reg_1021[7] & icmp_ln850_3_reg_1032;
assign and_ln850_fu_350_p2 = ret_V_19_reg_907[7] & icmp_ln850_reg_939;
assign overflow_fu_465_p2 = xor_ln785_fu_460_p2 & or_ln785_reg_1000;
assign ret_V_21_fu_299_p2 = op_3 & { op_2, 7'h00 };
assign xor_ln786_fu_470_p2 = ~ p_Result_8_reg_977;
assign xor_ln785_fu_460_p2 = ~ p_Result_7_reg_970;
assign xor_ln340_fu_485_p2 = ~ or_ln340_fu_480_p2;
assign xor_ln785_1_fu_510_p2 = ~ or_ln785_reg_1000;
assign xor_ln786_1_fu_505_p2 = ~ icmp_ln786_reg_989;
assign _060_ = ~ icmp_ln851_reg_874;
assign _061_ = ~ ap_start;
assign _062_ = ! op_3[6:0];
always @(posedge \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.clk )
\add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.bin_s1  <= _064_;
always @(posedge \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.clk )
\add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.ain_s1  <= _063_;
always @(posedge \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.clk )
\add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.sum_s1  <= _066_;
always @(posedge \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.clk )
\add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.carry_s1  <= _065_;
assign _064_ = \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.ce  ? \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.b [9:5] : \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.bin_s1 ;
assign _063_ = \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.ce  ? \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.a [9:5] : \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.ain_s1 ;
assign _065_ = \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.ce  ? \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.facout_s1  : \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.carry_s1 ;
assign _066_ = \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.ce  ? \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.fas_s1  : \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.sum_s1 ;
assign _067_ = \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.u1.a  + \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.u1.b ;
assign { \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.u1.cout , \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.u1.s  } = _067_ + \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.u1.cin ;
assign _068_ = \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.u2.a  + \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.u2.b ;
assign { \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.u2.cout , \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.u2.s  } = _068_ + \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.u2.cin ;
always @(posedge \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.clk )
\add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.bin_s1  <= _070_;
always @(posedge \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.clk )
\add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.ain_s1  <= _069_;
always @(posedge \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.clk )
\add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.sum_s1  <= _072_;
always @(posedge \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.clk )
\add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.carry_s1  <= _071_;
assign _070_ = \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.ce  ? \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.b [9:5] : \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.bin_s1 ;
assign _069_ = \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.ce  ? \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.a [9:5] : \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.ain_s1 ;
assign _071_ = \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.ce  ? \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.facout_s1  : \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.carry_s1 ;
assign _072_ = \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.ce  ? \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.fas_s1  : \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.sum_s1 ;
assign _073_ = \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.u1.a  + \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.u1.b ;
assign { \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.u1.cout , \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.u1.s  } = _073_ + \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.u1.cin ;
assign _074_ = \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.u2.a  + \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.u2.b ;
assign { \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.u2.cout , \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.u2.s  } = _074_ + \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.u2.cin ;
always @(posedge \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.clk )
\add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.bin_s1  <= _076_;
always @(posedge \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.clk )
\add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.ain_s1  <= _075_;
always @(posedge \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.clk )
\add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.sum_s1  <= _078_;
always @(posedge \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.clk )
\add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.carry_s1  <= _077_;
assign _076_ = \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.ce  ? \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.b [9:5] : \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.bin_s1 ;
assign _075_ = \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.ce  ? \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.a [9:5] : \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.ain_s1 ;
assign _077_ = \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.ce  ? \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.facout_s1  : \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.carry_s1 ;
assign _078_ = \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.ce  ? \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.fas_s1  : \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.sum_s1 ;
assign _079_ = \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.u1.a  + \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.u1.b ;
assign { \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.u1.cout , \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.u1.s  } = _079_ + \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.u1.cin ;
assign _080_ = \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.u2.a  + \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.u2.b ;
assign { \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.u2.cout , \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.u2.s  } = _080_ + \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.u2.cin ;
always @(posedge \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.clk )
\add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.bin_s1  <= _082_;
always @(posedge \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.clk )
\add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.ain_s1  <= _081_;
always @(posedge \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.clk )
\add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.sum_s1  <= _084_;
always @(posedge \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.clk )
\add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.carry_s1  <= _083_;
assign _082_ = \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.ce  ? \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.b [16:8] : \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.bin_s1 ;
assign _081_ = \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.ce  ? \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.a [16:8] : \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.ain_s1 ;
assign _083_ = \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.ce  ? \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.facout_s1  : \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.carry_s1 ;
assign _084_ = \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.ce  ? \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.fas_s1  : \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.sum_s1 ;
assign _085_ = \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.u1.a  + \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.u1.b ;
assign { \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.u1.cout , \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.u1.s  } = _085_ + \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.u1.cin ;
assign _086_ = \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.u2.a  + \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.u2.b ;
assign { \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.u2.cout , \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.u2.s  } = _086_ + \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.u2.cin ;
always @(posedge \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.clk )
\add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.bin_s1  <= _088_;
always @(posedge \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.clk )
\add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.ain_s1  <= _087_;
always @(posedge \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.clk )
\add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.sum_s1  <= _090_;
always @(posedge \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.clk )
\add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.carry_s1  <= _089_;
assign _088_ = \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.ce  ? \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.b [1] : \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.bin_s1 ;
assign _087_ = \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.ce  ? \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.a [1] : \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.ain_s1 ;
assign _089_ = \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.ce  ? \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.facout_s1  : \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.carry_s1 ;
assign _090_ = \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.ce  ? \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.fas_s1  : \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.sum_s1 ;
assign _091_ = \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.a  + \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.b ;
assign { \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.cout , \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.s  } = _091_ + \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.cin ;
assign _092_ = \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.a  + \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.b ;
assign { \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.cout , \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.s  } = _092_ + \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.cin ;
always @(posedge \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.clk )
\add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.bin_s1  <= _094_;
always @(posedge \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.clk )
\add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.ain_s1  <= _093_;
always @(posedge \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.clk )
\add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.sum_s1  <= _096_;
always @(posedge \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.clk )
\add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.carry_s1  <= _095_;
assign _094_ = \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.ce  ? \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.b [1] : \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.bin_s1 ;
assign _093_ = \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.ce  ? \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.a [1] : \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.ain_s1 ;
assign _095_ = \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.ce  ? \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.facout_s1  : \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.carry_s1 ;
assign _096_ = \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.ce  ? \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.fas_s1  : \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.sum_s1 ;
assign _097_ = \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.a  + \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.b ;
assign { \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.cout , \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.s  } = _097_ + \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.cin ;
assign _098_ = \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.a  + \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.b ;
assign { \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.cout , \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.s  } = _098_ + \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.cin ;
always @(posedge \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.clk )
\add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.bin_s1  <= _100_;
always @(posedge \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.clk )
\add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.ain_s1  <= _099_;
always @(posedge \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.clk )
\add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.sum_s1  <= _102_;
always @(posedge \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.clk )
\add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.carry_s1  <= _101_;
assign _100_ = \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.ce  ? \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.b [1] : \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.bin_s1 ;
assign _099_ = \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.ce  ? \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.a [1] : \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.ain_s1 ;
assign _101_ = \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.ce  ? \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.facout_s1  : \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.carry_s1 ;
assign _102_ = \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.ce  ? \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.fas_s1  : \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.sum_s1 ;
assign _103_ = \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.a  + \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.b ;
assign { \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.cout , \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.s  } = _103_ + \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.cin ;
assign _104_ = \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.a  + \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.b ;
assign { \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.cout , \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.s  } = _104_ + \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.cin ;
always @(posedge \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.clk )
\add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.bin_s1  <= _106_;
always @(posedge \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.clk )
\add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.ain_s1  <= _105_;
always @(posedge \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.clk )
\add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.sum_s1  <= _108_;
always @(posedge \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.clk )
\add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.carry_s1  <= _107_;
assign _106_ = \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.ce  ? \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.b [31:16] : \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.bin_s1 ;
assign _105_ = \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.ce  ? \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.a [31:16] : \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.ain_s1 ;
assign _107_ = \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.ce  ? \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.facout_s1  : \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.carry_s1 ;
assign _108_ = \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.ce  ? \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.fas_s1  : \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.sum_s1 ;
assign _109_ = \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.u1.a  + \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.u1.b ;
assign { \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.u1.cout , \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.u1.s  } = _109_ + \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.u1.cin ;
assign _110_ = \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.u2.a  + \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.u2.b ;
assign { \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.u2.cout , \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.u2.s  } = _110_ + \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.u2.cin ;
always @(posedge \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.clk )
\add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.bin_s1  <= _112_;
always @(posedge \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.clk )
\add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.ain_s1  <= _111_;
always @(posedge \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.clk )
\add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.sum_s1  <= _114_;
always @(posedge \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.clk )
\add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.carry_s1  <= _113_;
assign _112_ = \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.ce  ? \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.b [33:17] : \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.bin_s1 ;
assign _111_ = \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.ce  ? \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.a [33:17] : \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.ain_s1 ;
assign _113_ = \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.ce  ? \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.facout_s1  : \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.carry_s1 ;
assign _114_ = \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.ce  ? \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.fas_s1  : \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.sum_s1 ;
assign _115_ = \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.u1.a  + \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.u1.b ;
assign { \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.u1.cout , \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.u1.s  } = _115_ + \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.u1.cin ;
assign _116_ = \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.u2.a  + \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.u2.b ;
assign { \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.u2.cout , \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.u2.s  } = _116_ + \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.u2.cin ;
always @(posedge \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.clk )
\add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.bin_s1  <= _118_;
always @(posedge \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.clk )
\add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.ain_s1  <= _117_;
always @(posedge \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.clk )
\add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.sum_s1  <= _120_;
always @(posedge \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.clk )
\add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.carry_s1  <= _119_;
assign _118_ = \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.ce  ? \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.b [4:2] : \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.bin_s1 ;
assign _117_ = \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.ce  ? \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.a [4:2] : \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.ain_s1 ;
assign _119_ = \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.ce  ? \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.facout_s1  : \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.carry_s1 ;
assign _120_ = \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.ce  ? \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.fas_s1  : \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.sum_s1 ;
assign _121_ = \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.u1.a  + \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.u1.b ;
assign { \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.u1.cout , \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.u1.s  } = _121_ + \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.u1.cin ;
assign _122_ = \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.u2.a  + \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.u2.b ;
assign { \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.u2.cout , \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.u2.s  } = _122_ + \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.u2.cin ;
always @(posedge \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.clk )
\add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.bin_s1  <= _124_;
always @(posedge \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.clk )
\add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.ain_s1  <= _123_;
always @(posedge \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.clk )
\add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.sum_s1  <= _126_;
always @(posedge \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.clk )
\add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.carry_s1  <= _125_;
assign _124_ = \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.ce  ? \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.b [4:2] : \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.bin_s1 ;
assign _123_ = \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.ce  ? \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.a [4:2] : \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.ain_s1 ;
assign _125_ = \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.ce  ? \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.facout_s1  : \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.carry_s1 ;
assign _126_ = \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.ce  ? \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.fas_s1  : \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.sum_s1 ;
assign _127_ = \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.u1.a  + \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.u1.b ;
assign { \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.u1.cout , \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.u1.s  } = _127_ + \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.u1.cin ;
assign _128_ = \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.u2.a  + \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.u2.b ;
assign { \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.u2.cout , \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.u2.s  } = _128_ + \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.u2.cin ;
always @(posedge \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.clk )
\add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.bin_s1  <= _130_;
always @(posedge \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.clk )
\add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.ain_s1  <= _129_;
always @(posedge \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.clk )
\add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.sum_s1  <= _132_;
always @(posedge \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.clk )
\add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.carry_s1  <= _131_;
assign _130_ = \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.ce  ? \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.b [4:2] : \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.bin_s1 ;
assign _129_ = \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.ce  ? \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.a [4:2] : \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.ain_s1 ;
assign _131_ = \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.ce  ? \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.facout_s1  : \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.carry_s1 ;
assign _132_ = \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.ce  ? \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.fas_s1  : \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.sum_s1 ;
assign _133_ = \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.u1.a  + \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.u1.b ;
assign { \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.u1.cout , \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.u1.s  } = _133_ + \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.u1.cin ;
assign _134_ = \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.u2.a  + \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.u2.b ;
assign { \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.u2.cout , \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.u2.s  } = _134_ + \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.u2.cin ;
always @(posedge \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.clk )
\add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.bin_s1  <= _136_;
always @(posedge \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.clk )
\add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.ain_s1  <= _135_;
always @(posedge \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.clk )
\add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.sum_s1  <= _138_;
always @(posedge \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.clk )
\add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.carry_s1  <= _137_;
assign _136_ = \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.ce  ? \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.b [4:2] : \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.bin_s1 ;
assign _135_ = \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.ce  ? \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.a [4:2] : \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.ain_s1 ;
assign _137_ = \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.ce  ? \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.facout_s1  : \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.carry_s1 ;
assign _138_ = \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.ce  ? \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.fas_s1  : \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.sum_s1 ;
assign _139_ = \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.u1.a  + \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.u1.b ;
assign { \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.u1.cout , \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.u1.s  } = _139_ + \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.u1.cin ;
assign _140_ = \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.u2.a  + \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.u2.b ;
assign { \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.u2.cout , \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.u2.s  } = _140_ + \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.u2.cin ;
always @(posedge \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.clk )
\add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.bin_s1  <= _142_;
always @(posedge \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.clk )
\add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.ain_s1  <= _141_;
always @(posedge \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.clk )
\add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.sum_s1  <= _144_;
always @(posedge \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.clk )
\add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.carry_s1  <= _143_;
assign _142_ = \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.ce  ? \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.b [5:3] : \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.bin_s1 ;
assign _141_ = \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.ce  ? \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.a [5:3] : \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.ain_s1 ;
assign _143_ = \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.ce  ? \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.facout_s1  : \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.carry_s1 ;
assign _144_ = \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.ce  ? \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.fas_s1  : \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.sum_s1 ;
assign _145_ = \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.u1.a  + \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.u1.b ;
assign { \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.u1.cout , \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.u1.s  } = _145_ + \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.u1.cin ;
assign _146_ = \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.u2.a  + \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.u2.b ;
assign { \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.u2.cout , \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.u2.s  } = _146_ + \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.u2.cin ;
always @(posedge \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.clk )
\add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.bin_s1  <= _148_;
always @(posedge \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.clk )
\add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.ain_s1  <= _147_;
always @(posedge \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.clk )
\add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.sum_s1  <= _150_;
always @(posedge \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.clk )
\add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.carry_s1  <= _149_;
assign _148_ = \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.ce  ? \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.b [7:4] : \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.bin_s1 ;
assign _147_ = \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.ce  ? \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.a [7:4] : \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.ain_s1 ;
assign _149_ = \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.ce  ? \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.facout_s1  : \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.carry_s1 ;
assign _150_ = \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.ce  ? \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.fas_s1  : \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.sum_s1 ;
assign _151_ = \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.u1.a  + \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.u1.b ;
assign { \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.u1.cout , \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.u1.s  } = _151_ + \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.u1.cin ;
assign _152_ = \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.u2.a  + \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.u2.b ;
assign { \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.u2.cout , \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.u2.s  } = _152_ + \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.u2.cin ;
always @(posedge \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.clk )
\add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.bin_s1  <= _154_;
always @(posedge \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.clk )
\add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.ain_s1  <= _153_;
always @(posedge \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.clk )
\add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.sum_s1  <= _156_;
always @(posedge \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.clk )
\add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.carry_s1  <= _155_;
assign _154_ = \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.ce  ? \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.b [8:4] : \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.bin_s1 ;
assign _153_ = \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.ce  ? \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.a [8:4] : \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.ain_s1 ;
assign _155_ = \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.ce  ? \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.facout_s1  : \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.carry_s1 ;
assign _156_ = \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.ce  ? \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.fas_s1  : \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.sum_s1 ;
assign _157_ = \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.u1.a  + \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.u1.b ;
assign { \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.u1.cout , \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.u1.s  } = _157_ + \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.u1.cin ;
assign _158_ = \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.u2.a  + \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.u2.b ;
assign { \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.u2.cout , \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.u2.s  } = _158_ + \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.u2.cin ;
always @(posedge \shl_32s_8ns_32_7_1_U3.clk )
\shl_32s_8ns_32_7_1_U3.dout_array[5]  <= _170_;
always @(posedge \shl_32s_8ns_32_7_1_U3.clk )
\shl_32s_8ns_32_7_1_U3.din1_cast_array[5]  <= _164_;
always @(posedge \shl_32s_8ns_32_7_1_U3.clk )
\shl_32s_8ns_32_7_1_U3.dout_array[4]  <= _169_;
always @(posedge \shl_32s_8ns_32_7_1_U3.clk )
\shl_32s_8ns_32_7_1_U3.din1_cast_array[4]  <= _163_;
always @(posedge \shl_32s_8ns_32_7_1_U3.clk )
\shl_32s_8ns_32_7_1_U3.dout_array[3]  <= _168_;
always @(posedge \shl_32s_8ns_32_7_1_U3.clk )
\shl_32s_8ns_32_7_1_U3.din1_cast_array[3]  <= _162_;
always @(posedge \shl_32s_8ns_32_7_1_U3.clk )
\shl_32s_8ns_32_7_1_U3.dout_array[2]  <= _167_;
always @(posedge \shl_32s_8ns_32_7_1_U3.clk )
\shl_32s_8ns_32_7_1_U3.din1_cast_array[2]  <= _161_;
always @(posedge \shl_32s_8ns_32_7_1_U3.clk )
\shl_32s_8ns_32_7_1_U3.dout_array[1]  <= _166_;
always @(posedge \shl_32s_8ns_32_7_1_U3.clk )
\shl_32s_8ns_32_7_1_U3.din1_cast_array[1]  <= _160_;
always @(posedge \shl_32s_8ns_32_7_1_U3.clk )
\shl_32s_8ns_32_7_1_U3.dout_array[0]  <= _165_;
always @(posedge \shl_32s_8ns_32_7_1_U3.clk )
\shl_32s_8ns_32_7_1_U3.din1_cast_array[0]  <= _159_;
assign _171_ = \shl_32s_8ns_32_7_1_U3.ce  ? \shl_32s_8ns_32_7_1_U3.din1_cast_array[4]  : \shl_32s_8ns_32_7_1_U3.din1_cast_array[5] ;
assign _164_ = \shl_32s_8ns_32_7_1_U3.reset  ? 8'h00 : _171_;
assign _172_ = \shl_32s_8ns_32_7_1_U3.ce  ? _185_ : \shl_32s_8ns_32_7_1_U3.dout_array[5] ;
assign _170_ = \shl_32s_8ns_32_7_1_U3.reset  ? 32'd0 : _172_;
assign _173_ = \shl_32s_8ns_32_7_1_U3.ce  ? \shl_32s_8ns_32_7_1_U3.din1_cast_array[3]  : \shl_32s_8ns_32_7_1_U3.din1_cast_array[4] ;
assign _163_ = \shl_32s_8ns_32_7_1_U3.reset  ? 8'h00 : _173_;
assign _174_ = \shl_32s_8ns_32_7_1_U3.ce  ? _184_ : \shl_32s_8ns_32_7_1_U3.dout_array[4] ;
assign _169_ = \shl_32s_8ns_32_7_1_U3.reset  ? 32'd0 : _174_;
assign _175_ = \shl_32s_8ns_32_7_1_U3.ce  ? \shl_32s_8ns_32_7_1_U3.din1_cast_array[2]  : \shl_32s_8ns_32_7_1_U3.din1_cast_array[3] ;
assign _162_ = \shl_32s_8ns_32_7_1_U3.reset  ? 8'h00 : _175_;
assign _176_ = \shl_32s_8ns_32_7_1_U3.ce  ? _183_ : \shl_32s_8ns_32_7_1_U3.dout_array[3] ;
assign _168_ = \shl_32s_8ns_32_7_1_U3.reset  ? 32'd0 : _176_;
assign _177_ = \shl_32s_8ns_32_7_1_U3.ce  ? \shl_32s_8ns_32_7_1_U3.din1_cast_array[1]  : \shl_32s_8ns_32_7_1_U3.din1_cast_array[2] ;
assign _161_ = \shl_32s_8ns_32_7_1_U3.reset  ? 8'h00 : _177_;
assign _178_ = \shl_32s_8ns_32_7_1_U3.ce  ? \shl_32s_8ns_32_7_1_U3.dout_array[1]  : \shl_32s_8ns_32_7_1_U3.dout_array[2] ;
assign _167_ = \shl_32s_8ns_32_7_1_U3.reset  ? 32'd0 : _178_;
assign _179_ = \shl_32s_8ns_32_7_1_U3.ce  ? \shl_32s_8ns_32_7_1_U3.din1_cast_array[0]  : \shl_32s_8ns_32_7_1_U3.din1_cast_array[1] ;
assign _160_ = \shl_32s_8ns_32_7_1_U3.reset  ? 8'h00 : _179_;
assign _180_ = \shl_32s_8ns_32_7_1_U3.ce  ? \shl_32s_8ns_32_7_1_U3.dout_array[0]  : \shl_32s_8ns_32_7_1_U3.dout_array[1] ;
assign _166_ = \shl_32s_8ns_32_7_1_U3.reset  ? 32'd0 : _180_;
assign _181_ = \shl_32s_8ns_32_7_1_U3.ce  ? \shl_32s_8ns_32_7_1_U3.din1 [7:0] : \shl_32s_8ns_32_7_1_U3.din1_cast_array[0] ;
assign _159_ = \shl_32s_8ns_32_7_1_U3.reset  ? 8'h00 : _181_;
assign _182_ = \shl_32s_8ns_32_7_1_U3.ce  ? \shl_32s_8ns_32_7_1_U3.din0  : \shl_32s_8ns_32_7_1_U3.dout_array[0] ;
assign _165_ = \shl_32s_8ns_32_7_1_U3.reset  ? 32'd0 : _182_;
assign _183_ = \shl_32s_8ns_32_7_1_U3.dout_array[2]  << { \shl_32s_8ns_32_7_1_U3.din1_cast_array[2] [7:6], 6'h00 };
assign _184_ = \shl_32s_8ns_32_7_1_U3.dout_array[3]  << { \shl_32s_8ns_32_7_1_U3.din1_cast_array[3] [5:4], 4'h0 };
assign _185_ = \shl_32s_8ns_32_7_1_U3.dout_array[4]  << { \shl_32s_8ns_32_7_1_U3.din1_cast_array[4] [3:2], 2'h0 };
assign \shl_32s_8ns_32_7_1_U3.dout  = \shl_32s_8ns_32_7_1_U3.dout_array[5]  << \shl_32s_8ns_32_7_1_U3.din1_cast_array[5] [1:0];
assign \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.bin_s0  = ~ \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.b ;
always @(posedge \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.clk )
\sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.bin_s1  <= _187_;
always @(posedge \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.clk )
\sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.ain_s1  <= _186_;
always @(posedge \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.clk )
\sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.sum_s1  <= _189_;
always @(posedge \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.clk )
\sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.carry_s1  <= _188_;
assign _187_ = \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.ce  ? \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.bin_s0 [1] : \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.bin_s1 ;
assign _186_ = \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.ce  ? \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.a [1] : \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.ain_s1 ;
assign _188_ = \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.ce  ? \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.facout_s1  : \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.carry_s1 ;
assign _189_ = \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.ce  ? \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.fas_s1  : \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.sum_s1 ;
assign _190_ = \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.u1.a  + \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.u1.b ;
assign { \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.u1.cout , \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.u1.s  } = _190_ + \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.u1.cin ;
assign _191_ = \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.u2.a  + \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.u2.b ;
assign { \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.u2.cout , \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.u2.s  } = _191_ + \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.u2.cin ;
assign \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.bin_s0  = ~ \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.b ;
always @(posedge \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.clk )
\sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.bin_s1  <= _193_;
always @(posedge \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.clk )
\sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.ain_s1  <= _192_;
always @(posedge \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.clk )
\sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.sum_s1  <= _195_;
always @(posedge \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.clk )
\sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.carry_s1  <= _194_;
assign _193_ = \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.ce  ? \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.bin_s0 [3:2] : \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.bin_s1 ;
assign _192_ = \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.ce  ? \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.a [3:2] : \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.ain_s1 ;
assign _194_ = \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.ce  ? \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.facout_s1  : \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.carry_s1 ;
assign _195_ = \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.ce  ? \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.fas_s1  : \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.sum_s1 ;
assign _196_ = \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.u1.a  + \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.u1.b ;
assign { \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.u1.cout , \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.u1.s  } = _196_ + \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.u1.cin ;
assign _197_ = \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.u2.a  + \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.u2.b ;
assign { \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.u2.cout , \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.u2.s  } = _197_ + \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.u2.cin ;
assign _198_ = | op_0[15:3];
assign _199_ = op_0[15:3] != 13'h1fff;
assign _200_ = | trunc_ln851_1_reg_924;
assign _201_ = | ret_V_21_reg_918;
assign _202_ = | trunc_ln851_2_reg_1027;
assign _203_ = | trunc_ln851_reg_913;
assign _204_ = | op_10[9:0];
assign or_ln340_fu_480_p2 = p_Result_7_reg_970 | overflow_fu_465_p2;
assign or_ln785_1_fu_515_p2 = xor_ln785_1_fu_510_p2 | p_Result_7_reg_970;
assign or_ln785_fu_449_p2 = p_Result_8_reg_977 | icmp_ln768_reg_984;
assign or_ln786_fu_475_p2 = xor_ln786_fu_470_p2 | icmp_ln786_reg_989;
assign ret_V_19_fu_290_p2 = op_3 | { op_2, 7'h00 };
always @(posedge ap_clk)
select_ln703_reg_857[6:0] <= 7'h00;
always @(posedge ap_clk)
ret_V_21_reg_918[6:0] <= 7'h00;
always @(posedge ap_clk)
trunc_ln851_1_reg_924 <= 7'h00;
always @(posedge ap_clk)
select_ln1192_reg_960[4:2] <= 3'h0;
always @(posedge ap_clk)
p_Val2_s_reg_1006[0] <= 1'h0;
always @(posedge ap_clk)
select_ln340_reg_1011[0] <= 1'h0;
always @(posedge ap_clk)
op_1_V_reg_1016[0] <= 1'h0;
always @(posedge ap_clk)
select_ln703_reg_857[8:7] <= _047_;
always @(posedge ap_clk)
select_ln1347_reg_1082 <= _042_;
always @(posedge ap_clk)
select_ln1347_1_reg_1087 <= _041_;
always @(posedge ap_clk)
sext_ln850_reg_1092 <= _049_;
always @(posedge ap_clk)
select_ln69_2_reg_1099 <= _045_;
always @(posedge ap_clk)
ret_V_2_reg_891 <= _037_;
always @(posedge ap_clk)
ret_V_25_reg_1072 <= _034_;
always @(posedge ap_clk)
tmp_reg_1077 <= _051_;
always @(posedge ap_clk)
ret_V_24_reg_1042 <= _033_;
always @(posedge ap_clk)
select_ln69_reg_1047 <= _046_;
always @(posedge ap_clk)
ret_V_22_reg_954 <= _032_;
always @(posedge ap_clk)
select_ln1192_reg_960[1:0] <= _040_;
always @(posedge ap_clk)
ret_V_27_reg_1249 <= _036_;
always @(posedge ap_clk)
ret_V_21_cast_reg_1254 <= _030_;
always @(posedge ap_clk)
sext_ln353_reg_902 <= _048_;
always @(posedge ap_clk)
ret_V_19_reg_907 <= _029_;
always @(posedge ap_clk)
trunc_ln851_reg_913 <= _054_;
always @(posedge ap_clk)
ret_V_21_reg_918[7] <= _031_;
always @(posedge ap_clk)
ret_V_18_reg_896 <= _028_;
always @(posedge ap_clk)
ret_V_17_reg_879 <= _027_;
always @(posedge ap_clk)
ret_V_reg_884 <= _038_;
always @(posedge ap_clk)
p_Val2_s_reg_1006[3:1] <= _025_;
always @(posedge ap_clk)
select_ln340_reg_1011[3:1] <= _043_;
always @(posedge ap_clk)
or_ln785_reg_1000 <= _022_;
always @(posedge ap_clk)
op_30_V_reg_1229 <= _021_;
always @(posedge ap_clk)
op_21_V_reg_1052 <= _020_;
always @(posedge ap_clk)
op_1_V_reg_1016[3:1] <= _019_;
always @(posedge ap_clk)
shl_ln1299_reg_1021 <= _050_;
always @(posedge ap_clk)
trunc_ln851_2_reg_1027 <= _053_;
always @(posedge ap_clk)
icmp_ln851_reg_874 <= _017_;
always @(posedge ap_clk)
icmp_ln851_1_reg_1067 <= _016_;
always @(posedge ap_clk)
icmp_ln850_3_reg_1032 <= _014_;
always @(posedge ap_clk)
icmp_ln850_reg_939 <= _015_;
always @(posedge ap_clk)
icmp_ln850_1_reg_944 <= _012_;
always @(posedge ap_clk)
icmp_ln850_2_reg_949 <= _013_;
always @(posedge ap_clk)
trunc_ln703_reg_965 <= _052_;
always @(posedge ap_clk)
p_Result_7_reg_970 <= _023_;
always @(posedge ap_clk)
p_Result_8_reg_977 <= _024_;
always @(posedge ap_clk)
icmp_ln768_reg_984 <= _010_;
always @(posedge ap_clk)
icmp_ln786_reg_989 <= _011_;
always @(posedge ap_clk)
r_reg_995 <= _026_;
always @(posedge ap_clk)
op_14_V_reg_1124 <= _018_;
always @(posedge ap_clk)
ret_reg_1129 <= _039_;
always @(posedge ap_clk)
ret_V_26_reg_1134 <= _035_;
always @(posedge ap_clk)
select_ln69_1_reg_1139 <= _044_;
always @(posedge ap_clk)
add_ln69_4_reg_1144 <= _005_;
always @(posedge ap_clk)
add_ln69_2_reg_1214 <= _003_;
always @(posedge ap_clk)
add_ln69_6_reg_1219 <= _007_;
always @(posedge ap_clk)
add_ln69_reg_1179 <= _008_;
always @(posedge ap_clk)
add_ln69_1_reg_1184 <= _002_;
always @(posedge ap_clk)
add_ln69_3_reg_1189 <= _004_;
always @(posedge ap_clk)
add_ln69_5_reg_1194 <= _006_;
always @(posedge ap_clk)
add_ln691_reg_1114 <= _001_;
always @(posedge ap_clk)
add_ln691_1_reg_1261 <= _000_;
always @(posedge ap_clk)
ap_CS_fsm <= _009_;
assign _055_ = _059_ ? 2'h2 : 2'h1;
assign _205_ = ap_CS_fsm == 1'h1;
function [32:0] _592_;
input [32:0] a;
input [1088:0] b;
input [32:0] s;
case (s)
33'b000000000000000000000000000000001:
_592_ = b[32:0];
33'b000000000000000000000000000000010:
_592_ = b[65:33];
33'b000000000000000000000000000000100:
_592_ = b[98:66];
33'b000000000000000000000000000001000:
_592_ = b[131:99];
33'b000000000000000000000000000010000:
_592_ = b[164:132];
33'b000000000000000000000000000100000:
_592_ = b[197:165];
33'b000000000000000000000000001000000:
_592_ = b[230:198];
33'b000000000000000000000000010000000:
_592_ = b[263:231];
33'b000000000000000000000000100000000:
_592_ = b[296:264];
33'b000000000000000000000001000000000:
_592_ = b[329:297];
33'b000000000000000000000010000000000:
_592_ = b[362:330];
33'b000000000000000000000100000000000:
_592_ = b[395:363];
33'b000000000000000000001000000000000:
_592_ = b[428:396];
33'b000000000000000000010000000000000:
_592_ = b[461:429];
33'b000000000000000000100000000000000:
_592_ = b[494:462];
33'b000000000000000001000000000000000:
_592_ = b[527:495];
33'b000000000000000010000000000000000:
_592_ = b[560:528];
33'b000000000000000100000000000000000:
_592_ = b[593:561];
33'b000000000000001000000000000000000:
_592_ = b[626:594];
33'b000000000000010000000000000000000:
_592_ = b[659:627];
33'b000000000000100000000000000000000:
_592_ = b[692:660];
33'b000000000001000000000000000000000:
_592_ = b[725:693];
33'b000000000010000000000000000000000:
_592_ = b[758:726];
33'b000000000100000000000000000000000:
_592_ = b[791:759];
33'b000000001000000000000000000000000:
_592_ = b[824:792];
33'b000000010000000000000000000000000:
_592_ = b[857:825];
33'b000000100000000000000000000000000:
_592_ = b[890:858];
33'b000001000000000000000000000000000:
_592_ = b[923:891];
33'b000010000000000000000000000000000:
_592_ = b[956:924];
33'b000100000000000000000000000000000:
_592_ = b[989:957];
33'b001000000000000000000000000000000:
_592_ = b[1022:990];
33'b010000000000000000000000000000000:
_592_ = b[1055:1023];
33'b100000000000000000000000000000000:
_592_ = b[1088:1056];
33'b000000000000000000000000000000000:
_592_ = a;
default:
_592_ = 33'bx;
endcase
endfunction
assign ap_NS_fsm = _592_(33'hxxxxxxxxx, { 31'h00000000, _055_, 1056'h000000020000000200000002000000020000000200000002000000020000000200000002000000020000000200000002000000020000000200000002000000020000000200000002000000020000000200000002000000020000000200000002000000020000000200000002000000020000000200000002000000020000000000000001 }, { _205_, _237_, _236_, _235_, _234_, _233_, _232_, _231_, _230_, _229_, _228_, _227_, _226_, _225_, _224_, _223_, _222_, _221_, _220_, _219_, _218_, _217_, _216_, _215_, _214_, _213_, _212_, _211_, _210_, _209_, _208_, _207_, _206_ });
assign _206_ = ap_CS_fsm == 33'h100000000;
assign _207_ = ap_CS_fsm == 32'd2147483648;
assign _208_ = ap_CS_fsm == 31'h40000000;
assign _209_ = ap_CS_fsm == 30'h20000000;
assign _210_ = ap_CS_fsm == 29'h10000000;
assign _211_ = ap_CS_fsm == 28'h8000000;
assign _212_ = ap_CS_fsm == 27'h4000000;
assign _213_ = ap_CS_fsm == 26'h2000000;
assign _214_ = ap_CS_fsm == 25'h1000000;
assign _215_ = ap_CS_fsm == 24'h800000;
assign _216_ = ap_CS_fsm == 23'h400000;
assign _217_ = ap_CS_fsm == 22'h200000;
assign _218_ = ap_CS_fsm == 21'h100000;
assign _219_ = ap_CS_fsm == 20'h80000;
assign _220_ = ap_CS_fsm == 19'h40000;
assign _221_ = ap_CS_fsm == 18'h20000;
assign _222_ = ap_CS_fsm == 17'h10000;
assign _223_ = ap_CS_fsm == 16'h8000;
assign _224_ = ap_CS_fsm == 15'h4000;
assign _225_ = ap_CS_fsm == 14'h2000;
assign _226_ = ap_CS_fsm == 13'h1000;
assign _227_ = ap_CS_fsm == 12'h800;
assign _228_ = ap_CS_fsm == 11'h400;
assign _229_ = ap_CS_fsm == 10'h200;
assign _230_ = ap_CS_fsm == 9'h100;
assign _231_ = ap_CS_fsm == 8'h80;
assign _232_ = ap_CS_fsm == 7'h40;
assign _233_ = ap_CS_fsm == 6'h20;
assign _234_ = ap_CS_fsm == 5'h10;
assign _235_ = ap_CS_fsm == 4'h8;
assign _236_ = ap_CS_fsm == 3'h4;
assign _237_ = ap_CS_fsm == 2'h2;
assign op_31_ap_vld = ap_CS_fsm[32] ? 1'h1 : 1'h0;
assign ap_idle = _058_ ? 1'h1 : 1'h0;
assign _047_ = ap_CS_fsm[0] ? select_ln703_fu_219_p3[8:7] : select_ln703_reg_857[8:7];
assign _045_ = ap_CS_fsm[19] ? select_ln69_2_fu_655_p3 : select_ln69_2_reg_1099;
assign _049_ = ap_CS_fsm[19] ? { tmp_reg_1077[6], tmp_reg_1077 } : sext_ln850_reg_1092;
assign _041_ = ap_CS_fsm[19] ? select_ln1347_1_fu_639_p3 : select_ln1347_1_reg_1087;
assign _042_ = ap_CS_fsm[19] ? select_ln1347_fu_632_p3 : select_ln1347_reg_1082;
assign _037_ = _057_ ? grp_fu_256_p2 : ret_V_2_reg_891;
assign _051_ = ap_CS_fsm[18] ? grp_fu_606_p2[16:10] : tmp_reg_1077;
assign _034_ = ap_CS_fsm[18] ? grp_fu_606_p2 : ret_V_25_reg_1072;
assign _046_ = ap_CS_fsm[14] ? select_ln69_fu_579_p3 : select_ln69_reg_1047;
assign _033_ = ap_CS_fsm[14] ? grp_fu_549_p2 : ret_V_24_reg_1042;
assign _040_ = ap_CS_fsm[8] ? select_ln1192_fu_378_p3 : select_ln1192_reg_960[1:0];
assign _032_ = ap_CS_fsm[8] ? ret_V_22_fu_372_p2 : ret_V_22_reg_954;
assign _030_ = ap_CS_fsm[29] ? grp_fu_806_p2[32:1] : ret_V_21_cast_reg_1254;
assign _036_ = ap_CS_fsm[29] ? grp_fu_806_p2 : ret_V_27_reg_1249;
assign _031_ = ap_CS_fsm[6] ? ret_V_21_fu_299_p2[7] : ret_V_21_reg_918[7];
assign _054_ = ap_CS_fsm[6] ? ret_V_19_fu_290_p2[6:0] : trunc_ln851_reg_913;
assign _029_ = ap_CS_fsm[6] ? ret_V_19_fu_290_p2 : ret_V_19_reg_907;
assign _048_ = ap_CS_fsm[6] ? { ret_V_18_reg_896[1], ret_V_18_reg_896[1], ret_V_18_reg_896[1], ret_V_18_reg_896[1], ret_V_18_reg_896[1], ret_V_18_reg_896[1], ret_V_18_reg_896 } : sext_ln353_reg_902;
assign _028_ = ap_CS_fsm[5] ? ret_V_18_fu_273_p3 : ret_V_18_reg_896;
assign _038_ = ap_CS_fsm[2] ? grp_fu_235_p2[8:7] : ret_V_reg_884;
assign _027_ = ap_CS_fsm[2] ? grp_fu_235_p2 : ret_V_17_reg_879;
assign _043_ = ap_CS_fsm[11] ? select_ln340_fu_497_p3[3:1] : select_ln340_reg_1011[3:1];
assign _025_ = ap_CS_fsm[11] ? trunc_ln703_reg_965 : p_Val2_s_reg_1006[3:1];
assign _022_ = ap_CS_fsm[10] ? or_ln785_fu_449_p2 : or_ln785_reg_1000;
assign _021_ = ap_CS_fsm[27] ? grp_fu_786_p2 : op_30_V_reg_1229;
assign _020_ = ap_CS_fsm[16] ? grp_fu_587_p2 : op_21_V_reg_1052;
assign _053_ = ap_CS_fsm[12] ? grp_fu_315_p2[6:0] : trunc_ln851_2_reg_1027;
assign _050_ = ap_CS_fsm[12] ? grp_fu_315_p2 : shl_ln1299_reg_1021;
assign _019_ = ap_CS_fsm[12] ? op_1_V_fu_531_p3[3:1] : op_1_V_reg_1016[3:1];
assign _017_ = ap_CS_fsm[1] ? icmp_ln851_fu_240_p2 : icmp_ln851_reg_874;
assign _016_ = ap_CS_fsm[17] ? icmp_ln851_1_fu_616_p2 : icmp_ln851_1_reg_1067;
assign _014_ = ap_CS_fsm[13] ? icmp_ln850_3_fu_541_p2 : icmp_ln850_3_reg_1032;
assign _013_ = ap_CS_fsm[7] ? icmp_ln850_2_fu_331_p2 : icmp_ln850_2_reg_949;
assign _012_ = ap_CS_fsm[7] ? icmp_ln850_1_fu_326_p2 : icmp_ln850_1_reg_944;
assign _015_ = ap_CS_fsm[7] ? icmp_ln850_fu_321_p2 : icmp_ln850_reg_939;
assign _026_ = ap_CS_fsm[9] ? r_fu_443_p3 : r_reg_995;
assign _011_ = ap_CS_fsm[9] ? icmp_ln786_fu_422_p2 : icmp_ln786_reg_989;
assign _010_ = ap_CS_fsm[9] ? icmp_ln768_fu_416_p2 : icmp_ln768_reg_984;
assign _024_ = ap_CS_fsm[9] ? op_0[2] : p_Result_8_reg_977;
assign _023_ = ap_CS_fsm[9] ? op_0[15] : p_Result_7_reg_970;
assign _052_ = ap_CS_fsm[9] ? op_0[2:0] : trunc_ln703_reg_965;
assign _005_ = ap_CS_fsm[21] ? grp_fu_685_p2 : add_ln69_4_reg_1144;
assign _044_ = ap_CS_fsm[21] ? select_ln69_1_fu_709_p3 : select_ln69_1_reg_1139;
assign _035_ = ap_CS_fsm[21] ? ret_V_26_fu_702_p3 : ret_V_26_reg_1134;
assign _039_ = ap_CS_fsm[21] ? grp_fu_677_p2 : ret_reg_1129;
assign _018_ = ap_CS_fsm[21] ? grp_fu_671_p2 : op_14_V_reg_1124;
assign _007_ = ap_CS_fsm[25] ? grp_fu_777_p2 : add_ln69_6_reg_1219;
assign _003_ = ap_CS_fsm[25] ? grp_fu_766_p2 : add_ln69_2_reg_1214;
assign _006_ = ap_CS_fsm[23] ? grp_fu_759_p2 : add_ln69_5_reg_1194;
assign _004_ = ap_CS_fsm[23] ? grp_fu_753_p2 : add_ln69_3_reg_1189;
assign _002_ = ap_CS_fsm[23] ? grp_fu_747_p2 : add_ln69_1_reg_1184;
assign _008_ = ap_CS_fsm[23] ? grp_fu_741_p2 : add_ln69_reg_1179;
assign _001_ = _056_ ? grp_fu_649_p2 : add_ln691_reg_1114;
assign _000_ = ap_CS_fsm[31] ? grp_fu_822_p2 : add_ln691_1_reg_1261;
assign _009_ = ap_rst ? 33'h000000001 : ap_NS_fsm;
assign icmp_ln768_fu_416_p2 = _198_ ? 1'h1 : 1'h0;
assign icmp_ln786_fu_422_p2 = _199_ ? 1'h1 : 1'h0;
assign icmp_ln850_1_fu_326_p2 = _200_ ? 1'h1 : 1'h0;
assign icmp_ln850_2_fu_331_p2 = _201_ ? 1'h1 : 1'h0;
assign icmp_ln850_3_fu_541_p2 = _202_ ? 1'h1 : 1'h0;
assign icmp_ln850_fu_321_p2 = _203_ ? 1'h1 : 1'h0;
assign icmp_ln851_1_fu_616_p2 = _204_ ? 1'h1 : 1'h0;
assign icmp_ln851_fu_240_p2 = _062_ ? 1'h1 : 1'h0;
assign op_1_V_fu_531_p3 = and_ln785_1_fu_526_p2 ? p_Val2_s_reg_1006 : select_ln340_reg_1011;
assign op_31 = ret_V_27_reg_1249[33] ? select_ln850_2_fu_837_p3 : ret_V_21_cast_reg_1254;
assign r_fu_443_p3 = ret_V_22_reg_954 ? { 1'h0, select_ln850_4_fu_435_p3 } : sext_ln353_reg_902;
assign ret_V_18_fu_273_p3 = ret_V_17_reg_879[8] ? select_ln850_fu_268_p3 : ret_V_reg_884;
assign ret_V_26_fu_702_p3 = ret_V_25_reg_1072[16] ? select_ln850_1_fu_697_p3 : sext_ln850_reg_1092;
assign select_ln1192_fu_378_p3 = ret_V_20_fu_355_p2 ? 2'h3 : 2'h0;
assign select_ln1347_1_fu_639_p3 = ret_V_22_reg_954 ? 2'h3 : 2'h0;
assign select_ln1347_fu_632_p3 = op_2 ? 2'h3 : 2'h0;
assign select_ln340_fu_497_p3 = and_ln340_fu_491_p2 ? { trunc_ln703_reg_965, 1'h0 } : 4'h0;
assign select_ln69_1_fu_709_p3 = op_11 ? 2'h3 : 2'h0;
assign select_ln69_2_fu_655_p3 = op_18 ? 2'h3 : 2'h0;
assign select_ln69_fu_579_p3 = ret_V_23_fu_573_p2 ? 5'h1f : 5'h00;
assign select_ln703_fu_219_p3 = op_2 ? 9'h180 : 9'h000;
assign select_ln850_1_fu_697_p3 = icmp_ln851_1_reg_1067 ? add_ln691_reg_1114 : sext_ln850_reg_1092;
assign select_ln850_2_fu_837_p3 = op_19[0] ? add_ln691_1_reg_1261 : ret_V_21_cast_reg_1254;
assign select_ln850_4_fu_435_p3 = ret_V_18_reg_896[1] ? 7'h7f : 7'h00;
assign select_ln850_fu_268_p3 = icmp_ln851_reg_874 ? ret_V_reg_884 : ret_V_2_reg_891;
assign ret_V_20_fu_355_p2 = ret_V_19_reg_907[7] ^ and_ln850_fu_350_p2;
assign ret_V_22_fu_372_p2 = ret_V_21_reg_918[7] ^ and_ln850_1_fu_368_p2;
assign ret_V_23_fu_573_p2 = shl_ln1299_reg_1021[7] ^ and_ln850_2_fu_568_p2;
assign ap_CS_fsm_state1 = ap_CS_fsm[0];
assign ap_CS_fsm_state10 = ap_CS_fsm[9];
assign ap_CS_fsm_state11 = ap_CS_fsm[10];
assign ap_CS_fsm_state12 = ap_CS_fsm[11];
assign ap_CS_fsm_state13 = ap_CS_fsm[12];
assign ap_CS_fsm_state14 = ap_CS_fsm[13];
assign ap_CS_fsm_state15 = ap_CS_fsm[14];
assign ap_CS_fsm_state16 = ap_CS_fsm[15];
assign ap_CS_fsm_state17 = ap_CS_fsm[16];
assign ap_CS_fsm_state18 = ap_CS_fsm[17];
assign ap_CS_fsm_state19 = ap_CS_fsm[18];
assign ap_CS_fsm_state2 = ap_CS_fsm[1];
assign ap_CS_fsm_state20 = ap_CS_fsm[19];
assign ap_CS_fsm_state21 = ap_CS_fsm[20];
assign ap_CS_fsm_state22 = ap_CS_fsm[21];
assign ap_CS_fsm_state23 = ap_CS_fsm[22];
assign ap_CS_fsm_state24 = ap_CS_fsm[23];
assign ap_CS_fsm_state25 = ap_CS_fsm[24];
assign ap_CS_fsm_state26 = ap_CS_fsm[25];
assign ap_CS_fsm_state27 = ap_CS_fsm[26];
assign ap_CS_fsm_state28 = ap_CS_fsm[27];
assign ap_CS_fsm_state29 = ap_CS_fsm[28];
assign ap_CS_fsm_state3 = ap_CS_fsm[2];
assign ap_CS_fsm_state30 = ap_CS_fsm[29];
assign ap_CS_fsm_state31 = ap_CS_fsm[30];
assign ap_CS_fsm_state32 = ap_CS_fsm[31];
assign ap_CS_fsm_state33 = ap_CS_fsm[32];
assign ap_CS_fsm_state4 = ap_CS_fsm[3];
assign ap_CS_fsm_state5 = ap_CS_fsm[4];
assign ap_CS_fsm_state6 = ap_CS_fsm[5];
assign ap_CS_fsm_state7 = ap_CS_fsm[6];
assign ap_CS_fsm_state8 = ap_CS_fsm[7];
assign ap_CS_fsm_state9 = ap_CS_fsm[8];
assign ap_done = op_31_ap_vld;
assign ap_ready = op_31_ap_vld;
assign grp_fu_235_p1 = { op_3[7], op_3 };
assign grp_fu_315_p0 = { op_3[7], op_3[7], op_3[7], op_3[7], op_3[7], op_3[7], op_3[7], op_3[7], op_3[7], op_3[7], op_3[7], op_3[7], op_3[7], op_3[7], op_3[7], op_3[7], op_3[7], op_3[7], op_3[7], op_3[7], op_3[7], op_3[7], op_3[7], op_3[7], op_3 };
assign grp_fu_315_p1 = { 24'h000000, ret_V_18_reg_896[1], ret_V_18_reg_896[1], ret_V_18_reg_896[1], ret_V_18_reg_896[1], ret_V_18_reg_896[1], ret_V_18_reg_896[1], ret_V_18_reg_896 };
assign grp_fu_549_p1 = { op_1_V_reg_1016[3], op_1_V_reg_1016 };
assign grp_fu_606_p0 = { op_21_V_reg_1052[4], op_21_V_reg_1052[4], op_21_V_reg_1052, 10'h000 };
assign grp_fu_606_p1 = { op_10[15], op_10 };
assign grp_fu_649_p0 = { tmp_reg_1077[6], tmp_reg_1077 };
assign grp_fu_671_p0 = { op_6[1], op_6[1], op_6 };
assign grp_fu_671_p1 = op_7[3:0];
assign grp_fu_685_p1 = { 1'h0, op_12 };
assign grp_fu_741_p0 = { ret_V_26_reg_1134[7], ret_V_26_reg_1134[7], ret_V_26_reg_1134 };
assign grp_fu_741_p1 = { 2'h0, r_reg_995 };
assign grp_fu_747_p0 = { op_14_V_reg_1124[3], op_14_V_reg_1124 };
assign grp_fu_747_p1 = { op_16[3], op_16 };
assign grp_fu_753_p0 = { 1'h0, ret_reg_1129[1], ret_reg_1129[1], ret_reg_1129 };
assign grp_fu_753_p1 = { 3'h0, op_17 };
assign grp_fu_766_p0 = { add_ln69_1_reg_1184[4], add_ln69_1_reg_1184[4], add_ln69_1_reg_1184[4], add_ln69_1_reg_1184[4], add_ln69_1_reg_1184[4], add_ln69_1_reg_1184 };
assign grp_fu_777_p0 = { add_ln69_5_reg_1194[1], add_ln69_5_reg_1194[1], add_ln69_5_reg_1194[1], add_ln69_5_reg_1194[1], add_ln69_5_reg_1194 };
assign grp_fu_777_p1 = { 1'h0, add_ln69_3_reg_1189 };
assign grp_fu_786_p0 = { add_ln69_6_reg_1219[5], add_ln69_6_reg_1219[5], add_ln69_6_reg_1219[5], add_ln69_6_reg_1219[5], add_ln69_6_reg_1219 };
assign grp_fu_806_p0 = { op_30_V_reg_1229[9], op_30_V_reg_1229[9], op_30_V_reg_1229[9], op_30_V_reg_1229[9], op_30_V_reg_1229[9], op_30_V_reg_1229[9], op_30_V_reg_1229[9], op_30_V_reg_1229[9], op_30_V_reg_1229[9], op_30_V_reg_1229[9], op_30_V_reg_1229[9], op_30_V_reg_1229[9], op_30_V_reg_1229[9], op_30_V_reg_1229[9], op_30_V_reg_1229[9], op_30_V_reg_1229[9], op_30_V_reg_1229[9], op_30_V_reg_1229[9], op_30_V_reg_1229[9], op_30_V_reg_1229[9], op_30_V_reg_1229[9], op_30_V_reg_1229[9], op_30_V_reg_1229[9], op_30_V_reg_1229, 1'h0 };
assign grp_fu_806_p1 = { op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19 };
assign lhs_fu_283_p3 = { op_2, 7'h00 };
assign p_Result_1_fu_343_p3 = ret_V_19_reg_907[7];
assign p_Result_2_fu_561_p3 = shl_ln1299_reg_1021[7];
assign p_Result_5_fu_690_p3 = ret_V_25_reg_1072[16];
assign p_Result_6_fu_827_p3 = ret_V_27_reg_1249[33];
assign p_Result_s_12_fu_261_p3 = ret_V_17_reg_879[8];
assign p_Result_s_fu_406_p4 = op_0[15:3];
assign p_Val2_s_fu_453_p3 = { trunc_ln703_reg_965, 1'h0 };
assign ret_V_10_fu_554_p3 = shl_ln1299_reg_1021[7];
assign ret_V_19_fu_290_p1 = op_3;
assign ret_V_21_fu_299_p1 = op_3;
assign ret_V_5_fu_336_p3 = ret_V_19_reg_907[7];
assign ret_V_8_fu_361_p3 = ret_V_21_reg_918[7];
assign rhs_2_fu_595_p3 = { op_21_V_reg_1052, 10'h000 };
assign sext_ln1192_fu_591_p0 = op_10;
assign sext_ln1299_fu_312_p0 = op_3;
assign sext_ln353_fu_280_p1 = { ret_V_18_reg_896[1], ret_V_18_reg_896[1], ret_V_18_reg_896[1], ret_V_18_reg_896[1], ret_V_18_reg_896[1], ret_V_18_reg_896[1], ret_V_18_reg_896 };
assign sext_ln69_1_fu_720_p1 = { ret_reg_1129[1], ret_reg_1129[1], ret_reg_1129 };
assign sext_ln703_2_fu_791_p0 = op_19;
assign sext_ln703_fu_227_p0 = op_3;
assign sext_ln850_fu_646_p1 = { tmp_reg_1077[6], tmp_reg_1077 };
assign tmp_11_fu_795_p3 = { op_30_V_reg_1229, 1'h0 };
assign tmp_9_fu_428_p3 = ret_V_18_reg_896[1];
assign trunc_ln1192_fu_231_p0 = op_3;
assign trunc_ln1192_fu_231_p1 = op_3[6:0];
assign trunc_ln703_fu_386_p1 = op_0[2:0];
assign trunc_ln851_1_fu_304_p1 = ret_V_21_fu_299_p2[6:0];
assign trunc_ln851_2_fu_537_p1 = grp_fu_315_p2[6:0];
assign trunc_ln851_3_fu_612_p0 = op_10;
assign trunc_ln851_3_fu_612_p1 = op_10[9:0];
assign trunc_ln851_4_fu_834_p0 = op_19;
assign trunc_ln851_4_fu_834_p1 = op_19[0];
assign trunc_ln851_fu_295_p1 = ret_V_19_fu_290_p2[6:0];
assign \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.ain_s0  = \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.a ;
assign \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.s  = { \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.fas_s2 , \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.sum_s1  };
assign \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.u2.a  = \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.ain_s1 ;
assign \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.u2.b  = \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.bin_s1 ;
assign \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.u2.cin  = \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.carry_s1 ;
assign \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.facout_s2  = \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.u2.cout ;
assign \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.fas_s2  = \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.u2.s ;
assign \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.u1.a  = \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.a [1:0];
assign \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.u1.b  = \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.bin_s0 [1:0];
assign \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.u1.cin  = 1'h1;
assign \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.facout_s1  = \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.u1.cout ;
assign \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.fas_s1  = \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.u1.s ;
assign \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.a  = \sub_4s_4ns_4_2_1_U8.din0 ;
assign \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.b  = \sub_4s_4ns_4_2_1_U8.din1 ;
assign \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.ce  = \sub_4s_4ns_4_2_1_U8.ce ;
assign \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.clk  = \sub_4s_4ns_4_2_1_U8.clk ;
assign \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.reset  = \sub_4s_4ns_4_2_1_U8.reset ;
assign \sub_4s_4ns_4_2_1_U8.dout  = \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.s ;
assign \sub_4s_4ns_4_2_1_U8.ce  = 1'h1;
assign \sub_4s_4ns_4_2_1_U8.clk  = ap_clk;
assign \sub_4s_4ns_4_2_1_U8.din0  = { op_6[1], op_6[1], op_6 };
assign \sub_4s_4ns_4_2_1_U8.din1  = op_7[3:0];
assign grp_fu_671_p2 = \sub_4s_4ns_4_2_1_U8.dout ;
assign \sub_4s_4ns_4_2_1_U8.reset  = ap_rst;
assign \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.ain_s0  = \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.a ;
assign \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.s  = { \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.fas_s2 , \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.sum_s1  };
assign \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.u2.a  = \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.ain_s1 ;
assign \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.u2.b  = \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.bin_s1 ;
assign \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.u2.cin  = \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.carry_s1 ;
assign \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.facout_s2  = \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.u2.cout ;
assign \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.fas_s2  = \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.u2.s ;
assign \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.u1.a  = \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.a [0];
assign \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.u1.b  = \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.bin_s0 [0];
assign \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.u1.cin  = 1'h1;
assign \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.facout_s1  = \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.u1.cout ;
assign \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.fas_s1  = \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.u1.s ;
assign \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.a  = \sub_2ns_2ns_2_2_1_U9.din0 ;
assign \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.b  = \sub_2ns_2ns_2_2_1_U9.din1 ;
assign \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.ce  = \sub_2ns_2ns_2_2_1_U9.ce ;
assign \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.clk  = \sub_2ns_2ns_2_2_1_U9.clk ;
assign \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.reset  = \sub_2ns_2ns_2_2_1_U9.reset ;
assign \sub_2ns_2ns_2_2_1_U9.dout  = \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.s ;
assign \sub_2ns_2ns_2_2_1_U9.ce  = 1'h1;
assign \sub_2ns_2ns_2_2_1_U9.clk  = ap_clk;
assign \sub_2ns_2ns_2_2_1_U9.din0  = select_ln1347_reg_1082;
assign \sub_2ns_2ns_2_2_1_U9.din1  = select_ln1347_1_reg_1087;
assign grp_fu_677_p2 = \sub_2ns_2ns_2_2_1_U9.dout ;
assign \sub_2ns_2ns_2_2_1_U9.reset  = ap_rst;
assign \shl_32s_8ns_32_7_1_U3.din1_cast  = \shl_32s_8ns_32_7_1_U3.din1 [7:0];
assign \shl_32s_8ns_32_7_1_U3.din1_mask  = 8'h03;
assign \shl_32s_8ns_32_7_1_U3.ce  = 1'h1;
assign \shl_32s_8ns_32_7_1_U3.clk  = ap_clk;
assign \shl_32s_8ns_32_7_1_U3.din0  = { op_3[7], op_3[7], op_3[7], op_3[7], op_3[7], op_3[7], op_3[7], op_3[7], op_3[7], op_3[7], op_3[7], op_3[7], op_3[7], op_3[7], op_3[7], op_3[7], op_3[7], op_3[7], op_3[7], op_3[7], op_3[7], op_3[7], op_3[7], op_3[7], op_3 };
assign \shl_32s_8ns_32_7_1_U3.din1  = { 24'h000000, ret_V_18_reg_896[1], ret_V_18_reg_896[1], ret_V_18_reg_896[1], ret_V_18_reg_896[1], ret_V_18_reg_896[1], ret_V_18_reg_896[1], ret_V_18_reg_896 };
assign grp_fu_315_p2 = \shl_32s_8ns_32_7_1_U3.dout ;
assign \shl_32s_8ns_32_7_1_U3.reset  = ap_rst;
assign \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.ain_s0  = \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.a ;
assign \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.bin_s0  = \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.b ;
assign \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.s  = { \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.fas_s2 , \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.sum_s1  };
assign \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.u2.a  = \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.ain_s1 ;
assign \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.u2.b  = \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.bin_s1 ;
assign \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.u2.cin  = \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.carry_s1 ;
assign \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.facout_s2  = \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.u2.cout ;
assign \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.fas_s2  = \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.u2.s ;
assign \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.u1.a  = \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.a [3:0];
assign \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.u1.b  = \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.b [3:0];
assign \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.u1.cin  = 1'h0;
assign \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.facout_s1  = \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.u1.cout ;
assign \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.fas_s1  = \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.u1.s ;
assign \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.a  = \add_9ns_9s_9_2_1_U1.din0 ;
assign \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.b  = \add_9ns_9s_9_2_1_U1.din1 ;
assign \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.ce  = \add_9ns_9s_9_2_1_U1.ce ;
assign \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.clk  = \add_9ns_9s_9_2_1_U1.clk ;
assign \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.reset  = \add_9ns_9s_9_2_1_U1.reset ;
assign \add_9ns_9s_9_2_1_U1.dout  = \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.s ;
assign \add_9ns_9s_9_2_1_U1.ce  = 1'h1;
assign \add_9ns_9s_9_2_1_U1.clk  = ap_clk;
assign \add_9ns_9s_9_2_1_U1.din0  = select_ln703_reg_857;
assign \add_9ns_9s_9_2_1_U1.din1  = { op_3[7], op_3 };
assign grp_fu_235_p2 = \add_9ns_9s_9_2_1_U1.dout ;
assign \add_9ns_9s_9_2_1_U1.reset  = ap_rst;
assign \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.ain_s0  = \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.a ;
assign \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.bin_s0  = \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.b ;
assign \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.s  = { \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.fas_s2 , \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.sum_s1  };
assign \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.u2.a  = \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.ain_s1 ;
assign \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.u2.b  = \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.bin_s1 ;
assign \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.u2.cin  = \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.carry_s1 ;
assign \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.facout_s2  = \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.u2.cout ;
assign \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.fas_s2  = \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.u2.s ;
assign \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.u1.a  = \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.a [3:0];
assign \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.u1.b  = \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.b [3:0];
assign \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.u1.cin  = 1'h0;
assign \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.facout_s1  = \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.u1.cout ;
assign \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.fas_s1  = \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.u1.s ;
assign \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.a  = \add_8s_8ns_8_2_1_U7.din0 ;
assign \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.b  = \add_8s_8ns_8_2_1_U7.din1 ;
assign \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.ce  = \add_8s_8ns_8_2_1_U7.ce ;
assign \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.clk  = \add_8s_8ns_8_2_1_U7.clk ;
assign \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.reset  = \add_8s_8ns_8_2_1_U7.reset ;
assign \add_8s_8ns_8_2_1_U7.dout  = \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.s ;
assign \add_8s_8ns_8_2_1_U7.ce  = 1'h1;
assign \add_8s_8ns_8_2_1_U7.clk  = ap_clk;
assign \add_8s_8ns_8_2_1_U7.din0  = { tmp_reg_1077[6], tmp_reg_1077 };
assign \add_8s_8ns_8_2_1_U7.din1  = 8'h01;
assign grp_fu_649_p2 = \add_8s_8ns_8_2_1_U7.dout ;
assign \add_8s_8ns_8_2_1_U7.reset  = ap_rst;
assign \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.ain_s0  = \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.a ;
assign \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.bin_s0  = \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.b ;
assign \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.s  = { \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.fas_s2 , \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.sum_s1  };
assign \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.u2.a  = \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.ain_s1 ;
assign \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.u2.b  = \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.bin_s1 ;
assign \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.u2.cin  = \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.carry_s1 ;
assign \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.facout_s2  = \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.u2.cout ;
assign \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.fas_s2  = \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.u2.s ;
assign \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.u1.a  = \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.a [2:0];
assign \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.u1.b  = \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.b [2:0];
assign \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.u1.cin  = 1'h0;
assign \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.facout_s1  = \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.u1.cout ;
assign \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.fas_s1  = \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.u1.s ;
assign \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.a  = \add_6s_6ns_6_2_1_U16.din0 ;
assign \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.b  = \add_6s_6ns_6_2_1_U16.din1 ;
assign \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.ce  = \add_6s_6ns_6_2_1_U16.ce ;
assign \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.clk  = \add_6s_6ns_6_2_1_U16.clk ;
assign \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.reset  = \add_6s_6ns_6_2_1_U16.reset ;
assign \add_6s_6ns_6_2_1_U16.dout  = \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.s ;
assign \add_6s_6ns_6_2_1_U16.ce  = 1'h1;
assign \add_6s_6ns_6_2_1_U16.clk  = ap_clk;
assign \add_6s_6ns_6_2_1_U16.din0  = { add_ln69_5_reg_1194[1], add_ln69_5_reg_1194[1], add_ln69_5_reg_1194[1], add_ln69_5_reg_1194[1], add_ln69_5_reg_1194 };
assign \add_6s_6ns_6_2_1_U16.din1  = { 1'h0, add_ln69_3_reg_1189 };
assign grp_fu_777_p2 = \add_6s_6ns_6_2_1_U16.dout ;
assign \add_6s_6ns_6_2_1_U16.reset  = ap_rst;
assign \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.ain_s0  = \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.a ;
assign \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.bin_s0  = \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.b ;
assign \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.s  = { \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.fas_s2 , \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.sum_s1  };
assign \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.u2.a  = \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.ain_s1 ;
assign \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.u2.b  = \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.bin_s1 ;
assign \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.u2.cin  = \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.carry_s1 ;
assign \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.facout_s2  = \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.u2.cout ;
assign \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.fas_s2  = \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.u2.s ;
assign \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.u1.a  = \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.a [1:0];
assign \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.u1.b  = \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.b [1:0];
assign \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.u1.cin  = 1'h0;
assign \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.facout_s1  = \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.u1.cout ;
assign \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.fas_s1  = \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.u1.s ;
assign \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.a  = \add_5s_5s_5_2_1_U12.din0 ;
assign \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.b  = \add_5s_5s_5_2_1_U12.din1 ;
assign \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.ce  = \add_5s_5s_5_2_1_U12.ce ;
assign \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.clk  = \add_5s_5s_5_2_1_U12.clk ;
assign \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.reset  = \add_5s_5s_5_2_1_U12.reset ;
assign \add_5s_5s_5_2_1_U12.dout  = \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.s ;
assign \add_5s_5s_5_2_1_U12.ce  = 1'h1;
assign \add_5s_5s_5_2_1_U12.clk  = ap_clk;
assign \add_5s_5s_5_2_1_U12.din0  = { op_14_V_reg_1124[3], op_14_V_reg_1124 };
assign \add_5s_5s_5_2_1_U12.din1  = { op_16[3], op_16 };
assign grp_fu_747_p2 = \add_5s_5s_5_2_1_U12.dout ;
assign \add_5s_5s_5_2_1_U12.reset  = ap_rst;
assign \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.ain_s0  = \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.a ;
assign \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.bin_s0  = \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.b ;
assign \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.s  = { \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.fas_s2 , \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.sum_s1  };
assign \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.u2.a  = \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.ain_s1 ;
assign \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.u2.b  = \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.bin_s1 ;
assign \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.u2.cin  = \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.carry_s1 ;
assign \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.facout_s2  = \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.u2.cout ;
assign \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.fas_s2  = \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.u2.s ;
assign \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.u1.a  = \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.a [1:0];
assign \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.u1.b  = \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.b [1:0];
assign \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.u1.cin  = 1'h0;
assign \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.facout_s1  = \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.u1.cout ;
assign \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.fas_s1  = \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.u1.s ;
assign \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.a  = \add_5ns_5s_5_2_1_U4.din0 ;
assign \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.b  = \add_5ns_5s_5_2_1_U4.din1 ;
assign \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.ce  = \add_5ns_5s_5_2_1_U4.ce ;
assign \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.clk  = \add_5ns_5s_5_2_1_U4.clk ;
assign \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.reset  = \add_5ns_5s_5_2_1_U4.reset ;
assign \add_5ns_5s_5_2_1_U4.dout  = \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.s ;
assign \add_5ns_5s_5_2_1_U4.ce  = 1'h1;
assign \add_5ns_5s_5_2_1_U4.clk  = ap_clk;
assign \add_5ns_5s_5_2_1_U4.din0  = select_ln1192_reg_960;
assign \add_5ns_5s_5_2_1_U4.din1  = { op_1_V_reg_1016[3], op_1_V_reg_1016 };
assign grp_fu_549_p2 = \add_5ns_5s_5_2_1_U4.dout ;
assign \add_5ns_5s_5_2_1_U4.reset  = ap_rst;
assign \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.ain_s0  = \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.a ;
assign \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.bin_s0  = \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.b ;
assign \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.s  = { \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.fas_s2 , \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.sum_s1  };
assign \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.u2.a  = \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.ain_s1 ;
assign \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.u2.b  = \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.bin_s1 ;
assign \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.u2.cin  = \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.carry_s1 ;
assign \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.facout_s2  = \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.u2.cout ;
assign \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.fas_s2  = \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.u2.s ;
assign \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.u1.a  = \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.a [1:0];
assign \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.u1.b  = \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.b [1:0];
assign \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.u1.cin  = 1'h0;
assign \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.facout_s1  = \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.u1.cout ;
assign \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.fas_s1  = \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.u1.s ;
assign \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.a  = \add_5ns_5ns_5_2_1_U5.din0 ;
assign \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.b  = \add_5ns_5ns_5_2_1_U5.din1 ;
assign \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.ce  = \add_5ns_5ns_5_2_1_U5.ce ;
assign \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.clk  = \add_5ns_5ns_5_2_1_U5.clk ;
assign \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.reset  = \add_5ns_5ns_5_2_1_U5.reset ;
assign \add_5ns_5ns_5_2_1_U5.dout  = \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.s ;
assign \add_5ns_5ns_5_2_1_U5.ce  = 1'h1;
assign \add_5ns_5ns_5_2_1_U5.clk  = ap_clk;
assign \add_5ns_5ns_5_2_1_U5.din0  = ret_V_24_reg_1042;
assign \add_5ns_5ns_5_2_1_U5.din1  = select_ln69_reg_1047;
assign grp_fu_587_p2 = \add_5ns_5ns_5_2_1_U5.dout ;
assign \add_5ns_5ns_5_2_1_U5.reset  = ap_rst;
assign \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.ain_s0  = \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.a ;
assign \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.bin_s0  = \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.b ;
assign \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.s  = { \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.fas_s2 , \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.sum_s1  };
assign \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.u2.a  = \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.ain_s1 ;
assign \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.u2.b  = \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.bin_s1 ;
assign \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.u2.cin  = \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.carry_s1 ;
assign \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.facout_s2  = \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.u2.cout ;
assign \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.fas_s2  = \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.u2.s ;
assign \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.u1.a  = \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.a [1:0];
assign \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.u1.b  = \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.b [1:0];
assign \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.u1.cin  = 1'h0;
assign \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.facout_s1  = \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.u1.cout ;
assign \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.fas_s1  = \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.u1.s ;
assign \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.a  = \add_5ns_5ns_5_2_1_U13.din0 ;
assign \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.b  = \add_5ns_5ns_5_2_1_U13.din1 ;
assign \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.ce  = \add_5ns_5ns_5_2_1_U13.ce ;
assign \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.clk  = \add_5ns_5ns_5_2_1_U13.clk ;
assign \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.reset  = \add_5ns_5ns_5_2_1_U13.reset ;
assign \add_5ns_5ns_5_2_1_U13.dout  = \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.s ;
assign \add_5ns_5ns_5_2_1_U13.ce  = 1'h1;
assign \add_5ns_5ns_5_2_1_U13.clk  = ap_clk;
assign \add_5ns_5ns_5_2_1_U13.din0  = { 1'h0, ret_reg_1129[1], ret_reg_1129[1], ret_reg_1129 };
assign \add_5ns_5ns_5_2_1_U13.din1  = { 3'h0, op_17 };
assign grp_fu_753_p2 = \add_5ns_5ns_5_2_1_U13.dout ;
assign \add_5ns_5ns_5_2_1_U13.reset  = ap_rst;
assign \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.ain_s0  = \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.a ;
assign \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.bin_s0  = \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.b ;
assign \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.s  = { \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.fas_s2 , \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.sum_s1  };
assign \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.u2.a  = \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.ain_s1 ;
assign \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.u2.b  = \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.bin_s1 ;
assign \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.u2.cin  = \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.carry_s1 ;
assign \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.facout_s2  = \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.u2.cout ;
assign \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.fas_s2  = \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.u2.s ;
assign \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.u1.a  = \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.a [16:0];
assign \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.u1.b  = \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.b [16:0];
assign \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.u1.cin  = 1'h0;
assign \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.facout_s1  = \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.u1.cout ;
assign \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.fas_s1  = \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.u1.s ;
assign \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.a  = \add_34s_34s_34_2_1_U18.din0 ;
assign \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.b  = \add_34s_34s_34_2_1_U18.din1 ;
assign \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.ce  = \add_34s_34s_34_2_1_U18.ce ;
assign \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.clk  = \add_34s_34s_34_2_1_U18.clk ;
assign \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.reset  = \add_34s_34s_34_2_1_U18.reset ;
assign \add_34s_34s_34_2_1_U18.dout  = \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.s ;
assign \add_34s_34s_34_2_1_U18.ce  = 1'h1;
assign \add_34s_34s_34_2_1_U18.clk  = ap_clk;
assign \add_34s_34s_34_2_1_U18.din0  = { op_30_V_reg_1229[9], op_30_V_reg_1229[9], op_30_V_reg_1229[9], op_30_V_reg_1229[9], op_30_V_reg_1229[9], op_30_V_reg_1229[9], op_30_V_reg_1229[9], op_30_V_reg_1229[9], op_30_V_reg_1229[9], op_30_V_reg_1229[9], op_30_V_reg_1229[9], op_30_V_reg_1229[9], op_30_V_reg_1229[9], op_30_V_reg_1229[9], op_30_V_reg_1229[9], op_30_V_reg_1229[9], op_30_V_reg_1229[9], op_30_V_reg_1229[9], op_30_V_reg_1229[9], op_30_V_reg_1229[9], op_30_V_reg_1229[9], op_30_V_reg_1229[9], op_30_V_reg_1229[9], op_30_V_reg_1229, 1'h0 };
assign \add_34s_34s_34_2_1_U18.din1  = { op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19 };
assign grp_fu_806_p2 = \add_34s_34s_34_2_1_U18.dout ;
assign \add_34s_34s_34_2_1_U18.reset  = ap_rst;
assign \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.ain_s0  = \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.a ;
assign \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.bin_s0  = \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.b ;
assign \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.s  = { \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.fas_s2 , \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.sum_s1  };
assign \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.u2.a  = \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.ain_s1 ;
assign \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.u2.b  = \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.bin_s1 ;
assign \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.u2.cin  = \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.carry_s1 ;
assign \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.facout_s2  = \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.u2.cout ;
assign \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.fas_s2  = \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.u2.s ;
assign \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.u1.a  = \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.a [15:0];
assign \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.u1.b  = \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.b [15:0];
assign \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.u1.cin  = 1'h0;
assign \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.facout_s1  = \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.u1.cout ;
assign \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.fas_s1  = \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.u1.s ;
assign \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.a  = \add_32ns_32ns_32_2_1_U19.din0 ;
assign \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.b  = \add_32ns_32ns_32_2_1_U19.din1 ;
assign \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.ce  = \add_32ns_32ns_32_2_1_U19.ce ;
assign \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.clk  = \add_32ns_32ns_32_2_1_U19.clk ;
assign \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.reset  = \add_32ns_32ns_32_2_1_U19.reset ;
assign \add_32ns_32ns_32_2_1_U19.dout  = \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.s ;
assign \add_32ns_32ns_32_2_1_U19.ce  = 1'h1;
assign \add_32ns_32ns_32_2_1_U19.clk  = ap_clk;
assign \add_32ns_32ns_32_2_1_U19.din0  = ret_V_21_cast_reg_1254;
assign \add_32ns_32ns_32_2_1_U19.din1  = 32'd1;
assign grp_fu_822_p2 = \add_32ns_32ns_32_2_1_U19.dout ;
assign \add_32ns_32ns_32_2_1_U19.reset  = ap_rst;
assign \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.ain_s0  = \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.a ;
assign \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.bin_s0  = \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.b ;
assign \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.s  = { \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.fas_s2 , \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.sum_s1  };
assign \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.a  = \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.ain_s1 ;
assign \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.b  = \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.bin_s1 ;
assign \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.cin  = \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.carry_s1 ;
assign \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.facout_s2  = \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.cout ;
assign \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.fas_s2  = \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.s ;
assign \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.a  = \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.a [0];
assign \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.b  = \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.b [0];
assign \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.cin  = 1'h0;
assign \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.facout_s1  = \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.cout ;
assign \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.fas_s1  = \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.s ;
assign \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.a  = \add_2ns_2ns_2_2_1_U2.din0 ;
assign \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.b  = \add_2ns_2ns_2_2_1_U2.din1 ;
assign \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.ce  = \add_2ns_2ns_2_2_1_U2.ce ;
assign \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.clk  = \add_2ns_2ns_2_2_1_U2.clk ;
assign \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.reset  = \add_2ns_2ns_2_2_1_U2.reset ;
assign \add_2ns_2ns_2_2_1_U2.dout  = \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.s ;
assign \add_2ns_2ns_2_2_1_U2.ce  = 1'h1;
assign \add_2ns_2ns_2_2_1_U2.clk  = ap_clk;
assign \add_2ns_2ns_2_2_1_U2.din0  = ret_V_reg_884;
assign \add_2ns_2ns_2_2_1_U2.din1  = 2'h1;
assign grp_fu_256_p2 = \add_2ns_2ns_2_2_1_U2.dout ;
assign \add_2ns_2ns_2_2_1_U2.reset  = ap_rst;
assign \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.ain_s0  = \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.a ;
assign \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.bin_s0  = \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.b ;
assign \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.s  = { \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.fas_s2 , \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.sum_s1  };
assign \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.a  = \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.ain_s1 ;
assign \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.b  = \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.bin_s1 ;
assign \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.cin  = \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.carry_s1 ;
assign \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.facout_s2  = \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.cout ;
assign \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.fas_s2  = \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.s ;
assign \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.a  = \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.a [0];
assign \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.b  = \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.b [0];
assign \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.cin  = 1'h0;
assign \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.facout_s1  = \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.cout ;
assign \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.fas_s1  = \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.s ;
assign \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.a  = \add_2ns_2ns_2_2_1_U14.din0 ;
assign \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.b  = \add_2ns_2ns_2_2_1_U14.din1 ;
assign \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.ce  = \add_2ns_2ns_2_2_1_U14.ce ;
assign \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.clk  = \add_2ns_2ns_2_2_1_U14.clk ;
assign \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.reset  = \add_2ns_2ns_2_2_1_U14.reset ;
assign \add_2ns_2ns_2_2_1_U14.dout  = \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.s ;
assign \add_2ns_2ns_2_2_1_U14.ce  = 1'h1;
assign \add_2ns_2ns_2_2_1_U14.clk  = ap_clk;
assign \add_2ns_2ns_2_2_1_U14.din0  = add_ln69_4_reg_1144;
assign \add_2ns_2ns_2_2_1_U14.din1  = select_ln69_1_reg_1139;
assign grp_fu_759_p2 = \add_2ns_2ns_2_2_1_U14.dout ;
assign \add_2ns_2ns_2_2_1_U14.reset  = ap_rst;
assign \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.ain_s0  = \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.a ;
assign \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.bin_s0  = \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.b ;
assign \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.s  = { \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.fas_s2 , \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.sum_s1  };
assign \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.a  = \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.ain_s1 ;
assign \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.b  = \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.bin_s1 ;
assign \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.cin  = \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.carry_s1 ;
assign \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.facout_s2  = \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.cout ;
assign \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.fas_s2  = \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.s ;
assign \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.a  = \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.a [0];
assign \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.b  = \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.b [0];
assign \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.cin  = 1'h0;
assign \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.facout_s1  = \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.cout ;
assign \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.fas_s1  = \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.s ;
assign \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.a  = \add_2ns_2ns_2_2_1_U10.din0 ;
assign \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.b  = \add_2ns_2ns_2_2_1_U10.din1 ;
assign \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.ce  = \add_2ns_2ns_2_2_1_U10.ce ;
assign \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.clk  = \add_2ns_2ns_2_2_1_U10.clk ;
assign \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.reset  = \add_2ns_2ns_2_2_1_U10.reset ;
assign \add_2ns_2ns_2_2_1_U10.dout  = \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.s ;
assign \add_2ns_2ns_2_2_1_U10.ce  = 1'h1;
assign \add_2ns_2ns_2_2_1_U10.clk  = ap_clk;
assign \add_2ns_2ns_2_2_1_U10.din0  = select_ln69_2_reg_1099;
assign \add_2ns_2ns_2_2_1_U10.din1  = { 1'h0, op_12 };
assign grp_fu_685_p2 = \add_2ns_2ns_2_2_1_U10.dout ;
assign \add_2ns_2ns_2_2_1_U10.reset  = ap_rst;
assign \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.ain_s0  = \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.a ;
assign \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.bin_s0  = \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.b ;
assign \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.s  = { \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.fas_s2 , \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.sum_s1  };
assign \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.u2.a  = \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.ain_s1 ;
assign \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.u2.b  = \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.bin_s1 ;
assign \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.u2.cin  = \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.carry_s1 ;
assign \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.facout_s2  = \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.u2.cout ;
assign \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.fas_s2  = \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.u2.s ;
assign \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.u1.a  = \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.a [7:0];
assign \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.u1.b  = \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.b [7:0];
assign \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.u1.cin  = 1'h0;
assign \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.facout_s1  = \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.u1.cout ;
assign \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.fas_s1  = \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.u1.s ;
assign \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.a  = \add_17s_17s_17_2_1_U6.din0 ;
assign \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.b  = \add_17s_17s_17_2_1_U6.din1 ;
assign \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.ce  = \add_17s_17s_17_2_1_U6.ce ;
assign \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.clk  = \add_17s_17s_17_2_1_U6.clk ;
assign \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.reset  = \add_17s_17s_17_2_1_U6.reset ;
assign \add_17s_17s_17_2_1_U6.dout  = \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.s ;
assign \add_17s_17s_17_2_1_U6.ce  = 1'h1;
assign \add_17s_17s_17_2_1_U6.clk  = ap_clk;
assign \add_17s_17s_17_2_1_U6.din0  = { op_21_V_reg_1052[4], op_21_V_reg_1052[4], op_21_V_reg_1052, 10'h000 };
assign \add_17s_17s_17_2_1_U6.din1  = { op_10[15], op_10 };
assign grp_fu_606_p2 = \add_17s_17s_17_2_1_U6.dout ;
assign \add_17s_17s_17_2_1_U6.reset  = ap_rst;
assign \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.ain_s0  = \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.a ;
assign \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.bin_s0  = \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.b ;
assign \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.s  = { \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.fas_s2 , \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.sum_s1  };
assign \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.u2.a  = \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.ain_s1 ;
assign \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.u2.b  = \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.bin_s1 ;
assign \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.u2.cin  = \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.carry_s1 ;
assign \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.facout_s2  = \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.u2.cout ;
assign \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.fas_s2  = \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.u2.s ;
assign \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.u1.a  = \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.a [4:0];
assign \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.u1.b  = \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.b [4:0];
assign \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.u1.cin  = 1'h0;
assign \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.facout_s1  = \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.u1.cout ;
assign \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.fas_s1  = \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.u1.s ;
assign \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.a  = \add_10s_10ns_10_2_1_U17.din0 ;
assign \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.b  = \add_10s_10ns_10_2_1_U17.din1 ;
assign \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.ce  = \add_10s_10ns_10_2_1_U17.ce ;
assign \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.clk  = \add_10s_10ns_10_2_1_U17.clk ;
assign \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.reset  = \add_10s_10ns_10_2_1_U17.reset ;
assign \add_10s_10ns_10_2_1_U17.dout  = \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.s ;
assign \add_10s_10ns_10_2_1_U17.ce  = 1'h1;
assign \add_10s_10ns_10_2_1_U17.clk  = ap_clk;
assign \add_10s_10ns_10_2_1_U17.din0  = { add_ln69_6_reg_1219[5], add_ln69_6_reg_1219[5], add_ln69_6_reg_1219[5], add_ln69_6_reg_1219[5], add_ln69_6_reg_1219 };
assign \add_10s_10ns_10_2_1_U17.din1  = add_ln69_2_reg_1214;
assign grp_fu_786_p2 = \add_10s_10ns_10_2_1_U17.dout ;
assign \add_10s_10ns_10_2_1_U17.reset  = ap_rst;
assign \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.ain_s0  = \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.a ;
assign \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.bin_s0  = \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.b ;
assign \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.s  = { \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.fas_s2 , \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.sum_s1  };
assign \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.u2.a  = \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.ain_s1 ;
assign \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.u2.b  = \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.bin_s1 ;
assign \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.u2.cin  = \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.carry_s1 ;
assign \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.facout_s2  = \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.u2.cout ;
assign \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.fas_s2  = \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.u2.s ;
assign \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.u1.a  = \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.a [4:0];
assign \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.u1.b  = \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.b [4:0];
assign \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.u1.cin  = 1'h0;
assign \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.facout_s1  = \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.u1.cout ;
assign \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.fas_s1  = \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.u1.s ;
assign \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.a  = \add_10s_10ns_10_2_1_U15.din0 ;
assign \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.b  = \add_10s_10ns_10_2_1_U15.din1 ;
assign \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.ce  = \add_10s_10ns_10_2_1_U15.ce ;
assign \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.clk  = \add_10s_10ns_10_2_1_U15.clk ;
assign \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.reset  = \add_10s_10ns_10_2_1_U15.reset ;
assign \add_10s_10ns_10_2_1_U15.dout  = \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.s ;
assign \add_10s_10ns_10_2_1_U15.ce  = 1'h1;
assign \add_10s_10ns_10_2_1_U15.clk  = ap_clk;
assign \add_10s_10ns_10_2_1_U15.din0  = { add_ln69_1_reg_1184[4], add_ln69_1_reg_1184[4], add_ln69_1_reg_1184[4], add_ln69_1_reg_1184[4], add_ln69_1_reg_1184[4], add_ln69_1_reg_1184 };
assign \add_10s_10ns_10_2_1_U15.din1  = add_ln69_reg_1179;
assign grp_fu_766_p2 = \add_10s_10ns_10_2_1_U15.dout ;
assign \add_10s_10ns_10_2_1_U15.reset  = ap_rst;
assign \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.ain_s0  = \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.a ;
assign \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.bin_s0  = \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.b ;
assign \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.s  = { \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.fas_s2 , \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.sum_s1  };
assign \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.u2.a  = \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.ain_s1 ;
assign \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.u2.b  = \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.bin_s1 ;
assign \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.u2.cin  = \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.carry_s1 ;
assign \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.facout_s2  = \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.u2.cout ;
assign \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.fas_s2  = \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.u2.s ;
assign \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.u1.a  = \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.a [4:0];
assign \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.u1.b  = \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.b [4:0];
assign \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.u1.cin  = 1'h0;
assign \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.facout_s1  = \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.u1.cout ;
assign \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.fas_s1  = \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.u1.s ;
assign \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.a  = \add_10s_10ns_10_2_1_U11.din0 ;
assign \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.b  = \add_10s_10ns_10_2_1_U11.din1 ;
assign \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.ce  = \add_10s_10ns_10_2_1_U11.ce ;
assign \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.clk  = \add_10s_10ns_10_2_1_U11.clk ;
assign \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.reset  = \add_10s_10ns_10_2_1_U11.reset ;
assign \add_10s_10ns_10_2_1_U11.dout  = \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.s ;
assign \add_10s_10ns_10_2_1_U11.ce  = 1'h1;
assign \add_10s_10ns_10_2_1_U11.clk  = ap_clk;
assign \add_10s_10ns_10_2_1_U11.din0  = { ret_V_26_reg_1134[7], ret_V_26_reg_1134[7], ret_V_26_reg_1134 };
assign \add_10s_10ns_10_2_1_U11.din1  = { 2'h0, r_reg_995 };
assign grp_fu_741_p2 = \add_10s_10ns_10_2_1_U11.dout ;
assign \add_10s_10ns_10_2_1_U11.reset  = ap_rst;
endmodule


// Machine B:
// Processed by function `add_clk_enable_signal` in `verilog_tricks.py`.
// Processed by function `remove_reset_signal` in `verilog_tricks.py`.
module top_B (
  ap_clk,
  ap_start,
  ap_done,
  ap_idle,
  ap_ready,
  op_0,
  op_2,
  op_3,
  op_6,
  op_7,
  op_10,
  op_11,
  op_12,
  op_16,
  op_17,
  op_18,
  op_19,
  op_31,
  op_31_ap_vld,
clk_enable
);
input clk_enable;


input ap_clk;
wire ap_rst;
assign ap_rst = op_31_ap_vld;
input ap_start;
input [15:0] op_0;
input [15:0] op_10;
input op_11;
input op_12;
input [3:0] op_16;
input [1:0] op_17;
input op_18;
input [3:0] op_19;
input op_2;
input [7:0] op_3;
input [1:0] op_6;
input [31:0] op_7;
output ap_done;
output ap_idle;
output ap_ready;
output [31:0] op_31;
output op_31_ap_vld;


reg [4:0] \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.ain_s1 ;
reg [4:0] \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.bin_s1 ;
reg \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.carry_s1 ;
reg [4:0] \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.sum_s1 ;
reg [4:0] \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.ain_s1 ;
reg [4:0] \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.bin_s1 ;
reg \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.carry_s1 ;
reg [4:0] \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.sum_s1 ;
reg [4:0] \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.ain_s1 ;
reg [4:0] \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.bin_s1 ;
reg \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.carry_s1 ;
reg [4:0] \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.sum_s1 ;
reg [8:0] \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.ain_s1 ;
reg [8:0] \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.bin_s1 ;
reg \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.carry_s1 ;
reg [7:0] \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.sum_s1 ;
reg \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.ain_s1 ;
reg \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.bin_s1 ;
reg \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.carry_s1 ;
reg \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.sum_s1 ;
reg \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.ain_s1 ;
reg \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.bin_s1 ;
reg \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.carry_s1 ;
reg \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.sum_s1 ;
reg \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.ain_s1 ;
reg \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.bin_s1 ;
reg \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.carry_s1 ;
reg \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.sum_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.ain_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.bin_s1 ;
reg \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.carry_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.sum_s1 ;
reg [16:0] \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.ain_s1 ;
reg [16:0] \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.bin_s1 ;
reg \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.carry_s1 ;
reg [16:0] \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.sum_s1 ;
reg [2:0] \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.ain_s1 ;
reg [2:0] \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.bin_s1 ;
reg \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.carry_s1 ;
reg [1:0] \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.sum_s1 ;
reg [2:0] \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.ain_s1 ;
reg [2:0] \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.bin_s1 ;
reg \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.carry_s1 ;
reg [1:0] \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.sum_s1 ;
reg [2:0] \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.ain_s1 ;
reg [2:0] \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.bin_s1 ;
reg \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.carry_s1 ;
reg [1:0] \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.sum_s1 ;
reg [2:0] \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.ain_s1 ;
reg [2:0] \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.bin_s1 ;
reg \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.carry_s1 ;
reg [1:0] \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.sum_s1 ;
reg [2:0] \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.ain_s1 ;
reg [2:0] \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.bin_s1 ;
reg \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.carry_s1 ;
reg [2:0] \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.sum_s1 ;
reg [3:0] \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.ain_s1 ;
reg [3:0] \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.bin_s1 ;
reg \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.carry_s1 ;
reg [3:0] \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.sum_s1 ;
reg [4:0] \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.ain_s1 ;
reg [4:0] \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.bin_s1 ;
reg \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.carry_s1 ;
reg [3:0] \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.sum_s1 ;
reg [31:0] add_ln691_1_reg_1261;
reg [7:0] add_ln691_reg_1114;
reg [4:0] add_ln69_1_reg_1184;
reg [9:0] add_ln69_2_reg_1214;
reg [4:0] add_ln69_3_reg_1189;
reg [1:0] add_ln69_4_reg_1144;
reg [1:0] add_ln69_5_reg_1194;
reg [5:0] add_ln69_6_reg_1219;
reg [9:0] add_ln69_reg_1179;
reg [32:0] ap_CS_fsm = 33'h000000001;
reg icmp_ln768_reg_984;
reg icmp_ln786_reg_989;
reg icmp_ln850_1_reg_944;
reg icmp_ln850_2_reg_949;
reg icmp_ln850_3_reg_1032;
reg icmp_ln850_reg_939;
reg icmp_ln851_1_reg_1067;
reg icmp_ln851_reg_874;
reg [3:0] op_14_V_reg_1124;
reg [3:0] op_1_V_reg_1016;
reg [4:0] op_21_V_reg_1052;
reg [9:0] op_30_V_reg_1229;
reg or_ln785_reg_1000;
reg p_Result_7_reg_970;
reg p_Result_8_reg_977;
reg [3:0] p_Val2_s_reg_1006;
reg [7:0] r_reg_995;
reg [8:0] ret_V_17_reg_879;
reg [1:0] ret_V_18_reg_896;
reg [7:0] ret_V_19_reg_907;
reg [31:0] ret_V_21_cast_reg_1254;
reg [7:0] ret_V_21_reg_918;
reg ret_V_22_reg_954;
reg [4:0] ret_V_24_reg_1042;
reg [16:0] ret_V_25_reg_1072;
reg [7:0] ret_V_26_reg_1134;
reg [33:0] ret_V_27_reg_1249;
reg [1:0] ret_V_2_reg_891;
reg [1:0] ret_V_reg_884;
reg [1:0] ret_reg_1129;
reg [4:0] select_ln1192_reg_960;
reg [1:0] select_ln1347_1_reg_1087;
reg [1:0] select_ln1347_reg_1082;
reg [3:0] select_ln340_reg_1011;
reg [1:0] select_ln69_1_reg_1139;
reg [1:0] select_ln69_2_reg_1099;
reg [4:0] select_ln69_reg_1047;
reg [8:0] select_ln703_reg_857;
reg [7:0] sext_ln353_reg_902;
reg [7:0] sext_ln850_reg_1092;
reg [7:0] \shl_32s_8ns_32_7_1_U3.din1_cast_array[0] ;
reg [7:0] \shl_32s_8ns_32_7_1_U3.din1_cast_array[1] ;
reg [7:0] \shl_32s_8ns_32_7_1_U3.din1_cast_array[2] ;
reg [7:0] \shl_32s_8ns_32_7_1_U3.din1_cast_array[3] ;
reg [7:0] \shl_32s_8ns_32_7_1_U3.din1_cast_array[4] ;
reg [7:0] \shl_32s_8ns_32_7_1_U3.din1_cast_array[5] ;
reg [31:0] \shl_32s_8ns_32_7_1_U3.dout_array[0] ;
reg [31:0] \shl_32s_8ns_32_7_1_U3.dout_array[1] ;
reg [31:0] \shl_32s_8ns_32_7_1_U3.dout_array[2] ;
reg [31:0] \shl_32s_8ns_32_7_1_U3.dout_array[3] ;
reg [31:0] \shl_32s_8ns_32_7_1_U3.dout_array[4] ;
reg [31:0] \shl_32s_8ns_32_7_1_U3.dout_array[5] ;
reg [31:0] shl_ln1299_reg_1021;
reg \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.ain_s1 ;
reg \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.bin_s1 ;
reg \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.carry_s1 ;
reg \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.sum_s1 ;
reg [1:0] \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.ain_s1 ;
reg [1:0] \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.bin_s1 ;
reg \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.carry_s1 ;
reg [1:0] \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.sum_s1 ;
reg [6:0] tmp_reg_1077;
reg [2:0] trunc_ln703_reg_965;
reg [6:0] trunc_ln851_1_reg_924;
reg [6:0] trunc_ln851_2_reg_1027;
reg [6:0] trunc_ln851_reg_913;
wire [31:0] _000_;
wire [7:0] _001_;
wire [4:0] _002_;
wire [9:0] _003_;
wire [4:0] _004_;
wire [1:0] _005_;
wire [1:0] _006_;
wire [5:0] _007_;
wire [9:0] _008_;
wire [32:0] _009_;
wire _010_;
wire _011_;
wire _012_;
wire _013_;
wire _014_;
wire _015_;
wire _016_;
wire _017_;
wire [3:0] _018_;
wire [2:0] _019_;
wire [4:0] _020_;
wire [9:0] _021_;
wire _022_;
wire _023_;
wire _024_;
wire [2:0] _025_;
wire [7:0] _026_;
wire [8:0] _027_;
wire [1:0] _028_;
wire [7:0] _029_;
wire [31:0] _030_;
wire _031_;
wire _032_;
wire [4:0] _033_;
wire [16:0] _034_;
wire [7:0] _035_;
wire [33:0] _036_;
wire [1:0] _037_;
wire [1:0] _038_;
wire [1:0] _039_;
wire [1:0] _040_;
wire [1:0] _041_;
wire [1:0] _042_;
wire [2:0] _043_;
wire [1:0] _044_;
wire [1:0] _045_;
wire [4:0] _046_;
wire [1:0] _047_;
wire [7:0] _048_;
wire [7:0] _049_;
wire [31:0] _050_;
wire [6:0] _051_;
wire [2:0] _052_;
wire [6:0] _053_;
wire [6:0] _054_;
wire [1:0] _055_;
wire _056_;
wire _057_;
wire _058_;
wire _059_;
wire _060_;
wire _061_;
wire _062_;
wire [4:0] _063_;
wire [4:0] _064_;
wire _065_;
wire [4:0] _066_;
wire [5:0] _067_;
wire [5:0] _068_;
wire [4:0] _069_;
wire [4:0] _070_;
wire _071_;
wire [4:0] _072_;
wire [5:0] _073_;
wire [5:0] _074_;
wire [4:0] _075_;
wire [4:0] _076_;
wire _077_;
wire [4:0] _078_;
wire [5:0] _079_;
wire [5:0] _080_;
wire [8:0] _081_;
wire [8:0] _082_;
wire _083_;
wire [7:0] _084_;
wire [8:0] _085_;
wire [9:0] _086_;
wire _087_;
wire _088_;
wire _089_;
wire _090_;
wire [1:0] _091_;
wire [1:0] _092_;
wire _093_;
wire _094_;
wire _095_;
wire _096_;
wire [1:0] _097_;
wire [1:0] _098_;
wire _099_;
wire _100_;
wire _101_;
wire _102_;
wire [1:0] _103_;
wire [1:0] _104_;
wire [15:0] _105_;
wire [15:0] _106_;
wire _107_;
wire [15:0] _108_;
wire [16:0] _109_;
wire [16:0] _110_;
wire [16:0] _111_;
wire [16:0] _112_;
wire _113_;
wire [16:0] _114_;
wire [17:0] _115_;
wire [17:0] _116_;
wire [2:0] _117_;
wire [2:0] _118_;
wire _119_;
wire [1:0] _120_;
wire [2:0] _121_;
wire [3:0] _122_;
wire [2:0] _123_;
wire [2:0] _124_;
wire _125_;
wire [1:0] _126_;
wire [2:0] _127_;
wire [3:0] _128_;
wire [2:0] _129_;
wire [2:0] _130_;
wire _131_;
wire [1:0] _132_;
wire [2:0] _133_;
wire [3:0] _134_;
wire [2:0] _135_;
wire [2:0] _136_;
wire _137_;
wire [1:0] _138_;
wire [2:0] _139_;
wire [3:0] _140_;
wire [2:0] _141_;
wire [2:0] _142_;
wire _143_;
wire [2:0] _144_;
wire [3:0] _145_;
wire [3:0] _146_;
wire [3:0] _147_;
wire [3:0] _148_;
wire _149_;
wire [3:0] _150_;
wire [4:0] _151_;
wire [4:0] _152_;
wire [4:0] _153_;
wire [4:0] _154_;
wire _155_;
wire [3:0] _156_;
wire [4:0] _157_;
wire [5:0] _158_;
wire [7:0] _159_;
wire [7:0] _160_;
wire [7:0] _161_;
wire [7:0] _162_;
wire [7:0] _163_;
wire [7:0] _164_;
wire [31:0] _165_;
wire [31:0] _166_;
wire [31:0] _167_;
wire [31:0] _168_;
wire [31:0] _169_;
wire [31:0] _170_;
wire [7:0] _171_;
wire [31:0] _172_;
wire [7:0] _173_;
wire [31:0] _174_;
wire [7:0] _175_;
wire [31:0] _176_;
wire [7:0] _177_;
wire [31:0] _178_;
wire [7:0] _179_;
wire [31:0] _180_;
wire [7:0] _181_;
wire [31:0] _182_;
wire [31:0] _183_;
wire [31:0] _184_;
wire [31:0] _185_;
wire _186_;
wire _187_;
wire _188_;
wire _189_;
wire [1:0] _190_;
wire [1:0] _191_;
wire [1:0] _192_;
wire [1:0] _193_;
wire _194_;
wire [1:0] _195_;
wire [2:0] _196_;
wire [2:0] _197_;
wire _198_;
wire _199_;
wire _200_;
wire _201_;
wire _202_;
wire _203_;
wire _204_;
wire _205_;
wire _206_;
wire _207_;
wire _208_;
wire _209_;
wire _210_;
wire _211_;
wire _212_;
wire _213_;
wire _214_;
wire _215_;
wire _216_;
wire _217_;
wire _218_;
wire _219_;
wire _220_;
wire _221_;
wire _222_;
wire _223_;
wire _224_;
wire _225_;
wire _226_;
wire _227_;
wire _228_;
wire _229_;
wire _230_;
wire _231_;
wire _232_;
wire _233_;
wire _234_;
wire _235_;
wire _236_;
wire _237_;
wire \add_10s_10ns_10_2_1_U11.ce ;
wire \add_10s_10ns_10_2_1_U11.clk ;
wire [9:0] \add_10s_10ns_10_2_1_U11.din0 ;
wire [9:0] \add_10s_10ns_10_2_1_U11.din1 ;
wire [9:0] \add_10s_10ns_10_2_1_U11.dout ;
wire \add_10s_10ns_10_2_1_U11.reset ;
wire [9:0] \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.a ;
wire [9:0] \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.ain_s0 ;
wire [9:0] \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.b ;
wire [9:0] \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.bin_s0 ;
wire \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.ce ;
wire \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.clk ;
wire \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.facout_s1 ;
wire \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.facout_s2 ;
wire [4:0] \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.fas_s1 ;
wire [4:0] \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.fas_s2 ;
wire \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.reset ;
wire [9:0] \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.s ;
wire [4:0] \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.u1.a ;
wire [4:0] \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.u1.b ;
wire \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.u1.cin ;
wire \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.u1.cout ;
wire [4:0] \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.u1.s ;
wire [4:0] \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.u2.a ;
wire [4:0] \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.u2.b ;
wire \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.u2.cin ;
wire \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.u2.cout ;
wire [4:0] \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.u2.s ;
wire \add_10s_10ns_10_2_1_U15.ce ;
wire \add_10s_10ns_10_2_1_U15.clk ;
wire [9:0] \add_10s_10ns_10_2_1_U15.din0 ;
wire [9:0] \add_10s_10ns_10_2_1_U15.din1 ;
wire [9:0] \add_10s_10ns_10_2_1_U15.dout ;
wire \add_10s_10ns_10_2_1_U15.reset ;
wire [9:0] \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.a ;
wire [9:0] \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.ain_s0 ;
wire [9:0] \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.b ;
wire [9:0] \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.bin_s0 ;
wire \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.ce ;
wire \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.clk ;
wire \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.facout_s1 ;
wire \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.facout_s2 ;
wire [4:0] \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.fas_s1 ;
wire [4:0] \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.fas_s2 ;
wire \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.reset ;
wire [9:0] \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.s ;
wire [4:0] \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.u1.a ;
wire [4:0] \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.u1.b ;
wire \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.u1.cin ;
wire \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.u1.cout ;
wire [4:0] \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.u1.s ;
wire [4:0] \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.u2.a ;
wire [4:0] \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.u2.b ;
wire \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.u2.cin ;
wire \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.u2.cout ;
wire [4:0] \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.u2.s ;
wire \add_10s_10ns_10_2_1_U17.ce ;
wire \add_10s_10ns_10_2_1_U17.clk ;
wire [9:0] \add_10s_10ns_10_2_1_U17.din0 ;
wire [9:0] \add_10s_10ns_10_2_1_U17.din1 ;
wire [9:0] \add_10s_10ns_10_2_1_U17.dout ;
wire \add_10s_10ns_10_2_1_U17.reset ;
wire [9:0] \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.a ;
wire [9:0] \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.ain_s0 ;
wire [9:0] \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.b ;
wire [9:0] \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.bin_s0 ;
wire \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.ce ;
wire \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.clk ;
wire \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.facout_s1 ;
wire \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.facout_s2 ;
wire [4:0] \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.fas_s1 ;
wire [4:0] \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.fas_s2 ;
wire \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.reset ;
wire [9:0] \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.s ;
wire [4:0] \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.u1.a ;
wire [4:0] \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.u1.b ;
wire \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.u1.cin ;
wire \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.u1.cout ;
wire [4:0] \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.u1.s ;
wire [4:0] \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.u2.a ;
wire [4:0] \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.u2.b ;
wire \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.u2.cin ;
wire \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.u2.cout ;
wire [4:0] \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.u2.s ;
wire \add_17s_17s_17_2_1_U6.ce ;
wire \add_17s_17s_17_2_1_U6.clk ;
wire [16:0] \add_17s_17s_17_2_1_U6.din0 ;
wire [16:0] \add_17s_17s_17_2_1_U6.din1 ;
wire [16:0] \add_17s_17s_17_2_1_U6.dout ;
wire \add_17s_17s_17_2_1_U6.reset ;
wire [16:0] \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.a ;
wire [16:0] \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.ain_s0 ;
wire [16:0] \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.b ;
wire [16:0] \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.bin_s0 ;
wire \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.ce ;
wire \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.clk ;
wire \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.facout_s1 ;
wire \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.facout_s2 ;
wire [7:0] \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.fas_s1 ;
wire [8:0] \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.fas_s2 ;
wire \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.reset ;
wire [16:0] \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.s ;
wire [7:0] \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.u1.a ;
wire [7:0] \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.u1.b ;
wire \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.u1.cin ;
wire \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.u1.cout ;
wire [7:0] \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.u1.s ;
wire [8:0] \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.u2.a ;
wire [8:0] \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.u2.b ;
wire \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.u2.cin ;
wire \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.u2.cout ;
wire [8:0] \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.u2.s ;
wire \add_2ns_2ns_2_2_1_U10.ce ;
wire \add_2ns_2ns_2_2_1_U10.clk ;
wire [1:0] \add_2ns_2ns_2_2_1_U10.din0 ;
wire [1:0] \add_2ns_2ns_2_2_1_U10.din1 ;
wire [1:0] \add_2ns_2ns_2_2_1_U10.dout ;
wire \add_2ns_2ns_2_2_1_U10.reset ;
wire [1:0] \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.a ;
wire [1:0] \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.ain_s0 ;
wire [1:0] \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.b ;
wire [1:0] \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.bin_s0 ;
wire \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.ce ;
wire \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.clk ;
wire \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.facout_s1 ;
wire \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.facout_s2 ;
wire \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.fas_s1 ;
wire \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.fas_s2 ;
wire \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.reset ;
wire [1:0] \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.s ;
wire \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.a ;
wire \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.b ;
wire \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.cin ;
wire \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.cout ;
wire \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.s ;
wire \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.a ;
wire \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.b ;
wire \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.cin ;
wire \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.cout ;
wire \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.s ;
wire \add_2ns_2ns_2_2_1_U14.ce ;
wire \add_2ns_2ns_2_2_1_U14.clk ;
wire [1:0] \add_2ns_2ns_2_2_1_U14.din0 ;
wire [1:0] \add_2ns_2ns_2_2_1_U14.din1 ;
wire [1:0] \add_2ns_2ns_2_2_1_U14.dout ;
wire \add_2ns_2ns_2_2_1_U14.reset ;
wire [1:0] \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.a ;
wire [1:0] \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.ain_s0 ;
wire [1:0] \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.b ;
wire [1:0] \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.bin_s0 ;
wire \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.ce ;
wire \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.clk ;
wire \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.facout_s1 ;
wire \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.facout_s2 ;
wire \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.fas_s1 ;
wire \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.fas_s2 ;
wire \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.reset ;
wire [1:0] \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.s ;
wire \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.a ;
wire \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.b ;
wire \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.cin ;
wire \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.cout ;
wire \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.s ;
wire \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.a ;
wire \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.b ;
wire \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.cin ;
wire \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.cout ;
wire \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.s ;
wire \add_2ns_2ns_2_2_1_U2.ce ;
wire \add_2ns_2ns_2_2_1_U2.clk ;
wire [1:0] \add_2ns_2ns_2_2_1_U2.din0 ;
wire [1:0] \add_2ns_2ns_2_2_1_U2.din1 ;
wire [1:0] \add_2ns_2ns_2_2_1_U2.dout ;
wire \add_2ns_2ns_2_2_1_U2.reset ;
wire [1:0] \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.a ;
wire [1:0] \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.ain_s0 ;
wire [1:0] \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.b ;
wire [1:0] \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.bin_s0 ;
wire \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.ce ;
wire \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.clk ;
wire \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.facout_s1 ;
wire \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.facout_s2 ;
wire \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.fas_s1 ;
wire \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.fas_s2 ;
wire \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.reset ;
wire [1:0] \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.s ;
wire \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.a ;
wire \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.b ;
wire \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.cin ;
wire \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.cout ;
wire \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.s ;
wire \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.a ;
wire \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.b ;
wire \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.cin ;
wire \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.cout ;
wire \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.s ;
wire \add_32ns_32ns_32_2_1_U19.ce ;
wire \add_32ns_32ns_32_2_1_U19.clk ;
wire [31:0] \add_32ns_32ns_32_2_1_U19.din0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U19.din1 ;
wire [31:0] \add_32ns_32ns_32_2_1_U19.dout ;
wire \add_32ns_32ns_32_2_1_U19.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.a ;
wire [31:0] \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.ain_s0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.b ;
wire [31:0] \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.bin_s0 ;
wire \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.ce ;
wire \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.clk ;
wire \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.facout_s1 ;
wire \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.facout_s2 ;
wire [15:0] \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.fas_s1 ;
wire [15:0] \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.fas_s2 ;
wire \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.u1.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.u1.b ;
wire \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.u1.cin ;
wire \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.u1.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.u1.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.u2.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.u2.b ;
wire \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.u2.cin ;
wire \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.u2.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.u2.s ;
wire \add_34s_34s_34_2_1_U18.ce ;
wire \add_34s_34s_34_2_1_U18.clk ;
wire [33:0] \add_34s_34s_34_2_1_U18.din0 ;
wire [33:0] \add_34s_34s_34_2_1_U18.din1 ;
wire [33:0] \add_34s_34s_34_2_1_U18.dout ;
wire \add_34s_34s_34_2_1_U18.reset ;
wire [33:0] \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.a ;
wire [33:0] \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.ain_s0 ;
wire [33:0] \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.b ;
wire [33:0] \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.bin_s0 ;
wire \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.ce ;
wire \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.clk ;
wire \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.facout_s1 ;
wire \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.facout_s2 ;
wire [16:0] \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.fas_s1 ;
wire [16:0] \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.fas_s2 ;
wire \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.reset ;
wire [33:0] \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.s ;
wire [16:0] \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.u1.a ;
wire [16:0] \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.u1.b ;
wire \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.u1.cin ;
wire \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.u1.cout ;
wire [16:0] \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.u1.s ;
wire [16:0] \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.u2.a ;
wire [16:0] \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.u2.b ;
wire \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.u2.cin ;
wire \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.u2.cout ;
wire [16:0] \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.u2.s ;
wire \add_5ns_5ns_5_2_1_U13.ce ;
wire \add_5ns_5ns_5_2_1_U13.clk ;
wire [4:0] \add_5ns_5ns_5_2_1_U13.din0 ;
wire [4:0] \add_5ns_5ns_5_2_1_U13.din1 ;
wire [4:0] \add_5ns_5ns_5_2_1_U13.dout ;
wire \add_5ns_5ns_5_2_1_U13.reset ;
wire [4:0] \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.a ;
wire [4:0] \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.ain_s0 ;
wire [4:0] \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.b ;
wire [4:0] \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.bin_s0 ;
wire \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.ce ;
wire \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.clk ;
wire \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.facout_s1 ;
wire \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.facout_s2 ;
wire [1:0] \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.fas_s1 ;
wire [2:0] \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.fas_s2 ;
wire \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.reset ;
wire [4:0] \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.s ;
wire [1:0] \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.u1.a ;
wire [1:0] \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.u1.b ;
wire \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.u1.cin ;
wire \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.u1.cout ;
wire [1:0] \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.u1.s ;
wire [2:0] \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.u2.a ;
wire [2:0] \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.u2.b ;
wire \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.u2.cin ;
wire \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.u2.cout ;
wire [2:0] \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.u2.s ;
wire \add_5ns_5ns_5_2_1_U5.ce ;
wire \add_5ns_5ns_5_2_1_U5.clk ;
wire [4:0] \add_5ns_5ns_5_2_1_U5.din0 ;
wire [4:0] \add_5ns_5ns_5_2_1_U5.din1 ;
wire [4:0] \add_5ns_5ns_5_2_1_U5.dout ;
wire \add_5ns_5ns_5_2_1_U5.reset ;
wire [4:0] \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.a ;
wire [4:0] \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.ain_s0 ;
wire [4:0] \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.b ;
wire [4:0] \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.bin_s0 ;
wire \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.ce ;
wire \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.clk ;
wire \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.facout_s1 ;
wire \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.facout_s2 ;
wire [1:0] \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.fas_s1 ;
wire [2:0] \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.fas_s2 ;
wire \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.reset ;
wire [4:0] \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.s ;
wire [1:0] \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.u1.a ;
wire [1:0] \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.u1.b ;
wire \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.u1.cin ;
wire \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.u1.cout ;
wire [1:0] \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.u1.s ;
wire [2:0] \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.u2.a ;
wire [2:0] \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.u2.b ;
wire \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.u2.cin ;
wire \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.u2.cout ;
wire [2:0] \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.u2.s ;
wire \add_5ns_5s_5_2_1_U4.ce ;
wire \add_5ns_5s_5_2_1_U4.clk ;
wire [4:0] \add_5ns_5s_5_2_1_U4.din0 ;
wire [4:0] \add_5ns_5s_5_2_1_U4.din1 ;
wire [4:0] \add_5ns_5s_5_2_1_U4.dout ;
wire \add_5ns_5s_5_2_1_U4.reset ;
wire [4:0] \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.a ;
wire [4:0] \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.ain_s0 ;
wire [4:0] \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.b ;
wire [4:0] \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.bin_s0 ;
wire \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.ce ;
wire \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.clk ;
wire \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.facout_s1 ;
wire \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.facout_s2 ;
wire [1:0] \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.fas_s1 ;
wire [2:0] \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.fas_s2 ;
wire \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.reset ;
wire [4:0] \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.s ;
wire [1:0] \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.u1.a ;
wire [1:0] \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.u1.b ;
wire \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.u1.cin ;
wire \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.u1.cout ;
wire [1:0] \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.u1.s ;
wire [2:0] \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.u2.a ;
wire [2:0] \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.u2.b ;
wire \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.u2.cin ;
wire \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.u2.cout ;
wire [2:0] \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.u2.s ;
wire \add_5s_5s_5_2_1_U12.ce ;
wire \add_5s_5s_5_2_1_U12.clk ;
wire [4:0] \add_5s_5s_5_2_1_U12.din0 ;
wire [4:0] \add_5s_5s_5_2_1_U12.din1 ;
wire [4:0] \add_5s_5s_5_2_1_U12.dout ;
wire \add_5s_5s_5_2_1_U12.reset ;
wire [4:0] \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.a ;
wire [4:0] \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.ain_s0 ;
wire [4:0] \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.b ;
wire [4:0] \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.bin_s0 ;
wire \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.ce ;
wire \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.clk ;
wire \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.facout_s1 ;
wire \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.facout_s2 ;
wire [1:0] \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.fas_s1 ;
wire [2:0] \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.fas_s2 ;
wire \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.reset ;
wire [4:0] \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.s ;
wire [1:0] \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.u1.a ;
wire [1:0] \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.u1.b ;
wire \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.u1.cin ;
wire \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.u1.cout ;
wire [1:0] \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.u1.s ;
wire [2:0] \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.u2.a ;
wire [2:0] \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.u2.b ;
wire \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.u2.cin ;
wire \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.u2.cout ;
wire [2:0] \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.u2.s ;
wire \add_6s_6ns_6_2_1_U16.ce ;
wire \add_6s_6ns_6_2_1_U16.clk ;
wire [5:0] \add_6s_6ns_6_2_1_U16.din0 ;
wire [5:0] \add_6s_6ns_6_2_1_U16.din1 ;
wire [5:0] \add_6s_6ns_6_2_1_U16.dout ;
wire \add_6s_6ns_6_2_1_U16.reset ;
wire [5:0] \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.a ;
wire [5:0] \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.ain_s0 ;
wire [5:0] \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.b ;
wire [5:0] \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.bin_s0 ;
wire \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.ce ;
wire \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.clk ;
wire \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.facout_s1 ;
wire \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.facout_s2 ;
wire [2:0] \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.fas_s1 ;
wire [2:0] \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.fas_s2 ;
wire \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.reset ;
wire [5:0] \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.s ;
wire [2:0] \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.u1.a ;
wire [2:0] \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.u1.b ;
wire \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.u1.cin ;
wire \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.u1.cout ;
wire [2:0] \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.u1.s ;
wire [2:0] \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.u2.a ;
wire [2:0] \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.u2.b ;
wire \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.u2.cin ;
wire \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.u2.cout ;
wire [2:0] \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.u2.s ;
wire \add_8s_8ns_8_2_1_U7.ce ;
wire \add_8s_8ns_8_2_1_U7.clk ;
wire [7:0] \add_8s_8ns_8_2_1_U7.din0 ;
wire [7:0] \add_8s_8ns_8_2_1_U7.din1 ;
wire [7:0] \add_8s_8ns_8_2_1_U7.dout ;
wire \add_8s_8ns_8_2_1_U7.reset ;
wire [7:0] \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.a ;
wire [7:0] \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.ain_s0 ;
wire [7:0] \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.b ;
wire [7:0] \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.bin_s0 ;
wire \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.ce ;
wire \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.clk ;
wire \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.facout_s1 ;
wire \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.facout_s2 ;
wire [3:0] \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.fas_s1 ;
wire [3:0] \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.fas_s2 ;
wire \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.reset ;
wire [7:0] \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.s ;
wire [3:0] \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.u1.a ;
wire [3:0] \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.u1.b ;
wire \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.u1.cin ;
wire \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.u1.cout ;
wire [3:0] \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.u1.s ;
wire [3:0] \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.u2.a ;
wire [3:0] \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.u2.b ;
wire \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.u2.cin ;
wire \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.u2.cout ;
wire [3:0] \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.u2.s ;
wire \add_9ns_9s_9_2_1_U1.ce ;
wire \add_9ns_9s_9_2_1_U1.clk ;
wire [8:0] \add_9ns_9s_9_2_1_U1.din0 ;
wire [8:0] \add_9ns_9s_9_2_1_U1.din1 ;
wire [8:0] \add_9ns_9s_9_2_1_U1.dout ;
wire \add_9ns_9s_9_2_1_U1.reset ;
wire [8:0] \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.a ;
wire [8:0] \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.ain_s0 ;
wire [8:0] \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.b ;
wire [8:0] \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.bin_s0 ;
wire \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.ce ;
wire \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.clk ;
wire \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.facout_s1 ;
wire \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.facout_s2 ;
wire [3:0] \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.fas_s1 ;
wire [4:0] \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.fas_s2 ;
wire \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.reset ;
wire [8:0] \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.s ;
wire [3:0] \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.u1.a ;
wire [3:0] \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.u1.b ;
wire \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.u1.cin ;
wire \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.u1.cout ;
wire [3:0] \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.u1.s ;
wire [4:0] \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.u2.a ;
wire [4:0] \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.u2.b ;
wire \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.u2.cin ;
wire \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.u2.cout ;
wire [4:0] \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.u2.s ;
wire and_ln340_fu_491_p2;
wire and_ln785_1_fu_526_p2;
wire and_ln785_fu_520_p2;
wire and_ln850_1_fu_368_p2;
wire and_ln850_2_fu_568_p2;
wire and_ln850_fu_350_p2;
wire ap_CS_fsm_state1;
wire ap_CS_fsm_state10;
wire ap_CS_fsm_state11;
wire ap_CS_fsm_state12;
wire ap_CS_fsm_state13;
wire ap_CS_fsm_state14;
wire ap_CS_fsm_state15;
wire ap_CS_fsm_state16;
wire ap_CS_fsm_state17;
wire ap_CS_fsm_state18;
wire ap_CS_fsm_state19;
wire ap_CS_fsm_state2;
wire ap_CS_fsm_state20;
wire ap_CS_fsm_state21;
wire ap_CS_fsm_state22;
wire ap_CS_fsm_state23;
wire ap_CS_fsm_state24;
wire ap_CS_fsm_state25;
wire ap_CS_fsm_state26;
wire ap_CS_fsm_state27;
wire ap_CS_fsm_state28;
wire ap_CS_fsm_state29;
wire ap_CS_fsm_state3;
wire ap_CS_fsm_state30;
wire ap_CS_fsm_state31;
wire ap_CS_fsm_state32;
wire ap_CS_fsm_state33;
wire ap_CS_fsm_state4;
wire ap_CS_fsm_state5;
wire ap_CS_fsm_state6;
wire ap_CS_fsm_state7;
wire ap_CS_fsm_state8;
wire ap_CS_fsm_state9;
wire [32:0] ap_NS_fsm;
wire ap_clk;
wire ap_done;
wire ap_idle;
wire ap_ready;
wire ap_rst;
wire ap_start;
wire [8:0] grp_fu_235_p1;
wire [8:0] grp_fu_235_p2;
wire [1:0] grp_fu_256_p2;
wire [31:0] grp_fu_315_p0;
wire [31:0] grp_fu_315_p1;
wire [31:0] grp_fu_315_p2;
wire [4:0] grp_fu_549_p1;
wire [4:0] grp_fu_549_p2;
wire [4:0] grp_fu_587_p2;
wire [16:0] grp_fu_606_p0;
wire [16:0] grp_fu_606_p1;
wire [16:0] grp_fu_606_p2;
wire [7:0] grp_fu_649_p0;
wire [7:0] grp_fu_649_p2;
wire [3:0] grp_fu_671_p0;
wire [3:0] grp_fu_671_p1;
wire [3:0] grp_fu_671_p2;
wire [1:0] grp_fu_677_p2;
wire [1:0] grp_fu_685_p1;
wire [1:0] grp_fu_685_p2;
wire [9:0] grp_fu_741_p0;
wire [9:0] grp_fu_741_p1;
wire [9:0] grp_fu_741_p2;
wire [4:0] grp_fu_747_p0;
wire [4:0] grp_fu_747_p1;
wire [4:0] grp_fu_747_p2;
wire [4:0] grp_fu_753_p0;
wire [4:0] grp_fu_753_p1;
wire [4:0] grp_fu_753_p2;
wire [1:0] grp_fu_759_p2;
wire [9:0] grp_fu_766_p0;
wire [9:0] grp_fu_766_p2;
wire [5:0] grp_fu_777_p0;
wire [5:0] grp_fu_777_p1;
wire [5:0] grp_fu_777_p2;
wire [9:0] grp_fu_786_p0;
wire [9:0] grp_fu_786_p2;
wire [33:0] grp_fu_806_p0;
wire [33:0] grp_fu_806_p1;
wire [33:0] grp_fu_806_p2;
wire [31:0] grp_fu_822_p2;
wire icmp_ln768_fu_416_p2;
wire icmp_ln786_fu_422_p2;
wire icmp_ln850_1_fu_326_p2;
wire icmp_ln850_2_fu_331_p2;
wire icmp_ln850_3_fu_541_p2;
wire icmp_ln850_fu_321_p2;
wire icmp_ln851_1_fu_616_p2;
wire icmp_ln851_fu_240_p2;
wire [7:0] lhs_fu_283_p3;
wire [15:0] op_0;
wire [15:0] op_10;
wire op_11;
wire op_12;
wire [3:0] op_16;
wire [1:0] op_17;
wire op_18;
wire [3:0] op_19;
wire [3:0] op_1_V_fu_531_p3;
wire op_2;
wire [7:0] op_3;
wire [31:0] op_31;
wire op_31_ap_vld;
wire [1:0] op_6;
wire [31:0] op_7;
wire or_ln340_fu_480_p2;
wire or_ln785_1_fu_515_p2;
wire or_ln785_fu_449_p2;
wire or_ln786_fu_475_p2;
wire overflow_fu_465_p2;
wire p_Result_1_fu_343_p3;
wire p_Result_2_fu_561_p3;
wire p_Result_5_fu_690_p3;
wire p_Result_6_fu_827_p3;
wire p_Result_s_12_fu_261_p3;
wire [12:0] p_Result_s_fu_406_p4;
wire [3:0] p_Val2_s_fu_453_p3;
wire [7:0] r_fu_443_p3;
wire ret_V_10_fu_554_p3;
wire [1:0] ret_V_18_fu_273_p3;
wire [7:0] ret_V_19_fu_290_p1;
wire [7:0] ret_V_19_fu_290_p2;
wire ret_V_20_fu_355_p2;
wire [7:0] ret_V_21_fu_299_p1;
wire [7:0] ret_V_21_fu_299_p2;
wire ret_V_22_fu_372_p2;
wire ret_V_23_fu_573_p2;
wire [7:0] ret_V_26_fu_702_p3;
wire ret_V_5_fu_336_p3;
wire ret_V_8_fu_361_p3;
wire [14:0] rhs_2_fu_595_p3;
wire [1:0] select_ln1192_fu_378_p3;
wire [1:0] select_ln1347_1_fu_639_p3;
wire [1:0] select_ln1347_fu_632_p3;
wire [3:0] select_ln340_fu_497_p3;
wire [1:0] select_ln69_1_fu_709_p3;
wire [1:0] select_ln69_2_fu_655_p3;
wire [4:0] select_ln69_fu_579_p3;
wire [8:0] select_ln703_fu_219_p3;
wire [7:0] select_ln850_1_fu_697_p3;
wire [31:0] select_ln850_2_fu_837_p3;
wire [6:0] select_ln850_4_fu_435_p3;
wire [1:0] select_ln850_fu_268_p3;
wire [15:0] sext_ln1192_fu_591_p0;
wire [7:0] sext_ln1299_fu_312_p0;
wire [7:0] sext_ln353_fu_280_p1;
wire [3:0] sext_ln69_1_fu_720_p1;
wire [3:0] sext_ln703_2_fu_791_p0;
wire [7:0] sext_ln703_fu_227_p0;
wire [7:0] sext_ln850_fu_646_p1;
wire \shl_32s_8ns_32_7_1_U3.ce ;
wire \shl_32s_8ns_32_7_1_U3.clk ;
wire [31:0] \shl_32s_8ns_32_7_1_U3.din0 ;
wire [31:0] \shl_32s_8ns_32_7_1_U3.din1 ;
wire [7:0] \shl_32s_8ns_32_7_1_U3.din1_cast ;
wire [7:0] \shl_32s_8ns_32_7_1_U3.din1_mask ;
wire [31:0] \shl_32s_8ns_32_7_1_U3.dout ;
wire \shl_32s_8ns_32_7_1_U3.reset ;
wire \sub_2ns_2ns_2_2_1_U9.ce ;
wire \sub_2ns_2ns_2_2_1_U9.clk ;
wire [1:0] \sub_2ns_2ns_2_2_1_U9.din0 ;
wire [1:0] \sub_2ns_2ns_2_2_1_U9.din1 ;
wire [1:0] \sub_2ns_2ns_2_2_1_U9.dout ;
wire \sub_2ns_2ns_2_2_1_U9.reset ;
wire [1:0] \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.a ;
wire [1:0] \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.ain_s0 ;
wire [1:0] \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.b ;
wire [1:0] \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.bin_s0 ;
wire \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.ce ;
wire \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.clk ;
wire \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.facout_s1 ;
wire \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.facout_s2 ;
wire \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.fas_s1 ;
wire \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.fas_s2 ;
wire \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.reset ;
wire [1:0] \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.s ;
wire \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.u1.a ;
wire \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.u1.b ;
wire \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.u1.cin ;
wire \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.u1.cout ;
wire \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.u1.s ;
wire \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.u2.a ;
wire \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.u2.b ;
wire \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.u2.cin ;
wire \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.u2.cout ;
wire \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.u2.s ;
wire \sub_4s_4ns_4_2_1_U8.ce ;
wire \sub_4s_4ns_4_2_1_U8.clk ;
wire [3:0] \sub_4s_4ns_4_2_1_U8.din0 ;
wire [3:0] \sub_4s_4ns_4_2_1_U8.din1 ;
wire [3:0] \sub_4s_4ns_4_2_1_U8.dout ;
wire \sub_4s_4ns_4_2_1_U8.reset ;
wire [3:0] \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.a ;
wire [3:0] \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.ain_s0 ;
wire [3:0] \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.b ;
wire [3:0] \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.bin_s0 ;
wire \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.ce ;
wire \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.clk ;
wire \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.facout_s1 ;
wire \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.facout_s2 ;
wire [1:0] \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.fas_s1 ;
wire [1:0] \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.fas_s2 ;
wire \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.reset ;
wire [3:0] \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.s ;
wire [1:0] \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.u1.a ;
wire [1:0] \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.u1.b ;
wire \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.u1.cin ;
wire \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.u1.cout ;
wire [1:0] \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.u1.s ;
wire [1:0] \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.u2.a ;
wire [1:0] \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.u2.b ;
wire \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.u2.cin ;
wire \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.u2.cout ;
wire [1:0] \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.u2.s ;
wire [10:0] tmp_11_fu_795_p3;
wire tmp_9_fu_428_p3;
wire [7:0] trunc_ln1192_fu_231_p0;
wire [6:0] trunc_ln1192_fu_231_p1;
wire [2:0] trunc_ln703_fu_386_p1;
wire [6:0] trunc_ln851_1_fu_304_p1;
wire [6:0] trunc_ln851_2_fu_537_p1;
wire [15:0] trunc_ln851_3_fu_612_p0;
wire [9:0] trunc_ln851_3_fu_612_p1;
wire [3:0] trunc_ln851_4_fu_834_p0;
wire trunc_ln851_4_fu_834_p1;
wire [6:0] trunc_ln851_fu_295_p1;
wire xor_ln340_fu_485_p2;
wire xor_ln785_1_fu_510_p2;
wire xor_ln785_fu_460_p2;
wire xor_ln786_1_fu_505_p2;
wire xor_ln786_fu_470_p2;


assign _056_ = icmp_ln851_1_reg_1067 & ap_CS_fsm[20];
assign _057_ = _060_ & ap_CS_fsm[4];
assign _058_ = _061_ & ap_CS_fsm[0];
assign _059_ = ap_start & ap_CS_fsm[0];
assign and_ln340_fu_491_p2 = xor_ln340_fu_485_p2 & or_ln786_fu_475_p2;
assign and_ln785_1_fu_526_p2 = p_Result_8_reg_977 & and_ln785_fu_520_p2;
assign and_ln785_fu_520_p2 = xor_ln786_1_fu_505_p2 & or_ln785_1_fu_515_p2;
assign and_ln850_1_fu_368_p2 = icmp_ln850_2_reg_949 & icmp_ln850_1_reg_944;
assign and_ln850_2_fu_568_p2 = shl_ln1299_reg_1021[7] & icmp_ln850_3_reg_1032;
assign and_ln850_fu_350_p2 = ret_V_19_reg_907[7] & icmp_ln850_reg_939;
assign overflow_fu_465_p2 = xor_ln785_fu_460_p2 & or_ln785_reg_1000;
assign ret_V_21_fu_299_p2 = op_3 & { op_2, 7'h00 };
assign xor_ln786_fu_470_p2 = ~ p_Result_8_reg_977;
assign xor_ln785_fu_460_p2 = ~ p_Result_7_reg_970;
assign xor_ln340_fu_485_p2 = ~ or_ln340_fu_480_p2;
assign xor_ln785_1_fu_510_p2 = ~ or_ln785_reg_1000;
assign xor_ln786_1_fu_505_p2 = ~ icmp_ln786_reg_989;
assign _060_ = ~ icmp_ln851_reg_874;
assign _061_ = ~ ap_start;
assign _062_ = ! op_3[6:0];
always @(posedge \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.clk )
\add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.bin_s1  <= _064_;
always @(posedge \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.clk )
\add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.ain_s1  <= _063_;
always @(posedge \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.clk )
\add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.sum_s1  <= _066_;
always @(posedge \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.clk )
\add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.carry_s1  <= _065_;
assign _064_ = \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.ce  ? \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.b [9:5] : \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.bin_s1 ;
assign _063_ = \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.ce  ? \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.a [9:5] : \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.ain_s1 ;
assign _065_ = \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.ce  ? \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.facout_s1  : \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.carry_s1 ;
assign _066_ = \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.ce  ? \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.fas_s1  : \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.sum_s1 ;
assign _067_ = \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.u1.a  + \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.u1.b ;
assign { \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.u1.cout , \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.u1.s  } = _067_ + \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.u1.cin ;
assign _068_ = \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.u2.a  + \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.u2.b ;
assign { \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.u2.cout , \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.u2.s  } = _068_ + \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.u2.cin ;
always @(posedge \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.clk )
\add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.bin_s1  <= _070_;
always @(posedge \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.clk )
\add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.ain_s1  <= _069_;
always @(posedge \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.clk )
\add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.sum_s1  <= _072_;
always @(posedge \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.clk )
\add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.carry_s1  <= _071_;
assign _070_ = \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.ce  ? \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.b [9:5] : \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.bin_s1 ;
assign _069_ = \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.ce  ? \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.a [9:5] : \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.ain_s1 ;
assign _071_ = \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.ce  ? \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.facout_s1  : \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.carry_s1 ;
assign _072_ = \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.ce  ? \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.fas_s1  : \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.sum_s1 ;
assign _073_ = \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.u1.a  + \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.u1.b ;
assign { \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.u1.cout , \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.u1.s  } = _073_ + \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.u1.cin ;
assign _074_ = \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.u2.a  + \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.u2.b ;
assign { \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.u2.cout , \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.u2.s  } = _074_ + \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.u2.cin ;
always @(posedge \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.clk )
\add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.bin_s1  <= _076_;
always @(posedge \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.clk )
\add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.ain_s1  <= _075_;
always @(posedge \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.clk )
\add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.sum_s1  <= _078_;
always @(posedge \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.clk )
\add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.carry_s1  <= _077_;
assign _076_ = \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.ce  ? \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.b [9:5] : \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.bin_s1 ;
assign _075_ = \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.ce  ? \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.a [9:5] : \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.ain_s1 ;
assign _077_ = \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.ce  ? \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.facout_s1  : \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.carry_s1 ;
assign _078_ = \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.ce  ? \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.fas_s1  : \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.sum_s1 ;
assign _079_ = \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.u1.a  + \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.u1.b ;
assign { \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.u1.cout , \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.u1.s  } = _079_ + \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.u1.cin ;
assign _080_ = \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.u2.a  + \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.u2.b ;
assign { \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.u2.cout , \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.u2.s  } = _080_ + \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.u2.cin ;
always @(posedge \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.clk )
\add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.bin_s1  <= _082_;
always @(posedge \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.clk )
\add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.ain_s1  <= _081_;
always @(posedge \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.clk )
\add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.sum_s1  <= _084_;
always @(posedge \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.clk )
\add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.carry_s1  <= _083_;
assign _082_ = \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.ce  ? \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.b [16:8] : \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.bin_s1 ;
assign _081_ = \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.ce  ? \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.a [16:8] : \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.ain_s1 ;
assign _083_ = \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.ce  ? \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.facout_s1  : \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.carry_s1 ;
assign _084_ = \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.ce  ? \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.fas_s1  : \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.sum_s1 ;
assign _085_ = \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.u1.a  + \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.u1.b ;
assign { \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.u1.cout , \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.u1.s  } = _085_ + \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.u1.cin ;
assign _086_ = \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.u2.a  + \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.u2.b ;
assign { \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.u2.cout , \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.u2.s  } = _086_ + \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.u2.cin ;
always @(posedge \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.clk )
\add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.bin_s1  <= _088_;
always @(posedge \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.clk )
\add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.ain_s1  <= _087_;
always @(posedge \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.clk )
\add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.sum_s1  <= _090_;
always @(posedge \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.clk )
\add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.carry_s1  <= _089_;
assign _088_ = \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.ce  ? \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.b [1] : \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.bin_s1 ;
assign _087_ = \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.ce  ? \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.a [1] : \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.ain_s1 ;
assign _089_ = \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.ce  ? \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.facout_s1  : \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.carry_s1 ;
assign _090_ = \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.ce  ? \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.fas_s1  : \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.sum_s1 ;
assign _091_ = \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.a  + \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.b ;
assign { \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.cout , \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.s  } = _091_ + \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.cin ;
assign _092_ = \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.a  + \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.b ;
assign { \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.cout , \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.s  } = _092_ + \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.cin ;
always @(posedge \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.clk )
\add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.bin_s1  <= _094_;
always @(posedge \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.clk )
\add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.ain_s1  <= _093_;
always @(posedge \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.clk )
\add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.sum_s1  <= _096_;
always @(posedge \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.clk )
\add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.carry_s1  <= _095_;
assign _094_ = \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.ce  ? \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.b [1] : \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.bin_s1 ;
assign _093_ = \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.ce  ? \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.a [1] : \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.ain_s1 ;
assign _095_ = \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.ce  ? \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.facout_s1  : \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.carry_s1 ;
assign _096_ = \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.ce  ? \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.fas_s1  : \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.sum_s1 ;
assign _097_ = \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.a  + \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.b ;
assign { \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.cout , \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.s  } = _097_ + \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.cin ;
assign _098_ = \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.a  + \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.b ;
assign { \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.cout , \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.s  } = _098_ + \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.cin ;
always @(posedge \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.clk )
\add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.bin_s1  <= _100_;
always @(posedge \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.clk )
\add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.ain_s1  <= _099_;
always @(posedge \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.clk )
\add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.sum_s1  <= _102_;
always @(posedge \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.clk )
\add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.carry_s1  <= _101_;
assign _100_ = \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.ce  ? \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.b [1] : \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.bin_s1 ;
assign _099_ = \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.ce  ? \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.a [1] : \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.ain_s1 ;
assign _101_ = \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.ce  ? \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.facout_s1  : \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.carry_s1 ;
assign _102_ = \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.ce  ? \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.fas_s1  : \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.sum_s1 ;
assign _103_ = \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.a  + \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.b ;
assign { \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.cout , \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.s  } = _103_ + \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.cin ;
assign _104_ = \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.a  + \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.b ;
assign { \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.cout , \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.s  } = _104_ + \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.cin ;
always @(posedge \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.clk )
\add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.bin_s1  <= _106_;
always @(posedge \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.clk )
\add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.ain_s1  <= _105_;
always @(posedge \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.clk )
\add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.sum_s1  <= _108_;
always @(posedge \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.clk )
\add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.carry_s1  <= _107_;
assign _106_ = \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.ce  ? \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.b [31:16] : \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.bin_s1 ;
assign _105_ = \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.ce  ? \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.a [31:16] : \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.ain_s1 ;
assign _107_ = \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.ce  ? \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.facout_s1  : \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.carry_s1 ;
assign _108_ = \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.ce  ? \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.fas_s1  : \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.sum_s1 ;
assign _109_ = \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.u1.a  + \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.u1.b ;
assign { \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.u1.cout , \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.u1.s  } = _109_ + \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.u1.cin ;
assign _110_ = \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.u2.a  + \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.u2.b ;
assign { \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.u2.cout , \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.u2.s  } = _110_ + \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.u2.cin ;
always @(posedge \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.clk )
\add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.bin_s1  <= _112_;
always @(posedge \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.clk )
\add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.ain_s1  <= _111_;
always @(posedge \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.clk )
\add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.sum_s1  <= _114_;
always @(posedge \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.clk )
\add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.carry_s1  <= _113_;
assign _112_ = \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.ce  ? \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.b [33:17] : \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.bin_s1 ;
assign _111_ = \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.ce  ? \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.a [33:17] : \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.ain_s1 ;
assign _113_ = \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.ce  ? \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.facout_s1  : \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.carry_s1 ;
assign _114_ = \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.ce  ? \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.fas_s1  : \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.sum_s1 ;
assign _115_ = \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.u1.a  + \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.u1.b ;
assign { \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.u1.cout , \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.u1.s  } = _115_ + \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.u1.cin ;
assign _116_ = \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.u2.a  + \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.u2.b ;
assign { \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.u2.cout , \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.u2.s  } = _116_ + \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.u2.cin ;
always @(posedge \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.clk )
\add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.bin_s1  <= _118_;
always @(posedge \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.clk )
\add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.ain_s1  <= _117_;
always @(posedge \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.clk )
\add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.sum_s1  <= _120_;
always @(posedge \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.clk )
\add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.carry_s1  <= _119_;
assign _118_ = \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.ce  ? \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.b [4:2] : \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.bin_s1 ;
assign _117_ = \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.ce  ? \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.a [4:2] : \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.ain_s1 ;
assign _119_ = \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.ce  ? \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.facout_s1  : \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.carry_s1 ;
assign _120_ = \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.ce  ? \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.fas_s1  : \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.sum_s1 ;
assign _121_ = \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.u1.a  + \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.u1.b ;
assign { \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.u1.cout , \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.u1.s  } = _121_ + \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.u1.cin ;
assign _122_ = \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.u2.a  + \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.u2.b ;
assign { \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.u2.cout , \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.u2.s  } = _122_ + \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.u2.cin ;
always @(posedge \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.clk )
\add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.bin_s1  <= _124_;
always @(posedge \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.clk )
\add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.ain_s1  <= _123_;
always @(posedge \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.clk )
\add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.sum_s1  <= _126_;
always @(posedge \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.clk )
\add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.carry_s1  <= _125_;
assign _124_ = \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.ce  ? \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.b [4:2] : \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.bin_s1 ;
assign _123_ = \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.ce  ? \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.a [4:2] : \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.ain_s1 ;
assign _125_ = \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.ce  ? \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.facout_s1  : \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.carry_s1 ;
assign _126_ = \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.ce  ? \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.fas_s1  : \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.sum_s1 ;
assign _127_ = \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.u1.a  + \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.u1.b ;
assign { \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.u1.cout , \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.u1.s  } = _127_ + \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.u1.cin ;
assign _128_ = \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.u2.a  + \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.u2.b ;
assign { \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.u2.cout , \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.u2.s  } = _128_ + \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.u2.cin ;
always @(posedge \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.clk )
\add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.bin_s1  <= _130_;
always @(posedge \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.clk )
\add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.ain_s1  <= _129_;
always @(posedge \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.clk )
\add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.sum_s1  <= _132_;
always @(posedge \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.clk )
\add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.carry_s1  <= _131_;
assign _130_ = \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.ce  ? \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.b [4:2] : \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.bin_s1 ;
assign _129_ = \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.ce  ? \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.a [4:2] : \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.ain_s1 ;
assign _131_ = \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.ce  ? \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.facout_s1  : \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.carry_s1 ;
assign _132_ = \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.ce  ? \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.fas_s1  : \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.sum_s1 ;
assign _133_ = \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.u1.a  + \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.u1.b ;
assign { \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.u1.cout , \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.u1.s  } = _133_ + \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.u1.cin ;
assign _134_ = \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.u2.a  + \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.u2.b ;
assign { \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.u2.cout , \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.u2.s  } = _134_ + \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.u2.cin ;
always @(posedge \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.clk )
\add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.bin_s1  <= _136_;
always @(posedge \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.clk )
\add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.ain_s1  <= _135_;
always @(posedge \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.clk )
\add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.sum_s1  <= _138_;
always @(posedge \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.clk )
\add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.carry_s1  <= _137_;
assign _136_ = \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.ce  ? \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.b [4:2] : \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.bin_s1 ;
assign _135_ = \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.ce  ? \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.a [4:2] : \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.ain_s1 ;
assign _137_ = \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.ce  ? \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.facout_s1  : \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.carry_s1 ;
assign _138_ = \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.ce  ? \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.fas_s1  : \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.sum_s1 ;
assign _139_ = \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.u1.a  + \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.u1.b ;
assign { \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.u1.cout , \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.u1.s  } = _139_ + \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.u1.cin ;
assign _140_ = \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.u2.a  + \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.u2.b ;
assign { \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.u2.cout , \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.u2.s  } = _140_ + \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.u2.cin ;
always @(posedge \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.clk )
\add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.bin_s1  <= _142_;
always @(posedge \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.clk )
\add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.ain_s1  <= _141_;
always @(posedge \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.clk )
\add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.sum_s1  <= _144_;
always @(posedge \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.clk )
\add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.carry_s1  <= _143_;
assign _142_ = \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.ce  ? \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.b [5:3] : \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.bin_s1 ;
assign _141_ = \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.ce  ? \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.a [5:3] : \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.ain_s1 ;
assign _143_ = \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.ce  ? \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.facout_s1  : \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.carry_s1 ;
assign _144_ = \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.ce  ? \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.fas_s1  : \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.sum_s1 ;
assign _145_ = \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.u1.a  + \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.u1.b ;
assign { \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.u1.cout , \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.u1.s  } = _145_ + \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.u1.cin ;
assign _146_ = \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.u2.a  + \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.u2.b ;
assign { \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.u2.cout , \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.u2.s  } = _146_ + \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.u2.cin ;
always @(posedge \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.clk )
\add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.bin_s1  <= _148_;
always @(posedge \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.clk )
\add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.ain_s1  <= _147_;
always @(posedge \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.clk )
\add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.sum_s1  <= _150_;
always @(posedge \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.clk )
\add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.carry_s1  <= _149_;
assign _148_ = \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.ce  ? \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.b [7:4] : \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.bin_s1 ;
assign _147_ = \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.ce  ? \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.a [7:4] : \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.ain_s1 ;
assign _149_ = \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.ce  ? \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.facout_s1  : \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.carry_s1 ;
assign _150_ = \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.ce  ? \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.fas_s1  : \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.sum_s1 ;
assign _151_ = \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.u1.a  + \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.u1.b ;
assign { \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.u1.cout , \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.u1.s  } = _151_ + \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.u1.cin ;
assign _152_ = \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.u2.a  + \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.u2.b ;
assign { \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.u2.cout , \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.u2.s  } = _152_ + \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.u2.cin ;
always @(posedge \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.clk )
\add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.bin_s1  <= _154_;
always @(posedge \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.clk )
\add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.ain_s1  <= _153_;
always @(posedge \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.clk )
\add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.sum_s1  <= _156_;
always @(posedge \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.clk )
\add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.carry_s1  <= _155_;
assign _154_ = \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.ce  ? \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.b [8:4] : \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.bin_s1 ;
assign _153_ = \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.ce  ? \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.a [8:4] : \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.ain_s1 ;
assign _155_ = \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.ce  ? \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.facout_s1  : \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.carry_s1 ;
assign _156_ = \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.ce  ? \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.fas_s1  : \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.sum_s1 ;
assign _157_ = \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.u1.a  + \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.u1.b ;
assign { \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.u1.cout , \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.u1.s  } = _157_ + \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.u1.cin ;
assign _158_ = \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.u2.a  + \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.u2.b ;
assign { \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.u2.cout , \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.u2.s  } = _158_ + \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.u2.cin ;
always @(posedge \shl_32s_8ns_32_7_1_U3.clk )
\shl_32s_8ns_32_7_1_U3.dout_array[5]  <= _170_;
always @(posedge \shl_32s_8ns_32_7_1_U3.clk )
\shl_32s_8ns_32_7_1_U3.din1_cast_array[5]  <= _164_;
always @(posedge \shl_32s_8ns_32_7_1_U3.clk )
\shl_32s_8ns_32_7_1_U3.dout_array[4]  <= _169_;
always @(posedge \shl_32s_8ns_32_7_1_U3.clk )
\shl_32s_8ns_32_7_1_U3.din1_cast_array[4]  <= _163_;
always @(posedge \shl_32s_8ns_32_7_1_U3.clk )
\shl_32s_8ns_32_7_1_U3.dout_array[3]  <= _168_;
always @(posedge \shl_32s_8ns_32_7_1_U3.clk )
\shl_32s_8ns_32_7_1_U3.din1_cast_array[3]  <= _162_;
always @(posedge \shl_32s_8ns_32_7_1_U3.clk )
\shl_32s_8ns_32_7_1_U3.dout_array[2]  <= _167_;
always @(posedge \shl_32s_8ns_32_7_1_U3.clk )
\shl_32s_8ns_32_7_1_U3.din1_cast_array[2]  <= _161_;
always @(posedge \shl_32s_8ns_32_7_1_U3.clk )
\shl_32s_8ns_32_7_1_U3.dout_array[1]  <= _166_;
always @(posedge \shl_32s_8ns_32_7_1_U3.clk )
\shl_32s_8ns_32_7_1_U3.din1_cast_array[1]  <= _160_;
always @(posedge \shl_32s_8ns_32_7_1_U3.clk )
\shl_32s_8ns_32_7_1_U3.dout_array[0]  <= _165_;
always @(posedge \shl_32s_8ns_32_7_1_U3.clk )
\shl_32s_8ns_32_7_1_U3.din1_cast_array[0]  <= _159_;
assign _171_ = \shl_32s_8ns_32_7_1_U3.ce  ? \shl_32s_8ns_32_7_1_U3.din1_cast_array[4]  : \shl_32s_8ns_32_7_1_U3.din1_cast_array[5] ;
assign _164_ = \shl_32s_8ns_32_7_1_U3.reset  ? 8'h00 : _171_;
assign _172_ = \shl_32s_8ns_32_7_1_U3.ce  ? _185_ : \shl_32s_8ns_32_7_1_U3.dout_array[5] ;
assign _170_ = \shl_32s_8ns_32_7_1_U3.reset  ? 32'd0 : _172_;
assign _173_ = \shl_32s_8ns_32_7_1_U3.ce  ? \shl_32s_8ns_32_7_1_U3.din1_cast_array[3]  : \shl_32s_8ns_32_7_1_U3.din1_cast_array[4] ;
assign _163_ = \shl_32s_8ns_32_7_1_U3.reset  ? 8'h00 : _173_;
assign _174_ = \shl_32s_8ns_32_7_1_U3.ce  ? _184_ : \shl_32s_8ns_32_7_1_U3.dout_array[4] ;
assign _169_ = \shl_32s_8ns_32_7_1_U3.reset  ? 32'd0 : _174_;
assign _175_ = \shl_32s_8ns_32_7_1_U3.ce  ? \shl_32s_8ns_32_7_1_U3.din1_cast_array[2]  : \shl_32s_8ns_32_7_1_U3.din1_cast_array[3] ;
assign _162_ = \shl_32s_8ns_32_7_1_U3.reset  ? 8'h00 : _175_;
assign _176_ = \shl_32s_8ns_32_7_1_U3.ce  ? _183_ : \shl_32s_8ns_32_7_1_U3.dout_array[3] ;
assign _168_ = \shl_32s_8ns_32_7_1_U3.reset  ? 32'd0 : _176_;
assign _177_ = \shl_32s_8ns_32_7_1_U3.ce  ? \shl_32s_8ns_32_7_1_U3.din1_cast_array[1]  : \shl_32s_8ns_32_7_1_U3.din1_cast_array[2] ;
assign _161_ = \shl_32s_8ns_32_7_1_U3.reset  ? 8'h00 : _177_;
assign _178_ = \shl_32s_8ns_32_7_1_U3.ce  ? \shl_32s_8ns_32_7_1_U3.dout_array[1]  : \shl_32s_8ns_32_7_1_U3.dout_array[2] ;
assign _167_ = \shl_32s_8ns_32_7_1_U3.reset  ? 32'd0 : _178_;
assign _179_ = \shl_32s_8ns_32_7_1_U3.ce  ? \shl_32s_8ns_32_7_1_U3.din1_cast_array[0]  : \shl_32s_8ns_32_7_1_U3.din1_cast_array[1] ;
assign _160_ = \shl_32s_8ns_32_7_1_U3.reset  ? 8'h00 : _179_;
assign _180_ = \shl_32s_8ns_32_7_1_U3.ce  ? \shl_32s_8ns_32_7_1_U3.dout_array[0]  : \shl_32s_8ns_32_7_1_U3.dout_array[1] ;
assign _166_ = \shl_32s_8ns_32_7_1_U3.reset  ? 32'd0 : _180_;
assign _181_ = \shl_32s_8ns_32_7_1_U3.ce  ? \shl_32s_8ns_32_7_1_U3.din1 [7:0] : \shl_32s_8ns_32_7_1_U3.din1_cast_array[0] ;
assign _159_ = \shl_32s_8ns_32_7_1_U3.reset  ? 8'h00 : _181_;
assign _182_ = \shl_32s_8ns_32_7_1_U3.ce  ? \shl_32s_8ns_32_7_1_U3.din0  : \shl_32s_8ns_32_7_1_U3.dout_array[0] ;
assign _165_ = \shl_32s_8ns_32_7_1_U3.reset  ? 32'd0 : _182_;
assign _183_ = \shl_32s_8ns_32_7_1_U3.dout_array[2]  << { \shl_32s_8ns_32_7_1_U3.din1_cast_array[2] [7:6], 6'h00 };
assign _184_ = \shl_32s_8ns_32_7_1_U3.dout_array[3]  << { \shl_32s_8ns_32_7_1_U3.din1_cast_array[3] [5:4], 4'h0 };
assign _185_ = \shl_32s_8ns_32_7_1_U3.dout_array[4]  << { \shl_32s_8ns_32_7_1_U3.din1_cast_array[4] [3:2], 2'h0 };
assign \shl_32s_8ns_32_7_1_U3.dout  = \shl_32s_8ns_32_7_1_U3.dout_array[5]  << \shl_32s_8ns_32_7_1_U3.din1_cast_array[5] [1:0];
assign \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.bin_s0  = ~ \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.b ;
always @(posedge \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.clk )
\sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.bin_s1  <= _187_;
always @(posedge \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.clk )
\sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.ain_s1  <= _186_;
always @(posedge \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.clk )
\sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.sum_s1  <= _189_;
always @(posedge \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.clk )
\sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.carry_s1  <= _188_;
assign _187_ = \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.ce  ? \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.bin_s0 [1] : \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.bin_s1 ;
assign _186_ = \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.ce  ? \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.a [1] : \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.ain_s1 ;
assign _188_ = \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.ce  ? \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.facout_s1  : \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.carry_s1 ;
assign _189_ = \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.ce  ? \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.fas_s1  : \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.sum_s1 ;
assign _190_ = \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.u1.a  + \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.u1.b ;
assign { \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.u1.cout , \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.u1.s  } = _190_ + \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.u1.cin ;
assign _191_ = \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.u2.a  + \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.u2.b ;
assign { \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.u2.cout , \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.u2.s  } = _191_ + \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.u2.cin ;
assign \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.bin_s0  = ~ \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.b ;
always @(posedge \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.clk )
\sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.bin_s1  <= _193_;
always @(posedge \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.clk )
\sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.ain_s1  <= _192_;
always @(posedge \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.clk )
\sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.sum_s1  <= _195_;
always @(posedge \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.clk )
\sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.carry_s1  <= _194_;
assign _193_ = \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.ce  ? \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.bin_s0 [3:2] : \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.bin_s1 ;
assign _192_ = \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.ce  ? \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.a [3:2] : \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.ain_s1 ;
assign _194_ = \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.ce  ? \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.facout_s1  : \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.carry_s1 ;
assign _195_ = \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.ce  ? \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.fas_s1  : \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.sum_s1 ;
assign _196_ = \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.u1.a  + \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.u1.b ;
assign { \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.u1.cout , \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.u1.s  } = _196_ + \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.u1.cin ;
assign _197_ = \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.u2.a  + \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.u2.b ;
assign { \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.u2.cout , \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.u2.s  } = _197_ + \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.u2.cin ;
assign _198_ = | op_0[15:3];
assign _199_ = op_0[15:3] != 13'h1fff;
assign _200_ = | trunc_ln851_1_reg_924;
assign _201_ = | ret_V_21_reg_918;
assign _202_ = | trunc_ln851_2_reg_1027;
assign _203_ = | trunc_ln851_reg_913;
assign _204_ = | op_10[9:0];
assign or_ln340_fu_480_p2 = p_Result_7_reg_970 | overflow_fu_465_p2;
assign or_ln785_1_fu_515_p2 = xor_ln785_1_fu_510_p2 | p_Result_7_reg_970;
assign or_ln785_fu_449_p2 = p_Result_8_reg_977 | icmp_ln768_reg_984;
assign or_ln786_fu_475_p2 = xor_ln786_fu_470_p2 | icmp_ln786_reg_989;
assign ret_V_19_fu_290_p2 = op_3 | { op_2, 7'h00 };
always @(posedge ap_clk)
select_ln703_reg_857[6:0] <= 7'h00;
always @(posedge ap_clk)
ret_V_21_reg_918[6:0] <= 7'h00;
always @(posedge ap_clk)
trunc_ln851_1_reg_924 <= 7'h00;
always @(posedge ap_clk)
select_ln1192_reg_960[4:2] <= 3'h0;
always @(posedge ap_clk)
p_Val2_s_reg_1006[0] <= 1'h0;
always @(posedge ap_clk)
select_ln340_reg_1011[0] <= 1'h0;
always @(posedge ap_clk)
op_1_V_reg_1016[0] <= 1'h0;
always @(posedge ap_clk)
select_ln703_reg_857[8:7] <= _047_;
always @(posedge ap_clk)
select_ln1347_reg_1082 <= _042_;
always @(posedge ap_clk)
select_ln1347_1_reg_1087 <= _041_;
always @(posedge ap_clk)
sext_ln850_reg_1092 <= _049_;
always @(posedge ap_clk)
select_ln69_2_reg_1099 <= _045_;
always @(posedge ap_clk)
ret_V_2_reg_891 <= _037_;
always @(posedge ap_clk)
ret_V_25_reg_1072 <= _034_;
always @(posedge ap_clk)
tmp_reg_1077 <= _051_;
always @(posedge ap_clk)
ret_V_24_reg_1042 <= _033_;
always @(posedge ap_clk)
select_ln69_reg_1047 <= _046_;
always @(posedge ap_clk)
ret_V_22_reg_954 <= _032_;
always @(posedge ap_clk)
select_ln1192_reg_960[1:0] <= _040_;
always @(posedge ap_clk)
ret_V_27_reg_1249 <= _036_;
always @(posedge ap_clk)
ret_V_21_cast_reg_1254 <= _030_;
always @(posedge ap_clk)
sext_ln353_reg_902 <= _048_;
always @(posedge ap_clk)
ret_V_19_reg_907 <= _029_;
always @(posedge ap_clk)
trunc_ln851_reg_913 <= _054_;
always @(posedge ap_clk)
ret_V_21_reg_918[7] <= _031_;
always @(posedge ap_clk)
ret_V_18_reg_896 <= _028_;
always @(posedge ap_clk)
ret_V_17_reg_879 <= _027_;
always @(posedge ap_clk)
ret_V_reg_884 <= _038_;
always @(posedge ap_clk)
p_Val2_s_reg_1006[3:1] <= _025_;
always @(posedge ap_clk)
select_ln340_reg_1011[3:1] <= _043_;
always @(posedge ap_clk)
or_ln785_reg_1000 <= _022_;
always @(posedge ap_clk)
op_30_V_reg_1229 <= _021_;
always @(posedge ap_clk)
op_21_V_reg_1052 <= _020_;
always @(posedge ap_clk)
op_1_V_reg_1016[3:1] <= _019_;
always @(posedge ap_clk)
shl_ln1299_reg_1021 <= _050_;
always @(posedge ap_clk)
trunc_ln851_2_reg_1027 <= _053_;
always @(posedge ap_clk)
icmp_ln851_reg_874 <= _017_;
always @(posedge ap_clk)
icmp_ln851_1_reg_1067 <= _016_;
always @(posedge ap_clk)
icmp_ln850_3_reg_1032 <= _014_;
always @(posedge ap_clk)
icmp_ln850_reg_939 <= _015_;
always @(posedge ap_clk)
icmp_ln850_1_reg_944 <= _012_;
always @(posedge ap_clk)
icmp_ln850_2_reg_949 <= _013_;
always @(posedge ap_clk)
trunc_ln703_reg_965 <= _052_;
always @(posedge ap_clk)
p_Result_7_reg_970 <= _023_;
always @(posedge ap_clk)
p_Result_8_reg_977 <= _024_;
always @(posedge ap_clk)
icmp_ln768_reg_984 <= _010_;
always @(posedge ap_clk)
icmp_ln786_reg_989 <= _011_;
always @(posedge ap_clk)
r_reg_995 <= _026_;
always @(posedge ap_clk)
op_14_V_reg_1124 <= _018_;
always @(posedge ap_clk)
ret_reg_1129 <= _039_;
always @(posedge ap_clk)
ret_V_26_reg_1134 <= _035_;
always @(posedge ap_clk)
select_ln69_1_reg_1139 <= _044_;
always @(posedge ap_clk)
add_ln69_4_reg_1144 <= _005_;
always @(posedge ap_clk)
add_ln69_2_reg_1214 <= _003_;
always @(posedge ap_clk)
add_ln69_6_reg_1219 <= _007_;
always @(posedge ap_clk)
add_ln69_reg_1179 <= _008_;
always @(posedge ap_clk)
add_ln69_1_reg_1184 <= _002_;
always @(posedge ap_clk)
add_ln69_3_reg_1189 <= _004_;
always @(posedge ap_clk)
add_ln69_5_reg_1194 <= _006_;
always @(posedge ap_clk)
add_ln691_reg_1114 <= _001_;
always @(posedge ap_clk)
add_ln691_1_reg_1261 <= _000_;
always @(posedge ap_clk)
ap_CS_fsm <= _009_;
assign _055_ = _059_ ? 2'h2 : 2'h1;
assign _205_ = ap_CS_fsm == 1'h1;
function [32:0] _592_;
input [32:0] a;
input [1088:0] b;
input [32:0] s;
case (s)
33'b000000000000000000000000000000001:
_592_ = b[32:0];
33'b000000000000000000000000000000010:
_592_ = b[65:33];
33'b000000000000000000000000000000100:
_592_ = b[98:66];
33'b000000000000000000000000000001000:
_592_ = b[131:99];
33'b000000000000000000000000000010000:
_592_ = b[164:132];
33'b000000000000000000000000000100000:
_592_ = b[197:165];
33'b000000000000000000000000001000000:
_592_ = b[230:198];
33'b000000000000000000000000010000000:
_592_ = b[263:231];
33'b000000000000000000000000100000000:
_592_ = b[296:264];
33'b000000000000000000000001000000000:
_592_ = b[329:297];
33'b000000000000000000000010000000000:
_592_ = b[362:330];
33'b000000000000000000000100000000000:
_592_ = b[395:363];
33'b000000000000000000001000000000000:
_592_ = b[428:396];
33'b000000000000000000010000000000000:
_592_ = b[461:429];
33'b000000000000000000100000000000000:
_592_ = b[494:462];
33'b000000000000000001000000000000000:
_592_ = b[527:495];
33'b000000000000000010000000000000000:
_592_ = b[560:528];
33'b000000000000000100000000000000000:
_592_ = b[593:561];
33'b000000000000001000000000000000000:
_592_ = b[626:594];
33'b000000000000010000000000000000000:
_592_ = b[659:627];
33'b000000000000100000000000000000000:
_592_ = b[692:660];
33'b000000000001000000000000000000000:
_592_ = b[725:693];
33'b000000000010000000000000000000000:
_592_ = b[758:726];
33'b000000000100000000000000000000000:
_592_ = b[791:759];
33'b000000001000000000000000000000000:
_592_ = b[824:792];
33'b000000010000000000000000000000000:
_592_ = b[857:825];
33'b000000100000000000000000000000000:
_592_ = b[890:858];
33'b000001000000000000000000000000000:
_592_ = b[923:891];
33'b000010000000000000000000000000000:
_592_ = b[956:924];
33'b000100000000000000000000000000000:
_592_ = b[989:957];
33'b001000000000000000000000000000000:
_592_ = b[1022:990];
33'b010000000000000000000000000000000:
_592_ = b[1055:1023];
33'b100000000000000000000000000000000:
_592_ = b[1088:1056];
33'b000000000000000000000000000000000:
_592_ = a;
default:
_592_ = 33'bx;
endcase
endfunction
assign ap_NS_fsm = _592_(33'hxxxxxxxxx, { 31'h00000000, _055_, 1056'h000000020000000200000002000000020000000200000002000000020000000200000002000000020000000200000002000000020000000200000002000000020000000200000002000000020000000200000002000000020000000200000002000000020000000200000002000000020000000200000002000000020000000000000001 }, { _205_, _237_, _236_, _235_, _234_, _233_, _232_, _231_, _230_, _229_, _228_, _227_, _226_, _225_, _224_, _223_, _222_, _221_, _220_, _219_, _218_, _217_, _216_, _215_, _214_, _213_, _212_, _211_, _210_, _209_, _208_, _207_, _206_ });
assign _206_ = ap_CS_fsm == 33'h100000000;
assign _207_ = ap_CS_fsm == 32'd2147483648;
assign _208_ = ap_CS_fsm == 31'h40000000;
assign _209_ = ap_CS_fsm == 30'h20000000;
assign _210_ = ap_CS_fsm == 29'h10000000;
assign _211_ = ap_CS_fsm == 28'h8000000;
assign _212_ = ap_CS_fsm == 27'h4000000;
assign _213_ = ap_CS_fsm == 26'h2000000;
assign _214_ = ap_CS_fsm == 25'h1000000;
assign _215_ = ap_CS_fsm == 24'h800000;
assign _216_ = ap_CS_fsm == 23'h400000;
assign _217_ = ap_CS_fsm == 22'h200000;
assign _218_ = ap_CS_fsm == 21'h100000;
assign _219_ = ap_CS_fsm == 20'h80000;
assign _220_ = ap_CS_fsm == 19'h40000;
assign _221_ = ap_CS_fsm == 18'h20000;
assign _222_ = ap_CS_fsm == 17'h10000;
assign _223_ = ap_CS_fsm == 16'h8000;
assign _224_ = ap_CS_fsm == 15'h4000;
assign _225_ = ap_CS_fsm == 14'h2000;
assign _226_ = ap_CS_fsm == 13'h1000;
assign _227_ = ap_CS_fsm == 12'h800;
assign _228_ = ap_CS_fsm == 11'h400;
assign _229_ = ap_CS_fsm == 10'h200;
assign _230_ = ap_CS_fsm == 9'h100;
assign _231_ = ap_CS_fsm == 8'h80;
assign _232_ = ap_CS_fsm == 7'h40;
assign _233_ = ap_CS_fsm == 6'h20;
assign _234_ = ap_CS_fsm == 5'h10;
assign _235_ = ap_CS_fsm == 4'h8;
assign _236_ = ap_CS_fsm == 3'h4;
assign _237_ = ap_CS_fsm == 2'h2;
assign op_31_ap_vld = ap_CS_fsm[32] ? 1'h1 : 1'h0;
assign ap_idle = _058_ ? 1'h1 : 1'h0;
assign _047_ = ap_CS_fsm[0] ? select_ln703_fu_219_p3[8:7] : select_ln703_reg_857[8:7];
assign _045_ = ap_CS_fsm[19] ? select_ln69_2_fu_655_p3 : select_ln69_2_reg_1099;
assign _049_ = ap_CS_fsm[19] ? { tmp_reg_1077[6], tmp_reg_1077 } : sext_ln850_reg_1092;
assign _041_ = ap_CS_fsm[19] ? select_ln1347_1_fu_639_p3 : select_ln1347_1_reg_1087;
assign _042_ = ap_CS_fsm[19] ? select_ln1347_fu_632_p3 : select_ln1347_reg_1082;
assign _037_ = _057_ ? grp_fu_256_p2 : ret_V_2_reg_891;
assign _051_ = ap_CS_fsm[18] ? grp_fu_606_p2[16:10] : tmp_reg_1077;
assign _034_ = ap_CS_fsm[18] ? grp_fu_606_p2 : ret_V_25_reg_1072;
assign _046_ = ap_CS_fsm[14] ? select_ln69_fu_579_p3 : select_ln69_reg_1047;
assign _033_ = ap_CS_fsm[14] ? grp_fu_549_p2 : ret_V_24_reg_1042;
assign _040_ = ap_CS_fsm[8] ? select_ln1192_fu_378_p3 : select_ln1192_reg_960[1:0];
assign _032_ = ap_CS_fsm[8] ? ret_V_22_fu_372_p2 : ret_V_22_reg_954;
assign _030_ = ap_CS_fsm[29] ? grp_fu_806_p2[32:1] : ret_V_21_cast_reg_1254;
assign _036_ = ap_CS_fsm[29] ? grp_fu_806_p2 : ret_V_27_reg_1249;
assign _031_ = ap_CS_fsm[6] ? ret_V_21_fu_299_p2[7] : ret_V_21_reg_918[7];
assign _054_ = ap_CS_fsm[6] ? ret_V_19_fu_290_p2[6:0] : trunc_ln851_reg_913;
assign _029_ = ap_CS_fsm[6] ? ret_V_19_fu_290_p2 : ret_V_19_reg_907;
assign _048_ = ap_CS_fsm[6] ? { ret_V_18_reg_896[1], ret_V_18_reg_896[1], ret_V_18_reg_896[1], ret_V_18_reg_896[1], ret_V_18_reg_896[1], ret_V_18_reg_896[1], ret_V_18_reg_896 } : sext_ln353_reg_902;
assign _028_ = ap_CS_fsm[5] ? ret_V_18_fu_273_p3 : ret_V_18_reg_896;
assign _038_ = ap_CS_fsm[2] ? grp_fu_235_p2[8:7] : ret_V_reg_884;
assign _027_ = ap_CS_fsm[2] ? grp_fu_235_p2 : ret_V_17_reg_879;
assign _043_ = ap_CS_fsm[11] ? select_ln340_fu_497_p3[3:1] : select_ln340_reg_1011[3:1];
assign _025_ = ap_CS_fsm[11] ? trunc_ln703_reg_965 : p_Val2_s_reg_1006[3:1];
assign _022_ = ap_CS_fsm[10] ? or_ln785_fu_449_p2 : or_ln785_reg_1000;
assign _021_ = ap_CS_fsm[27] ? grp_fu_786_p2 : op_30_V_reg_1229;
assign _020_ = ap_CS_fsm[16] ? grp_fu_587_p2 : op_21_V_reg_1052;
assign _053_ = ap_CS_fsm[12] ? grp_fu_315_p2[6:0] : trunc_ln851_2_reg_1027;
assign _050_ = ap_CS_fsm[12] ? grp_fu_315_p2 : shl_ln1299_reg_1021;
assign _019_ = ap_CS_fsm[12] ? op_1_V_fu_531_p3[3:1] : op_1_V_reg_1016[3:1];
assign _017_ = ap_CS_fsm[1] ? icmp_ln851_fu_240_p2 : icmp_ln851_reg_874;
assign _016_ = ap_CS_fsm[17] ? icmp_ln851_1_fu_616_p2 : icmp_ln851_1_reg_1067;
assign _014_ = ap_CS_fsm[13] ? icmp_ln850_3_fu_541_p2 : icmp_ln850_3_reg_1032;
assign _013_ = ap_CS_fsm[7] ? icmp_ln850_2_fu_331_p2 : icmp_ln850_2_reg_949;
assign _012_ = ap_CS_fsm[7] ? icmp_ln850_1_fu_326_p2 : icmp_ln850_1_reg_944;
assign _015_ = ap_CS_fsm[7] ? icmp_ln850_fu_321_p2 : icmp_ln850_reg_939;
assign _026_ = ap_CS_fsm[9] ? r_fu_443_p3 : r_reg_995;
assign _011_ = ap_CS_fsm[9] ? icmp_ln786_fu_422_p2 : icmp_ln786_reg_989;
assign _010_ = ap_CS_fsm[9] ? icmp_ln768_fu_416_p2 : icmp_ln768_reg_984;
assign _024_ = ap_CS_fsm[9] ? op_0[2] : p_Result_8_reg_977;
assign _023_ = ap_CS_fsm[9] ? op_0[15] : p_Result_7_reg_970;
assign _052_ = ap_CS_fsm[9] ? op_0[2:0] : trunc_ln703_reg_965;
assign _005_ = ap_CS_fsm[21] ? grp_fu_685_p2 : add_ln69_4_reg_1144;
assign _044_ = ap_CS_fsm[21] ? select_ln69_1_fu_709_p3 : select_ln69_1_reg_1139;
assign _035_ = ap_CS_fsm[21] ? ret_V_26_fu_702_p3 : ret_V_26_reg_1134;
assign _039_ = ap_CS_fsm[21] ? grp_fu_677_p2 : ret_reg_1129;
assign _018_ = ap_CS_fsm[21] ? grp_fu_671_p2 : op_14_V_reg_1124;
assign _007_ = ap_CS_fsm[25] ? grp_fu_777_p2 : add_ln69_6_reg_1219;
assign _003_ = ap_CS_fsm[25] ? grp_fu_766_p2 : add_ln69_2_reg_1214;
assign _006_ = ap_CS_fsm[23] ? grp_fu_759_p2 : add_ln69_5_reg_1194;
assign _004_ = ap_CS_fsm[23] ? grp_fu_753_p2 : add_ln69_3_reg_1189;
assign _002_ = ap_CS_fsm[23] ? grp_fu_747_p2 : add_ln69_1_reg_1184;
assign _008_ = ap_CS_fsm[23] ? grp_fu_741_p2 : add_ln69_reg_1179;
assign _001_ = _056_ ? grp_fu_649_p2 : add_ln691_reg_1114;
assign _000_ = ap_CS_fsm[31] ? grp_fu_822_p2 : add_ln691_1_reg_1261;
assign _009_ = ap_rst ? 33'h000000001 : ap_NS_fsm;
assign icmp_ln768_fu_416_p2 = _198_ ? 1'h1 : 1'h0;
assign icmp_ln786_fu_422_p2 = _199_ ? 1'h1 : 1'h0;
assign icmp_ln850_1_fu_326_p2 = _200_ ? 1'h1 : 1'h0;
assign icmp_ln850_2_fu_331_p2 = _201_ ? 1'h1 : 1'h0;
assign icmp_ln850_3_fu_541_p2 = _202_ ? 1'h1 : 1'h0;
assign icmp_ln850_fu_321_p2 = _203_ ? 1'h1 : 1'h0;
assign icmp_ln851_1_fu_616_p2 = _204_ ? 1'h1 : 1'h0;
assign icmp_ln851_fu_240_p2 = _062_ ? 1'h1 : 1'h0;
assign op_1_V_fu_531_p3 = and_ln785_1_fu_526_p2 ? p_Val2_s_reg_1006 : select_ln340_reg_1011;
assign op_31 = ret_V_27_reg_1249[33] ? select_ln850_2_fu_837_p3 : ret_V_21_cast_reg_1254;
assign r_fu_443_p3 = ret_V_22_reg_954 ? { 1'h0, select_ln850_4_fu_435_p3 } : sext_ln353_reg_902;
assign ret_V_18_fu_273_p3 = ret_V_17_reg_879[8] ? select_ln850_fu_268_p3 : ret_V_reg_884;
assign ret_V_26_fu_702_p3 = ret_V_25_reg_1072[16] ? select_ln850_1_fu_697_p3 : sext_ln850_reg_1092;
assign select_ln1192_fu_378_p3 = ret_V_20_fu_355_p2 ? 2'h3 : 2'h0;
assign select_ln1347_1_fu_639_p3 = ret_V_22_reg_954 ? 2'h3 : 2'h0;
assign select_ln1347_fu_632_p3 = op_2 ? 2'h3 : 2'h0;
assign select_ln340_fu_497_p3 = and_ln340_fu_491_p2 ? { trunc_ln703_reg_965, 1'h0 } : 4'h0;
assign select_ln69_1_fu_709_p3 = op_11 ? 2'h3 : 2'h0;
assign select_ln69_2_fu_655_p3 = op_18 ? 2'h3 : 2'h0;
assign select_ln69_fu_579_p3 = ret_V_23_fu_573_p2 ? 5'h1f : 5'h00;
assign select_ln703_fu_219_p3 = op_2 ? 9'h180 : 9'h000;
assign select_ln850_1_fu_697_p3 = icmp_ln851_1_reg_1067 ? add_ln691_reg_1114 : sext_ln850_reg_1092;
assign select_ln850_2_fu_837_p3 = op_19[0] ? add_ln691_1_reg_1261 : ret_V_21_cast_reg_1254;
assign select_ln850_4_fu_435_p3 = ret_V_18_reg_896[1] ? 7'h7f : 7'h00;
assign select_ln850_fu_268_p3 = icmp_ln851_reg_874 ? ret_V_reg_884 : ret_V_2_reg_891;
assign ret_V_20_fu_355_p2 = ret_V_19_reg_907[7] ^ and_ln850_fu_350_p2;
assign ret_V_22_fu_372_p2 = ret_V_21_reg_918[7] ^ and_ln850_1_fu_368_p2;
assign ret_V_23_fu_573_p2 = shl_ln1299_reg_1021[7] ^ and_ln850_2_fu_568_p2;
assign ap_CS_fsm_state1 = ap_CS_fsm[0];
assign ap_CS_fsm_state10 = ap_CS_fsm[9];
assign ap_CS_fsm_state11 = ap_CS_fsm[10];
assign ap_CS_fsm_state12 = ap_CS_fsm[11];
assign ap_CS_fsm_state13 = ap_CS_fsm[12];
assign ap_CS_fsm_state14 = ap_CS_fsm[13];
assign ap_CS_fsm_state15 = ap_CS_fsm[14];
assign ap_CS_fsm_state16 = ap_CS_fsm[15];
assign ap_CS_fsm_state17 = ap_CS_fsm[16];
assign ap_CS_fsm_state18 = ap_CS_fsm[17];
assign ap_CS_fsm_state19 = ap_CS_fsm[18];
assign ap_CS_fsm_state2 = ap_CS_fsm[1];
assign ap_CS_fsm_state20 = ap_CS_fsm[19];
assign ap_CS_fsm_state21 = ap_CS_fsm[20];
assign ap_CS_fsm_state22 = ap_CS_fsm[21];
assign ap_CS_fsm_state23 = ap_CS_fsm[22];
assign ap_CS_fsm_state24 = ap_CS_fsm[23];
assign ap_CS_fsm_state25 = ap_CS_fsm[24];
assign ap_CS_fsm_state26 = ap_CS_fsm[25];
assign ap_CS_fsm_state27 = ap_CS_fsm[26];
assign ap_CS_fsm_state28 = ap_CS_fsm[27];
assign ap_CS_fsm_state29 = ap_CS_fsm[28];
assign ap_CS_fsm_state3 = ap_CS_fsm[2];
assign ap_CS_fsm_state30 = ap_CS_fsm[29];
assign ap_CS_fsm_state31 = ap_CS_fsm[30];
assign ap_CS_fsm_state32 = ap_CS_fsm[31];
assign ap_CS_fsm_state33 = ap_CS_fsm[32];
assign ap_CS_fsm_state4 = ap_CS_fsm[3];
assign ap_CS_fsm_state5 = ap_CS_fsm[4];
assign ap_CS_fsm_state6 = ap_CS_fsm[5];
assign ap_CS_fsm_state7 = ap_CS_fsm[6];
assign ap_CS_fsm_state8 = ap_CS_fsm[7];
assign ap_CS_fsm_state9 = ap_CS_fsm[8];
assign ap_done = op_31_ap_vld;
assign ap_ready = op_31_ap_vld;
assign grp_fu_235_p1 = { op_3[7], op_3 };
assign grp_fu_315_p0 = { op_3[7], op_3[7], op_3[7], op_3[7], op_3[7], op_3[7], op_3[7], op_3[7], op_3[7], op_3[7], op_3[7], op_3[7], op_3[7], op_3[7], op_3[7], op_3[7], op_3[7], op_3[7], op_3[7], op_3[7], op_3[7], op_3[7], op_3[7], op_3[7], op_3 };
assign grp_fu_315_p1 = { 24'h000000, ret_V_18_reg_896[1], ret_V_18_reg_896[1], ret_V_18_reg_896[1], ret_V_18_reg_896[1], ret_V_18_reg_896[1], ret_V_18_reg_896[1], ret_V_18_reg_896 };
assign grp_fu_549_p1 = { op_1_V_reg_1016[3], op_1_V_reg_1016 };
assign grp_fu_606_p0 = { op_21_V_reg_1052[4], op_21_V_reg_1052[4], op_21_V_reg_1052, 10'h000 };
assign grp_fu_606_p1 = { op_10[15], op_10 };
assign grp_fu_649_p0 = { tmp_reg_1077[6], tmp_reg_1077 };
assign grp_fu_671_p0 = { op_6[1], op_6[1], op_6 };
assign grp_fu_671_p1 = op_7[3:0];
assign grp_fu_685_p1 = { 1'h0, op_12 };
assign grp_fu_741_p0 = { ret_V_26_reg_1134[7], ret_V_26_reg_1134[7], ret_V_26_reg_1134 };
assign grp_fu_741_p1 = { 2'h0, r_reg_995 };
assign grp_fu_747_p0 = { op_14_V_reg_1124[3], op_14_V_reg_1124 };
assign grp_fu_747_p1 = { op_16[3], op_16 };
assign grp_fu_753_p0 = { 1'h0, ret_reg_1129[1], ret_reg_1129[1], ret_reg_1129 };
assign grp_fu_753_p1 = { 3'h0, op_17 };
assign grp_fu_766_p0 = { add_ln69_1_reg_1184[4], add_ln69_1_reg_1184[4], add_ln69_1_reg_1184[4], add_ln69_1_reg_1184[4], add_ln69_1_reg_1184[4], add_ln69_1_reg_1184 };
assign grp_fu_777_p0 = { add_ln69_5_reg_1194[1], add_ln69_5_reg_1194[1], add_ln69_5_reg_1194[1], add_ln69_5_reg_1194[1], add_ln69_5_reg_1194 };
assign grp_fu_777_p1 = { 1'h0, add_ln69_3_reg_1189 };
assign grp_fu_786_p0 = { add_ln69_6_reg_1219[5], add_ln69_6_reg_1219[5], add_ln69_6_reg_1219[5], add_ln69_6_reg_1219[5], add_ln69_6_reg_1219 };
assign grp_fu_806_p0 = { op_30_V_reg_1229[9], op_30_V_reg_1229[9], op_30_V_reg_1229[9], op_30_V_reg_1229[9], op_30_V_reg_1229[9], op_30_V_reg_1229[9], op_30_V_reg_1229[9], op_30_V_reg_1229[9], op_30_V_reg_1229[9], op_30_V_reg_1229[9], op_30_V_reg_1229[9], op_30_V_reg_1229[9], op_30_V_reg_1229[9], op_30_V_reg_1229[9], op_30_V_reg_1229[9], op_30_V_reg_1229[9], op_30_V_reg_1229[9], op_30_V_reg_1229[9], op_30_V_reg_1229[9], op_30_V_reg_1229[9], op_30_V_reg_1229[9], op_30_V_reg_1229[9], op_30_V_reg_1229[9], op_30_V_reg_1229, 1'h0 };
assign grp_fu_806_p1 = { op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19 };
assign lhs_fu_283_p3 = { op_2, 7'h00 };
assign p_Result_1_fu_343_p3 = ret_V_19_reg_907[7];
assign p_Result_2_fu_561_p3 = shl_ln1299_reg_1021[7];
assign p_Result_5_fu_690_p3 = ret_V_25_reg_1072[16];
assign p_Result_6_fu_827_p3 = ret_V_27_reg_1249[33];
assign p_Result_s_12_fu_261_p3 = ret_V_17_reg_879[8];
assign p_Result_s_fu_406_p4 = op_0[15:3];
assign p_Val2_s_fu_453_p3 = { trunc_ln703_reg_965, 1'h0 };
assign ret_V_10_fu_554_p3 = shl_ln1299_reg_1021[7];
assign ret_V_19_fu_290_p1 = op_3;
assign ret_V_21_fu_299_p1 = op_3;
assign ret_V_5_fu_336_p3 = ret_V_19_reg_907[7];
assign ret_V_8_fu_361_p3 = ret_V_21_reg_918[7];
assign rhs_2_fu_595_p3 = { op_21_V_reg_1052, 10'h000 };
assign sext_ln1192_fu_591_p0 = op_10;
assign sext_ln1299_fu_312_p0 = op_3;
assign sext_ln353_fu_280_p1 = { ret_V_18_reg_896[1], ret_V_18_reg_896[1], ret_V_18_reg_896[1], ret_V_18_reg_896[1], ret_V_18_reg_896[1], ret_V_18_reg_896[1], ret_V_18_reg_896 };
assign sext_ln69_1_fu_720_p1 = { ret_reg_1129[1], ret_reg_1129[1], ret_reg_1129 };
assign sext_ln703_2_fu_791_p0 = op_19;
assign sext_ln703_fu_227_p0 = op_3;
assign sext_ln850_fu_646_p1 = { tmp_reg_1077[6], tmp_reg_1077 };
assign tmp_11_fu_795_p3 = { op_30_V_reg_1229, 1'h0 };
assign tmp_9_fu_428_p3 = ret_V_18_reg_896[1];
assign trunc_ln1192_fu_231_p0 = op_3;
assign trunc_ln1192_fu_231_p1 = op_3[6:0];
assign trunc_ln703_fu_386_p1 = op_0[2:0];
assign trunc_ln851_1_fu_304_p1 = ret_V_21_fu_299_p2[6:0];
assign trunc_ln851_2_fu_537_p1 = grp_fu_315_p2[6:0];
assign trunc_ln851_3_fu_612_p0 = op_10;
assign trunc_ln851_3_fu_612_p1 = op_10[9:0];
assign trunc_ln851_4_fu_834_p0 = op_19;
assign trunc_ln851_4_fu_834_p1 = op_19[0];
assign trunc_ln851_fu_295_p1 = ret_V_19_fu_290_p2[6:0];
assign \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.ain_s0  = \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.a ;
assign \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.s  = { \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.fas_s2 , \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.sum_s1  };
assign \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.u2.a  = \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.ain_s1 ;
assign \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.u2.b  = \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.bin_s1 ;
assign \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.u2.cin  = \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.carry_s1 ;
assign \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.facout_s2  = \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.u2.cout ;
assign \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.fas_s2  = \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.u2.s ;
assign \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.u1.a  = \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.a [1:0];
assign \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.u1.b  = \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.bin_s0 [1:0];
assign \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.u1.cin  = 1'h1;
assign \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.facout_s1  = \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.u1.cout ;
assign \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.fas_s1  = \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.u1.s ;
assign \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.a  = \sub_4s_4ns_4_2_1_U8.din0 ;
assign \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.b  = \sub_4s_4ns_4_2_1_U8.din1 ;
assign \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.ce  = \sub_4s_4ns_4_2_1_U8.ce ;
assign \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.clk  = \sub_4s_4ns_4_2_1_U8.clk ;
assign \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.reset  = \sub_4s_4ns_4_2_1_U8.reset ;
assign \sub_4s_4ns_4_2_1_U8.dout  = \sub_4s_4ns_4_2_1_U8.top_sub_4s_4ns_4_2_1_Adder_6_U.s ;
assign \sub_4s_4ns_4_2_1_U8.ce  = 1'h1;
assign \sub_4s_4ns_4_2_1_U8.clk  = ap_clk;
assign \sub_4s_4ns_4_2_1_U8.din0  = { op_6[1], op_6[1], op_6 };
assign \sub_4s_4ns_4_2_1_U8.din1  = op_7[3:0];
assign grp_fu_671_p2 = \sub_4s_4ns_4_2_1_U8.dout ;
assign \sub_4s_4ns_4_2_1_U8.reset  = ap_rst;
assign \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.ain_s0  = \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.a ;
assign \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.s  = { \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.fas_s2 , \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.sum_s1  };
assign \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.u2.a  = \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.ain_s1 ;
assign \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.u2.b  = \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.bin_s1 ;
assign \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.u2.cin  = \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.carry_s1 ;
assign \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.facout_s2  = \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.u2.cout ;
assign \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.fas_s2  = \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.u2.s ;
assign \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.u1.a  = \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.a [0];
assign \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.u1.b  = \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.bin_s0 [0];
assign \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.u1.cin  = 1'h1;
assign \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.facout_s1  = \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.u1.cout ;
assign \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.fas_s1  = \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.u1.s ;
assign \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.a  = \sub_2ns_2ns_2_2_1_U9.din0 ;
assign \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.b  = \sub_2ns_2ns_2_2_1_U9.din1 ;
assign \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.ce  = \sub_2ns_2ns_2_2_1_U9.ce ;
assign \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.clk  = \sub_2ns_2ns_2_2_1_U9.clk ;
assign \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.reset  = \sub_2ns_2ns_2_2_1_U9.reset ;
assign \sub_2ns_2ns_2_2_1_U9.dout  = \sub_2ns_2ns_2_2_1_U9.top_sub_2ns_2ns_2_2_1_Adder_7_U.s ;
assign \sub_2ns_2ns_2_2_1_U9.ce  = 1'h1;
assign \sub_2ns_2ns_2_2_1_U9.clk  = ap_clk;
assign \sub_2ns_2ns_2_2_1_U9.din0  = select_ln1347_reg_1082;
assign \sub_2ns_2ns_2_2_1_U9.din1  = select_ln1347_1_reg_1087;
assign grp_fu_677_p2 = \sub_2ns_2ns_2_2_1_U9.dout ;
assign \sub_2ns_2ns_2_2_1_U9.reset  = ap_rst;
assign \shl_32s_8ns_32_7_1_U3.din1_cast  = \shl_32s_8ns_32_7_1_U3.din1 [7:0];
assign \shl_32s_8ns_32_7_1_U3.din1_mask  = 8'h03;
assign \shl_32s_8ns_32_7_1_U3.ce  = 1'h1;
assign \shl_32s_8ns_32_7_1_U3.clk  = ap_clk;
assign \shl_32s_8ns_32_7_1_U3.din0  = { op_3[7], op_3[7], op_3[7], op_3[7], op_3[7], op_3[7], op_3[7], op_3[7], op_3[7], op_3[7], op_3[7], op_3[7], op_3[7], op_3[7], op_3[7], op_3[7], op_3[7], op_3[7], op_3[7], op_3[7], op_3[7], op_3[7], op_3[7], op_3[7], op_3 };
assign \shl_32s_8ns_32_7_1_U3.din1  = { 24'h000000, ret_V_18_reg_896[1], ret_V_18_reg_896[1], ret_V_18_reg_896[1], ret_V_18_reg_896[1], ret_V_18_reg_896[1], ret_V_18_reg_896[1], ret_V_18_reg_896 };
assign grp_fu_315_p2 = \shl_32s_8ns_32_7_1_U3.dout ;
assign \shl_32s_8ns_32_7_1_U3.reset  = ap_rst;
assign \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.ain_s0  = \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.a ;
assign \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.bin_s0  = \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.b ;
assign \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.s  = { \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.fas_s2 , \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.sum_s1  };
assign \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.u2.a  = \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.ain_s1 ;
assign \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.u2.b  = \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.bin_s1 ;
assign \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.u2.cin  = \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.carry_s1 ;
assign \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.facout_s2  = \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.u2.cout ;
assign \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.fas_s2  = \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.u2.s ;
assign \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.u1.a  = \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.a [3:0];
assign \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.u1.b  = \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.b [3:0];
assign \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.u1.cin  = 1'h0;
assign \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.facout_s1  = \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.u1.cout ;
assign \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.fas_s1  = \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.u1.s ;
assign \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.a  = \add_9ns_9s_9_2_1_U1.din0 ;
assign \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.b  = \add_9ns_9s_9_2_1_U1.din1 ;
assign \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.ce  = \add_9ns_9s_9_2_1_U1.ce ;
assign \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.clk  = \add_9ns_9s_9_2_1_U1.clk ;
assign \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.reset  = \add_9ns_9s_9_2_1_U1.reset ;
assign \add_9ns_9s_9_2_1_U1.dout  = \add_9ns_9s_9_2_1_U1.top_add_9ns_9s_9_2_1_Adder_0_U.s ;
assign \add_9ns_9s_9_2_1_U1.ce  = 1'h1;
assign \add_9ns_9s_9_2_1_U1.clk  = ap_clk;
assign \add_9ns_9s_9_2_1_U1.din0  = select_ln703_reg_857;
assign \add_9ns_9s_9_2_1_U1.din1  = { op_3[7], op_3 };
assign grp_fu_235_p2 = \add_9ns_9s_9_2_1_U1.dout ;
assign \add_9ns_9s_9_2_1_U1.reset  = ap_rst;
assign \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.ain_s0  = \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.a ;
assign \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.bin_s0  = \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.b ;
assign \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.s  = { \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.fas_s2 , \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.sum_s1  };
assign \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.u2.a  = \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.ain_s1 ;
assign \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.u2.b  = \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.bin_s1 ;
assign \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.u2.cin  = \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.carry_s1 ;
assign \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.facout_s2  = \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.u2.cout ;
assign \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.fas_s2  = \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.u2.s ;
assign \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.u1.a  = \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.a [3:0];
assign \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.u1.b  = \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.b [3:0];
assign \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.u1.cin  = 1'h0;
assign \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.facout_s1  = \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.u1.cout ;
assign \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.fas_s1  = \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.u1.s ;
assign \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.a  = \add_8s_8ns_8_2_1_U7.din0 ;
assign \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.b  = \add_8s_8ns_8_2_1_U7.din1 ;
assign \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.ce  = \add_8s_8ns_8_2_1_U7.ce ;
assign \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.clk  = \add_8s_8ns_8_2_1_U7.clk ;
assign \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.reset  = \add_8s_8ns_8_2_1_U7.reset ;
assign \add_8s_8ns_8_2_1_U7.dout  = \add_8s_8ns_8_2_1_U7.top_add_8s_8ns_8_2_1_Adder_5_U.s ;
assign \add_8s_8ns_8_2_1_U7.ce  = 1'h1;
assign \add_8s_8ns_8_2_1_U7.clk  = ap_clk;
assign \add_8s_8ns_8_2_1_U7.din0  = { tmp_reg_1077[6], tmp_reg_1077 };
assign \add_8s_8ns_8_2_1_U7.din1  = 8'h01;
assign grp_fu_649_p2 = \add_8s_8ns_8_2_1_U7.dout ;
assign \add_8s_8ns_8_2_1_U7.reset  = ap_rst;
assign \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.ain_s0  = \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.a ;
assign \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.bin_s0  = \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.b ;
assign \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.s  = { \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.fas_s2 , \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.sum_s1  };
assign \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.u2.a  = \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.ain_s1 ;
assign \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.u2.b  = \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.bin_s1 ;
assign \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.u2.cin  = \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.carry_s1 ;
assign \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.facout_s2  = \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.u2.cout ;
assign \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.fas_s2  = \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.u2.s ;
assign \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.u1.a  = \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.a [2:0];
assign \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.u1.b  = \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.b [2:0];
assign \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.u1.cin  = 1'h0;
assign \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.facout_s1  = \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.u1.cout ;
assign \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.fas_s1  = \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.u1.s ;
assign \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.a  = \add_6s_6ns_6_2_1_U16.din0 ;
assign \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.b  = \add_6s_6ns_6_2_1_U16.din1 ;
assign \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.ce  = \add_6s_6ns_6_2_1_U16.ce ;
assign \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.clk  = \add_6s_6ns_6_2_1_U16.clk ;
assign \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.reset  = \add_6s_6ns_6_2_1_U16.reset ;
assign \add_6s_6ns_6_2_1_U16.dout  = \add_6s_6ns_6_2_1_U16.top_add_6s_6ns_6_2_1_Adder_10_U.s ;
assign \add_6s_6ns_6_2_1_U16.ce  = 1'h1;
assign \add_6s_6ns_6_2_1_U16.clk  = ap_clk;
assign \add_6s_6ns_6_2_1_U16.din0  = { add_ln69_5_reg_1194[1], add_ln69_5_reg_1194[1], add_ln69_5_reg_1194[1], add_ln69_5_reg_1194[1], add_ln69_5_reg_1194 };
assign \add_6s_6ns_6_2_1_U16.din1  = { 1'h0, add_ln69_3_reg_1189 };
assign grp_fu_777_p2 = \add_6s_6ns_6_2_1_U16.dout ;
assign \add_6s_6ns_6_2_1_U16.reset  = ap_rst;
assign \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.ain_s0  = \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.a ;
assign \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.bin_s0  = \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.b ;
assign \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.s  = { \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.fas_s2 , \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.sum_s1  };
assign \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.u2.a  = \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.ain_s1 ;
assign \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.u2.b  = \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.bin_s1 ;
assign \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.u2.cin  = \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.carry_s1 ;
assign \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.facout_s2  = \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.u2.cout ;
assign \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.fas_s2  = \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.u2.s ;
assign \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.u1.a  = \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.a [1:0];
assign \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.u1.b  = \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.b [1:0];
assign \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.u1.cin  = 1'h0;
assign \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.facout_s1  = \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.u1.cout ;
assign \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.fas_s1  = \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.u1.s ;
assign \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.a  = \add_5s_5s_5_2_1_U12.din0 ;
assign \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.b  = \add_5s_5s_5_2_1_U12.din1 ;
assign \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.ce  = \add_5s_5s_5_2_1_U12.ce ;
assign \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.clk  = \add_5s_5s_5_2_1_U12.clk ;
assign \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.reset  = \add_5s_5s_5_2_1_U12.reset ;
assign \add_5s_5s_5_2_1_U12.dout  = \add_5s_5s_5_2_1_U12.top_add_5s_5s_5_2_1_Adder_9_U.s ;
assign \add_5s_5s_5_2_1_U12.ce  = 1'h1;
assign \add_5s_5s_5_2_1_U12.clk  = ap_clk;
assign \add_5s_5s_5_2_1_U12.din0  = { op_14_V_reg_1124[3], op_14_V_reg_1124 };
assign \add_5s_5s_5_2_1_U12.din1  = { op_16[3], op_16 };
assign grp_fu_747_p2 = \add_5s_5s_5_2_1_U12.dout ;
assign \add_5s_5s_5_2_1_U12.reset  = ap_rst;
assign \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.ain_s0  = \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.a ;
assign \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.bin_s0  = \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.b ;
assign \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.s  = { \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.fas_s2 , \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.sum_s1  };
assign \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.u2.a  = \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.ain_s1 ;
assign \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.u2.b  = \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.bin_s1 ;
assign \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.u2.cin  = \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.carry_s1 ;
assign \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.facout_s2  = \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.u2.cout ;
assign \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.fas_s2  = \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.u2.s ;
assign \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.u1.a  = \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.a [1:0];
assign \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.u1.b  = \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.b [1:0];
assign \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.u1.cin  = 1'h0;
assign \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.facout_s1  = \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.u1.cout ;
assign \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.fas_s1  = \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.u1.s ;
assign \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.a  = \add_5ns_5s_5_2_1_U4.din0 ;
assign \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.b  = \add_5ns_5s_5_2_1_U4.din1 ;
assign \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.ce  = \add_5ns_5s_5_2_1_U4.ce ;
assign \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.clk  = \add_5ns_5s_5_2_1_U4.clk ;
assign \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.reset  = \add_5ns_5s_5_2_1_U4.reset ;
assign \add_5ns_5s_5_2_1_U4.dout  = \add_5ns_5s_5_2_1_U4.top_add_5ns_5s_5_2_1_Adder_2_U.s ;
assign \add_5ns_5s_5_2_1_U4.ce  = 1'h1;
assign \add_5ns_5s_5_2_1_U4.clk  = ap_clk;
assign \add_5ns_5s_5_2_1_U4.din0  = select_ln1192_reg_960;
assign \add_5ns_5s_5_2_1_U4.din1  = { op_1_V_reg_1016[3], op_1_V_reg_1016 };
assign grp_fu_549_p2 = \add_5ns_5s_5_2_1_U4.dout ;
assign \add_5ns_5s_5_2_1_U4.reset  = ap_rst;
assign \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.ain_s0  = \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.a ;
assign \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.bin_s0  = \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.b ;
assign \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.s  = { \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.fas_s2 , \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.sum_s1  };
assign \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.u2.a  = \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.ain_s1 ;
assign \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.u2.b  = \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.bin_s1 ;
assign \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.u2.cin  = \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.carry_s1 ;
assign \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.facout_s2  = \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.u2.cout ;
assign \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.fas_s2  = \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.u2.s ;
assign \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.u1.a  = \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.a [1:0];
assign \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.u1.b  = \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.b [1:0];
assign \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.u1.cin  = 1'h0;
assign \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.facout_s1  = \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.u1.cout ;
assign \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.fas_s1  = \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.u1.s ;
assign \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.a  = \add_5ns_5ns_5_2_1_U5.din0 ;
assign \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.b  = \add_5ns_5ns_5_2_1_U5.din1 ;
assign \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.ce  = \add_5ns_5ns_5_2_1_U5.ce ;
assign \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.clk  = \add_5ns_5ns_5_2_1_U5.clk ;
assign \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.reset  = \add_5ns_5ns_5_2_1_U5.reset ;
assign \add_5ns_5ns_5_2_1_U5.dout  = \add_5ns_5ns_5_2_1_U5.top_add_5ns_5ns_5_2_1_Adder_3_U.s ;
assign \add_5ns_5ns_5_2_1_U5.ce  = 1'h1;
assign \add_5ns_5ns_5_2_1_U5.clk  = ap_clk;
assign \add_5ns_5ns_5_2_1_U5.din0  = ret_V_24_reg_1042;
assign \add_5ns_5ns_5_2_1_U5.din1  = select_ln69_reg_1047;
assign grp_fu_587_p2 = \add_5ns_5ns_5_2_1_U5.dout ;
assign \add_5ns_5ns_5_2_1_U5.reset  = ap_rst;
assign \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.ain_s0  = \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.a ;
assign \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.bin_s0  = \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.b ;
assign \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.s  = { \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.fas_s2 , \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.sum_s1  };
assign \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.u2.a  = \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.ain_s1 ;
assign \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.u2.b  = \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.bin_s1 ;
assign \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.u2.cin  = \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.carry_s1 ;
assign \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.facout_s2  = \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.u2.cout ;
assign \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.fas_s2  = \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.u2.s ;
assign \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.u1.a  = \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.a [1:0];
assign \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.u1.b  = \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.b [1:0];
assign \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.u1.cin  = 1'h0;
assign \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.facout_s1  = \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.u1.cout ;
assign \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.fas_s1  = \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.u1.s ;
assign \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.a  = \add_5ns_5ns_5_2_1_U13.din0 ;
assign \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.b  = \add_5ns_5ns_5_2_1_U13.din1 ;
assign \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.ce  = \add_5ns_5ns_5_2_1_U13.ce ;
assign \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.clk  = \add_5ns_5ns_5_2_1_U13.clk ;
assign \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.reset  = \add_5ns_5ns_5_2_1_U13.reset ;
assign \add_5ns_5ns_5_2_1_U13.dout  = \add_5ns_5ns_5_2_1_U13.top_add_5ns_5ns_5_2_1_Adder_3_U.s ;
assign \add_5ns_5ns_5_2_1_U13.ce  = 1'h1;
assign \add_5ns_5ns_5_2_1_U13.clk  = ap_clk;
assign \add_5ns_5ns_5_2_1_U13.din0  = { 1'h0, ret_reg_1129[1], ret_reg_1129[1], ret_reg_1129 };
assign \add_5ns_5ns_5_2_1_U13.din1  = { 3'h0, op_17 };
assign grp_fu_753_p2 = \add_5ns_5ns_5_2_1_U13.dout ;
assign \add_5ns_5ns_5_2_1_U13.reset  = ap_rst;
assign \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.ain_s0  = \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.a ;
assign \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.bin_s0  = \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.b ;
assign \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.s  = { \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.fas_s2 , \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.sum_s1  };
assign \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.u2.a  = \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.ain_s1 ;
assign \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.u2.b  = \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.bin_s1 ;
assign \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.u2.cin  = \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.carry_s1 ;
assign \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.facout_s2  = \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.u2.cout ;
assign \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.fas_s2  = \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.u2.s ;
assign \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.u1.a  = \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.a [16:0];
assign \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.u1.b  = \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.b [16:0];
assign \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.u1.cin  = 1'h0;
assign \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.facout_s1  = \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.u1.cout ;
assign \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.fas_s1  = \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.u1.s ;
assign \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.a  = \add_34s_34s_34_2_1_U18.din0 ;
assign \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.b  = \add_34s_34s_34_2_1_U18.din1 ;
assign \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.ce  = \add_34s_34s_34_2_1_U18.ce ;
assign \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.clk  = \add_34s_34s_34_2_1_U18.clk ;
assign \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.reset  = \add_34s_34s_34_2_1_U18.reset ;
assign \add_34s_34s_34_2_1_U18.dout  = \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_11_U.s ;
assign \add_34s_34s_34_2_1_U18.ce  = 1'h1;
assign \add_34s_34s_34_2_1_U18.clk  = ap_clk;
assign \add_34s_34s_34_2_1_U18.din0  = { op_30_V_reg_1229[9], op_30_V_reg_1229[9], op_30_V_reg_1229[9], op_30_V_reg_1229[9], op_30_V_reg_1229[9], op_30_V_reg_1229[9], op_30_V_reg_1229[9], op_30_V_reg_1229[9], op_30_V_reg_1229[9], op_30_V_reg_1229[9], op_30_V_reg_1229[9], op_30_V_reg_1229[9], op_30_V_reg_1229[9], op_30_V_reg_1229[9], op_30_V_reg_1229[9], op_30_V_reg_1229[9], op_30_V_reg_1229[9], op_30_V_reg_1229[9], op_30_V_reg_1229[9], op_30_V_reg_1229[9], op_30_V_reg_1229[9], op_30_V_reg_1229[9], op_30_V_reg_1229[9], op_30_V_reg_1229, 1'h0 };
assign \add_34s_34s_34_2_1_U18.din1  = { op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19 };
assign grp_fu_806_p2 = \add_34s_34s_34_2_1_U18.dout ;
assign \add_34s_34s_34_2_1_U18.reset  = ap_rst;
assign \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.ain_s0  = \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.a ;
assign \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.bin_s0  = \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.b ;
assign \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.s  = { \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.fas_s2 , \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.sum_s1  };
assign \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.u2.a  = \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.ain_s1 ;
assign \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.u2.b  = \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.bin_s1 ;
assign \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.u2.cin  = \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.carry_s1 ;
assign \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.facout_s2  = \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.u2.cout ;
assign \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.fas_s2  = \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.u2.s ;
assign \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.u1.a  = \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.a [15:0];
assign \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.u1.b  = \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.b [15:0];
assign \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.u1.cin  = 1'h0;
assign \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.facout_s1  = \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.u1.cout ;
assign \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.fas_s1  = \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.u1.s ;
assign \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.a  = \add_32ns_32ns_32_2_1_U19.din0 ;
assign \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.b  = \add_32ns_32ns_32_2_1_U19.din1 ;
assign \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.ce  = \add_32ns_32ns_32_2_1_U19.ce ;
assign \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.clk  = \add_32ns_32ns_32_2_1_U19.clk ;
assign \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.reset  = \add_32ns_32ns_32_2_1_U19.reset ;
assign \add_32ns_32ns_32_2_1_U19.dout  = \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_12_U.s ;
assign \add_32ns_32ns_32_2_1_U19.ce  = 1'h1;
assign \add_32ns_32ns_32_2_1_U19.clk  = ap_clk;
assign \add_32ns_32ns_32_2_1_U19.din0  = ret_V_21_cast_reg_1254;
assign \add_32ns_32ns_32_2_1_U19.din1  = 32'd1;
assign grp_fu_822_p2 = \add_32ns_32ns_32_2_1_U19.dout ;
assign \add_32ns_32ns_32_2_1_U19.reset  = ap_rst;
assign \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.ain_s0  = \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.a ;
assign \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.bin_s0  = \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.b ;
assign \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.s  = { \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.fas_s2 , \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.sum_s1  };
assign \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.a  = \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.ain_s1 ;
assign \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.b  = \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.bin_s1 ;
assign \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.cin  = \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.carry_s1 ;
assign \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.facout_s2  = \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.cout ;
assign \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.fas_s2  = \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.s ;
assign \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.a  = \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.a [0];
assign \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.b  = \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.b [0];
assign \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.cin  = 1'h0;
assign \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.facout_s1  = \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.cout ;
assign \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.fas_s1  = \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.s ;
assign \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.a  = \add_2ns_2ns_2_2_1_U2.din0 ;
assign \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.b  = \add_2ns_2ns_2_2_1_U2.din1 ;
assign \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.ce  = \add_2ns_2ns_2_2_1_U2.ce ;
assign \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.clk  = \add_2ns_2ns_2_2_1_U2.clk ;
assign \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.reset  = \add_2ns_2ns_2_2_1_U2.reset ;
assign \add_2ns_2ns_2_2_1_U2.dout  = \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.s ;
assign \add_2ns_2ns_2_2_1_U2.ce  = 1'h1;
assign \add_2ns_2ns_2_2_1_U2.clk  = ap_clk;
assign \add_2ns_2ns_2_2_1_U2.din0  = ret_V_reg_884;
assign \add_2ns_2ns_2_2_1_U2.din1  = 2'h1;
assign grp_fu_256_p2 = \add_2ns_2ns_2_2_1_U2.dout ;
assign \add_2ns_2ns_2_2_1_U2.reset  = ap_rst;
assign \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.ain_s0  = \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.a ;
assign \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.bin_s0  = \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.b ;
assign \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.s  = { \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.fas_s2 , \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.sum_s1  };
assign \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.a  = \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.ain_s1 ;
assign \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.b  = \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.bin_s1 ;
assign \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.cin  = \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.carry_s1 ;
assign \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.facout_s2  = \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.cout ;
assign \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.fas_s2  = \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.s ;
assign \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.a  = \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.a [0];
assign \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.b  = \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.b [0];
assign \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.cin  = 1'h0;
assign \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.facout_s1  = \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.cout ;
assign \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.fas_s1  = \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.s ;
assign \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.a  = \add_2ns_2ns_2_2_1_U14.din0 ;
assign \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.b  = \add_2ns_2ns_2_2_1_U14.din1 ;
assign \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.ce  = \add_2ns_2ns_2_2_1_U14.ce ;
assign \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.clk  = \add_2ns_2ns_2_2_1_U14.clk ;
assign \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.reset  = \add_2ns_2ns_2_2_1_U14.reset ;
assign \add_2ns_2ns_2_2_1_U14.dout  = \add_2ns_2ns_2_2_1_U14.top_add_2ns_2ns_2_2_1_Adder_1_U.s ;
assign \add_2ns_2ns_2_2_1_U14.ce  = 1'h1;
assign \add_2ns_2ns_2_2_1_U14.clk  = ap_clk;
assign \add_2ns_2ns_2_2_1_U14.din0  = add_ln69_4_reg_1144;
assign \add_2ns_2ns_2_2_1_U14.din1  = select_ln69_1_reg_1139;
assign grp_fu_759_p2 = \add_2ns_2ns_2_2_1_U14.dout ;
assign \add_2ns_2ns_2_2_1_U14.reset  = ap_rst;
assign \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.ain_s0  = \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.a ;
assign \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.bin_s0  = \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.b ;
assign \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.s  = { \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.fas_s2 , \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.sum_s1  };
assign \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.a  = \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.ain_s1 ;
assign \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.b  = \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.bin_s1 ;
assign \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.cin  = \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.carry_s1 ;
assign \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.facout_s2  = \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.cout ;
assign \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.fas_s2  = \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.s ;
assign \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.a  = \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.a [0];
assign \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.b  = \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.b [0];
assign \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.cin  = 1'h0;
assign \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.facout_s1  = \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.cout ;
assign \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.fas_s1  = \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.s ;
assign \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.a  = \add_2ns_2ns_2_2_1_U10.din0 ;
assign \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.b  = \add_2ns_2ns_2_2_1_U10.din1 ;
assign \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.ce  = \add_2ns_2ns_2_2_1_U10.ce ;
assign \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.clk  = \add_2ns_2ns_2_2_1_U10.clk ;
assign \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.reset  = \add_2ns_2ns_2_2_1_U10.reset ;
assign \add_2ns_2ns_2_2_1_U10.dout  = \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_1_U.s ;
assign \add_2ns_2ns_2_2_1_U10.ce  = 1'h1;
assign \add_2ns_2ns_2_2_1_U10.clk  = ap_clk;
assign \add_2ns_2ns_2_2_1_U10.din0  = select_ln69_2_reg_1099;
assign \add_2ns_2ns_2_2_1_U10.din1  = { 1'h0, op_12 };
assign grp_fu_685_p2 = \add_2ns_2ns_2_2_1_U10.dout ;
assign \add_2ns_2ns_2_2_1_U10.reset  = ap_rst;
assign \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.ain_s0  = \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.a ;
assign \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.bin_s0  = \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.b ;
assign \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.s  = { \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.fas_s2 , \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.sum_s1  };
assign \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.u2.a  = \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.ain_s1 ;
assign \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.u2.b  = \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.bin_s1 ;
assign \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.u2.cin  = \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.carry_s1 ;
assign \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.facout_s2  = \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.u2.cout ;
assign \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.fas_s2  = \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.u2.s ;
assign \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.u1.a  = \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.a [7:0];
assign \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.u1.b  = \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.b [7:0];
assign \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.u1.cin  = 1'h0;
assign \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.facout_s1  = \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.u1.cout ;
assign \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.fas_s1  = \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.u1.s ;
assign \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.a  = \add_17s_17s_17_2_1_U6.din0 ;
assign \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.b  = \add_17s_17s_17_2_1_U6.din1 ;
assign \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.ce  = \add_17s_17s_17_2_1_U6.ce ;
assign \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.clk  = \add_17s_17s_17_2_1_U6.clk ;
assign \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.reset  = \add_17s_17s_17_2_1_U6.reset ;
assign \add_17s_17s_17_2_1_U6.dout  = \add_17s_17s_17_2_1_U6.top_add_17s_17s_17_2_1_Adder_4_U.s ;
assign \add_17s_17s_17_2_1_U6.ce  = 1'h1;
assign \add_17s_17s_17_2_1_U6.clk  = ap_clk;
assign \add_17s_17s_17_2_1_U6.din0  = { op_21_V_reg_1052[4], op_21_V_reg_1052[4], op_21_V_reg_1052, 10'h000 };
assign \add_17s_17s_17_2_1_U6.din1  = { op_10[15], op_10 };
assign grp_fu_606_p2 = \add_17s_17s_17_2_1_U6.dout ;
assign \add_17s_17s_17_2_1_U6.reset  = ap_rst;
assign \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.ain_s0  = \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.a ;
assign \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.bin_s0  = \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.b ;
assign \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.s  = { \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.fas_s2 , \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.sum_s1  };
assign \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.u2.a  = \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.ain_s1 ;
assign \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.u2.b  = \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.bin_s1 ;
assign \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.u2.cin  = \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.carry_s1 ;
assign \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.facout_s2  = \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.u2.cout ;
assign \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.fas_s2  = \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.u2.s ;
assign \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.u1.a  = \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.a [4:0];
assign \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.u1.b  = \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.b [4:0];
assign \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.u1.cin  = 1'h0;
assign \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.facout_s1  = \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.u1.cout ;
assign \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.fas_s1  = \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.u1.s ;
assign \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.a  = \add_10s_10ns_10_2_1_U17.din0 ;
assign \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.b  = \add_10s_10ns_10_2_1_U17.din1 ;
assign \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.ce  = \add_10s_10ns_10_2_1_U17.ce ;
assign \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.clk  = \add_10s_10ns_10_2_1_U17.clk ;
assign \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.reset  = \add_10s_10ns_10_2_1_U17.reset ;
assign \add_10s_10ns_10_2_1_U17.dout  = \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_8_U.s ;
assign \add_10s_10ns_10_2_1_U17.ce  = 1'h1;
assign \add_10s_10ns_10_2_1_U17.clk  = ap_clk;
assign \add_10s_10ns_10_2_1_U17.din0  = { add_ln69_6_reg_1219[5], add_ln69_6_reg_1219[5], add_ln69_6_reg_1219[5], add_ln69_6_reg_1219[5], add_ln69_6_reg_1219 };
assign \add_10s_10ns_10_2_1_U17.din1  = add_ln69_2_reg_1214;
assign grp_fu_786_p2 = \add_10s_10ns_10_2_1_U17.dout ;
assign \add_10s_10ns_10_2_1_U17.reset  = ap_rst;
assign \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.ain_s0  = \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.a ;
assign \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.bin_s0  = \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.b ;
assign \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.s  = { \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.fas_s2 , \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.sum_s1  };
assign \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.u2.a  = \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.ain_s1 ;
assign \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.u2.b  = \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.bin_s1 ;
assign \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.u2.cin  = \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.carry_s1 ;
assign \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.facout_s2  = \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.u2.cout ;
assign \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.fas_s2  = \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.u2.s ;
assign \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.u1.a  = \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.a [4:0];
assign \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.u1.b  = \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.b [4:0];
assign \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.u1.cin  = 1'h0;
assign \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.facout_s1  = \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.u1.cout ;
assign \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.fas_s1  = \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.u1.s ;
assign \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.a  = \add_10s_10ns_10_2_1_U15.din0 ;
assign \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.b  = \add_10s_10ns_10_2_1_U15.din1 ;
assign \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.ce  = \add_10s_10ns_10_2_1_U15.ce ;
assign \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.clk  = \add_10s_10ns_10_2_1_U15.clk ;
assign \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.reset  = \add_10s_10ns_10_2_1_U15.reset ;
assign \add_10s_10ns_10_2_1_U15.dout  = \add_10s_10ns_10_2_1_U15.top_add_10s_10ns_10_2_1_Adder_8_U.s ;
assign \add_10s_10ns_10_2_1_U15.ce  = 1'h1;
assign \add_10s_10ns_10_2_1_U15.clk  = ap_clk;
assign \add_10s_10ns_10_2_1_U15.din0  = { add_ln69_1_reg_1184[4], add_ln69_1_reg_1184[4], add_ln69_1_reg_1184[4], add_ln69_1_reg_1184[4], add_ln69_1_reg_1184[4], add_ln69_1_reg_1184 };
assign \add_10s_10ns_10_2_1_U15.din1  = add_ln69_reg_1179;
assign grp_fu_766_p2 = \add_10s_10ns_10_2_1_U15.dout ;
assign \add_10s_10ns_10_2_1_U15.reset  = ap_rst;
assign \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.ain_s0  = \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.a ;
assign \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.bin_s0  = \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.b ;
assign \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.s  = { \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.fas_s2 , \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.sum_s1  };
assign \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.u2.a  = \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.ain_s1 ;
assign \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.u2.b  = \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.bin_s1 ;
assign \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.u2.cin  = \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.carry_s1 ;
assign \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.facout_s2  = \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.u2.cout ;
assign \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.fas_s2  = \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.u2.s ;
assign \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.u1.a  = \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.a [4:0];
assign \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.u1.b  = \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.b [4:0];
assign \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.u1.cin  = 1'h0;
assign \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.facout_s1  = \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.u1.cout ;
assign \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.fas_s1  = \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.u1.s ;
assign \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.a  = \add_10s_10ns_10_2_1_U11.din0 ;
assign \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.b  = \add_10s_10ns_10_2_1_U11.din1 ;
assign \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.ce  = \add_10s_10ns_10_2_1_U11.ce ;
assign \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.clk  = \add_10s_10ns_10_2_1_U11.clk ;
assign \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.reset  = \add_10s_10ns_10_2_1_U11.reset ;
assign \add_10s_10ns_10_2_1_U11.dout  = \add_10s_10ns_10_2_1_U11.top_add_10s_10ns_10_2_1_Adder_8_U.s ;
assign \add_10s_10ns_10_2_1_U11.ce  = 1'h1;
assign \add_10s_10ns_10_2_1_U11.clk  = ap_clk;
assign \add_10s_10ns_10_2_1_U11.din0  = { ret_V_26_reg_1134[7], ret_V_26_reg_1134[7], ret_V_26_reg_1134 };
assign \add_10s_10ns_10_2_1_U11.din1  = { 2'h0, r_reg_995 };
assign grp_fu_741_p2 = \add_10s_10ns_10_2_1_U11.dout ;
assign \add_10s_10ns_10_2_1_U11.reset  = ap_rst;
endmodule


// Product machine:
module top_A_times_top_B (ap_start, op_0, op_10, op_11, op_12, op_16, op_17, op_18, op_19, op_2, op_3, op_6, op_7, ap_clk, unsafe_signal);
input ap_start;
input [15:0] op_0;
input [15:0] op_10;
input op_11;
input op_12;
input [3:0] op_16;
input [1:0] op_17;
input op_18;
input [3:0] op_19;
input op_2;
input [7:0] op_3;
input [1:0] op_6;
input [31:0] op_7;
input ap_clk;
output unsafe_signal;
reg _setup;
initial _setup = 1'b0;
always @ (posedge ap_clk) _setup <= 1'b1;
reg ap_start_internal;
always @ (posedge ap_clk) if (!_setup) ap_start_internal <= ap_start;
reg [15:0] op_0_internal;
always @ (posedge ap_clk) if (!_setup) op_0_internal <= op_0;
reg [15:0] op_10_internal;
always @ (posedge ap_clk) if (!_setup) op_10_internal <= op_10;
reg op_11_internal;
always @ (posedge ap_clk) if (!_setup) op_11_internal <= op_11;
reg op_12_internal;
always @ (posedge ap_clk) if (!_setup) op_12_internal <= op_12;
reg [3:0] op_16_internal;
always @ (posedge ap_clk) if (!_setup) op_16_internal <= op_16;
reg [1:0] op_17_internal;
always @ (posedge ap_clk) if (!_setup) op_17_internal <= op_17;
reg op_18_internal;
always @ (posedge ap_clk) if (!_setup) op_18_internal <= op_18;
reg [3:0] op_19_internal;
always @ (posedge ap_clk) if (!_setup) op_19_internal <= op_19;
reg op_2_internal;
always @ (posedge ap_clk) if (!_setup) op_2_internal <= op_2;
reg [7:0] op_3_internal;
always @ (posedge ap_clk) if (!_setup) op_3_internal <= op_3;
reg [1:0] op_6_internal;
always @ (posedge ap_clk) if (!_setup) op_6_internal <= op_6;
reg [31:0] op_7_internal;
always @ (posedge ap_clk) if (!_setup) op_7_internal <= op_7;
wire ap_done_A;
wire ap_done_B;
wire ap_done_eq;
assign ap_done_eq = ap_done_A == ap_done_B;
wire ap_idle_A;
wire ap_idle_B;
wire ap_idle_eq;
assign ap_idle_eq = ap_idle_A == ap_idle_B;
wire ap_ready_A;
wire ap_ready_B;
wire ap_ready_eq;
assign ap_ready_eq = ap_ready_A == ap_ready_B;
wire [31:0] op_31_A;
wire [31:0] op_31_B;
wire op_31_eq;
assign op_31_eq = op_31_A == op_31_B;
wire op_31_ap_vld_A;
wire op_31_ap_vld_B;
wire clk_enable_A;
wire clk_enable_B;
assign clk_enable_A = _setup & (~op_31_ap_vld_A | op_31_ap_vld_B);
assign clk_enable_B = _setup;
wire divergent;
assign divergent = ~(ap_done_eq & ap_idle_eq & ap_ready_eq & op_31_eq);
assign unsafe_signal = op_31_ap_vld_A & op_31_ap_vld_B & divergent;
top_A instance_A (
    .ap_clk(ap_clk),
    .clk_enable(clk_enable_A),
    .ap_start(ap_start_internal),
    .op_0(op_0_internal),
    .op_10(op_10_internal),
    .op_11(op_11_internal),
    .op_12(op_12_internal),
    .op_16(op_16_internal),
    .op_17(op_17_internal),
    .op_18(op_18_internal),
    .op_19(op_19_internal),
    .op_2(op_2_internal),
    .op_3(op_3_internal),
    .op_6(op_6_internal),
    .op_7(op_7_internal),
    .ap_done(ap_done_A),
    .ap_idle(ap_idle_A),
    .ap_ready(ap_ready_A),
    .op_31(op_31_A),
    .op_31_ap_vld(op_31_ap_vld_A)
);
top_B instance_B (
    .ap_clk(ap_clk),
    .clk_enable(clk_enable_B),
    .ap_start(ap_start_internal),
    .op_0(op_0_internal),
    .op_10(op_10_internal),
    .op_11(op_11_internal),
    .op_12(op_12_internal),
    .op_16(op_16_internal),
    .op_17(op_17_internal),
    .op_18(op_18_internal),
    .op_19(op_19_internal),
    .op_2(op_2_internal),
    .op_3(op_3_internal),
    .op_6(op_6_internal),
    .op_7(op_7_internal),
    .ap_done(ap_done_B),
    .ap_idle(ap_idle_B),
    .ap_ready(ap_ready_B),
    .op_31(op_31_B),
    .op_31_ap_vld(op_31_ap_vld_B)
);
endmodule
