// Processed by function `construct_kairos` in `verilog_tricks.py`.
// Machine A:
// Processed by function `add_clk_enable_signal` in `verilog_tricks.py`.
// Processed by function `remove_reset_signal` in `verilog_tricks.py`.
module top_A (
  ap_clk,
  ap_start,
  ap_done,
  ap_idle,
  ap_ready,
  op_0,
  op_1,
  op_3,
  op_4,
  op_7,
  op_9,
  op_11,
  op_14,
  op_15,
  op_16,
  op_17,
  op_18,
  op_19,
  op_30,
  op_30_ap_vld,
clk_enable
);
input clk_enable;


input ap_clk;
wire ap_rst;
assign ap_rst = op_30_ap_vld;
input ap_start;
input [3:0] op_0;
input [1:0] op_1;
input [15:0] op_11;
input [3:0] op_14;
input op_15;
input [7:0] op_16;
input [31:0] op_17;
input [7:0] op_18;
input op_19;
input [7:0] op_3;
input [15:0] op_4;
input [3:0] op_7;
input [7:0] op_9;
output ap_done;
output ap_idle;
output ap_ready;
output [31:0] op_30;
output op_30_ap_vld;


reg [31:0] add_ln691_1_reg_1220;
reg [31:0] add_ln691_2_reg_1242;
reg [1:0] add_ln69_3_reg_1174;
reg [10:0] ap_CS_fsm = 11'h001;
reg icmp_ln851_1_reg_1136;
reg icmp_ln851_2_reg_1098;
reg icmp_ln851_3_reg_1189;
reg icmp_ln851_4_reg_1215;
reg icmp_ln851_5_reg_1237;
reg icmp_ln851_6_reg_1259;
reg [3:0] op_12_V_reg_1179;
reg [17:0] op_22_V_reg_1184;
reg [18:0] op_26_V_reg_1199;
reg [1:0] op_2_V_reg_1103;
reg p_Result_11_reg_1151;
reg [1:0] p_Result_s_20_reg_1163;
reg [9:0] r_V_reg_1081;
reg [3:0] r_reg_1146;
reg [6:0] ret_V_18_reg_1108;
reg [31:0] ret_V_19_cast_reg_1209;
reg [8:0] ret_V_19_reg_1125;
reg [31:0] ret_V_22_cast_reg_1230;
reg [1:0] ret_V_24_reg_1169;
reg [31:0] ret_V_25_cast_reg_1252;
reg [18:0] ret_V_26_reg_1194;
reg [36:0] ret_V_27_reg_1204;
reg [56:0] ret_V_28_reg_1225;
reg [34:0] ret_V_29_reg_1247;
reg [5:0] ret_V_4_reg_1130;
reg [5:0] ret_V_5_reg_1141;
reg [6:0] ret_V_reg_1086;
reg [2:0] ret_reg_1115;
reg [7:0] sh_V_1_reg_1120;
reg tmp_5_reg_1157;
reg [2:0] trunc_ln851_reg_1093;
wire [31:0] _000_;
wire [31:0] _001_;
wire [1:0] _002_;
wire [10:0] _003_;
wire _004_;
wire _005_;
wire _006_;
wire _007_;
wire _008_;
wire _009_;
wire [3:0] _010_;
wire [17:0] _011_;
wire [18:0] _012_;
wire [1:0] _013_;
wire _014_;
wire [1:0] _015_;
wire [9:0] _016_;
wire [3:0] _017_;
wire [6:0] _018_;
wire [31:0] _019_;
wire [8:0] _020_;
wire [31:0] _021_;
wire [1:0] _022_;
wire [31:0] _023_;
wire [18:0] _024_;
wire [36:0] _025_;
wire [56:0] _026_;
wire [34:0] _027_;
wire [5:0] _028_;
wire [5:0] _029_;
wire [6:0] _030_;
wire [2:0] _031_;
wire [7:0] _032_;
wire _033_;
wire [2:0] _034_;
wire [1:0] _035_;
wire _036_;
wire _037_;
wire _038_;
wire _039_;
wire _040_;
wire _041_;
wire _042_;
wire _043_;
wire _044_;
wire _045_;
wire _046_;
wire _047_;
wire _048_;
wire _049_;
wire _050_;
wire _051_;
wire _052_;
wire _053_;
wire _054_;
wire _055_;
wire _056_;
wire _057_;
wire _058_;
wire _059_;
wire _060_;
wire _061_;
wire [31:0] add_ln691_1_fu_896_p2;
wire [31:0] add_ln691_2_fu_963_p2;
wire [31:0] add_ln691_3_fu_1036_p2;
wire [18:0] add_ln691_fu_816_p2;
wire [18:0] add_ln69_2_fu_841_p2;
wire [1:0] add_ln69_3_fu_635_p2;
wire [6:0] add_ln69_fu_752_p2;
wire and_ln353_fu_469_p2;
wire [3:0] and_ln_fu_669_p3;
wire ap_CS_fsm_state1;
wire ap_CS_fsm_state10;
wire ap_CS_fsm_state11;
wire ap_CS_fsm_state2;
wire ap_CS_fsm_state3;
wire ap_CS_fsm_state4;
wire ap_CS_fsm_state5;
wire ap_CS_fsm_state6;
wire ap_CS_fsm_state7;
wire ap_CS_fsm_state8;
wire ap_CS_fsm_state9;
wire [10:0] ap_NS_fsm;
wire ap_clk;
wire ap_done;
wire ap_idle;
wire ap_ready;
wire ap_rst;
wire ap_start;
wire [31:0] ashr_ln799_fu_498_p2;
wire icmp_ln785_fu_684_p2;
wire icmp_ln786_1_fu_707_p2;
wire icmp_ln786_fu_701_p2;
wire icmp_ln850_fu_463_p2;
wire icmp_ln851_1_fu_398_p2;
wire icmp_ln851_2_fu_293_p2;
wire icmp_ln851_3_fu_772_p2;
wire icmp_ln851_4_fu_890_p2;
wire icmp_ln851_5_fu_957_p2;
wire icmp_ln851_6_fu_1023_p2;
wire icmp_ln851_fu_315_p2;
wire [6:0] lhs_fu_362_p3;
wire [7:0] \mul_8s_2s_10_1_1_U1.din0 ;
wire [1:0] \mul_8s_2s_10_1_1_U1.din1 ;
wire [9:0] \mul_8s_2s_10_1_1_U1.dout ;
wire [7:0] \mul_8s_2s_10_1_1_U1.top_mul_8s_2s_10_1_1_Multiplier_0_U.a ;
wire [1:0] \mul_8s_2s_10_1_1_U1.top_mul_8s_2s_10_1_1_Multiplier_0_U.b ;
wire [9:0] \mul_8s_2s_10_1_1_U1.top_mul_8s_2s_10_1_1_Multiplier_0_U.p ;
wire [3:0] op_0;
wire [1:0] op_1;
wire [15:0] op_11;
wire [3:0] op_12_V_fu_737_p3;
wire [3:0] op_14;
wire op_15;
wire [7:0] op_16;
wire [31:0] op_17;
wire [7:0] op_18;
wire op_19;
wire [17:0] op_22_V_fu_762_p2;
wire [18:0] op_26_V_fu_849_p2;
wire [1:0] op_2_V_fu_303_p1;
wire [1:0] op_2_V_fu_303_p2;
wire [7:0] op_3;
wire [31:0] op_30;
wire op_30_ap_vld;
wire [15:0] op_4;
wire [3:0] op_7;
wire [7:0] op_8_V_fu_417_p2;
wire [7:0] op_9;
wire or_ln384_fu_731_p2;
wire or_ln786_fu_712_p2;
wire [3:0] or_ln_fu_676_p4;
wire overflow_fu_695_p2;
wire p_Result_10_fu_481_p3;
wire p_Result_1_fu_641_p3;
wire p_Result_2_fu_451_p3;
wire p_Result_5_fu_594_p3;
wire p_Result_6_fu_808_p3;
wire p_Result_7_fu_902_p3;
wire p_Result_8_fu_968_p3;
wire p_Result_9_fu_1029_p3;
wire p_Result_s_fu_308_p3;
wire [3:0] p_Val2_5_fu_664_p2;
wire [9:0] r_V_fu_269_p2;
wire [3:0] r_fu_529_p3;
wire [1:0] ret_V_10_fu_602_p2;
wire [1:0] ret_V_12_cast_fu_584_p4;
wire [6:0] ret_V_18_fu_332_p3;
wire [31:0] ret_V_19_cast_fu_876_p4;
wire [8:0] ret_V_19_fu_378_p2;
wire [6:0] ret_V_1_fu_320_p2;
wire [5:0] ret_V_20_fu_653_p3;
wire [10:0] ret_V_21_fu_437_p2;
wire ret_V_22_fu_475_p2;
wire [11:0] ret_V_23_fu_578_p2;
wire [1:0] ret_V_24_fu_615_p3;
wire [19:0] ret_V_25_fu_788_p2;
wire [18:0] ret_V_26_fu_829_p3;
wire [36:0] ret_V_27_fu_870_p2;
wire [56:0] ret_V_28_fu_937_p2;
wire [34:0] ret_V_29_fu_1003_p2;
wire [31:0] ret_V_30_fu_1047_p3;
wire [5:0] ret_V_4_fu_384_p4;
wire [5:0] ret_V_5_fu_404_p2;
wire [2:0] ret_fu_350_p2;
wire [9:0] rhs_2_fu_426_p3;
wire [10:0] rhs_4_fu_566_p3;
wire [19:0] rhs_6_fu_781_p3;
wire [55:0] rhs_8_fu_925_p3;
wire [33:0] rhs_9_fu_991_p3;
wire [31:0] select_ln353_1_fu_984_p3;
wire [31:0] select_ln353_fu_918_p3;
wire [3:0] select_ln384_fu_723_p3;
wire [31:0] select_ln69_1_fu_1054_p3;
wire [1:0] select_ln69_fu_627_p3;
wire [5:0] select_ln850_1_fu_648_p3;
wire [1:0] select_ln850_3_fu_608_p3;
wire [18:0] select_ln850_4_fu_822_p3;
wire [31:0] select_ln850_6_fu_913_p3;
wire [31:0] select_ln850_7_fu_1041_p3;
wire [31:0] select_ln850_8_fu_979_p3;
wire [6:0] select_ln850_fu_325_p3;
wire [19:0] sext_ln1192_1_fu_778_p1;
wire [36:0] sext_ln1192_2_fu_866_p1;
wire [56:0] sext_ln1192_3_fu_933_p1;
wire [34:0] sext_ln1192_4_fu_999_p1;
wire [11:0] sext_ln1192_fu_574_p1;
wire [10:0] sext_ln1193_1_fu_433_p1;
wire [7:0] sext_ln1193_fu_423_p0;
wire [10:0] sext_ln1193_fu_423_p1;
wire [7:0] sext_ln1349_fu_410_p1;
wire [7:0] sext_ln15_fu_339_p1;
wire [6:0] sext_ln20_fu_660_p1;
wire [2:0] sext_ln215_1_fu_346_p1;
wire [1:0] sext_ln215_fu_343_p0;
wire [2:0] sext_ln215_fu_343_p1;
wire [3:0] sext_ln546_1_fu_508_p1;
wire [15:0] sext_ln546_2_fu_512_p1;
wire [15:0] sext_ln546_fu_491_p1;
wire [17:0] sext_ln69_1_fu_758_p1;
wire [18:0] sext_ln69_2_fu_837_p1;
wire [18:0] sext_ln69_4_fu_846_p1;
wire [6:0] sext_ln69_fu_745_p1;
wire [7:0] sext_ln703_1_fu_563_p0;
wire [11:0] sext_ln703_1_fu_563_p1;
wire [7:0] sext_ln703_2_fu_855_p0;
wire [36:0] sext_ln703_2_fu_855_p1;
wire [31:0] sext_ln703_3_fu_909_p0;
wire [56:0] sext_ln703_3_fu_909_p1;
wire [7:0] sext_ln703_4_fu_975_p0;
wire [34:0] sext_ln703_4_fu_975_p1;
wire [7:0] sext_ln703_fu_374_p0;
wire [8:0] sext_ln703_fu_374_p1;
wire [31:0] sext_ln781_fu_488_p1;
wire [18:0] sext_ln850_fu_804_p1;
wire [7:0] sh_V_1_fu_356_p2;
wire [31:0] shl_ln781_fu_519_p2;
wire [17:0] tmp_1_fu_794_p4;
wire [22:0] tmp_8_fu_859_p3;
wire tmp_fu_443_p3;
wire [7:0] trunc_ln1349_fu_413_p1;
wire [2:0] trunc_ln546_fu_504_p1;
wire [1:0] trunc_ln69_fu_299_p1;
wire [3:0] trunc_ln769_fu_525_p1;
wire [7:0] trunc_ln851_1_fu_394_p0;
wire [2:0] trunc_ln851_1_fu_394_p1;
wire [2:0] trunc_ln851_2_fu_459_p1;
wire [7:0] trunc_ln851_3_fu_289_p0;
wire [2:0] trunc_ln851_3_fu_289_p1;
wire [1:0] trunc_ln851_4_fu_768_p1;
wire [7:0] trunc_ln851_5_fu_886_p0;
wire [3:0] trunc_ln851_5_fu_886_p1;
wire [31:0] trunc_ln851_6_fu_953_p0;
wire [23:0] trunc_ln851_6_fu_953_p1;
wire [7:0] trunc_ln851_7_fu_1019_p0;
wire [1:0] trunc_ln851_7_fu_1019_p1;
wire [2:0] trunc_ln851_fu_285_p1;
wire underflow_fu_718_p2;
wire xor_ln785_fu_690_p2;
wire [8:0] zext_ln1192_fu_370_p1;
wire [31:0] zext_ln546_1_fu_515_p1;
wire [31:0] zext_ln546_fu_494_p1;
wire [1:0] zext_ln69_1_fu_623_p1;
wire [17:0] zext_ln69_fu_748_p1;


assign add_ln691_1_fu_896_p2 = { ret_V_27_fu_870_p2[36], ret_V_27_fu_870_p2[36], ret_V_27_fu_870_p2[36], ret_V_27_fu_870_p2[36], ret_V_27_fu_870_p2[36], ret_V_27_fu_870_p2[36], ret_V_27_fu_870_p2[36], ret_V_27_fu_870_p2[36], ret_V_27_fu_870_p2[36], ret_V_27_fu_870_p2[36], ret_V_27_fu_870_p2[36], ret_V_27_fu_870_p2[36], ret_V_27_fu_870_p2[36], ret_V_27_fu_870_p2[22:4] } + 1'h1;
assign add_ln691_2_fu_963_p2 = ret_V_22_cast_reg_1230 + 1'h1;
assign add_ln691_3_fu_1036_p2 = ret_V_25_cast_reg_1252 + 1'h1;
assign add_ln691_fu_816_p2 = $signed(ret_V_25_fu_788_p2[19:2]) + $signed(2'h1);
assign add_ln69_2_fu_841_p2 = $signed(ret_V_26_reg_1194) + $signed(op_14);
assign add_ln69_3_fu_635_p2 = select_ln69_fu_627_p3 + ret_V_22_fu_475_p2;
assign add_ln69_fu_752_p2 = $signed(ret_V_20_fu_653_p3) + $signed(ret_V_24_reg_1169);
assign op_22_V_fu_762_p2 = $signed(add_ln69_fu_752_p2) + $signed({ 1'h0, op_11 });
assign op_26_V_fu_849_p2 = $signed(add_ln69_3_reg_1174) + $signed(add_ln69_2_fu_841_p2);
assign op_2_V_fu_303_p2 = $signed(op_0[1:0]) + $signed(op_1);
assign op_30 = ret_V_30_fu_1047_p3 + select_ln69_1_fu_1054_p3;
assign ret_V_10_fu_602_p2 = ret_V_23_fu_578_p2[4:3] + 1'h1;
assign ret_V_19_fu_378_p2 = $signed({ 1'h0, op_7, 3'h0 }) + $signed(op_9);
assign ret_V_1_fu_320_p2 = ret_V_reg_1086 + 1'h1;
assign ret_V_23_fu_578_p2 = $signed({ op_8_V_fu_417_p2, 3'h0 }) + $signed(op_3);
assign ret_V_25_fu_788_p2 = $signed({ op_22_V_reg_1184, 2'h0 }) + $signed(op_12_V_reg_1179);
assign { ret_V_27_fu_870_p2[36], ret_V_27_fu_870_p2[22:0] } = $signed({ op_26_V_reg_1199, 4'h0 }) + $signed(op_16);
assign ret_V_28_fu_937_p2 = $signed({ select_ln353_fu_918_p3, 24'h000000 }) + $signed(op_17);
assign ret_V_29_fu_1003_p2 = $signed({ select_ln353_1_fu_984_p3, 2'h0 }) + $signed(op_18);
assign ret_V_5_fu_404_p2 = ret_V_19_fu_378_p2[8:3] + 1'h1;
assign ret_fu_350_p2 = $signed(op_2_V_fu_303_p2) + $signed(op_1);
assign _036_ = ap_CS_fsm[8] & icmp_ln851_5_reg_1237;
assign _037_ = ap_CS_fsm[0] & _039_;
assign _038_ = ap_CS_fsm[0] & ap_start;
assign and_ln353_fu_469_p2 = ret_V_21_fu_437_p2[10] & icmp_ln850_fu_463_p2;
assign overflow_fu_695_p2 = xor_ln785_fu_690_p2 & icmp_ln785_fu_684_p2;
assign underflow_fu_718_p2 = p_Result_11_reg_1151 & or_ln786_fu_712_p2;
assign xor_ln785_fu_690_p2 = ~ p_Result_11_reg_1151;
assign _039_ = ~ ap_start;
assign _040_ = ! { tmp_5_reg_1157, 3'h0 };
assign _041_ = ! op_9[2:0];
assign _042_ = ! op_3[2:0];
assign _043_ = ! trunc_ln851_reg_1093;
assign \mul_8s_2s_10_1_1_U1.top_mul_8s_2s_10_1_1_Multiplier_0_U.p  = $signed(\mul_8s_2s_10_1_1_U1.top_mul_8s_2s_10_1_1_Multiplier_0_U.a ) * $signed(\mul_8s_2s_10_1_1_U1.top_mul_8s_2s_10_1_1_Multiplier_0_U.b );
assign _044_ = | { tmp_5_reg_1157, 1'h0, p_Result_s_20_reg_1163 };
assign _045_ = p_Result_s_20_reg_1163 != 2'h3;
assign _046_ = | ret_V_21_fu_437_p2[2:0];
assign _047_ = | op_12_V_fu_737_p3[1:0];
assign _048_ = | op_16[3:0];
assign _049_ = | op_17[23:0];
assign _050_ = | op_18[1:0];
assign op_8_V_fu_417_p2 = op_4[7:0] | { op_2_V_reg_1103[1], op_2_V_reg_1103[1], op_2_V_reg_1103[1], op_2_V_reg_1103[1], op_2_V_reg_1103[1], op_2_V_reg_1103[1], op_2_V_reg_1103 };
assign or_ln384_fu_731_p2 = underflow_fu_718_p2 | overflow_fu_695_p2;
assign or_ln786_fu_712_p2 = icmp_ln786_fu_701_p2 | icmp_ln786_1_fu_707_p2;
always @(posedge ap_clk)
ret_V_26_reg_1194 <= _024_;
always @(posedge ap_clk)
op_2_V_reg_1103 <= _013_;
always @(posedge ap_clk)
ret_V_18_reg_1108 <= _018_;
always @(posedge ap_clk)
ret_reg_1115 <= _031_;
always @(posedge ap_clk)
sh_V_1_reg_1120 <= _032_;
always @(posedge ap_clk)
op_26_V_reg_1199 <= _012_;
always @(posedge ap_clk)
ret_V_29_reg_1247 <= _027_;
always @(posedge ap_clk)
ret_V_25_cast_reg_1252 <= _023_;
always @(posedge ap_clk)
icmp_ln851_6_reg_1259 <= _009_;
always @(posedge ap_clk)
ret_V_28_reg_1225 <= _026_;
always @(posedge ap_clk)
ret_V_22_cast_reg_1230 <= _021_;
always @(posedge ap_clk)
icmp_ln851_5_reg_1237 <= _008_;
always @(posedge ap_clk)
op_12_V_reg_1179 <= _010_;
always @(posedge ap_clk)
op_22_V_reg_1184 <= _011_;
always @(posedge ap_clk)
icmp_ln851_3_reg_1189 <= _006_;
always @(posedge ap_clk)
r_V_reg_1081 <= _016_;
always @(posedge ap_clk)
ret_V_reg_1086 <= _030_;
always @(posedge ap_clk)
trunc_ln851_reg_1093 <= _034_;
always @(posedge ap_clk)
icmp_ln851_2_reg_1098 <= _005_;
always @(posedge ap_clk)
ret_V_19_reg_1125 <= _020_;
always @(posedge ap_clk)
ret_V_4_reg_1130 <= _028_;
always @(posedge ap_clk)
icmp_ln851_1_reg_1136 <= _004_;
always @(posedge ap_clk)
ret_V_5_reg_1141 <= _029_;
always @(posedge ap_clk)
r_reg_1146 <= _017_;
always @(posedge ap_clk)
p_Result_11_reg_1151 <= _014_;
always @(posedge ap_clk)
tmp_5_reg_1157 <= _033_;
always @(posedge ap_clk)
p_Result_s_20_reg_1163 <= _015_;
always @(posedge ap_clk)
ret_V_24_reg_1169 <= _022_;
always @(posedge ap_clk)
add_ln69_3_reg_1174 <= _002_;
always @(posedge ap_clk)
add_ln691_2_reg_1242 <= _001_;
always @(posedge ap_clk)
ret_V_27_reg_1204 <= _025_;
always @(posedge ap_clk)
ret_V_19_cast_reg_1209 <= _019_;
always @(posedge ap_clk)
icmp_ln851_4_reg_1215 <= _007_;
always @(posedge ap_clk)
add_ln691_1_reg_1220 <= _000_;
always @(posedge ap_clk)
ap_CS_fsm <= _003_;
assign _035_ = _038_ ? 2'h2 : 2'h1;
assign _051_ = ap_CS_fsm == 1'h1;
function [10:0] _143_;
input [10:0] a;
input [120:0] b;
input [10:0] s;
case (s)
11'b00000000001:
_143_ = b[10:0];
11'b00000000010:
_143_ = b[21:11];
11'b00000000100:
_143_ = b[32:22];
11'b00000001000:
_143_ = b[43:33];
11'b00000010000:
_143_ = b[54:44];
11'b00000100000:
_143_ = b[65:55];
11'b00001000000:
_143_ = b[76:66];
11'b00010000000:
_143_ = b[87:77];
11'b00100000000:
_143_ = b[98:88];
11'b01000000000:
_143_ = b[109:99];
11'b10000000000:
_143_ = b[120:110];
11'b00000000000:
_143_ = a;
default:
_143_ = 11'bx;
endcase
endfunction
assign ap_NS_fsm = _143_(11'hxxx, { 9'h000, _035_, 110'h0020080200802008020080200001 }, { _051_, _061_, _060_, _059_, _058_, _057_, _056_, _055_, _054_, _053_, _052_ });
assign _052_ = ap_CS_fsm == 11'h400;
assign _053_ = ap_CS_fsm == 10'h200;
assign _054_ = ap_CS_fsm == 9'h100;
assign _055_ = ap_CS_fsm == 8'h80;
assign _056_ = ap_CS_fsm == 7'h40;
assign _057_ = ap_CS_fsm == 6'h20;
assign _058_ = ap_CS_fsm == 5'h10;
assign _059_ = ap_CS_fsm == 4'h8;
assign _060_ = ap_CS_fsm == 3'h4;
assign _061_ = ap_CS_fsm == 2'h2;
assign op_30_ap_vld = ap_CS_fsm[10] ? 1'h1 : 1'h0;
assign ap_idle = _037_ ? 1'h1 : 1'h0;
assign _024_ = ap_CS_fsm[4] ? ret_V_26_fu_829_p3 : ret_V_26_reg_1194;
assign _032_ = ap_CS_fsm[1] ? sh_V_1_fu_356_p2 : sh_V_1_reg_1120;
assign _031_ = ap_CS_fsm[1] ? ret_fu_350_p2 : ret_reg_1115;
assign _018_ = ap_CS_fsm[1] ? ret_V_18_fu_332_p3 : ret_V_18_reg_1108;
assign _013_ = ap_CS_fsm[1] ? op_2_V_fu_303_p2 : op_2_V_reg_1103;
assign _012_ = ap_CS_fsm[5] ? op_26_V_fu_849_p2 : op_26_V_reg_1199;
assign _009_ = ap_CS_fsm[9] ? icmp_ln851_6_fu_1023_p2 : icmp_ln851_6_reg_1259;
assign _023_ = ap_CS_fsm[9] ? ret_V_29_fu_1003_p2[33:2] : ret_V_25_cast_reg_1252;
assign _027_ = ap_CS_fsm[9] ? ret_V_29_fu_1003_p2 : ret_V_29_reg_1247;
assign _008_ = ap_CS_fsm[7] ? icmp_ln851_5_fu_957_p2 : icmp_ln851_5_reg_1237;
assign _021_ = ap_CS_fsm[7] ? ret_V_28_fu_937_p2[55:24] : ret_V_22_cast_reg_1230;
assign _026_ = ap_CS_fsm[7] ? ret_V_28_fu_937_p2 : ret_V_28_reg_1225;
assign _006_ = ap_CS_fsm[3] ? icmp_ln851_3_fu_772_p2 : icmp_ln851_3_reg_1189;
assign _011_ = ap_CS_fsm[3] ? op_22_V_fu_762_p2 : op_22_V_reg_1184;
assign _010_ = ap_CS_fsm[3] ? op_12_V_fu_737_p3 : op_12_V_reg_1179;
assign _005_ = ap_CS_fsm[0] ? icmp_ln851_2_fu_293_p2 : icmp_ln851_2_reg_1098;
assign _034_ = ap_CS_fsm[0] ? r_V_fu_269_p2[2:0] : trunc_ln851_reg_1093;
assign _030_ = ap_CS_fsm[0] ? r_V_fu_269_p2[9:3] : ret_V_reg_1086;
assign _016_ = ap_CS_fsm[0] ? r_V_fu_269_p2 : r_V_reg_1081;
assign _002_ = ap_CS_fsm[2] ? add_ln69_3_fu_635_p2 : add_ln69_3_reg_1174;
assign _022_ = ap_CS_fsm[2] ? ret_V_24_fu_615_p3 : ret_V_24_reg_1169;
assign _015_ = ap_CS_fsm[2] ? r_fu_529_p3[3:2] : p_Result_s_20_reg_1163;
assign _033_ = ap_CS_fsm[2] ? r_fu_529_p3[1] : tmp_5_reg_1157;
assign _014_ = ap_CS_fsm[2] ? r_fu_529_p3[3] : p_Result_11_reg_1151;
assign _017_ = ap_CS_fsm[2] ? r_fu_529_p3 : r_reg_1146;
assign _029_ = ap_CS_fsm[2] ? ret_V_5_fu_404_p2 : ret_V_5_reg_1141;
assign _004_ = ap_CS_fsm[2] ? icmp_ln851_1_fu_398_p2 : icmp_ln851_1_reg_1136;
assign _028_ = ap_CS_fsm[2] ? ret_V_19_fu_378_p2[8:3] : ret_V_4_reg_1130;
assign _020_ = ap_CS_fsm[2] ? ret_V_19_fu_378_p2 : ret_V_19_reg_1125;
assign _001_ = _036_ ? add_ln691_2_fu_963_p2 : add_ln691_2_reg_1242;
assign _000_ = ap_CS_fsm[6] ? add_ln691_1_fu_896_p2 : add_ln691_1_reg_1220;
assign _007_ = ap_CS_fsm[6] ? icmp_ln851_4_fu_890_p2 : icmp_ln851_4_reg_1215;
assign _019_ = ap_CS_fsm[6] ? { ret_V_27_fu_870_p2[36], ret_V_27_fu_870_p2[36], ret_V_27_fu_870_p2[36], ret_V_27_fu_870_p2[36], ret_V_27_fu_870_p2[36], ret_V_27_fu_870_p2[36], ret_V_27_fu_870_p2[36], ret_V_27_fu_870_p2[36], ret_V_27_fu_870_p2[36], ret_V_27_fu_870_p2[36], ret_V_27_fu_870_p2[36], ret_V_27_fu_870_p2[36], ret_V_27_fu_870_p2[36], ret_V_27_fu_870_p2[22:4] } : ret_V_19_cast_reg_1209;
assign _025_ = ap_CS_fsm[6] ? { ret_V_27_fu_870_p2[36], ret_V_27_fu_870_p2[36], ret_V_27_fu_870_p2[36], ret_V_27_fu_870_p2[36], ret_V_27_fu_870_p2[36], ret_V_27_fu_870_p2[36], ret_V_27_fu_870_p2[36], ret_V_27_fu_870_p2[36], ret_V_27_fu_870_p2[36], ret_V_27_fu_870_p2[36], ret_V_27_fu_870_p2[36], ret_V_27_fu_870_p2[36], ret_V_27_fu_870_p2[36], ret_V_27_fu_870_p2[36], ret_V_27_fu_870_p2[22:0] } : ret_V_27_reg_1204;
assign _003_ = ap_rst ? 11'h001 : ap_NS_fsm;
assign trunc_ln769_fu_525_p1 = $signed(ret_reg_1115) << { ret_V_18_reg_1108[6], ret_V_18_reg_1108[6], ret_V_18_reg_1108[6], ret_V_18_reg_1108[6], ret_V_18_reg_1108[6], ret_V_18_reg_1108[6], ret_V_18_reg_1108[6], ret_V_18_reg_1108[6], ret_V_18_reg_1108[6], ret_V_18_reg_1108 };
assign trunc_ln546_fu_504_p1 = $signed(ret_reg_1115) >>> { sh_V_1_reg_1120[7], sh_V_1_reg_1120[7], sh_V_1_reg_1120[7], sh_V_1_reg_1120[7], sh_V_1_reg_1120[7], sh_V_1_reg_1120[7], sh_V_1_reg_1120[7], sh_V_1_reg_1120[7], sh_V_1_reg_1120 };
assign ret_V_21_fu_437_p2 = $signed(op_3) - $signed({ ret_V_18_reg_1108, 3'h0 });
assign sh_V_1_fu_356_p2 = $signed(1'h0) - $signed(ret_V_18_fu_332_p3);
assign icmp_ln785_fu_684_p2 = _044_ ? 1'h1 : 1'h0;
assign icmp_ln786_1_fu_707_p2 = _045_ ? 1'h1 : 1'h0;
assign icmp_ln786_fu_701_p2 = _040_ ? 1'h1 : 1'h0;
assign icmp_ln850_fu_463_p2 = _046_ ? 1'h1 : 1'h0;
assign icmp_ln851_1_fu_398_p2 = _041_ ? 1'h1 : 1'h0;
assign icmp_ln851_2_fu_293_p2 = _042_ ? 1'h1 : 1'h0;
assign icmp_ln851_3_fu_772_p2 = _047_ ? 1'h1 : 1'h0;
assign icmp_ln851_4_fu_890_p2 = _048_ ? 1'h1 : 1'h0;
assign icmp_ln851_5_fu_957_p2 = _049_ ? 1'h1 : 1'h0;
assign icmp_ln851_6_fu_1023_p2 = _050_ ? 1'h1 : 1'h0;
assign icmp_ln851_fu_315_p2 = _043_ ? 1'h1 : 1'h0;
assign op_12_V_fu_737_p3 = or_ln384_fu_731_p2 ? select_ln384_fu_723_p3 : { r_reg_1146[1:0], 2'h0 };
assign r_fu_529_p3 = ret_V_18_reg_1108[6] ? { trunc_ln546_fu_504_p1[2], trunc_ln546_fu_504_p1 } : trunc_ln769_fu_525_p1;
assign ret_V_18_fu_332_p3 = r_V_reg_1081[9] ? select_ln850_fu_325_p3 : ret_V_reg_1086;
assign ret_V_20_fu_653_p3 = ret_V_19_reg_1125[8] ? select_ln850_1_fu_648_p3 : ret_V_4_reg_1130;
assign ret_V_24_fu_615_p3 = ret_V_23_fu_578_p2[11] ? select_ln850_3_fu_608_p3 : ret_V_23_fu_578_p2[4:3];
assign ret_V_26_fu_829_p3 = ret_V_25_fu_788_p2[19] ? select_ln850_4_fu_822_p3 : { 2'h0, ret_V_25_fu_788_p2[18:2] };
assign ret_V_30_fu_1047_p3 = ret_V_29_reg_1247[34] ? select_ln850_7_fu_1041_p3 : ret_V_25_cast_reg_1252;
assign select_ln353_1_fu_984_p3 = ret_V_28_reg_1225[56] ? select_ln850_8_fu_979_p3 : ret_V_22_cast_reg_1230;
assign select_ln353_fu_918_p3 = ret_V_27_reg_1204[36] ? select_ln850_6_fu_913_p3 : ret_V_19_cast_reg_1209;
assign select_ln384_fu_723_p3 = overflow_fu_695_p2 ? 4'h7 : 4'h8;
assign select_ln69_1_fu_1054_p3 = op_19 ? 32'd4294967295 : 32'd0;
assign select_ln69_fu_627_p3 = op_15 ? 2'h3 : 2'h0;
assign select_ln850_1_fu_648_p3 = icmp_ln851_1_reg_1136 ? ret_V_4_reg_1130 : ret_V_5_reg_1141;
assign select_ln850_3_fu_608_p3 = icmp_ln851_2_reg_1098 ? ret_V_23_fu_578_p2[4:3] : ret_V_10_fu_602_p2;
assign select_ln850_4_fu_822_p3 = icmp_ln851_3_reg_1189 ? add_ln691_fu_816_p2 : { 2'h3, ret_V_25_fu_788_p2[18:2] };
assign select_ln850_6_fu_913_p3 = icmp_ln851_4_reg_1215 ? add_ln691_1_reg_1220 : ret_V_19_cast_reg_1209;
assign select_ln850_7_fu_1041_p3 = icmp_ln851_6_reg_1259 ? add_ln691_3_fu_1036_p2 : ret_V_25_cast_reg_1252;
assign select_ln850_8_fu_979_p3 = icmp_ln851_5_reg_1237 ? add_ln691_2_reg_1242 : ret_V_22_cast_reg_1230;
assign select_ln850_fu_325_p3 = icmp_ln851_fu_315_p2 ? ret_V_reg_1086 : ret_V_1_fu_320_p2;
assign ret_V_22_fu_475_p2 = ret_V_21_fu_437_p2[3] ^ and_ln353_fu_469_p2;
assign and_ln_fu_669_p3 = { tmp_5_reg_1157, 3'h0 };
assign ap_CS_fsm_state1 = ap_CS_fsm[0];
assign ap_CS_fsm_state10 = ap_CS_fsm[9];
assign ap_CS_fsm_state11 = ap_CS_fsm[10];
assign ap_CS_fsm_state2 = ap_CS_fsm[1];
assign ap_CS_fsm_state3 = ap_CS_fsm[2];
assign ap_CS_fsm_state4 = ap_CS_fsm[3];
assign ap_CS_fsm_state5 = ap_CS_fsm[4];
assign ap_CS_fsm_state6 = ap_CS_fsm[5];
assign ap_CS_fsm_state7 = ap_CS_fsm[6];
assign ap_CS_fsm_state8 = ap_CS_fsm[7];
assign ap_CS_fsm_state9 = ap_CS_fsm[8];
assign ap_done = op_30_ap_vld;
assign ap_ready = op_30_ap_vld;
assign ashr_ln799_fu_498_p2[2:0] = trunc_ln546_fu_504_p1;
assign lhs_fu_362_p3 = { op_7, 3'h0 };
assign op_2_V_fu_303_p1 = op_1;
assign or_ln_fu_676_p4 = { tmp_5_reg_1157, 1'h0, p_Result_s_20_reg_1163 };
assign p_Result_10_fu_481_p3 = ret_V_18_reg_1108[6];
assign p_Result_1_fu_641_p3 = ret_V_19_reg_1125[8];
assign p_Result_2_fu_451_p3 = ret_V_21_fu_437_p2[10];
assign p_Result_5_fu_594_p3 = ret_V_23_fu_578_p2[11];
assign p_Result_6_fu_808_p3 = ret_V_25_fu_788_p2[19];
assign p_Result_7_fu_902_p3 = ret_V_27_reg_1204[36];
assign p_Result_8_fu_968_p3 = ret_V_28_reg_1225[56];
assign p_Result_9_fu_1029_p3 = ret_V_29_reg_1247[34];
assign p_Result_s_fu_308_p3 = r_V_reg_1081[9];
assign p_Val2_5_fu_664_p2 = { r_reg_1146[1:0], 2'h0 };
assign ret_V_12_cast_fu_584_p4 = ret_V_23_fu_578_p2[4:3];
assign ret_V_19_cast_fu_876_p4 = { ret_V_27_fu_870_p2[36], ret_V_27_fu_870_p2[36], ret_V_27_fu_870_p2[36], ret_V_27_fu_870_p2[36], ret_V_27_fu_870_p2[36], ret_V_27_fu_870_p2[36], ret_V_27_fu_870_p2[36], ret_V_27_fu_870_p2[36], ret_V_27_fu_870_p2[36], ret_V_27_fu_870_p2[36], ret_V_27_fu_870_p2[36], ret_V_27_fu_870_p2[36], ret_V_27_fu_870_p2[36], ret_V_27_fu_870_p2[22:4] };
assign ret_V_27_fu_870_p2[35:23] = { ret_V_27_fu_870_p2[36], ret_V_27_fu_870_p2[36], ret_V_27_fu_870_p2[36], ret_V_27_fu_870_p2[36], ret_V_27_fu_870_p2[36], ret_V_27_fu_870_p2[36], ret_V_27_fu_870_p2[36], ret_V_27_fu_870_p2[36], ret_V_27_fu_870_p2[36], ret_V_27_fu_870_p2[36], ret_V_27_fu_870_p2[36], ret_V_27_fu_870_p2[36], ret_V_27_fu_870_p2[36] };
assign ret_V_4_fu_384_p4 = ret_V_19_fu_378_p2[8:3];
assign rhs_2_fu_426_p3 = { ret_V_18_reg_1108, 3'h0 };
assign rhs_4_fu_566_p3 = { op_8_V_fu_417_p2, 3'h0 };
assign rhs_6_fu_781_p3 = { op_22_V_reg_1184, 2'h0 };
assign rhs_8_fu_925_p3 = { select_ln353_fu_918_p3, 24'h000000 };
assign rhs_9_fu_991_p3 = { select_ln353_1_fu_984_p3, 2'h0 };
assign sext_ln1192_1_fu_778_p1 = { op_12_V_reg_1179[3], op_12_V_reg_1179[3], op_12_V_reg_1179[3], op_12_V_reg_1179[3], op_12_V_reg_1179[3], op_12_V_reg_1179[3], op_12_V_reg_1179[3], op_12_V_reg_1179[3], op_12_V_reg_1179[3], op_12_V_reg_1179[3], op_12_V_reg_1179[3], op_12_V_reg_1179[3], op_12_V_reg_1179[3], op_12_V_reg_1179[3], op_12_V_reg_1179[3], op_12_V_reg_1179[3], op_12_V_reg_1179 };
assign sext_ln1192_2_fu_866_p1 = { op_26_V_reg_1199[18], op_26_V_reg_1199[18], op_26_V_reg_1199[18], op_26_V_reg_1199[18], op_26_V_reg_1199[18], op_26_V_reg_1199[18], op_26_V_reg_1199[18], op_26_V_reg_1199[18], op_26_V_reg_1199[18], op_26_V_reg_1199[18], op_26_V_reg_1199[18], op_26_V_reg_1199[18], op_26_V_reg_1199[18], op_26_V_reg_1199[18], op_26_V_reg_1199, 4'h0 };
assign sext_ln1192_3_fu_933_p1 = { select_ln353_fu_918_p3[31], select_ln353_fu_918_p3, 24'h000000 };
assign sext_ln1192_4_fu_999_p1 = { select_ln353_1_fu_984_p3[31], select_ln353_1_fu_984_p3, 2'h0 };
assign sext_ln1192_fu_574_p1 = { op_8_V_fu_417_p2[7], op_8_V_fu_417_p2, 3'h0 };
assign sext_ln1193_1_fu_433_p1 = { ret_V_18_reg_1108[6], ret_V_18_reg_1108, 3'h0 };
assign sext_ln1193_fu_423_p0 = op_3;
assign sext_ln1193_fu_423_p1 = { op_3[7], op_3[7], op_3[7], op_3 };
assign sext_ln1349_fu_410_p1 = { op_2_V_reg_1103[1], op_2_V_reg_1103[1], op_2_V_reg_1103[1], op_2_V_reg_1103[1], op_2_V_reg_1103[1], op_2_V_reg_1103[1], op_2_V_reg_1103 };
assign sext_ln15_fu_339_p1 = { ret_V_18_fu_332_p3[6], ret_V_18_fu_332_p3 };
assign sext_ln20_fu_660_p1 = { ret_V_20_fu_653_p3[5], ret_V_20_fu_653_p3 };
assign sext_ln215_1_fu_346_p1 = { op_2_V_fu_303_p2[1], op_2_V_fu_303_p2 };
assign sext_ln215_fu_343_p0 = op_1;
assign sext_ln215_fu_343_p1 = { op_1[1], op_1 };
assign sext_ln546_1_fu_508_p1 = { trunc_ln546_fu_504_p1[2], trunc_ln546_fu_504_p1 };
assign sext_ln546_2_fu_512_p1 = { ret_V_18_reg_1108[6], ret_V_18_reg_1108[6], ret_V_18_reg_1108[6], ret_V_18_reg_1108[6], ret_V_18_reg_1108[6], ret_V_18_reg_1108[6], ret_V_18_reg_1108[6], ret_V_18_reg_1108[6], ret_V_18_reg_1108[6], ret_V_18_reg_1108 };
assign sext_ln546_fu_491_p1 = { sh_V_1_reg_1120[7], sh_V_1_reg_1120[7], sh_V_1_reg_1120[7], sh_V_1_reg_1120[7], sh_V_1_reg_1120[7], sh_V_1_reg_1120[7], sh_V_1_reg_1120[7], sh_V_1_reg_1120[7], sh_V_1_reg_1120 };
assign sext_ln69_1_fu_758_p1 = { add_ln69_fu_752_p2[6], add_ln69_fu_752_p2[6], add_ln69_fu_752_p2[6], add_ln69_fu_752_p2[6], add_ln69_fu_752_p2[6], add_ln69_fu_752_p2[6], add_ln69_fu_752_p2[6], add_ln69_fu_752_p2[6], add_ln69_fu_752_p2[6], add_ln69_fu_752_p2[6], add_ln69_fu_752_p2[6], add_ln69_fu_752_p2 };
assign sext_ln69_2_fu_837_p1 = { op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14 };
assign sext_ln69_4_fu_846_p1 = { add_ln69_3_reg_1174[1], add_ln69_3_reg_1174[1], add_ln69_3_reg_1174[1], add_ln69_3_reg_1174[1], add_ln69_3_reg_1174[1], add_ln69_3_reg_1174[1], add_ln69_3_reg_1174[1], add_ln69_3_reg_1174[1], add_ln69_3_reg_1174[1], add_ln69_3_reg_1174[1], add_ln69_3_reg_1174[1], add_ln69_3_reg_1174[1], add_ln69_3_reg_1174[1], add_ln69_3_reg_1174[1], add_ln69_3_reg_1174[1], add_ln69_3_reg_1174[1], add_ln69_3_reg_1174[1], add_ln69_3_reg_1174 };
assign sext_ln69_fu_745_p1 = { ret_V_24_reg_1169[1], ret_V_24_reg_1169[1], ret_V_24_reg_1169[1], ret_V_24_reg_1169[1], ret_V_24_reg_1169[1], ret_V_24_reg_1169 };
assign sext_ln703_1_fu_563_p0 = op_3;
assign sext_ln703_1_fu_563_p1 = { op_3[7], op_3[7], op_3[7], op_3[7], op_3 };
assign sext_ln703_2_fu_855_p0 = op_16;
assign sext_ln703_2_fu_855_p1 = { op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16 };
assign sext_ln703_3_fu_909_p0 = op_17;
assign sext_ln703_3_fu_909_p1 = { op_17[31], op_17[31], op_17[31], op_17[31], op_17[31], op_17[31], op_17[31], op_17[31], op_17[31], op_17[31], op_17[31], op_17[31], op_17[31], op_17[31], op_17[31], op_17[31], op_17[31], op_17[31], op_17[31], op_17[31], op_17[31], op_17[31], op_17[31], op_17[31], op_17[31], op_17 };
assign sext_ln703_4_fu_975_p0 = op_18;
assign sext_ln703_4_fu_975_p1 = { op_18[7], op_18[7], op_18[7], op_18[7], op_18[7], op_18[7], op_18[7], op_18[7], op_18[7], op_18[7], op_18[7], op_18[7], op_18[7], op_18[7], op_18[7], op_18[7], op_18[7], op_18[7], op_18[7], op_18[7], op_18[7], op_18[7], op_18[7], op_18[7], op_18[7], op_18[7], op_18[7], op_18 };
assign sext_ln703_fu_374_p0 = op_9;
assign sext_ln703_fu_374_p1 = { op_9[7], op_9 };
assign sext_ln781_fu_488_p1 = { ret_reg_1115[2], ret_reg_1115[2], ret_reg_1115[2], ret_reg_1115[2], ret_reg_1115[2], ret_reg_1115[2], ret_reg_1115[2], ret_reg_1115[2], ret_reg_1115[2], ret_reg_1115[2], ret_reg_1115[2], ret_reg_1115[2], ret_reg_1115[2], ret_reg_1115[2], ret_reg_1115[2], ret_reg_1115[2], ret_reg_1115[2], ret_reg_1115[2], ret_reg_1115[2], ret_reg_1115[2], ret_reg_1115[2], ret_reg_1115[2], ret_reg_1115[2], ret_reg_1115[2], ret_reg_1115[2], ret_reg_1115[2], ret_reg_1115[2], ret_reg_1115[2], ret_reg_1115[2], ret_reg_1115 };
assign sext_ln850_fu_804_p1 = { ret_V_25_fu_788_p2[19], ret_V_25_fu_788_p2[19:2] };
assign shl_ln781_fu_519_p2[3:0] = trunc_ln769_fu_525_p1;
assign tmp_1_fu_794_p4 = ret_V_25_fu_788_p2[19:2];
assign tmp_8_fu_859_p3 = { op_26_V_reg_1199, 4'h0 };
assign tmp_fu_443_p3 = ret_V_21_fu_437_p2[3];
assign trunc_ln1349_fu_413_p1 = op_4[7:0];
assign trunc_ln69_fu_299_p1 = op_0[1:0];
assign trunc_ln851_1_fu_394_p0 = op_9;
assign trunc_ln851_1_fu_394_p1 = op_9[2:0];
assign trunc_ln851_2_fu_459_p1 = ret_V_21_fu_437_p2[2:0];
assign trunc_ln851_3_fu_289_p0 = op_3;
assign trunc_ln851_3_fu_289_p1 = op_3[2:0];
assign trunc_ln851_4_fu_768_p1 = op_12_V_fu_737_p3[1:0];
assign trunc_ln851_5_fu_886_p0 = op_16;
assign trunc_ln851_5_fu_886_p1 = op_16[3:0];
assign trunc_ln851_6_fu_953_p0 = op_17;
assign trunc_ln851_6_fu_953_p1 = op_17[23:0];
assign trunc_ln851_7_fu_1019_p0 = op_18;
assign trunc_ln851_7_fu_1019_p1 = op_18[1:0];
assign trunc_ln851_fu_285_p1 = r_V_fu_269_p2[2:0];
assign zext_ln1192_fu_370_p1 = { 2'h0, op_7, 3'h0 };
assign zext_ln546_1_fu_515_p1 = { 16'h0000, ret_V_18_reg_1108[6], ret_V_18_reg_1108[6], ret_V_18_reg_1108[6], ret_V_18_reg_1108[6], ret_V_18_reg_1108[6], ret_V_18_reg_1108[6], ret_V_18_reg_1108[6], ret_V_18_reg_1108[6], ret_V_18_reg_1108[6], ret_V_18_reg_1108 };
assign zext_ln546_fu_494_p1 = { 16'h0000, sh_V_1_reg_1120[7], sh_V_1_reg_1120[7], sh_V_1_reg_1120[7], sh_V_1_reg_1120[7], sh_V_1_reg_1120[7], sh_V_1_reg_1120[7], sh_V_1_reg_1120[7], sh_V_1_reg_1120[7], sh_V_1_reg_1120 };
assign zext_ln69_1_fu_623_p1 = { 1'h0, ret_V_22_fu_475_p2 };
assign zext_ln69_fu_748_p1 = { 2'h0, op_11 };
assign \mul_8s_2s_10_1_1_U1.top_mul_8s_2s_10_1_1_Multiplier_0_U.a  = \mul_8s_2s_10_1_1_U1.din0 ;
assign \mul_8s_2s_10_1_1_U1.top_mul_8s_2s_10_1_1_Multiplier_0_U.b  = \mul_8s_2s_10_1_1_U1.din1 ;
assign \mul_8s_2s_10_1_1_U1.dout  = \mul_8s_2s_10_1_1_U1.top_mul_8s_2s_10_1_1_Multiplier_0_U.p ;
assign \mul_8s_2s_10_1_1_U1.din0  = op_3;
assign \mul_8s_2s_10_1_1_U1.din1  = op_1;
assign r_V_fu_269_p2 = \mul_8s_2s_10_1_1_U1.dout ;
endmodule


// Machine B:
// Processed by function `add_clk_enable_signal` in `verilog_tricks.py`.
// Processed by function `remove_reset_signal` in `verilog_tricks.py`.
module top_B (
  ap_clk,
  ap_start,
  ap_done,
  ap_idle,
  ap_ready,
  op_0,
  op_1,
  op_3,
  op_4,
  op_7,
  op_9,
  op_11,
  op_14,
  op_15,
  op_16,
  op_17,
  op_18,
  op_19,
  op_30,
  op_30_ap_vld,
clk_enable
);
input clk_enable;


input ap_clk;
wire ap_rst;
assign ap_rst = op_30_ap_vld;
input ap_start;
input [3:0] op_0;
input [1:0] op_1;
input [15:0] op_11;
input [3:0] op_14;
input op_15;
input [7:0] op_16;
input [31:0] op_17;
input [7:0] op_18;
input op_19;
input [7:0] op_3;
input [15:0] op_4;
input [3:0] op_7;
input [7:0] op_9;
output ap_done;
output ap_idle;
output ap_ready;
output [31:0] op_30;
output op_30_ap_vld;


reg [5:0] \add_12s_12s_12_2_1_U7.top_add_12s_12s_12_2_1_Adder_5_U.ain_s1 ;
reg [5:0] \add_12s_12s_12_2_1_U7.top_add_12s_12s_12_2_1_Adder_5_U.bin_s1 ;
reg \add_12s_12s_12_2_1_U7.top_add_12s_12s_12_2_1_Adder_5_U.carry_s1 ;
reg [5:0] \add_12s_12s_12_2_1_U7.top_add_12s_12s_12_2_1_Adder_5_U.sum_s1 ;
reg [8:0] \add_18s_18ns_18_2_1_U14.top_add_18s_18ns_18_2_1_Adder_10_U.ain_s1 ;
reg [8:0] \add_18s_18ns_18_2_1_U14.top_add_18s_18ns_18_2_1_Adder_10_U.bin_s1 ;
reg \add_18s_18ns_18_2_1_U14.top_add_18s_18ns_18_2_1_Adder_10_U.carry_s1 ;
reg [8:0] \add_18s_18ns_18_2_1_U14.top_add_18s_18ns_18_2_1_Adder_10_U.sum_s1 ;
reg [9:0] \add_19ns_19s_19_2_1_U17.top_add_19ns_19s_19_2_1_Adder_13_U.ain_s1 ;
reg [9:0] \add_19ns_19s_19_2_1_U17.top_add_19ns_19s_19_2_1_Adder_13_U.bin_s1 ;
reg \add_19ns_19s_19_2_1_U17.top_add_19ns_19s_19_2_1_Adder_13_U.carry_s1 ;
reg [8:0] \add_19ns_19s_19_2_1_U17.top_add_19ns_19s_19_2_1_Adder_13_U.sum_s1 ;
reg [9:0] \add_19s_19ns_19_2_1_U16.top_add_19s_19ns_19_2_1_Adder_12_U.ain_s1 ;
reg [9:0] \add_19s_19ns_19_2_1_U16.top_add_19s_19ns_19_2_1_Adder_12_U.bin_s1 ;
reg \add_19s_19ns_19_2_1_U16.top_add_19s_19ns_19_2_1_Adder_12_U.carry_s1 ;
reg [8:0] \add_19s_19ns_19_2_1_U16.top_add_19s_19ns_19_2_1_Adder_12_U.sum_s1 ;
reg [9:0] \add_19s_19ns_19_2_1_U19.top_add_19s_19ns_19_2_1_Adder_12_U.ain_s1 ;
reg [9:0] \add_19s_19ns_19_2_1_U19.top_add_19s_19ns_19_2_1_Adder_12_U.bin_s1 ;
reg \add_19s_19ns_19_2_1_U19.top_add_19s_19ns_19_2_1_Adder_12_U.carry_s1 ;
reg [8:0] \add_19s_19ns_19_2_1_U19.top_add_19s_19ns_19_2_1_Adder_12_U.sum_s1 ;
reg [9:0] \add_20ns_20s_20_2_1_U15.top_add_20ns_20s_20_2_1_Adder_11_U.ain_s1 ;
reg [9:0] \add_20ns_20s_20_2_1_U15.top_add_20ns_20s_20_2_1_Adder_11_U.bin_s1 ;
reg \add_20ns_20s_20_2_1_U15.top_add_20ns_20s_20_2_1_Adder_11_U.carry_s1 ;
reg [9:0] \add_20ns_20s_20_2_1_U15.top_add_20ns_20s_20_2_1_Adder_11_U.sum_s1 ;
reg \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_6_U.ain_s1 ;
reg \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_6_U.bin_s1 ;
reg \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_6_U.carry_s1 ;
reg \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_6_U.sum_s1 ;
reg \add_2ns_2ns_2_2_1_U18.top_add_2ns_2ns_2_2_1_Adder_6_U.ain_s1 ;
reg \add_2ns_2ns_2_2_1_U18.top_add_2ns_2ns_2_2_1_Adder_6_U.bin_s1 ;
reg \add_2ns_2ns_2_2_1_U18.top_add_2ns_2ns_2_2_1_Adder_6_U.carry_s1 ;
reg \add_2ns_2ns_2_2_1_U18.top_add_2ns_2ns_2_2_1_Adder_6_U.sum_s1 ;
reg \add_2ns_2s_2_2_1_U2.top_add_2ns_2s_2_2_1_Adder_0_U.ain_s1 ;
reg \add_2ns_2s_2_2_1_U2.top_add_2ns_2s_2_2_1_Adder_0_U.bin_s1 ;
reg \add_2ns_2s_2_2_1_U2.top_add_2ns_2s_2_2_1_Adder_0_U.carry_s1 ;
reg \add_2ns_2s_2_2_1_U2.top_add_2ns_2s_2_2_1_Adder_0_U.sum_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.ain_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.bin_s1 ;
reg \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.carry_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.sum_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.ain_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.bin_s1 ;
reg \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.carry_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.sum_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.ain_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.bin_s1 ;
reg \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.carry_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.sum_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U26.top_add_32ns_32ns_32_2_1_Adder_15_U.ain_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U26.top_add_32ns_32ns_32_2_1_Adder_15_U.bin_s1 ;
reg \add_32ns_32ns_32_2_1_U26.top_add_32ns_32ns_32_2_1_Adder_15_U.carry_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U26.top_add_32ns_32ns_32_2_1_Adder_15_U.sum_s1 ;
reg [17:0] \add_35s_35s_35_2_1_U24.top_add_35s_35s_35_2_1_Adder_17_U.ain_s1 ;
reg [17:0] \add_35s_35s_35_2_1_U24.top_add_35s_35s_35_2_1_Adder_17_U.bin_s1 ;
reg \add_35s_35s_35_2_1_U24.top_add_35s_35s_35_2_1_Adder_17_U.carry_s1 ;
reg [16:0] \add_35s_35s_35_2_1_U24.top_add_35s_35s_35_2_1_Adder_17_U.sum_s1 ;
reg [18:0] \add_37s_37s_37_2_1_U20.top_add_37s_37s_37_2_1_Adder_14_U.ain_s1 ;
reg [18:0] \add_37s_37s_37_2_1_U20.top_add_37s_37s_37_2_1_Adder_14_U.bin_s1 ;
reg \add_37s_37s_37_2_1_U20.top_add_37s_37s_37_2_1_Adder_14_U.carry_s1 ;
reg [17:0] \add_37s_37s_37_2_1_U20.top_add_37s_37s_37_2_1_Adder_14_U.sum_s1 ;
reg [1:0] \add_3s_3s_3_2_1_U4.top_add_3s_3s_3_2_1_Adder_2_U.ain_s1 ;
reg [1:0] \add_3s_3s_3_2_1_U4.top_add_3s_3s_3_2_1_Adder_2_U.bin_s1 ;
reg \add_3s_3s_3_2_1_U4.top_add_3s_3s_3_2_1_Adder_2_U.carry_s1 ;
reg \add_3s_3s_3_2_1_U4.top_add_3s_3s_3_2_1_Adder_2_U.sum_s1 ;
reg [28:0] \add_57s_57s_57_2_1_U22.top_add_57s_57s_57_2_1_Adder_16_U.ain_s1 ;
reg [28:0] \add_57s_57s_57_2_1_U22.top_add_57s_57s_57_2_1_Adder_16_U.bin_s1 ;
reg \add_57s_57s_57_2_1_U22.top_add_57s_57s_57_2_1_Adder_16_U.carry_s1 ;
reg [27:0] \add_57s_57s_57_2_1_U22.top_add_57s_57s_57_2_1_Adder_16_U.sum_s1 ;
reg [2:0] \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_8_U.ain_s1 ;
reg [2:0] \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_8_U.bin_s1 ;
reg \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_8_U.carry_s1 ;
reg [2:0] \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_8_U.sum_s1 ;
reg [3:0] \add_7ns_7ns_7_2_1_U3.top_add_7ns_7ns_7_2_1_Adder_1_U.ain_s1 ;
reg [3:0] \add_7ns_7ns_7_2_1_U3.top_add_7ns_7ns_7_2_1_Adder_1_U.bin_s1 ;
reg \add_7ns_7ns_7_2_1_U3.top_add_7ns_7ns_7_2_1_Adder_1_U.carry_s1 ;
reg [2:0] \add_7ns_7ns_7_2_1_U3.top_add_7ns_7ns_7_2_1_Adder_1_U.sum_s1 ;
reg [3:0] \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_9_U.ain_s1 ;
reg [3:0] \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_9_U.bin_s1 ;
reg \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_9_U.carry_s1 ;
reg [2:0] \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_9_U.sum_s1 ;
reg [4:0] \add_9ns_9s_9_2_1_U11.top_add_9ns_9s_9_2_1_Adder_7_U.ain_s1 ;
reg [4:0] \add_9ns_9s_9_2_1_U11.top_add_9ns_9s_9_2_1_Adder_7_U.bin_s1 ;
reg \add_9ns_9s_9_2_1_U11.top_add_9ns_9s_9_2_1_Adder_7_U.carry_s1 ;
reg [3:0] \add_9ns_9s_9_2_1_U11.top_add_9ns_9s_9_2_1_Adder_7_U.sum_s1 ;
reg [31:0] add_ln691_1_reg_1451;
reg [31:0] add_ln691_2_reg_1488;
reg [31:0] add_ln691_3_reg_1525;
reg [18:0] add_ln691_reg_1379;
reg [18:0] add_ln69_2_reg_1404;
reg [1:0] add_ln69_3_reg_1409;
reg [6:0] add_ln69_reg_1306;
reg [48:0] ap_CS_fsm = 49'h0000000000001;
reg [15:0] \ashr_32s_16ns_32_7_1_U8.din1_cast_array[0] ;
reg [15:0] \ashr_32s_16ns_32_7_1_U8.din1_cast_array[1] ;
reg [15:0] \ashr_32s_16ns_32_7_1_U8.din1_cast_array[2] ;
reg [15:0] \ashr_32s_16ns_32_7_1_U8.din1_cast_array[3] ;
reg [15:0] \ashr_32s_16ns_32_7_1_U8.din1_cast_array[4] ;
reg [15:0] \ashr_32s_16ns_32_7_1_U8.din1_cast_array[5] ;
reg [31:0] \ashr_32s_16ns_32_7_1_U8.dout_array[0] ;
reg [31:0] \ashr_32s_16ns_32_7_1_U8.dout_array[1] ;
reg [31:0] \ashr_32s_16ns_32_7_1_U8.dout_array[2] ;
reg [31:0] \ashr_32s_16ns_32_7_1_U8.dout_array[3] ;
reg [31:0] \ashr_32s_16ns_32_7_1_U8.dout_array[4] ;
reg [31:0] \ashr_32s_16ns_32_7_1_U8.dout_array[5] ;
reg icmp_ln785_reg_1296;
reg icmp_ln786_1_reg_1301;
reg icmp_ln786_reg_1317;
reg icmp_ln850_reg_1180;
reg icmp_ln851_1_reg_1221;
reg icmp_ln851_2_reg_1052;
reg icmp_ln851_3_reg_1357;
reg icmp_ln851_4_reg_1434;
reg icmp_ln851_5_reg_1471;
reg icmp_ln851_6_reg_1508;
reg icmp_ln851_reg_1079;
reg [7:0] \mul_8s_2s_10_7_1_U1.top_mul_8s_2s_10_7_1_Mul_DSP_0_U.a_reg0 ;
reg [1:0] \mul_8s_2s_10_7_1_U1.top_mul_8s_2s_10_7_1_Mul_DSP_0_U.b_reg0 ;
reg [9:0] \mul_8s_2s_10_7_1_U1.top_mul_8s_2s_10_7_1_Mul_DSP_0_U.buff0 ;
reg [9:0] \mul_8s_2s_10_7_1_U1.top_mul_8s_2s_10_7_1_Mul_DSP_0_U.buff1 ;
reg [9:0] \mul_8s_2s_10_7_1_U1.top_mul_8s_2s_10_7_1_Mul_DSP_0_U.buff2 ;
reg [9:0] \mul_8s_2s_10_7_1_U1.top_mul_8s_2s_10_7_1_Mul_DSP_0_U.buff3 ;
reg [9:0] \mul_8s_2s_10_7_1_U1.top_mul_8s_2s_10_7_1_Mul_DSP_0_U.buff4 ;
reg [3:0] op_12_V_reg_1332;
reg [17:0] op_22_V_reg_1337;
reg [18:0] op_26_V_reg_1419;
reg [1:0] op_2_V_reg_1084;
reg [7:0] op_8_V_reg_1112;
reg overflow_reg_1311;
reg p_Result_10_reg_1117;
reg p_Result_11_reg_1273;
reg [1:0] p_Result_s_20_reg_1285;
reg [9:0] r_V_reg_1057;
reg [3:0] r_reg_1268;
reg [1:0] ret_V_10_reg_1206;
reg [1:0] ret_V_12_cast_reg_1173;
reg [6:0] ret_V_18_reg_1095;
reg [31:0] ret_V_19_cast_reg_1444;
reg [8:0] ret_V_19_reg_1231;
reg [6:0] ret_V_1_reg_1090;
reg [5:0] ret_V_20_reg_1248;
reg [10:0] ret_V_21_reg_1152;
reg [31:0] ret_V_22_cast_reg_1481;
reg ret_V_22_reg_1201;
reg [11:0] ret_V_23_reg_1168;
reg [1:0] ret_V_24_reg_1226;
reg [31:0] ret_V_25_cast_reg_1518;
reg [19:0] ret_V_25_reg_1362;
reg [18:0] ret_V_26_reg_1384;
reg [36:0] ret_V_27_reg_1439;
reg [56:0] ret_V_28_reg_1476;
reg [34:0] ret_V_29_reg_1513;
reg [31:0] ret_V_30_reg_1530;
reg [5:0] ret_V_4_reg_1236;
reg [5:0] ret_V_5_reg_1243;
reg [6:0] ret_V_reg_1062;
reg [2:0] ret_reg_1127;
reg [31:0] select_ln353_1_reg_1493;
reg [31:0] select_ln353_reg_1456;
reg [31:0] select_ln69_1_reg_1535;
reg [1:0] select_ln69_reg_1389;
reg [18:0] sext_ln850_reg_1372;
reg [7:0] sh_V_1_reg_1163;
reg [15:0] \shl_32s_16ns_32_7_1_U9.din1_cast_array[0] ;
reg [15:0] \shl_32s_16ns_32_7_1_U9.din1_cast_array[1] ;
reg [15:0] \shl_32s_16ns_32_7_1_U9.din1_cast_array[2] ;
reg [15:0] \shl_32s_16ns_32_7_1_U9.din1_cast_array[3] ;
reg [15:0] \shl_32s_16ns_32_7_1_U9.din1_cast_array[4] ;
reg [15:0] \shl_32s_16ns_32_7_1_U9.din1_cast_array[5] ;
reg [31:0] \shl_32s_16ns_32_7_1_U9.dout_array[0] ;
reg [31:0] \shl_32s_16ns_32_7_1_U9.dout_array[1] ;
reg [31:0] \shl_32s_16ns_32_7_1_U9.dout_array[2] ;
reg [31:0] \shl_32s_16ns_32_7_1_U9.dout_array[3] ;
reg [31:0] \shl_32s_16ns_32_7_1_U9.dout_array[4] ;
reg [31:0] \shl_32s_16ns_32_7_1_U9.dout_array[5] ;
reg [5:0] \sub_11s_11s_11_2_1_U5.top_sub_11s_11s_11_2_1_Adder_3_U.ain_s1 ;
reg [5:0] \sub_11s_11s_11_2_1_U5.top_sub_11s_11s_11_2_1_Adder_3_U.bin_s1 ;
reg \sub_11s_11s_11_2_1_U5.top_sub_11s_11s_11_2_1_Adder_3_U.carry_s1 ;
reg [4:0] \sub_11s_11s_11_2_1_U5.top_sub_11s_11s_11_2_1_Adder_3_U.sum_s1 ;
reg [3:0] \sub_8ns_8s_8_2_1_U6.top_sub_8ns_8s_8_2_1_Adder_4_U.ain_s1 ;
reg [3:0] \sub_8ns_8s_8_2_1_U6.top_sub_8ns_8s_8_2_1_Adder_4_U.bin_s1 ;
reg \sub_8ns_8s_8_2_1_U6.top_sub_8ns_8s_8_2_1_Adder_4_U.carry_s1 ;
reg [3:0] \sub_8ns_8s_8_2_1_U6.top_sub_8ns_8s_8_2_1_Adder_4_U.sum_s1 ;
reg [17:0] tmp_1_reg_1367;
reg tmp_5_reg_1279;
reg [2:0] trunc_ln546_reg_1253;
reg [3:0] trunc_ln769_reg_1258;
reg [2:0] trunc_ln851_2_reg_1158;
reg [1:0] trunc_ln851_4_reg_1342;
reg [2:0] trunc_ln851_reg_1069;
wire [31:0] _000_;
wire [31:0] _001_;
wire [31:0] _002_;
wire [18:0] _003_;
wire [18:0] _004_;
wire [1:0] _005_;
wire [6:0] _006_;
wire [48:0] _007_;
wire _008_;
wire _009_;
wire _010_;
wire _011_;
wire _012_;
wire _013_;
wire _014_;
wire _015_;
wire _016_;
wire _017_;
wire _018_;
wire [3:0] _019_;
wire [17:0] _020_;
wire [18:0] _021_;
wire [1:0] _022_;
wire [7:0] _023_;
wire _024_;
wire _025_;
wire _026_;
wire [1:0] _027_;
wire [9:0] _028_;
wire [3:0] _029_;
wire [1:0] _030_;
wire [1:0] _031_;
wire [6:0] _032_;
wire [31:0] _033_;
wire [8:0] _034_;
wire [6:0] _035_;
wire [5:0] _036_;
wire [10:0] _037_;
wire [31:0] _038_;
wire _039_;
wire [11:0] _040_;
wire [1:0] _041_;
wire [31:0] _042_;
wire [19:0] _043_;
wire [18:0] _044_;
wire [36:0] _045_;
wire [56:0] _046_;
wire [34:0] _047_;
wire [31:0] _048_;
wire [5:0] _049_;
wire [5:0] _050_;
wire [6:0] _051_;
wire [2:0] _052_;
wire [31:0] _053_;
wire [31:0] _054_;
wire [31:0] _055_;
wire [1:0] _056_;
wire [18:0] _057_;
wire [7:0] _058_;
wire [17:0] _059_;
wire _060_;
wire [2:0] _061_;
wire [3:0] _062_;
wire [2:0] _063_;
wire [1:0] _064_;
wire [2:0] _065_;
wire [1:0] _066_;
wire _067_;
wire _068_;
wire _069_;
wire _070_;
wire _071_;
wire _072_;
wire _073_;
wire _074_;
wire _075_;
wire _076_;
wire _077_;
wire _078_;
wire _079_;
wire _080_;
wire _081_;
wire _082_;
wire _083_;
wire _084_;
wire _085_;
wire [5:0] _086_;
wire [5:0] _087_;
wire _088_;
wire [5:0] _089_;
wire [6:0] _090_;
wire [6:0] _091_;
wire [8:0] _092_;
wire [8:0] _093_;
wire _094_;
wire [8:0] _095_;
wire [9:0] _096_;
wire [9:0] _097_;
wire [9:0] _098_;
wire [9:0] _099_;
wire _100_;
wire [8:0] _101_;
wire [9:0] _102_;
wire [10:0] _103_;
wire [9:0] _104_;
wire [9:0] _105_;
wire _106_;
wire [8:0] _107_;
wire [9:0] _108_;
wire [10:0] _109_;
wire [9:0] _110_;
wire [9:0] _111_;
wire _112_;
wire [8:0] _113_;
wire [9:0] _114_;
wire [10:0] _115_;
wire [9:0] _116_;
wire [9:0] _117_;
wire _118_;
wire [9:0] _119_;
wire [10:0] _120_;
wire [10:0] _121_;
wire _122_;
wire _123_;
wire _124_;
wire _125_;
wire [1:0] _126_;
wire [1:0] _127_;
wire _128_;
wire _129_;
wire _130_;
wire _131_;
wire [1:0] _132_;
wire [1:0] _133_;
wire _134_;
wire _135_;
wire _136_;
wire _137_;
wire [1:0] _138_;
wire [1:0] _139_;
wire [15:0] _140_;
wire [15:0] _141_;
wire _142_;
wire [15:0] _143_;
wire [16:0] _144_;
wire [16:0] _145_;
wire [15:0] _146_;
wire [15:0] _147_;
wire _148_;
wire [15:0] _149_;
wire [16:0] _150_;
wire [16:0] _151_;
wire [15:0] _152_;
wire [15:0] _153_;
wire _154_;
wire [15:0] _155_;
wire [16:0] _156_;
wire [16:0] _157_;
wire [15:0] _158_;
wire [15:0] _159_;
wire _160_;
wire [15:0] _161_;
wire [16:0] _162_;
wire [16:0] _163_;
wire [17:0] _164_;
wire [17:0] _165_;
wire _166_;
wire [16:0] _167_;
wire [17:0] _168_;
wire [18:0] _169_;
wire [18:0] _170_;
wire [18:0] _171_;
wire _172_;
wire [17:0] _173_;
wire [18:0] _174_;
wire [19:0] _175_;
wire [1:0] _176_;
wire [1:0] _177_;
wire _178_;
wire _179_;
wire [1:0] _180_;
wire [2:0] _181_;
wire [28:0] _182_;
wire [28:0] _183_;
wire _184_;
wire [27:0] _185_;
wire [28:0] _186_;
wire [29:0] _187_;
wire [2:0] _188_;
wire [2:0] _189_;
wire _190_;
wire [2:0] _191_;
wire [3:0] _192_;
wire [3:0] _193_;
wire [3:0] _194_;
wire [3:0] _195_;
wire _196_;
wire [2:0] _197_;
wire [3:0] _198_;
wire [4:0] _199_;
wire [3:0] _200_;
wire [3:0] _201_;
wire _202_;
wire [2:0] _203_;
wire [3:0] _204_;
wire [4:0] _205_;
wire [4:0] _206_;
wire [4:0] _207_;
wire _208_;
wire [3:0] _209_;
wire [4:0] _210_;
wire [5:0] _211_;
wire [15:0] _212_;
wire [15:0] _213_;
wire [15:0] _214_;
wire [15:0] _215_;
wire [15:0] _216_;
wire [15:0] _217_;
wire [31:0] _218_;
wire [31:0] _219_;
wire [31:0] _220_;
wire [31:0] _221_;
wire [31:0] _222_;
wire [31:0] _223_;
wire [15:0] _224_;
wire [31:0] _225_;
wire [15:0] _226_;
wire [31:0] _227_;
wire [15:0] _228_;
wire [31:0] _229_;
wire [15:0] _230_;
wire [31:0] _231_;
wire [15:0] _232_;
wire [31:0] _233_;
wire [15:0] _234_;
wire [31:0] _235_;
wire [31:0] _236_;
wire [31:0] _237_;
wire [31:0] _238_;
wire [31:0] _239_;
wire [31:0] _240_;
wire [7:0] _241_;
wire [1:0] _242_;
wire [9:0] _243_;
wire [9:0] _244_;
wire [9:0] _245_;
wire [9:0] _246_;
wire [9:0] _247_;
wire [15:0] _248_;
wire [15:0] _249_;
wire [15:0] _250_;
wire [15:0] _251_;
wire [15:0] _252_;
wire [15:0] _253_;
wire [31:0] _254_;
wire [31:0] _255_;
wire [31:0] _256_;
wire [31:0] _257_;
wire [31:0] _258_;
wire [31:0] _259_;
wire [15:0] _260_;
wire [31:0] _261_;
wire [15:0] _262_;
wire [31:0] _263_;
wire [15:0] _264_;
wire [31:0] _265_;
wire [15:0] _266_;
wire [31:0] _267_;
wire [15:0] _268_;
wire [31:0] _269_;
wire [15:0] _270_;
wire [31:0] _271_;
wire [31:0] _272_;
wire [31:0] _273_;
wire [31:0] _274_;
wire [31:0] _275_;
wire [31:0] _276_;
wire [5:0] _277_;
wire [5:0] _278_;
wire _279_;
wire [4:0] _280_;
wire [5:0] _281_;
wire [6:0] _282_;
wire [3:0] _283_;
wire [3:0] _284_;
wire _285_;
wire [3:0] _286_;
wire [4:0] _287_;
wire [4:0] _288_;
wire _289_;
wire _290_;
wire _291_;
wire _292_;
wire _293_;
wire _294_;
wire _295_;
wire _296_;
wire _297_;
wire _298_;
wire _299_;
wire _300_;
wire _301_;
wire _302_;
wire _303_;
wire _304_;
wire _305_;
wire _306_;
wire _307_;
wire _308_;
wire _309_;
wire _310_;
wire _311_;
wire _312_;
wire _313_;
wire _314_;
wire _315_;
wire _316_;
wire _317_;
wire _318_;
wire _319_;
wire _320_;
wire _321_;
wire _322_;
wire _323_;
wire _324_;
wire _325_;
wire _326_;
wire _327_;
wire _328_;
wire _329_;
wire _330_;
wire _331_;
wire _332_;
wire _333_;
wire _334_;
wire _335_;
wire _336_;
wire _337_;
wire _338_;
wire _339_;
wire _340_;
wire _341_;
wire _342_;
wire _343_;
wire _344_;
wire \add_12s_12s_12_2_1_U7.ce ;
wire \add_12s_12s_12_2_1_U7.clk ;
wire [11:0] \add_12s_12s_12_2_1_U7.din0 ;
wire [11:0] \add_12s_12s_12_2_1_U7.din1 ;
wire [11:0] \add_12s_12s_12_2_1_U7.dout ;
wire \add_12s_12s_12_2_1_U7.reset ;
wire [11:0] \add_12s_12s_12_2_1_U7.top_add_12s_12s_12_2_1_Adder_5_U.a ;
wire [11:0] \add_12s_12s_12_2_1_U7.top_add_12s_12s_12_2_1_Adder_5_U.ain_s0 ;
wire [11:0] \add_12s_12s_12_2_1_U7.top_add_12s_12s_12_2_1_Adder_5_U.b ;
wire [11:0] \add_12s_12s_12_2_1_U7.top_add_12s_12s_12_2_1_Adder_5_U.bin_s0 ;
wire \add_12s_12s_12_2_1_U7.top_add_12s_12s_12_2_1_Adder_5_U.ce ;
wire \add_12s_12s_12_2_1_U7.top_add_12s_12s_12_2_1_Adder_5_U.clk ;
wire \add_12s_12s_12_2_1_U7.top_add_12s_12s_12_2_1_Adder_5_U.facout_s1 ;
wire \add_12s_12s_12_2_1_U7.top_add_12s_12s_12_2_1_Adder_5_U.facout_s2 ;
wire [5:0] \add_12s_12s_12_2_1_U7.top_add_12s_12s_12_2_1_Adder_5_U.fas_s1 ;
wire [5:0] \add_12s_12s_12_2_1_U7.top_add_12s_12s_12_2_1_Adder_5_U.fas_s2 ;
wire \add_12s_12s_12_2_1_U7.top_add_12s_12s_12_2_1_Adder_5_U.reset ;
wire [11:0] \add_12s_12s_12_2_1_U7.top_add_12s_12s_12_2_1_Adder_5_U.s ;
wire [5:0] \add_12s_12s_12_2_1_U7.top_add_12s_12s_12_2_1_Adder_5_U.u1.a ;
wire [5:0] \add_12s_12s_12_2_1_U7.top_add_12s_12s_12_2_1_Adder_5_U.u1.b ;
wire \add_12s_12s_12_2_1_U7.top_add_12s_12s_12_2_1_Adder_5_U.u1.cin ;
wire \add_12s_12s_12_2_1_U7.top_add_12s_12s_12_2_1_Adder_5_U.u1.cout ;
wire [5:0] \add_12s_12s_12_2_1_U7.top_add_12s_12s_12_2_1_Adder_5_U.u1.s ;
wire [5:0] \add_12s_12s_12_2_1_U7.top_add_12s_12s_12_2_1_Adder_5_U.u2.a ;
wire [5:0] \add_12s_12s_12_2_1_U7.top_add_12s_12s_12_2_1_Adder_5_U.u2.b ;
wire \add_12s_12s_12_2_1_U7.top_add_12s_12s_12_2_1_Adder_5_U.u2.cin ;
wire \add_12s_12s_12_2_1_U7.top_add_12s_12s_12_2_1_Adder_5_U.u2.cout ;
wire [5:0] \add_12s_12s_12_2_1_U7.top_add_12s_12s_12_2_1_Adder_5_U.u2.s ;
wire \add_18s_18ns_18_2_1_U14.ce ;
wire \add_18s_18ns_18_2_1_U14.clk ;
wire [17:0] \add_18s_18ns_18_2_1_U14.din0 ;
wire [17:0] \add_18s_18ns_18_2_1_U14.din1 ;
wire [17:0] \add_18s_18ns_18_2_1_U14.dout ;
wire \add_18s_18ns_18_2_1_U14.reset ;
wire [17:0] \add_18s_18ns_18_2_1_U14.top_add_18s_18ns_18_2_1_Adder_10_U.a ;
wire [17:0] \add_18s_18ns_18_2_1_U14.top_add_18s_18ns_18_2_1_Adder_10_U.ain_s0 ;
wire [17:0] \add_18s_18ns_18_2_1_U14.top_add_18s_18ns_18_2_1_Adder_10_U.b ;
wire [17:0] \add_18s_18ns_18_2_1_U14.top_add_18s_18ns_18_2_1_Adder_10_U.bin_s0 ;
wire \add_18s_18ns_18_2_1_U14.top_add_18s_18ns_18_2_1_Adder_10_U.ce ;
wire \add_18s_18ns_18_2_1_U14.top_add_18s_18ns_18_2_1_Adder_10_U.clk ;
wire \add_18s_18ns_18_2_1_U14.top_add_18s_18ns_18_2_1_Adder_10_U.facout_s1 ;
wire \add_18s_18ns_18_2_1_U14.top_add_18s_18ns_18_2_1_Adder_10_U.facout_s2 ;
wire [8:0] \add_18s_18ns_18_2_1_U14.top_add_18s_18ns_18_2_1_Adder_10_U.fas_s1 ;
wire [8:0] \add_18s_18ns_18_2_1_U14.top_add_18s_18ns_18_2_1_Adder_10_U.fas_s2 ;
wire \add_18s_18ns_18_2_1_U14.top_add_18s_18ns_18_2_1_Adder_10_U.reset ;
wire [17:0] \add_18s_18ns_18_2_1_U14.top_add_18s_18ns_18_2_1_Adder_10_U.s ;
wire [8:0] \add_18s_18ns_18_2_1_U14.top_add_18s_18ns_18_2_1_Adder_10_U.u1.a ;
wire [8:0] \add_18s_18ns_18_2_1_U14.top_add_18s_18ns_18_2_1_Adder_10_U.u1.b ;
wire \add_18s_18ns_18_2_1_U14.top_add_18s_18ns_18_2_1_Adder_10_U.u1.cin ;
wire \add_18s_18ns_18_2_1_U14.top_add_18s_18ns_18_2_1_Adder_10_U.u1.cout ;
wire [8:0] \add_18s_18ns_18_2_1_U14.top_add_18s_18ns_18_2_1_Adder_10_U.u1.s ;
wire [8:0] \add_18s_18ns_18_2_1_U14.top_add_18s_18ns_18_2_1_Adder_10_U.u2.a ;
wire [8:0] \add_18s_18ns_18_2_1_U14.top_add_18s_18ns_18_2_1_Adder_10_U.u2.b ;
wire \add_18s_18ns_18_2_1_U14.top_add_18s_18ns_18_2_1_Adder_10_U.u2.cin ;
wire \add_18s_18ns_18_2_1_U14.top_add_18s_18ns_18_2_1_Adder_10_U.u2.cout ;
wire [8:0] \add_18s_18ns_18_2_1_U14.top_add_18s_18ns_18_2_1_Adder_10_U.u2.s ;
wire \add_19ns_19s_19_2_1_U17.ce ;
wire \add_19ns_19s_19_2_1_U17.clk ;
wire [18:0] \add_19ns_19s_19_2_1_U17.din0 ;
wire [18:0] \add_19ns_19s_19_2_1_U17.din1 ;
wire [18:0] \add_19ns_19s_19_2_1_U17.dout ;
wire \add_19ns_19s_19_2_1_U17.reset ;
wire [18:0] \add_19ns_19s_19_2_1_U17.top_add_19ns_19s_19_2_1_Adder_13_U.a ;
wire [18:0] \add_19ns_19s_19_2_1_U17.top_add_19ns_19s_19_2_1_Adder_13_U.ain_s0 ;
wire [18:0] \add_19ns_19s_19_2_1_U17.top_add_19ns_19s_19_2_1_Adder_13_U.b ;
wire [18:0] \add_19ns_19s_19_2_1_U17.top_add_19ns_19s_19_2_1_Adder_13_U.bin_s0 ;
wire \add_19ns_19s_19_2_1_U17.top_add_19ns_19s_19_2_1_Adder_13_U.ce ;
wire \add_19ns_19s_19_2_1_U17.top_add_19ns_19s_19_2_1_Adder_13_U.clk ;
wire \add_19ns_19s_19_2_1_U17.top_add_19ns_19s_19_2_1_Adder_13_U.facout_s1 ;
wire \add_19ns_19s_19_2_1_U17.top_add_19ns_19s_19_2_1_Adder_13_U.facout_s2 ;
wire [8:0] \add_19ns_19s_19_2_1_U17.top_add_19ns_19s_19_2_1_Adder_13_U.fas_s1 ;
wire [9:0] \add_19ns_19s_19_2_1_U17.top_add_19ns_19s_19_2_1_Adder_13_U.fas_s2 ;
wire \add_19ns_19s_19_2_1_U17.top_add_19ns_19s_19_2_1_Adder_13_U.reset ;
wire [18:0] \add_19ns_19s_19_2_1_U17.top_add_19ns_19s_19_2_1_Adder_13_U.s ;
wire [8:0] \add_19ns_19s_19_2_1_U17.top_add_19ns_19s_19_2_1_Adder_13_U.u1.a ;
wire [8:0] \add_19ns_19s_19_2_1_U17.top_add_19ns_19s_19_2_1_Adder_13_U.u1.b ;
wire \add_19ns_19s_19_2_1_U17.top_add_19ns_19s_19_2_1_Adder_13_U.u1.cin ;
wire \add_19ns_19s_19_2_1_U17.top_add_19ns_19s_19_2_1_Adder_13_U.u1.cout ;
wire [8:0] \add_19ns_19s_19_2_1_U17.top_add_19ns_19s_19_2_1_Adder_13_U.u1.s ;
wire [9:0] \add_19ns_19s_19_2_1_U17.top_add_19ns_19s_19_2_1_Adder_13_U.u2.a ;
wire [9:0] \add_19ns_19s_19_2_1_U17.top_add_19ns_19s_19_2_1_Adder_13_U.u2.b ;
wire \add_19ns_19s_19_2_1_U17.top_add_19ns_19s_19_2_1_Adder_13_U.u2.cin ;
wire \add_19ns_19s_19_2_1_U17.top_add_19ns_19s_19_2_1_Adder_13_U.u2.cout ;
wire [9:0] \add_19ns_19s_19_2_1_U17.top_add_19ns_19s_19_2_1_Adder_13_U.u2.s ;
wire \add_19s_19ns_19_2_1_U16.ce ;
wire \add_19s_19ns_19_2_1_U16.clk ;
wire [18:0] \add_19s_19ns_19_2_1_U16.din0 ;
wire [18:0] \add_19s_19ns_19_2_1_U16.din1 ;
wire [18:0] \add_19s_19ns_19_2_1_U16.dout ;
wire \add_19s_19ns_19_2_1_U16.reset ;
wire [18:0] \add_19s_19ns_19_2_1_U16.top_add_19s_19ns_19_2_1_Adder_12_U.a ;
wire [18:0] \add_19s_19ns_19_2_1_U16.top_add_19s_19ns_19_2_1_Adder_12_U.ain_s0 ;
wire [18:0] \add_19s_19ns_19_2_1_U16.top_add_19s_19ns_19_2_1_Adder_12_U.b ;
wire [18:0] \add_19s_19ns_19_2_1_U16.top_add_19s_19ns_19_2_1_Adder_12_U.bin_s0 ;
wire \add_19s_19ns_19_2_1_U16.top_add_19s_19ns_19_2_1_Adder_12_U.ce ;
wire \add_19s_19ns_19_2_1_U16.top_add_19s_19ns_19_2_1_Adder_12_U.clk ;
wire \add_19s_19ns_19_2_1_U16.top_add_19s_19ns_19_2_1_Adder_12_U.facout_s1 ;
wire \add_19s_19ns_19_2_1_U16.top_add_19s_19ns_19_2_1_Adder_12_U.facout_s2 ;
wire [8:0] \add_19s_19ns_19_2_1_U16.top_add_19s_19ns_19_2_1_Adder_12_U.fas_s1 ;
wire [9:0] \add_19s_19ns_19_2_1_U16.top_add_19s_19ns_19_2_1_Adder_12_U.fas_s2 ;
wire \add_19s_19ns_19_2_1_U16.top_add_19s_19ns_19_2_1_Adder_12_U.reset ;
wire [18:0] \add_19s_19ns_19_2_1_U16.top_add_19s_19ns_19_2_1_Adder_12_U.s ;
wire [8:0] \add_19s_19ns_19_2_1_U16.top_add_19s_19ns_19_2_1_Adder_12_U.u1.a ;
wire [8:0] \add_19s_19ns_19_2_1_U16.top_add_19s_19ns_19_2_1_Adder_12_U.u1.b ;
wire \add_19s_19ns_19_2_1_U16.top_add_19s_19ns_19_2_1_Adder_12_U.u1.cin ;
wire \add_19s_19ns_19_2_1_U16.top_add_19s_19ns_19_2_1_Adder_12_U.u1.cout ;
wire [8:0] \add_19s_19ns_19_2_1_U16.top_add_19s_19ns_19_2_1_Adder_12_U.u1.s ;
wire [9:0] \add_19s_19ns_19_2_1_U16.top_add_19s_19ns_19_2_1_Adder_12_U.u2.a ;
wire [9:0] \add_19s_19ns_19_2_1_U16.top_add_19s_19ns_19_2_1_Adder_12_U.u2.b ;
wire \add_19s_19ns_19_2_1_U16.top_add_19s_19ns_19_2_1_Adder_12_U.u2.cin ;
wire \add_19s_19ns_19_2_1_U16.top_add_19s_19ns_19_2_1_Adder_12_U.u2.cout ;
wire [9:0] \add_19s_19ns_19_2_1_U16.top_add_19s_19ns_19_2_1_Adder_12_U.u2.s ;
wire \add_19s_19ns_19_2_1_U19.ce ;
wire \add_19s_19ns_19_2_1_U19.clk ;
wire [18:0] \add_19s_19ns_19_2_1_U19.din0 ;
wire [18:0] \add_19s_19ns_19_2_1_U19.din1 ;
wire [18:0] \add_19s_19ns_19_2_1_U19.dout ;
wire \add_19s_19ns_19_2_1_U19.reset ;
wire [18:0] \add_19s_19ns_19_2_1_U19.top_add_19s_19ns_19_2_1_Adder_12_U.a ;
wire [18:0] \add_19s_19ns_19_2_1_U19.top_add_19s_19ns_19_2_1_Adder_12_U.ain_s0 ;
wire [18:0] \add_19s_19ns_19_2_1_U19.top_add_19s_19ns_19_2_1_Adder_12_U.b ;
wire [18:0] \add_19s_19ns_19_2_1_U19.top_add_19s_19ns_19_2_1_Adder_12_U.bin_s0 ;
wire \add_19s_19ns_19_2_1_U19.top_add_19s_19ns_19_2_1_Adder_12_U.ce ;
wire \add_19s_19ns_19_2_1_U19.top_add_19s_19ns_19_2_1_Adder_12_U.clk ;
wire \add_19s_19ns_19_2_1_U19.top_add_19s_19ns_19_2_1_Adder_12_U.facout_s1 ;
wire \add_19s_19ns_19_2_1_U19.top_add_19s_19ns_19_2_1_Adder_12_U.facout_s2 ;
wire [8:0] \add_19s_19ns_19_2_1_U19.top_add_19s_19ns_19_2_1_Adder_12_U.fas_s1 ;
wire [9:0] \add_19s_19ns_19_2_1_U19.top_add_19s_19ns_19_2_1_Adder_12_U.fas_s2 ;
wire \add_19s_19ns_19_2_1_U19.top_add_19s_19ns_19_2_1_Adder_12_U.reset ;
wire [18:0] \add_19s_19ns_19_2_1_U19.top_add_19s_19ns_19_2_1_Adder_12_U.s ;
wire [8:0] \add_19s_19ns_19_2_1_U19.top_add_19s_19ns_19_2_1_Adder_12_U.u1.a ;
wire [8:0] \add_19s_19ns_19_2_1_U19.top_add_19s_19ns_19_2_1_Adder_12_U.u1.b ;
wire \add_19s_19ns_19_2_1_U19.top_add_19s_19ns_19_2_1_Adder_12_U.u1.cin ;
wire \add_19s_19ns_19_2_1_U19.top_add_19s_19ns_19_2_1_Adder_12_U.u1.cout ;
wire [8:0] \add_19s_19ns_19_2_1_U19.top_add_19s_19ns_19_2_1_Adder_12_U.u1.s ;
wire [9:0] \add_19s_19ns_19_2_1_U19.top_add_19s_19ns_19_2_1_Adder_12_U.u2.a ;
wire [9:0] \add_19s_19ns_19_2_1_U19.top_add_19s_19ns_19_2_1_Adder_12_U.u2.b ;
wire \add_19s_19ns_19_2_1_U19.top_add_19s_19ns_19_2_1_Adder_12_U.u2.cin ;
wire \add_19s_19ns_19_2_1_U19.top_add_19s_19ns_19_2_1_Adder_12_U.u2.cout ;
wire [9:0] \add_19s_19ns_19_2_1_U19.top_add_19s_19ns_19_2_1_Adder_12_U.u2.s ;
wire \add_20ns_20s_20_2_1_U15.ce ;
wire \add_20ns_20s_20_2_1_U15.clk ;
wire [19:0] \add_20ns_20s_20_2_1_U15.din0 ;
wire [19:0] \add_20ns_20s_20_2_1_U15.din1 ;
wire [19:0] \add_20ns_20s_20_2_1_U15.dout ;
wire \add_20ns_20s_20_2_1_U15.reset ;
wire [19:0] \add_20ns_20s_20_2_1_U15.top_add_20ns_20s_20_2_1_Adder_11_U.a ;
wire [19:0] \add_20ns_20s_20_2_1_U15.top_add_20ns_20s_20_2_1_Adder_11_U.ain_s0 ;
wire [19:0] \add_20ns_20s_20_2_1_U15.top_add_20ns_20s_20_2_1_Adder_11_U.b ;
wire [19:0] \add_20ns_20s_20_2_1_U15.top_add_20ns_20s_20_2_1_Adder_11_U.bin_s0 ;
wire \add_20ns_20s_20_2_1_U15.top_add_20ns_20s_20_2_1_Adder_11_U.ce ;
wire \add_20ns_20s_20_2_1_U15.top_add_20ns_20s_20_2_1_Adder_11_U.clk ;
wire \add_20ns_20s_20_2_1_U15.top_add_20ns_20s_20_2_1_Adder_11_U.facout_s1 ;
wire \add_20ns_20s_20_2_1_U15.top_add_20ns_20s_20_2_1_Adder_11_U.facout_s2 ;
wire [9:0] \add_20ns_20s_20_2_1_U15.top_add_20ns_20s_20_2_1_Adder_11_U.fas_s1 ;
wire [9:0] \add_20ns_20s_20_2_1_U15.top_add_20ns_20s_20_2_1_Adder_11_U.fas_s2 ;
wire \add_20ns_20s_20_2_1_U15.top_add_20ns_20s_20_2_1_Adder_11_U.reset ;
wire [19:0] \add_20ns_20s_20_2_1_U15.top_add_20ns_20s_20_2_1_Adder_11_U.s ;
wire [9:0] \add_20ns_20s_20_2_1_U15.top_add_20ns_20s_20_2_1_Adder_11_U.u1.a ;
wire [9:0] \add_20ns_20s_20_2_1_U15.top_add_20ns_20s_20_2_1_Adder_11_U.u1.b ;
wire \add_20ns_20s_20_2_1_U15.top_add_20ns_20s_20_2_1_Adder_11_U.u1.cin ;
wire \add_20ns_20s_20_2_1_U15.top_add_20ns_20s_20_2_1_Adder_11_U.u1.cout ;
wire [9:0] \add_20ns_20s_20_2_1_U15.top_add_20ns_20s_20_2_1_Adder_11_U.u1.s ;
wire [9:0] \add_20ns_20s_20_2_1_U15.top_add_20ns_20s_20_2_1_Adder_11_U.u2.a ;
wire [9:0] \add_20ns_20s_20_2_1_U15.top_add_20ns_20s_20_2_1_Adder_11_U.u2.b ;
wire \add_20ns_20s_20_2_1_U15.top_add_20ns_20s_20_2_1_Adder_11_U.u2.cin ;
wire \add_20ns_20s_20_2_1_U15.top_add_20ns_20s_20_2_1_Adder_11_U.u2.cout ;
wire [9:0] \add_20ns_20s_20_2_1_U15.top_add_20ns_20s_20_2_1_Adder_11_U.u2.s ;
wire \add_2ns_2ns_2_2_1_U10.ce ;
wire \add_2ns_2ns_2_2_1_U10.clk ;
wire [1:0] \add_2ns_2ns_2_2_1_U10.din0 ;
wire [1:0] \add_2ns_2ns_2_2_1_U10.din1 ;
wire [1:0] \add_2ns_2ns_2_2_1_U10.dout ;
wire \add_2ns_2ns_2_2_1_U10.reset ;
wire [1:0] \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_6_U.a ;
wire [1:0] \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_6_U.ain_s0 ;
wire [1:0] \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_6_U.b ;
wire [1:0] \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_6_U.bin_s0 ;
wire \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_6_U.ce ;
wire \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_6_U.clk ;
wire \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_6_U.facout_s1 ;
wire \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_6_U.facout_s2 ;
wire \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_6_U.fas_s1 ;
wire \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_6_U.fas_s2 ;
wire \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_6_U.reset ;
wire [1:0] \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_6_U.s ;
wire \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_6_U.u1.a ;
wire \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_6_U.u1.b ;
wire \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_6_U.u1.cin ;
wire \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_6_U.u1.cout ;
wire \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_6_U.u1.s ;
wire \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_6_U.u2.a ;
wire \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_6_U.u2.b ;
wire \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_6_U.u2.cin ;
wire \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_6_U.u2.cout ;
wire \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_6_U.u2.s ;
wire \add_2ns_2ns_2_2_1_U18.ce ;
wire \add_2ns_2ns_2_2_1_U18.clk ;
wire [1:0] \add_2ns_2ns_2_2_1_U18.din0 ;
wire [1:0] \add_2ns_2ns_2_2_1_U18.din1 ;
wire [1:0] \add_2ns_2ns_2_2_1_U18.dout ;
wire \add_2ns_2ns_2_2_1_U18.reset ;
wire [1:0] \add_2ns_2ns_2_2_1_U18.top_add_2ns_2ns_2_2_1_Adder_6_U.a ;
wire [1:0] \add_2ns_2ns_2_2_1_U18.top_add_2ns_2ns_2_2_1_Adder_6_U.ain_s0 ;
wire [1:0] \add_2ns_2ns_2_2_1_U18.top_add_2ns_2ns_2_2_1_Adder_6_U.b ;
wire [1:0] \add_2ns_2ns_2_2_1_U18.top_add_2ns_2ns_2_2_1_Adder_6_U.bin_s0 ;
wire \add_2ns_2ns_2_2_1_U18.top_add_2ns_2ns_2_2_1_Adder_6_U.ce ;
wire \add_2ns_2ns_2_2_1_U18.top_add_2ns_2ns_2_2_1_Adder_6_U.clk ;
wire \add_2ns_2ns_2_2_1_U18.top_add_2ns_2ns_2_2_1_Adder_6_U.facout_s1 ;
wire \add_2ns_2ns_2_2_1_U18.top_add_2ns_2ns_2_2_1_Adder_6_U.facout_s2 ;
wire \add_2ns_2ns_2_2_1_U18.top_add_2ns_2ns_2_2_1_Adder_6_U.fas_s1 ;
wire \add_2ns_2ns_2_2_1_U18.top_add_2ns_2ns_2_2_1_Adder_6_U.fas_s2 ;
wire \add_2ns_2ns_2_2_1_U18.top_add_2ns_2ns_2_2_1_Adder_6_U.reset ;
wire [1:0] \add_2ns_2ns_2_2_1_U18.top_add_2ns_2ns_2_2_1_Adder_6_U.s ;
wire \add_2ns_2ns_2_2_1_U18.top_add_2ns_2ns_2_2_1_Adder_6_U.u1.a ;
wire \add_2ns_2ns_2_2_1_U18.top_add_2ns_2ns_2_2_1_Adder_6_U.u1.b ;
wire \add_2ns_2ns_2_2_1_U18.top_add_2ns_2ns_2_2_1_Adder_6_U.u1.cin ;
wire \add_2ns_2ns_2_2_1_U18.top_add_2ns_2ns_2_2_1_Adder_6_U.u1.cout ;
wire \add_2ns_2ns_2_2_1_U18.top_add_2ns_2ns_2_2_1_Adder_6_U.u1.s ;
wire \add_2ns_2ns_2_2_1_U18.top_add_2ns_2ns_2_2_1_Adder_6_U.u2.a ;
wire \add_2ns_2ns_2_2_1_U18.top_add_2ns_2ns_2_2_1_Adder_6_U.u2.b ;
wire \add_2ns_2ns_2_2_1_U18.top_add_2ns_2ns_2_2_1_Adder_6_U.u2.cin ;
wire \add_2ns_2ns_2_2_1_U18.top_add_2ns_2ns_2_2_1_Adder_6_U.u2.cout ;
wire \add_2ns_2ns_2_2_1_U18.top_add_2ns_2ns_2_2_1_Adder_6_U.u2.s ;
wire \add_2ns_2s_2_2_1_U2.ce ;
wire \add_2ns_2s_2_2_1_U2.clk ;
wire [1:0] \add_2ns_2s_2_2_1_U2.din0 ;
wire [1:0] \add_2ns_2s_2_2_1_U2.din1 ;
wire [1:0] \add_2ns_2s_2_2_1_U2.dout ;
wire \add_2ns_2s_2_2_1_U2.reset ;
wire [1:0] \add_2ns_2s_2_2_1_U2.top_add_2ns_2s_2_2_1_Adder_0_U.a ;
wire [1:0] \add_2ns_2s_2_2_1_U2.top_add_2ns_2s_2_2_1_Adder_0_U.ain_s0 ;
wire [1:0] \add_2ns_2s_2_2_1_U2.top_add_2ns_2s_2_2_1_Adder_0_U.b ;
wire [1:0] \add_2ns_2s_2_2_1_U2.top_add_2ns_2s_2_2_1_Adder_0_U.bin_s0 ;
wire \add_2ns_2s_2_2_1_U2.top_add_2ns_2s_2_2_1_Adder_0_U.ce ;
wire \add_2ns_2s_2_2_1_U2.top_add_2ns_2s_2_2_1_Adder_0_U.clk ;
wire \add_2ns_2s_2_2_1_U2.top_add_2ns_2s_2_2_1_Adder_0_U.facout_s1 ;
wire \add_2ns_2s_2_2_1_U2.top_add_2ns_2s_2_2_1_Adder_0_U.facout_s2 ;
wire \add_2ns_2s_2_2_1_U2.top_add_2ns_2s_2_2_1_Adder_0_U.fas_s1 ;
wire \add_2ns_2s_2_2_1_U2.top_add_2ns_2s_2_2_1_Adder_0_U.fas_s2 ;
wire \add_2ns_2s_2_2_1_U2.top_add_2ns_2s_2_2_1_Adder_0_U.reset ;
wire [1:0] \add_2ns_2s_2_2_1_U2.top_add_2ns_2s_2_2_1_Adder_0_U.s ;
wire \add_2ns_2s_2_2_1_U2.top_add_2ns_2s_2_2_1_Adder_0_U.u1.a ;
wire \add_2ns_2s_2_2_1_U2.top_add_2ns_2s_2_2_1_Adder_0_U.u1.b ;
wire \add_2ns_2s_2_2_1_U2.top_add_2ns_2s_2_2_1_Adder_0_U.u1.cin ;
wire \add_2ns_2s_2_2_1_U2.top_add_2ns_2s_2_2_1_Adder_0_U.u1.cout ;
wire \add_2ns_2s_2_2_1_U2.top_add_2ns_2s_2_2_1_Adder_0_U.u1.s ;
wire \add_2ns_2s_2_2_1_U2.top_add_2ns_2s_2_2_1_Adder_0_U.u2.a ;
wire \add_2ns_2s_2_2_1_U2.top_add_2ns_2s_2_2_1_Adder_0_U.u2.b ;
wire \add_2ns_2s_2_2_1_U2.top_add_2ns_2s_2_2_1_Adder_0_U.u2.cin ;
wire \add_2ns_2s_2_2_1_U2.top_add_2ns_2s_2_2_1_Adder_0_U.u2.cout ;
wire \add_2ns_2s_2_2_1_U2.top_add_2ns_2s_2_2_1_Adder_0_U.u2.s ;
wire \add_32ns_32ns_32_2_1_U21.ce ;
wire \add_32ns_32ns_32_2_1_U21.clk ;
wire [31:0] \add_32ns_32ns_32_2_1_U21.din0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U21.din1 ;
wire [31:0] \add_32ns_32ns_32_2_1_U21.dout ;
wire \add_32ns_32ns_32_2_1_U21.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.a ;
wire [31:0] \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.ain_s0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.b ;
wire [31:0] \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.bin_s0 ;
wire \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.ce ;
wire \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.clk ;
wire \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.facout_s1 ;
wire \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.facout_s2 ;
wire [15:0] \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.fas_s1 ;
wire [15:0] \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.fas_s2 ;
wire \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.b ;
wire \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.cin ;
wire \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.b ;
wire \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.cin ;
wire \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.s ;
wire \add_32ns_32ns_32_2_1_U23.ce ;
wire \add_32ns_32ns_32_2_1_U23.clk ;
wire [31:0] \add_32ns_32ns_32_2_1_U23.din0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U23.din1 ;
wire [31:0] \add_32ns_32ns_32_2_1_U23.dout ;
wire \add_32ns_32ns_32_2_1_U23.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.a ;
wire [31:0] \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.ain_s0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.b ;
wire [31:0] \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.bin_s0 ;
wire \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.ce ;
wire \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.clk ;
wire \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.facout_s1 ;
wire \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.facout_s2 ;
wire [15:0] \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.fas_s1 ;
wire [15:0] \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.fas_s2 ;
wire \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.b ;
wire \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.cin ;
wire \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.b ;
wire \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.cin ;
wire \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.s ;
wire \add_32ns_32ns_32_2_1_U25.ce ;
wire \add_32ns_32ns_32_2_1_U25.clk ;
wire [31:0] \add_32ns_32ns_32_2_1_U25.din0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U25.din1 ;
wire [31:0] \add_32ns_32ns_32_2_1_U25.dout ;
wire \add_32ns_32ns_32_2_1_U25.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.a ;
wire [31:0] \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.ain_s0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.b ;
wire [31:0] \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.bin_s0 ;
wire \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.ce ;
wire \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.clk ;
wire \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.facout_s1 ;
wire \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.facout_s2 ;
wire [15:0] \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.fas_s1 ;
wire [15:0] \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.fas_s2 ;
wire \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.b ;
wire \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.cin ;
wire \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.b ;
wire \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.cin ;
wire \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.s ;
wire \add_32ns_32ns_32_2_1_U26.ce ;
wire \add_32ns_32ns_32_2_1_U26.clk ;
wire [31:0] \add_32ns_32ns_32_2_1_U26.din0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U26.din1 ;
wire [31:0] \add_32ns_32ns_32_2_1_U26.dout ;
wire \add_32ns_32ns_32_2_1_U26.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U26.top_add_32ns_32ns_32_2_1_Adder_15_U.a ;
wire [31:0] \add_32ns_32ns_32_2_1_U26.top_add_32ns_32ns_32_2_1_Adder_15_U.ain_s0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U26.top_add_32ns_32ns_32_2_1_Adder_15_U.b ;
wire [31:0] \add_32ns_32ns_32_2_1_U26.top_add_32ns_32ns_32_2_1_Adder_15_U.bin_s0 ;
wire \add_32ns_32ns_32_2_1_U26.top_add_32ns_32ns_32_2_1_Adder_15_U.ce ;
wire \add_32ns_32ns_32_2_1_U26.top_add_32ns_32ns_32_2_1_Adder_15_U.clk ;
wire \add_32ns_32ns_32_2_1_U26.top_add_32ns_32ns_32_2_1_Adder_15_U.facout_s1 ;
wire \add_32ns_32ns_32_2_1_U26.top_add_32ns_32ns_32_2_1_Adder_15_U.facout_s2 ;
wire [15:0] \add_32ns_32ns_32_2_1_U26.top_add_32ns_32ns_32_2_1_Adder_15_U.fas_s1 ;
wire [15:0] \add_32ns_32ns_32_2_1_U26.top_add_32ns_32ns_32_2_1_Adder_15_U.fas_s2 ;
wire \add_32ns_32ns_32_2_1_U26.top_add_32ns_32ns_32_2_1_Adder_15_U.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U26.top_add_32ns_32ns_32_2_1_Adder_15_U.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U26.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U26.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.b ;
wire \add_32ns_32ns_32_2_1_U26.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.cin ;
wire \add_32ns_32ns_32_2_1_U26.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U26.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U26.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U26.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.b ;
wire \add_32ns_32ns_32_2_1_U26.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.cin ;
wire \add_32ns_32ns_32_2_1_U26.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U26.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.s ;
wire \add_35s_35s_35_2_1_U24.ce ;
wire \add_35s_35s_35_2_1_U24.clk ;
wire [34:0] \add_35s_35s_35_2_1_U24.din0 ;
wire [34:0] \add_35s_35s_35_2_1_U24.din1 ;
wire [34:0] \add_35s_35s_35_2_1_U24.dout ;
wire \add_35s_35s_35_2_1_U24.reset ;
wire [34:0] \add_35s_35s_35_2_1_U24.top_add_35s_35s_35_2_1_Adder_17_U.a ;
wire [34:0] \add_35s_35s_35_2_1_U24.top_add_35s_35s_35_2_1_Adder_17_U.ain_s0 ;
wire [34:0] \add_35s_35s_35_2_1_U24.top_add_35s_35s_35_2_1_Adder_17_U.b ;
wire [34:0] \add_35s_35s_35_2_1_U24.top_add_35s_35s_35_2_1_Adder_17_U.bin_s0 ;
wire \add_35s_35s_35_2_1_U24.top_add_35s_35s_35_2_1_Adder_17_U.ce ;
wire \add_35s_35s_35_2_1_U24.top_add_35s_35s_35_2_1_Adder_17_U.clk ;
wire \add_35s_35s_35_2_1_U24.top_add_35s_35s_35_2_1_Adder_17_U.facout_s1 ;
wire \add_35s_35s_35_2_1_U24.top_add_35s_35s_35_2_1_Adder_17_U.facout_s2 ;
wire [16:0] \add_35s_35s_35_2_1_U24.top_add_35s_35s_35_2_1_Adder_17_U.fas_s1 ;
wire [17:0] \add_35s_35s_35_2_1_U24.top_add_35s_35s_35_2_1_Adder_17_U.fas_s2 ;
wire \add_35s_35s_35_2_1_U24.top_add_35s_35s_35_2_1_Adder_17_U.reset ;
wire [34:0] \add_35s_35s_35_2_1_U24.top_add_35s_35s_35_2_1_Adder_17_U.s ;
wire [16:0] \add_35s_35s_35_2_1_U24.top_add_35s_35s_35_2_1_Adder_17_U.u1.a ;
wire [16:0] \add_35s_35s_35_2_1_U24.top_add_35s_35s_35_2_1_Adder_17_U.u1.b ;
wire \add_35s_35s_35_2_1_U24.top_add_35s_35s_35_2_1_Adder_17_U.u1.cin ;
wire \add_35s_35s_35_2_1_U24.top_add_35s_35s_35_2_1_Adder_17_U.u1.cout ;
wire [16:0] \add_35s_35s_35_2_1_U24.top_add_35s_35s_35_2_1_Adder_17_U.u1.s ;
wire [17:0] \add_35s_35s_35_2_1_U24.top_add_35s_35s_35_2_1_Adder_17_U.u2.a ;
wire [17:0] \add_35s_35s_35_2_1_U24.top_add_35s_35s_35_2_1_Adder_17_U.u2.b ;
wire \add_35s_35s_35_2_1_U24.top_add_35s_35s_35_2_1_Adder_17_U.u2.cin ;
wire \add_35s_35s_35_2_1_U24.top_add_35s_35s_35_2_1_Adder_17_U.u2.cout ;
wire [17:0] \add_35s_35s_35_2_1_U24.top_add_35s_35s_35_2_1_Adder_17_U.u2.s ;
wire \add_37s_37s_37_2_1_U20.ce ;
wire \add_37s_37s_37_2_1_U20.clk ;
wire [36:0] \add_37s_37s_37_2_1_U20.din0 ;
wire [36:0] \add_37s_37s_37_2_1_U20.din1 ;
wire [36:0] \add_37s_37s_37_2_1_U20.dout ;
wire \add_37s_37s_37_2_1_U20.reset ;
wire [36:0] \add_37s_37s_37_2_1_U20.top_add_37s_37s_37_2_1_Adder_14_U.a ;
wire [36:0] \add_37s_37s_37_2_1_U20.top_add_37s_37s_37_2_1_Adder_14_U.ain_s0 ;
wire [36:0] \add_37s_37s_37_2_1_U20.top_add_37s_37s_37_2_1_Adder_14_U.b ;
wire [36:0] \add_37s_37s_37_2_1_U20.top_add_37s_37s_37_2_1_Adder_14_U.bin_s0 ;
wire \add_37s_37s_37_2_1_U20.top_add_37s_37s_37_2_1_Adder_14_U.ce ;
wire \add_37s_37s_37_2_1_U20.top_add_37s_37s_37_2_1_Adder_14_U.clk ;
wire \add_37s_37s_37_2_1_U20.top_add_37s_37s_37_2_1_Adder_14_U.facout_s1 ;
wire \add_37s_37s_37_2_1_U20.top_add_37s_37s_37_2_1_Adder_14_U.facout_s2 ;
wire [17:0] \add_37s_37s_37_2_1_U20.top_add_37s_37s_37_2_1_Adder_14_U.fas_s1 ;
wire [18:0] \add_37s_37s_37_2_1_U20.top_add_37s_37s_37_2_1_Adder_14_U.fas_s2 ;
wire \add_37s_37s_37_2_1_U20.top_add_37s_37s_37_2_1_Adder_14_U.reset ;
wire [36:0] \add_37s_37s_37_2_1_U20.top_add_37s_37s_37_2_1_Adder_14_U.s ;
wire [17:0] \add_37s_37s_37_2_1_U20.top_add_37s_37s_37_2_1_Adder_14_U.u1.a ;
wire [17:0] \add_37s_37s_37_2_1_U20.top_add_37s_37s_37_2_1_Adder_14_U.u1.b ;
wire \add_37s_37s_37_2_1_U20.top_add_37s_37s_37_2_1_Adder_14_U.u1.cin ;
wire \add_37s_37s_37_2_1_U20.top_add_37s_37s_37_2_1_Adder_14_U.u1.cout ;
wire [17:0] \add_37s_37s_37_2_1_U20.top_add_37s_37s_37_2_1_Adder_14_U.u1.s ;
wire [18:0] \add_37s_37s_37_2_1_U20.top_add_37s_37s_37_2_1_Adder_14_U.u2.a ;
wire [18:0] \add_37s_37s_37_2_1_U20.top_add_37s_37s_37_2_1_Adder_14_U.u2.b ;
wire \add_37s_37s_37_2_1_U20.top_add_37s_37s_37_2_1_Adder_14_U.u2.cin ;
wire \add_37s_37s_37_2_1_U20.top_add_37s_37s_37_2_1_Adder_14_U.u2.cout ;
wire [18:0] \add_37s_37s_37_2_1_U20.top_add_37s_37s_37_2_1_Adder_14_U.u2.s ;
wire \add_3s_3s_3_2_1_U4.ce ;
wire \add_3s_3s_3_2_1_U4.clk ;
wire [2:0] \add_3s_3s_3_2_1_U4.din0 ;
wire [2:0] \add_3s_3s_3_2_1_U4.din1 ;
wire [2:0] \add_3s_3s_3_2_1_U4.dout ;
wire \add_3s_3s_3_2_1_U4.reset ;
wire [2:0] \add_3s_3s_3_2_1_U4.top_add_3s_3s_3_2_1_Adder_2_U.a ;
wire [2:0] \add_3s_3s_3_2_1_U4.top_add_3s_3s_3_2_1_Adder_2_U.ain_s0 ;
wire [2:0] \add_3s_3s_3_2_1_U4.top_add_3s_3s_3_2_1_Adder_2_U.b ;
wire [2:0] \add_3s_3s_3_2_1_U4.top_add_3s_3s_3_2_1_Adder_2_U.bin_s0 ;
wire \add_3s_3s_3_2_1_U4.top_add_3s_3s_3_2_1_Adder_2_U.ce ;
wire \add_3s_3s_3_2_1_U4.top_add_3s_3s_3_2_1_Adder_2_U.clk ;
wire \add_3s_3s_3_2_1_U4.top_add_3s_3s_3_2_1_Adder_2_U.facout_s1 ;
wire \add_3s_3s_3_2_1_U4.top_add_3s_3s_3_2_1_Adder_2_U.facout_s2 ;
wire \add_3s_3s_3_2_1_U4.top_add_3s_3s_3_2_1_Adder_2_U.fas_s1 ;
wire [1:0] \add_3s_3s_3_2_1_U4.top_add_3s_3s_3_2_1_Adder_2_U.fas_s2 ;
wire \add_3s_3s_3_2_1_U4.top_add_3s_3s_3_2_1_Adder_2_U.reset ;
wire [2:0] \add_3s_3s_3_2_1_U4.top_add_3s_3s_3_2_1_Adder_2_U.s ;
wire \add_3s_3s_3_2_1_U4.top_add_3s_3s_3_2_1_Adder_2_U.u1.a ;
wire \add_3s_3s_3_2_1_U4.top_add_3s_3s_3_2_1_Adder_2_U.u1.b ;
wire \add_3s_3s_3_2_1_U4.top_add_3s_3s_3_2_1_Adder_2_U.u1.cin ;
wire \add_3s_3s_3_2_1_U4.top_add_3s_3s_3_2_1_Adder_2_U.u1.cout ;
wire \add_3s_3s_3_2_1_U4.top_add_3s_3s_3_2_1_Adder_2_U.u1.s ;
wire [1:0] \add_3s_3s_3_2_1_U4.top_add_3s_3s_3_2_1_Adder_2_U.u2.a ;
wire [1:0] \add_3s_3s_3_2_1_U4.top_add_3s_3s_3_2_1_Adder_2_U.u2.b ;
wire \add_3s_3s_3_2_1_U4.top_add_3s_3s_3_2_1_Adder_2_U.u2.cin ;
wire \add_3s_3s_3_2_1_U4.top_add_3s_3s_3_2_1_Adder_2_U.u2.cout ;
wire [1:0] \add_3s_3s_3_2_1_U4.top_add_3s_3s_3_2_1_Adder_2_U.u2.s ;
wire \add_57s_57s_57_2_1_U22.ce ;
wire \add_57s_57s_57_2_1_U22.clk ;
wire [56:0] \add_57s_57s_57_2_1_U22.din0 ;
wire [56:0] \add_57s_57s_57_2_1_U22.din1 ;
wire [56:0] \add_57s_57s_57_2_1_U22.dout ;
wire \add_57s_57s_57_2_1_U22.reset ;
wire [56:0] \add_57s_57s_57_2_1_U22.top_add_57s_57s_57_2_1_Adder_16_U.a ;
wire [56:0] \add_57s_57s_57_2_1_U22.top_add_57s_57s_57_2_1_Adder_16_U.ain_s0 ;
wire [56:0] \add_57s_57s_57_2_1_U22.top_add_57s_57s_57_2_1_Adder_16_U.b ;
wire [56:0] \add_57s_57s_57_2_1_U22.top_add_57s_57s_57_2_1_Adder_16_U.bin_s0 ;
wire \add_57s_57s_57_2_1_U22.top_add_57s_57s_57_2_1_Adder_16_U.ce ;
wire \add_57s_57s_57_2_1_U22.top_add_57s_57s_57_2_1_Adder_16_U.clk ;
wire \add_57s_57s_57_2_1_U22.top_add_57s_57s_57_2_1_Adder_16_U.facout_s1 ;
wire \add_57s_57s_57_2_1_U22.top_add_57s_57s_57_2_1_Adder_16_U.facout_s2 ;
wire [27:0] \add_57s_57s_57_2_1_U22.top_add_57s_57s_57_2_1_Adder_16_U.fas_s1 ;
wire [28:0] \add_57s_57s_57_2_1_U22.top_add_57s_57s_57_2_1_Adder_16_U.fas_s2 ;
wire \add_57s_57s_57_2_1_U22.top_add_57s_57s_57_2_1_Adder_16_U.reset ;
wire [56:0] \add_57s_57s_57_2_1_U22.top_add_57s_57s_57_2_1_Adder_16_U.s ;
wire [27:0] \add_57s_57s_57_2_1_U22.top_add_57s_57s_57_2_1_Adder_16_U.u1.a ;
wire [27:0] \add_57s_57s_57_2_1_U22.top_add_57s_57s_57_2_1_Adder_16_U.u1.b ;
wire \add_57s_57s_57_2_1_U22.top_add_57s_57s_57_2_1_Adder_16_U.u1.cin ;
wire \add_57s_57s_57_2_1_U22.top_add_57s_57s_57_2_1_Adder_16_U.u1.cout ;
wire [27:0] \add_57s_57s_57_2_1_U22.top_add_57s_57s_57_2_1_Adder_16_U.u1.s ;
wire [28:0] \add_57s_57s_57_2_1_U22.top_add_57s_57s_57_2_1_Adder_16_U.u2.a ;
wire [28:0] \add_57s_57s_57_2_1_U22.top_add_57s_57s_57_2_1_Adder_16_U.u2.b ;
wire \add_57s_57s_57_2_1_U22.top_add_57s_57s_57_2_1_Adder_16_U.u2.cin ;
wire \add_57s_57s_57_2_1_U22.top_add_57s_57s_57_2_1_Adder_16_U.u2.cout ;
wire [28:0] \add_57s_57s_57_2_1_U22.top_add_57s_57s_57_2_1_Adder_16_U.u2.s ;
wire \add_6ns_6ns_6_2_1_U12.ce ;
wire \add_6ns_6ns_6_2_1_U12.clk ;
wire [5:0] \add_6ns_6ns_6_2_1_U12.din0 ;
wire [5:0] \add_6ns_6ns_6_2_1_U12.din1 ;
wire [5:0] \add_6ns_6ns_6_2_1_U12.dout ;
wire \add_6ns_6ns_6_2_1_U12.reset ;
wire [5:0] \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_8_U.a ;
wire [5:0] \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_8_U.ain_s0 ;
wire [5:0] \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_8_U.b ;
wire [5:0] \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_8_U.bin_s0 ;
wire \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_8_U.ce ;
wire \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_8_U.clk ;
wire \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_8_U.facout_s1 ;
wire \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_8_U.facout_s2 ;
wire [2:0] \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_8_U.fas_s1 ;
wire [2:0] \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_8_U.fas_s2 ;
wire \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_8_U.reset ;
wire [5:0] \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_8_U.s ;
wire [2:0] \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_8_U.u1.a ;
wire [2:0] \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_8_U.u1.b ;
wire \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_8_U.u1.cin ;
wire \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_8_U.u1.cout ;
wire [2:0] \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_8_U.u1.s ;
wire [2:0] \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_8_U.u2.a ;
wire [2:0] \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_8_U.u2.b ;
wire \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_8_U.u2.cin ;
wire \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_8_U.u2.cout ;
wire [2:0] \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_8_U.u2.s ;
wire \add_7ns_7ns_7_2_1_U3.ce ;
wire \add_7ns_7ns_7_2_1_U3.clk ;
wire [6:0] \add_7ns_7ns_7_2_1_U3.din0 ;
wire [6:0] \add_7ns_7ns_7_2_1_U3.din1 ;
wire [6:0] \add_7ns_7ns_7_2_1_U3.dout ;
wire \add_7ns_7ns_7_2_1_U3.reset ;
wire [6:0] \add_7ns_7ns_7_2_1_U3.top_add_7ns_7ns_7_2_1_Adder_1_U.a ;
wire [6:0] \add_7ns_7ns_7_2_1_U3.top_add_7ns_7ns_7_2_1_Adder_1_U.ain_s0 ;
wire [6:0] \add_7ns_7ns_7_2_1_U3.top_add_7ns_7ns_7_2_1_Adder_1_U.b ;
wire [6:0] \add_7ns_7ns_7_2_1_U3.top_add_7ns_7ns_7_2_1_Adder_1_U.bin_s0 ;
wire \add_7ns_7ns_7_2_1_U3.top_add_7ns_7ns_7_2_1_Adder_1_U.ce ;
wire \add_7ns_7ns_7_2_1_U3.top_add_7ns_7ns_7_2_1_Adder_1_U.clk ;
wire \add_7ns_7ns_7_2_1_U3.top_add_7ns_7ns_7_2_1_Adder_1_U.facout_s1 ;
wire \add_7ns_7ns_7_2_1_U3.top_add_7ns_7ns_7_2_1_Adder_1_U.facout_s2 ;
wire [2:0] \add_7ns_7ns_7_2_1_U3.top_add_7ns_7ns_7_2_1_Adder_1_U.fas_s1 ;
wire [3:0] \add_7ns_7ns_7_2_1_U3.top_add_7ns_7ns_7_2_1_Adder_1_U.fas_s2 ;
wire \add_7ns_7ns_7_2_1_U3.top_add_7ns_7ns_7_2_1_Adder_1_U.reset ;
wire [6:0] \add_7ns_7ns_7_2_1_U3.top_add_7ns_7ns_7_2_1_Adder_1_U.s ;
wire [2:0] \add_7ns_7ns_7_2_1_U3.top_add_7ns_7ns_7_2_1_Adder_1_U.u1.a ;
wire [2:0] \add_7ns_7ns_7_2_1_U3.top_add_7ns_7ns_7_2_1_Adder_1_U.u1.b ;
wire \add_7ns_7ns_7_2_1_U3.top_add_7ns_7ns_7_2_1_Adder_1_U.u1.cin ;
wire \add_7ns_7ns_7_2_1_U3.top_add_7ns_7ns_7_2_1_Adder_1_U.u1.cout ;
wire [2:0] \add_7ns_7ns_7_2_1_U3.top_add_7ns_7ns_7_2_1_Adder_1_U.u1.s ;
wire [3:0] \add_7ns_7ns_7_2_1_U3.top_add_7ns_7ns_7_2_1_Adder_1_U.u2.a ;
wire [3:0] \add_7ns_7ns_7_2_1_U3.top_add_7ns_7ns_7_2_1_Adder_1_U.u2.b ;
wire \add_7ns_7ns_7_2_1_U3.top_add_7ns_7ns_7_2_1_Adder_1_U.u2.cin ;
wire \add_7ns_7ns_7_2_1_U3.top_add_7ns_7ns_7_2_1_Adder_1_U.u2.cout ;
wire [3:0] \add_7ns_7ns_7_2_1_U3.top_add_7ns_7ns_7_2_1_Adder_1_U.u2.s ;
wire \add_7s_7s_7_2_1_U13.ce ;
wire \add_7s_7s_7_2_1_U13.clk ;
wire [6:0] \add_7s_7s_7_2_1_U13.din0 ;
wire [6:0] \add_7s_7s_7_2_1_U13.din1 ;
wire [6:0] \add_7s_7s_7_2_1_U13.dout ;
wire \add_7s_7s_7_2_1_U13.reset ;
wire [6:0] \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_9_U.a ;
wire [6:0] \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_9_U.ain_s0 ;
wire [6:0] \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_9_U.b ;
wire [6:0] \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_9_U.bin_s0 ;
wire \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_9_U.ce ;
wire \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_9_U.clk ;
wire \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_9_U.facout_s1 ;
wire \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_9_U.facout_s2 ;
wire [2:0] \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_9_U.fas_s1 ;
wire [3:0] \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_9_U.fas_s2 ;
wire \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_9_U.reset ;
wire [6:0] \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_9_U.s ;
wire [2:0] \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_9_U.u1.a ;
wire [2:0] \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_9_U.u1.b ;
wire \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_9_U.u1.cin ;
wire \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_9_U.u1.cout ;
wire [2:0] \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_9_U.u1.s ;
wire [3:0] \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_9_U.u2.a ;
wire [3:0] \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_9_U.u2.b ;
wire \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_9_U.u2.cin ;
wire \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_9_U.u2.cout ;
wire [3:0] \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_9_U.u2.s ;
wire \add_9ns_9s_9_2_1_U11.ce ;
wire \add_9ns_9s_9_2_1_U11.clk ;
wire [8:0] \add_9ns_9s_9_2_1_U11.din0 ;
wire [8:0] \add_9ns_9s_9_2_1_U11.din1 ;
wire [8:0] \add_9ns_9s_9_2_1_U11.dout ;
wire \add_9ns_9s_9_2_1_U11.reset ;
wire [8:0] \add_9ns_9s_9_2_1_U11.top_add_9ns_9s_9_2_1_Adder_7_U.a ;
wire [8:0] \add_9ns_9s_9_2_1_U11.top_add_9ns_9s_9_2_1_Adder_7_U.ain_s0 ;
wire [8:0] \add_9ns_9s_9_2_1_U11.top_add_9ns_9s_9_2_1_Adder_7_U.b ;
wire [8:0] \add_9ns_9s_9_2_1_U11.top_add_9ns_9s_9_2_1_Adder_7_U.bin_s0 ;
wire \add_9ns_9s_9_2_1_U11.top_add_9ns_9s_9_2_1_Adder_7_U.ce ;
wire \add_9ns_9s_9_2_1_U11.top_add_9ns_9s_9_2_1_Adder_7_U.clk ;
wire \add_9ns_9s_9_2_1_U11.top_add_9ns_9s_9_2_1_Adder_7_U.facout_s1 ;
wire \add_9ns_9s_9_2_1_U11.top_add_9ns_9s_9_2_1_Adder_7_U.facout_s2 ;
wire [3:0] \add_9ns_9s_9_2_1_U11.top_add_9ns_9s_9_2_1_Adder_7_U.fas_s1 ;
wire [4:0] \add_9ns_9s_9_2_1_U11.top_add_9ns_9s_9_2_1_Adder_7_U.fas_s2 ;
wire \add_9ns_9s_9_2_1_U11.top_add_9ns_9s_9_2_1_Adder_7_U.reset ;
wire [8:0] \add_9ns_9s_9_2_1_U11.top_add_9ns_9s_9_2_1_Adder_7_U.s ;
wire [3:0] \add_9ns_9s_9_2_1_U11.top_add_9ns_9s_9_2_1_Adder_7_U.u1.a ;
wire [3:0] \add_9ns_9s_9_2_1_U11.top_add_9ns_9s_9_2_1_Adder_7_U.u1.b ;
wire \add_9ns_9s_9_2_1_U11.top_add_9ns_9s_9_2_1_Adder_7_U.u1.cin ;
wire \add_9ns_9s_9_2_1_U11.top_add_9ns_9s_9_2_1_Adder_7_U.u1.cout ;
wire [3:0] \add_9ns_9s_9_2_1_U11.top_add_9ns_9s_9_2_1_Adder_7_U.u1.s ;
wire [4:0] \add_9ns_9s_9_2_1_U11.top_add_9ns_9s_9_2_1_Adder_7_U.u2.a ;
wire [4:0] \add_9ns_9s_9_2_1_U11.top_add_9ns_9s_9_2_1_Adder_7_U.u2.b ;
wire \add_9ns_9s_9_2_1_U11.top_add_9ns_9s_9_2_1_Adder_7_U.u2.cin ;
wire \add_9ns_9s_9_2_1_U11.top_add_9ns_9s_9_2_1_Adder_7_U.u2.cout ;
wire [4:0] \add_9ns_9s_9_2_1_U11.top_add_9ns_9s_9_2_1_Adder_7_U.u2.s ;
wire and_ln353_fu_486_p2;
wire [3:0] and_ln_fu_656_p3;
wire ap_CS_fsm_state1;
wire ap_CS_fsm_state10;
wire ap_CS_fsm_state11;
wire ap_CS_fsm_state12;
wire ap_CS_fsm_state13;
wire ap_CS_fsm_state14;
wire ap_CS_fsm_state15;
wire ap_CS_fsm_state16;
wire ap_CS_fsm_state17;
wire ap_CS_fsm_state18;
wire ap_CS_fsm_state19;
wire ap_CS_fsm_state20;
wire ap_CS_fsm_state21;
wire ap_CS_fsm_state22;
wire ap_CS_fsm_state23;
wire ap_CS_fsm_state24;
wire ap_CS_fsm_state25;
wire ap_CS_fsm_state26;
wire ap_CS_fsm_state27;
wire ap_CS_fsm_state28;
wire ap_CS_fsm_state29;
wire ap_CS_fsm_state30;
wire ap_CS_fsm_state31;
wire ap_CS_fsm_state32;
wire ap_CS_fsm_state33;
wire ap_CS_fsm_state34;
wire ap_CS_fsm_state35;
wire ap_CS_fsm_state36;
wire ap_CS_fsm_state37;
wire ap_CS_fsm_state38;
wire ap_CS_fsm_state39;
wire ap_CS_fsm_state40;
wire ap_CS_fsm_state41;
wire ap_CS_fsm_state42;
wire ap_CS_fsm_state43;
wire ap_CS_fsm_state44;
wire ap_CS_fsm_state45;
wire ap_CS_fsm_state46;
wire ap_CS_fsm_state47;
wire ap_CS_fsm_state48;
wire ap_CS_fsm_state49;
wire ap_CS_fsm_state7;
wire ap_CS_fsm_state8;
wire ap_CS_fsm_state9;
wire [48:0] ap_NS_fsm;
wire ap_clk;
wire ap_done;
wire ap_idle;
wire ap_ready;
wire ap_rst;
wire ap_start;
wire \ashr_32s_16ns_32_7_1_U8.ce ;
wire \ashr_32s_16ns_32_7_1_U8.clk ;
wire [31:0] \ashr_32s_16ns_32_7_1_U8.din0 ;
wire [31:0] \ashr_32s_16ns_32_7_1_U8.din1 ;
wire [15:0] \ashr_32s_16ns_32_7_1_U8.din1_cast ;
wire [15:0] \ashr_32s_16ns_32_7_1_U8.din1_mask ;
wire [31:0] \ashr_32s_16ns_32_7_1_U8.dout ;
wire \ashr_32s_16ns_32_7_1_U8.reset ;
wire [31:0] grp_fu_1025_p2;
wire [9:0] grp_fu_269_p2;
wire [1:0] grp_fu_303_p0;
wire [1:0] grp_fu_303_p2;
wire [6:0] grp_fu_313_p2;
wire [2:0] grp_fu_343_p0;
wire [2:0] grp_fu_343_p1;
wire [2:0] grp_fu_343_p2;
wire [10:0] grp_fu_387_p0;
wire [10:0] grp_fu_387_p1;
wire [10:0] grp_fu_387_p2;
wire [7:0] grp_fu_393_p1;
wire [7:0] grp_fu_393_p2;
wire [11:0] grp_fu_413_p0;
wire [11:0] grp_fu_413_p1;
wire [11:0] grp_fu_413_p2;
wire [31:0] grp_fu_448_p1;
wire [31:0] grp_fu_448_p2;
wire [31:0] grp_fu_461_p1;
wire [31:0] grp_fu_461_p2;
wire [1:0] grp_fu_467_p2;
wire [8:0] grp_fu_513_p0;
wire [8:0] grp_fu_513_p1;
wire [8:0] grp_fu_513_p2;
wire [5:0] grp_fu_558_p2;
wire [6:0] grp_fu_631_p0;
wire [6:0] grp_fu_631_p1;
wire [6:0] grp_fu_631_p2;
wire [17:0] grp_fu_686_p0;
wire [17:0] grp_fu_686_p1;
wire [17:0] grp_fu_686_p2;
wire [19:0] grp_fu_740_p0;
wire [19:0] grp_fu_740_p1;
wire [19:0] grp_fu_740_p2;
wire [18:0] grp_fu_764_p0;
wire [18:0] grp_fu_764_p2;
wire [18:0] grp_fu_804_p1;
wire [18:0] grp_fu_804_p2;
wire [1:0] grp_fu_809_p1;
wire [1:0] grp_fu_809_p2;
wire [18:0] grp_fu_817_p0;
wire [18:0] grp_fu_817_p2;
wire [36:0] grp_fu_837_p0;
wire [36:0] grp_fu_837_p1;
wire [36:0] grp_fu_837_p2;
wire [31:0] grp_fu_863_p2;
wire [56:0] grp_fu_902_p0;
wire [56:0] grp_fu_902_p1;
wire [56:0] grp_fu_902_p2;
wire [31:0] grp_fu_928_p2;
wire [34:0] grp_fu_967_p0;
wire [34:0] grp_fu_967_p1;
wire [34:0] grp_fu_967_p2;
wire [31:0] grp_fu_993_p2;
wire icmp_ln785_fu_645_p2;
wire icmp_ln786_1_fu_651_p2;
wire icmp_ln786_fu_673_p2;
wire icmp_ln850_fu_433_p2;
wire icmp_ln851_1_fu_523_p2;
wire icmp_ln851_2_fu_279_p2;
wire icmp_ln851_3_fu_746_p2;
wire icmp_ln851_4_fu_847_p2;
wire icmp_ln851_5_fu_912_p2;
wire icmp_ln851_6_fu_977_p2;
wire icmp_ln851_fu_308_p2;
wire [6:0] lhs_fu_497_p3;
wire \mul_8s_2s_10_7_1_U1.ce ;
wire \mul_8s_2s_10_7_1_U1.clk ;
wire [7:0] \mul_8s_2s_10_7_1_U1.din0 ;
wire [1:0] \mul_8s_2s_10_7_1_U1.din1 ;
wire [9:0] \mul_8s_2s_10_7_1_U1.dout ;
wire \mul_8s_2s_10_7_1_U1.reset ;
wire [7:0] \mul_8s_2s_10_7_1_U1.top_mul_8s_2s_10_7_1_Mul_DSP_0_U.a ;
wire [1:0] \mul_8s_2s_10_7_1_U1.top_mul_8s_2s_10_7_1_Mul_DSP_0_U.b ;
wire \mul_8s_2s_10_7_1_U1.top_mul_8s_2s_10_7_1_Mul_DSP_0_U.ce ;
wire \mul_8s_2s_10_7_1_U1.top_mul_8s_2s_10_7_1_Mul_DSP_0_U.clk ;
wire [9:0] \mul_8s_2s_10_7_1_U1.top_mul_8s_2s_10_7_1_Mul_DSP_0_U.p ;
wire [9:0] \mul_8s_2s_10_7_1_U1.top_mul_8s_2s_10_7_1_Mul_DSP_0_U.tmp_product ;
wire [3:0] op_0;
wire [1:0] op_1;
wire [15:0] op_11;
wire [3:0] op_12_V_fu_718_p3;
wire [3:0] op_14;
wire op_15;
wire [7:0] op_16;
wire [31:0] op_17;
wire [7:0] op_18;
wire op_19;
wire [7:0] op_3;
wire [31:0] op_30;
wire op_30_ap_vld;
wire [15:0] op_4;
wire [3:0] op_7;
wire [7:0] op_8_V_fu_356_p2;
wire [7:0] op_9;
wire or_ln384_fu_713_p2;
wire or_ln786_fu_697_p2;
wire [3:0] or_ln_fu_637_p4;
wire overflow_fu_668_p2;
wire p_Result_1_fu_563_p3;
wire p_Result_2_fu_479_p3;
wire p_Result_5_fu_529_p3;
wire p_Result_6_fu_770_p3;
wire p_Result_7_fu_868_p3;
wire p_Result_8_fu_933_p3;
wire p_Result_9_fu_998_p3;
wire p_Result_s_fu_318_p3;
wire [3:0] p_Val2_5_fu_692_p2;
wire [3:0] r_fu_596_p3;
wire [6:0] ret_V_18_fu_330_p3;
wire [5:0] ret_V_20_fu_575_p3;
wire ret_V_22_fu_491_p2;
wire [1:0] ret_V_24_fu_541_p3;
wire [18:0] ret_V_26_fu_782_p3;
wire [31:0] ret_V_30_fu_1010_p3;
wire [9:0] rhs_2_fu_376_p3;
wire [10:0] rhs_4_fu_402_p3;
wire [55:0] rhs_8_fu_891_p3;
wire [33:0] rhs_9_fu_956_p3;
wire [31:0] select_ln353_1_fu_945_p3;
wire [31:0] select_ln353_fu_880_p3;
wire [3:0] select_ln384_fu_706_p3;
wire [31:0] select_ln69_1_fu_1017_p3;
wire [1:0] select_ln69_fu_789_p3;
wire [5:0] select_ln850_1_fu_570_p3;
wire [1:0] select_ln850_3_fu_536_p3;
wire [18:0] select_ln850_4_fu_777_p3;
wire [31:0] select_ln850_6_fu_875_p3;
wire [31:0] select_ln850_7_fu_1005_p3;
wire [31:0] select_ln850_8_fu_940_p3;
wire [6:0] select_ln850_fu_325_p3;
wire [7:0] sext_ln1193_fu_373_p0;
wire [7:0] sext_ln1349_fu_349_p1;
wire [1:0] sext_ln215_fu_337_p0;
wire [3:0] sext_ln546_1_fu_593_p1;
wire [15:0] sext_ln546_2_fu_454_p1;
wire [15:0] sext_ln546_fu_441_p1;
wire [7:0] sext_ln703_1_fu_399_p0;
wire [7:0] sext_ln703_2_fu_822_p0;
wire [31:0] sext_ln703_3_fu_887_p0;
wire [7:0] sext_ln703_4_fu_952_p0;
wire [7:0] sext_ln703_fu_509_p0;
wire [31:0] sext_ln781_fu_438_p1;
wire [18:0] sext_ln850_fu_761_p1;
wire \shl_32s_16ns_32_7_1_U9.ce ;
wire \shl_32s_16ns_32_7_1_U9.clk ;
wire [31:0] \shl_32s_16ns_32_7_1_U9.din0 ;
wire [31:0] \shl_32s_16ns_32_7_1_U9.din1 ;
wire [15:0] \shl_32s_16ns_32_7_1_U9.din1_cast ;
wire [15:0] \shl_32s_16ns_32_7_1_U9.din1_mask ;
wire [31:0] \shl_32s_16ns_32_7_1_U9.dout ;
wire \shl_32s_16ns_32_7_1_U9.reset ;
wire \sub_11s_11s_11_2_1_U5.ce ;
wire \sub_11s_11s_11_2_1_U5.clk ;
wire [10:0] \sub_11s_11s_11_2_1_U5.din0 ;
wire [10:0] \sub_11s_11s_11_2_1_U5.din1 ;
wire [10:0] \sub_11s_11s_11_2_1_U5.dout ;
wire \sub_11s_11s_11_2_1_U5.reset ;
wire [10:0] \sub_11s_11s_11_2_1_U5.top_sub_11s_11s_11_2_1_Adder_3_U.a ;
wire [10:0] \sub_11s_11s_11_2_1_U5.top_sub_11s_11s_11_2_1_Adder_3_U.ain_s0 ;
wire [10:0] \sub_11s_11s_11_2_1_U5.top_sub_11s_11s_11_2_1_Adder_3_U.b ;
wire [10:0] \sub_11s_11s_11_2_1_U5.top_sub_11s_11s_11_2_1_Adder_3_U.bin_s0 ;
wire \sub_11s_11s_11_2_1_U5.top_sub_11s_11s_11_2_1_Adder_3_U.ce ;
wire \sub_11s_11s_11_2_1_U5.top_sub_11s_11s_11_2_1_Adder_3_U.clk ;
wire \sub_11s_11s_11_2_1_U5.top_sub_11s_11s_11_2_1_Adder_3_U.facout_s1 ;
wire \sub_11s_11s_11_2_1_U5.top_sub_11s_11s_11_2_1_Adder_3_U.facout_s2 ;
wire [4:0] \sub_11s_11s_11_2_1_U5.top_sub_11s_11s_11_2_1_Adder_3_U.fas_s1 ;
wire [5:0] \sub_11s_11s_11_2_1_U5.top_sub_11s_11s_11_2_1_Adder_3_U.fas_s2 ;
wire \sub_11s_11s_11_2_1_U5.top_sub_11s_11s_11_2_1_Adder_3_U.reset ;
wire [10:0] \sub_11s_11s_11_2_1_U5.top_sub_11s_11s_11_2_1_Adder_3_U.s ;
wire [4:0] \sub_11s_11s_11_2_1_U5.top_sub_11s_11s_11_2_1_Adder_3_U.u1.a ;
wire [4:0] \sub_11s_11s_11_2_1_U5.top_sub_11s_11s_11_2_1_Adder_3_U.u1.b ;
wire \sub_11s_11s_11_2_1_U5.top_sub_11s_11s_11_2_1_Adder_3_U.u1.cin ;
wire \sub_11s_11s_11_2_1_U5.top_sub_11s_11s_11_2_1_Adder_3_U.u1.cout ;
wire [4:0] \sub_11s_11s_11_2_1_U5.top_sub_11s_11s_11_2_1_Adder_3_U.u1.s ;
wire [5:0] \sub_11s_11s_11_2_1_U5.top_sub_11s_11s_11_2_1_Adder_3_U.u2.a ;
wire [5:0] \sub_11s_11s_11_2_1_U5.top_sub_11s_11s_11_2_1_Adder_3_U.u2.b ;
wire \sub_11s_11s_11_2_1_U5.top_sub_11s_11s_11_2_1_Adder_3_U.u2.cin ;
wire \sub_11s_11s_11_2_1_U5.top_sub_11s_11s_11_2_1_Adder_3_U.u2.cout ;
wire [5:0] \sub_11s_11s_11_2_1_U5.top_sub_11s_11s_11_2_1_Adder_3_U.u2.s ;
wire \sub_8ns_8s_8_2_1_U6.ce ;
wire \sub_8ns_8s_8_2_1_U6.clk ;
wire [7:0] \sub_8ns_8s_8_2_1_U6.din0 ;
wire [7:0] \sub_8ns_8s_8_2_1_U6.din1 ;
wire [7:0] \sub_8ns_8s_8_2_1_U6.dout ;
wire \sub_8ns_8s_8_2_1_U6.reset ;
wire [7:0] \sub_8ns_8s_8_2_1_U6.top_sub_8ns_8s_8_2_1_Adder_4_U.a ;
wire [7:0] \sub_8ns_8s_8_2_1_U6.top_sub_8ns_8s_8_2_1_Adder_4_U.ain_s0 ;
wire [7:0] \sub_8ns_8s_8_2_1_U6.top_sub_8ns_8s_8_2_1_Adder_4_U.b ;
wire [7:0] \sub_8ns_8s_8_2_1_U6.top_sub_8ns_8s_8_2_1_Adder_4_U.bin_s0 ;
wire \sub_8ns_8s_8_2_1_U6.top_sub_8ns_8s_8_2_1_Adder_4_U.ce ;
wire \sub_8ns_8s_8_2_1_U6.top_sub_8ns_8s_8_2_1_Adder_4_U.clk ;
wire \sub_8ns_8s_8_2_1_U6.top_sub_8ns_8s_8_2_1_Adder_4_U.facout_s1 ;
wire \sub_8ns_8s_8_2_1_U6.top_sub_8ns_8s_8_2_1_Adder_4_U.facout_s2 ;
wire [3:0] \sub_8ns_8s_8_2_1_U6.top_sub_8ns_8s_8_2_1_Adder_4_U.fas_s1 ;
wire [3:0] \sub_8ns_8s_8_2_1_U6.top_sub_8ns_8s_8_2_1_Adder_4_U.fas_s2 ;
wire \sub_8ns_8s_8_2_1_U6.top_sub_8ns_8s_8_2_1_Adder_4_U.reset ;
wire [7:0] \sub_8ns_8s_8_2_1_U6.top_sub_8ns_8s_8_2_1_Adder_4_U.s ;
wire [3:0] \sub_8ns_8s_8_2_1_U6.top_sub_8ns_8s_8_2_1_Adder_4_U.u1.a ;
wire [3:0] \sub_8ns_8s_8_2_1_U6.top_sub_8ns_8s_8_2_1_Adder_4_U.u1.b ;
wire \sub_8ns_8s_8_2_1_U6.top_sub_8ns_8s_8_2_1_Adder_4_U.u1.cin ;
wire \sub_8ns_8s_8_2_1_U6.top_sub_8ns_8s_8_2_1_Adder_4_U.u1.cout ;
wire [3:0] \sub_8ns_8s_8_2_1_U6.top_sub_8ns_8s_8_2_1_Adder_4_U.u1.s ;
wire [3:0] \sub_8ns_8s_8_2_1_U6.top_sub_8ns_8s_8_2_1_Adder_4_U.u2.a ;
wire [3:0] \sub_8ns_8s_8_2_1_U6.top_sub_8ns_8s_8_2_1_Adder_4_U.u2.b ;
wire \sub_8ns_8s_8_2_1_U6.top_sub_8ns_8s_8_2_1_Adder_4_U.u2.cin ;
wire \sub_8ns_8s_8_2_1_U6.top_sub_8ns_8s_8_2_1_Adder_4_U.u2.cout ;
wire [3:0] \sub_8ns_8s_8_2_1_U6.top_sub_8ns_8s_8_2_1_Adder_4_U.u2.s ;
wire [22:0] tmp_8_fu_826_p3;
wire tmp_fu_472_p3;
wire [7:0] trunc_ln1349_fu_352_p1;
wire [2:0] trunc_ln546_fu_582_p1;
wire [3:0] trunc_ln769_fu_586_p1;
wire [7:0] trunc_ln851_1_fu_519_p0;
wire [2:0] trunc_ln851_1_fu_519_p1;
wire [2:0] trunc_ln851_2_fu_419_p1;
wire [7:0] trunc_ln851_3_fu_275_p0;
wire [2:0] trunc_ln851_3_fu_275_p1;
wire [1:0] trunc_ln851_4_fu_726_p1;
wire [7:0] trunc_ln851_5_fu_843_p0;
wire [3:0] trunc_ln851_5_fu_843_p1;
wire [31:0] trunc_ln851_6_fu_908_p0;
wire [23:0] trunc_ln851_6_fu_908_p1;
wire [7:0] trunc_ln851_7_fu_973_p0;
wire [1:0] trunc_ln851_7_fu_973_p1;
wire [2:0] trunc_ln851_fu_295_p1;
wire underflow_fu_701_p2;
wire xor_ln785_fu_663_p2;


assign _067_ = icmp_ln851_4_reg_1434 & ap_CS_fsm[35];
assign _068_ = icmp_ln851_5_reg_1471 & ap_CS_fsm[40];
assign _069_ = icmp_ln851_6_reg_1508 & ap_CS_fsm[45];
assign _070_ = icmp_ln851_3_reg_1357 & ap_CS_fsm[26];
assign _071_ = _078_ & ap_CS_fsm[13];
assign _072_ = _079_ & ap_CS_fsm[17];
assign _073_ = ap_CS_fsm[11] & p_Result_10_reg_1117;
assign _074_ = ap_CS_fsm[18] & p_Result_10_reg_1117;
assign _075_ = ap_CS_fsm[18] & _080_;
assign _076_ = _081_ & ap_CS_fsm[0];
assign _077_ = ap_start & ap_CS_fsm[0];
assign and_ln353_fu_486_p2 = ret_V_21_reg_1152[10] & icmp_ln850_reg_1180;
assign overflow_fu_668_p2 = xor_ln785_fu_663_p2 & icmp_ln785_reg_1296;
assign underflow_fu_701_p2 = p_Result_11_reg_1273 & or_ln786_fu_697_p2;
assign xor_ln785_fu_663_p2 = ~ p_Result_11_reg_1273;
assign _078_ = ~ icmp_ln851_2_reg_1052;
assign _079_ = ~ icmp_ln851_1_reg_1221;
assign _080_ = ~ p_Result_10_reg_1117;
assign _081_ = ~ ap_start;
assign _082_ = ! { tmp_5_reg_1279, 3'h0 };
assign _083_ = ! op_9[2:0];
assign _084_ = ! op_3[2:0];
assign _085_ = ! trunc_ln851_reg_1069;
always @(posedge \add_12s_12s_12_2_1_U7.top_add_12s_12s_12_2_1_Adder_5_U.clk )
\add_12s_12s_12_2_1_U7.top_add_12s_12s_12_2_1_Adder_5_U.bin_s1  <= _087_;
always @(posedge \add_12s_12s_12_2_1_U7.top_add_12s_12s_12_2_1_Adder_5_U.clk )
\add_12s_12s_12_2_1_U7.top_add_12s_12s_12_2_1_Adder_5_U.ain_s1  <= _086_;
always @(posedge \add_12s_12s_12_2_1_U7.top_add_12s_12s_12_2_1_Adder_5_U.clk )
\add_12s_12s_12_2_1_U7.top_add_12s_12s_12_2_1_Adder_5_U.sum_s1  <= _089_;
always @(posedge \add_12s_12s_12_2_1_U7.top_add_12s_12s_12_2_1_Adder_5_U.clk )
\add_12s_12s_12_2_1_U7.top_add_12s_12s_12_2_1_Adder_5_U.carry_s1  <= _088_;
assign _087_ = \add_12s_12s_12_2_1_U7.top_add_12s_12s_12_2_1_Adder_5_U.ce  ? \add_12s_12s_12_2_1_U7.top_add_12s_12s_12_2_1_Adder_5_U.b [11:6] : \add_12s_12s_12_2_1_U7.top_add_12s_12s_12_2_1_Adder_5_U.bin_s1 ;
assign _086_ = \add_12s_12s_12_2_1_U7.top_add_12s_12s_12_2_1_Adder_5_U.ce  ? \add_12s_12s_12_2_1_U7.top_add_12s_12s_12_2_1_Adder_5_U.a [11:6] : \add_12s_12s_12_2_1_U7.top_add_12s_12s_12_2_1_Adder_5_U.ain_s1 ;
assign _088_ = \add_12s_12s_12_2_1_U7.top_add_12s_12s_12_2_1_Adder_5_U.ce  ? \add_12s_12s_12_2_1_U7.top_add_12s_12s_12_2_1_Adder_5_U.facout_s1  : \add_12s_12s_12_2_1_U7.top_add_12s_12s_12_2_1_Adder_5_U.carry_s1 ;
assign _089_ = \add_12s_12s_12_2_1_U7.top_add_12s_12s_12_2_1_Adder_5_U.ce  ? \add_12s_12s_12_2_1_U7.top_add_12s_12s_12_2_1_Adder_5_U.fas_s1  : \add_12s_12s_12_2_1_U7.top_add_12s_12s_12_2_1_Adder_5_U.sum_s1 ;
assign _090_ = \add_12s_12s_12_2_1_U7.top_add_12s_12s_12_2_1_Adder_5_U.u1.a  + \add_12s_12s_12_2_1_U7.top_add_12s_12s_12_2_1_Adder_5_U.u1.b ;
assign { \add_12s_12s_12_2_1_U7.top_add_12s_12s_12_2_1_Adder_5_U.u1.cout , \add_12s_12s_12_2_1_U7.top_add_12s_12s_12_2_1_Adder_5_U.u1.s  } = _090_ + \add_12s_12s_12_2_1_U7.top_add_12s_12s_12_2_1_Adder_5_U.u1.cin ;
assign _091_ = \add_12s_12s_12_2_1_U7.top_add_12s_12s_12_2_1_Adder_5_U.u2.a  + \add_12s_12s_12_2_1_U7.top_add_12s_12s_12_2_1_Adder_5_U.u2.b ;
assign { \add_12s_12s_12_2_1_U7.top_add_12s_12s_12_2_1_Adder_5_U.u2.cout , \add_12s_12s_12_2_1_U7.top_add_12s_12s_12_2_1_Adder_5_U.u2.s  } = _091_ + \add_12s_12s_12_2_1_U7.top_add_12s_12s_12_2_1_Adder_5_U.u2.cin ;
always @(posedge \add_18s_18ns_18_2_1_U14.top_add_18s_18ns_18_2_1_Adder_10_U.clk )
\add_18s_18ns_18_2_1_U14.top_add_18s_18ns_18_2_1_Adder_10_U.bin_s1  <= _093_;
always @(posedge \add_18s_18ns_18_2_1_U14.top_add_18s_18ns_18_2_1_Adder_10_U.clk )
\add_18s_18ns_18_2_1_U14.top_add_18s_18ns_18_2_1_Adder_10_U.ain_s1  <= _092_;
always @(posedge \add_18s_18ns_18_2_1_U14.top_add_18s_18ns_18_2_1_Adder_10_U.clk )
\add_18s_18ns_18_2_1_U14.top_add_18s_18ns_18_2_1_Adder_10_U.sum_s1  <= _095_;
always @(posedge \add_18s_18ns_18_2_1_U14.top_add_18s_18ns_18_2_1_Adder_10_U.clk )
\add_18s_18ns_18_2_1_U14.top_add_18s_18ns_18_2_1_Adder_10_U.carry_s1  <= _094_;
assign _093_ = \add_18s_18ns_18_2_1_U14.top_add_18s_18ns_18_2_1_Adder_10_U.ce  ? \add_18s_18ns_18_2_1_U14.top_add_18s_18ns_18_2_1_Adder_10_U.b [17:9] : \add_18s_18ns_18_2_1_U14.top_add_18s_18ns_18_2_1_Adder_10_U.bin_s1 ;
assign _092_ = \add_18s_18ns_18_2_1_U14.top_add_18s_18ns_18_2_1_Adder_10_U.ce  ? \add_18s_18ns_18_2_1_U14.top_add_18s_18ns_18_2_1_Adder_10_U.a [17:9] : \add_18s_18ns_18_2_1_U14.top_add_18s_18ns_18_2_1_Adder_10_U.ain_s1 ;
assign _094_ = \add_18s_18ns_18_2_1_U14.top_add_18s_18ns_18_2_1_Adder_10_U.ce  ? \add_18s_18ns_18_2_1_U14.top_add_18s_18ns_18_2_1_Adder_10_U.facout_s1  : \add_18s_18ns_18_2_1_U14.top_add_18s_18ns_18_2_1_Adder_10_U.carry_s1 ;
assign _095_ = \add_18s_18ns_18_2_1_U14.top_add_18s_18ns_18_2_1_Adder_10_U.ce  ? \add_18s_18ns_18_2_1_U14.top_add_18s_18ns_18_2_1_Adder_10_U.fas_s1  : \add_18s_18ns_18_2_1_U14.top_add_18s_18ns_18_2_1_Adder_10_U.sum_s1 ;
assign _096_ = \add_18s_18ns_18_2_1_U14.top_add_18s_18ns_18_2_1_Adder_10_U.u1.a  + \add_18s_18ns_18_2_1_U14.top_add_18s_18ns_18_2_1_Adder_10_U.u1.b ;
assign { \add_18s_18ns_18_2_1_U14.top_add_18s_18ns_18_2_1_Adder_10_U.u1.cout , \add_18s_18ns_18_2_1_U14.top_add_18s_18ns_18_2_1_Adder_10_U.u1.s  } = _096_ + \add_18s_18ns_18_2_1_U14.top_add_18s_18ns_18_2_1_Adder_10_U.u1.cin ;
assign _097_ = \add_18s_18ns_18_2_1_U14.top_add_18s_18ns_18_2_1_Adder_10_U.u2.a  + \add_18s_18ns_18_2_1_U14.top_add_18s_18ns_18_2_1_Adder_10_U.u2.b ;
assign { \add_18s_18ns_18_2_1_U14.top_add_18s_18ns_18_2_1_Adder_10_U.u2.cout , \add_18s_18ns_18_2_1_U14.top_add_18s_18ns_18_2_1_Adder_10_U.u2.s  } = _097_ + \add_18s_18ns_18_2_1_U14.top_add_18s_18ns_18_2_1_Adder_10_U.u2.cin ;
always @(posedge \add_19ns_19s_19_2_1_U17.top_add_19ns_19s_19_2_1_Adder_13_U.clk )
\add_19ns_19s_19_2_1_U17.top_add_19ns_19s_19_2_1_Adder_13_U.bin_s1  <= _099_;
always @(posedge \add_19ns_19s_19_2_1_U17.top_add_19ns_19s_19_2_1_Adder_13_U.clk )
\add_19ns_19s_19_2_1_U17.top_add_19ns_19s_19_2_1_Adder_13_U.ain_s1  <= _098_;
always @(posedge \add_19ns_19s_19_2_1_U17.top_add_19ns_19s_19_2_1_Adder_13_U.clk )
\add_19ns_19s_19_2_1_U17.top_add_19ns_19s_19_2_1_Adder_13_U.sum_s1  <= _101_;
always @(posedge \add_19ns_19s_19_2_1_U17.top_add_19ns_19s_19_2_1_Adder_13_U.clk )
\add_19ns_19s_19_2_1_U17.top_add_19ns_19s_19_2_1_Adder_13_U.carry_s1  <= _100_;
assign _099_ = \add_19ns_19s_19_2_1_U17.top_add_19ns_19s_19_2_1_Adder_13_U.ce  ? \add_19ns_19s_19_2_1_U17.top_add_19ns_19s_19_2_1_Adder_13_U.b [18:9] : \add_19ns_19s_19_2_1_U17.top_add_19ns_19s_19_2_1_Adder_13_U.bin_s1 ;
assign _098_ = \add_19ns_19s_19_2_1_U17.top_add_19ns_19s_19_2_1_Adder_13_U.ce  ? \add_19ns_19s_19_2_1_U17.top_add_19ns_19s_19_2_1_Adder_13_U.a [18:9] : \add_19ns_19s_19_2_1_U17.top_add_19ns_19s_19_2_1_Adder_13_U.ain_s1 ;
assign _100_ = \add_19ns_19s_19_2_1_U17.top_add_19ns_19s_19_2_1_Adder_13_U.ce  ? \add_19ns_19s_19_2_1_U17.top_add_19ns_19s_19_2_1_Adder_13_U.facout_s1  : \add_19ns_19s_19_2_1_U17.top_add_19ns_19s_19_2_1_Adder_13_U.carry_s1 ;
assign _101_ = \add_19ns_19s_19_2_1_U17.top_add_19ns_19s_19_2_1_Adder_13_U.ce  ? \add_19ns_19s_19_2_1_U17.top_add_19ns_19s_19_2_1_Adder_13_U.fas_s1  : \add_19ns_19s_19_2_1_U17.top_add_19ns_19s_19_2_1_Adder_13_U.sum_s1 ;
assign _102_ = \add_19ns_19s_19_2_1_U17.top_add_19ns_19s_19_2_1_Adder_13_U.u1.a  + \add_19ns_19s_19_2_1_U17.top_add_19ns_19s_19_2_1_Adder_13_U.u1.b ;
assign { \add_19ns_19s_19_2_1_U17.top_add_19ns_19s_19_2_1_Adder_13_U.u1.cout , \add_19ns_19s_19_2_1_U17.top_add_19ns_19s_19_2_1_Adder_13_U.u1.s  } = _102_ + \add_19ns_19s_19_2_1_U17.top_add_19ns_19s_19_2_1_Adder_13_U.u1.cin ;
assign _103_ = \add_19ns_19s_19_2_1_U17.top_add_19ns_19s_19_2_1_Adder_13_U.u2.a  + \add_19ns_19s_19_2_1_U17.top_add_19ns_19s_19_2_1_Adder_13_U.u2.b ;
assign { \add_19ns_19s_19_2_1_U17.top_add_19ns_19s_19_2_1_Adder_13_U.u2.cout , \add_19ns_19s_19_2_1_U17.top_add_19ns_19s_19_2_1_Adder_13_U.u2.s  } = _103_ + \add_19ns_19s_19_2_1_U17.top_add_19ns_19s_19_2_1_Adder_13_U.u2.cin ;
always @(posedge \add_19s_19ns_19_2_1_U16.top_add_19s_19ns_19_2_1_Adder_12_U.clk )
\add_19s_19ns_19_2_1_U16.top_add_19s_19ns_19_2_1_Adder_12_U.bin_s1  <= _105_;
always @(posedge \add_19s_19ns_19_2_1_U16.top_add_19s_19ns_19_2_1_Adder_12_U.clk )
\add_19s_19ns_19_2_1_U16.top_add_19s_19ns_19_2_1_Adder_12_U.ain_s1  <= _104_;
always @(posedge \add_19s_19ns_19_2_1_U16.top_add_19s_19ns_19_2_1_Adder_12_U.clk )
\add_19s_19ns_19_2_1_U16.top_add_19s_19ns_19_2_1_Adder_12_U.sum_s1  <= _107_;
always @(posedge \add_19s_19ns_19_2_1_U16.top_add_19s_19ns_19_2_1_Adder_12_U.clk )
\add_19s_19ns_19_2_1_U16.top_add_19s_19ns_19_2_1_Adder_12_U.carry_s1  <= _106_;
assign _105_ = \add_19s_19ns_19_2_1_U16.top_add_19s_19ns_19_2_1_Adder_12_U.ce  ? \add_19s_19ns_19_2_1_U16.top_add_19s_19ns_19_2_1_Adder_12_U.b [18:9] : \add_19s_19ns_19_2_1_U16.top_add_19s_19ns_19_2_1_Adder_12_U.bin_s1 ;
assign _104_ = \add_19s_19ns_19_2_1_U16.top_add_19s_19ns_19_2_1_Adder_12_U.ce  ? \add_19s_19ns_19_2_1_U16.top_add_19s_19ns_19_2_1_Adder_12_U.a [18:9] : \add_19s_19ns_19_2_1_U16.top_add_19s_19ns_19_2_1_Adder_12_U.ain_s1 ;
assign _106_ = \add_19s_19ns_19_2_1_U16.top_add_19s_19ns_19_2_1_Adder_12_U.ce  ? \add_19s_19ns_19_2_1_U16.top_add_19s_19ns_19_2_1_Adder_12_U.facout_s1  : \add_19s_19ns_19_2_1_U16.top_add_19s_19ns_19_2_1_Adder_12_U.carry_s1 ;
assign _107_ = \add_19s_19ns_19_2_1_U16.top_add_19s_19ns_19_2_1_Adder_12_U.ce  ? \add_19s_19ns_19_2_1_U16.top_add_19s_19ns_19_2_1_Adder_12_U.fas_s1  : \add_19s_19ns_19_2_1_U16.top_add_19s_19ns_19_2_1_Adder_12_U.sum_s1 ;
assign _108_ = \add_19s_19ns_19_2_1_U16.top_add_19s_19ns_19_2_1_Adder_12_U.u1.a  + \add_19s_19ns_19_2_1_U16.top_add_19s_19ns_19_2_1_Adder_12_U.u1.b ;
assign { \add_19s_19ns_19_2_1_U16.top_add_19s_19ns_19_2_1_Adder_12_U.u1.cout , \add_19s_19ns_19_2_1_U16.top_add_19s_19ns_19_2_1_Adder_12_U.u1.s  } = _108_ + \add_19s_19ns_19_2_1_U16.top_add_19s_19ns_19_2_1_Adder_12_U.u1.cin ;
assign _109_ = \add_19s_19ns_19_2_1_U16.top_add_19s_19ns_19_2_1_Adder_12_U.u2.a  + \add_19s_19ns_19_2_1_U16.top_add_19s_19ns_19_2_1_Adder_12_U.u2.b ;
assign { \add_19s_19ns_19_2_1_U16.top_add_19s_19ns_19_2_1_Adder_12_U.u2.cout , \add_19s_19ns_19_2_1_U16.top_add_19s_19ns_19_2_1_Adder_12_U.u2.s  } = _109_ + \add_19s_19ns_19_2_1_U16.top_add_19s_19ns_19_2_1_Adder_12_U.u2.cin ;
always @(posedge \add_19s_19ns_19_2_1_U19.top_add_19s_19ns_19_2_1_Adder_12_U.clk )
\add_19s_19ns_19_2_1_U19.top_add_19s_19ns_19_2_1_Adder_12_U.bin_s1  <= _111_;
always @(posedge \add_19s_19ns_19_2_1_U19.top_add_19s_19ns_19_2_1_Adder_12_U.clk )
\add_19s_19ns_19_2_1_U19.top_add_19s_19ns_19_2_1_Adder_12_U.ain_s1  <= _110_;
always @(posedge \add_19s_19ns_19_2_1_U19.top_add_19s_19ns_19_2_1_Adder_12_U.clk )
\add_19s_19ns_19_2_1_U19.top_add_19s_19ns_19_2_1_Adder_12_U.sum_s1  <= _113_;
always @(posedge \add_19s_19ns_19_2_1_U19.top_add_19s_19ns_19_2_1_Adder_12_U.clk )
\add_19s_19ns_19_2_1_U19.top_add_19s_19ns_19_2_1_Adder_12_U.carry_s1  <= _112_;
assign _111_ = \add_19s_19ns_19_2_1_U19.top_add_19s_19ns_19_2_1_Adder_12_U.ce  ? \add_19s_19ns_19_2_1_U19.top_add_19s_19ns_19_2_1_Adder_12_U.b [18:9] : \add_19s_19ns_19_2_1_U19.top_add_19s_19ns_19_2_1_Adder_12_U.bin_s1 ;
assign _110_ = \add_19s_19ns_19_2_1_U19.top_add_19s_19ns_19_2_1_Adder_12_U.ce  ? \add_19s_19ns_19_2_1_U19.top_add_19s_19ns_19_2_1_Adder_12_U.a [18:9] : \add_19s_19ns_19_2_1_U19.top_add_19s_19ns_19_2_1_Adder_12_U.ain_s1 ;
assign _112_ = \add_19s_19ns_19_2_1_U19.top_add_19s_19ns_19_2_1_Adder_12_U.ce  ? \add_19s_19ns_19_2_1_U19.top_add_19s_19ns_19_2_1_Adder_12_U.facout_s1  : \add_19s_19ns_19_2_1_U19.top_add_19s_19ns_19_2_1_Adder_12_U.carry_s1 ;
assign _113_ = \add_19s_19ns_19_2_1_U19.top_add_19s_19ns_19_2_1_Adder_12_U.ce  ? \add_19s_19ns_19_2_1_U19.top_add_19s_19ns_19_2_1_Adder_12_U.fas_s1  : \add_19s_19ns_19_2_1_U19.top_add_19s_19ns_19_2_1_Adder_12_U.sum_s1 ;
assign _114_ = \add_19s_19ns_19_2_1_U19.top_add_19s_19ns_19_2_1_Adder_12_U.u1.a  + \add_19s_19ns_19_2_1_U19.top_add_19s_19ns_19_2_1_Adder_12_U.u1.b ;
assign { \add_19s_19ns_19_2_1_U19.top_add_19s_19ns_19_2_1_Adder_12_U.u1.cout , \add_19s_19ns_19_2_1_U19.top_add_19s_19ns_19_2_1_Adder_12_U.u1.s  } = _114_ + \add_19s_19ns_19_2_1_U19.top_add_19s_19ns_19_2_1_Adder_12_U.u1.cin ;
assign _115_ = \add_19s_19ns_19_2_1_U19.top_add_19s_19ns_19_2_1_Adder_12_U.u2.a  + \add_19s_19ns_19_2_1_U19.top_add_19s_19ns_19_2_1_Adder_12_U.u2.b ;
assign { \add_19s_19ns_19_2_1_U19.top_add_19s_19ns_19_2_1_Adder_12_U.u2.cout , \add_19s_19ns_19_2_1_U19.top_add_19s_19ns_19_2_1_Adder_12_U.u2.s  } = _115_ + \add_19s_19ns_19_2_1_U19.top_add_19s_19ns_19_2_1_Adder_12_U.u2.cin ;
always @(posedge \add_20ns_20s_20_2_1_U15.top_add_20ns_20s_20_2_1_Adder_11_U.clk )
\add_20ns_20s_20_2_1_U15.top_add_20ns_20s_20_2_1_Adder_11_U.bin_s1  <= _117_;
always @(posedge \add_20ns_20s_20_2_1_U15.top_add_20ns_20s_20_2_1_Adder_11_U.clk )
\add_20ns_20s_20_2_1_U15.top_add_20ns_20s_20_2_1_Adder_11_U.ain_s1  <= _116_;
always @(posedge \add_20ns_20s_20_2_1_U15.top_add_20ns_20s_20_2_1_Adder_11_U.clk )
\add_20ns_20s_20_2_1_U15.top_add_20ns_20s_20_2_1_Adder_11_U.sum_s1  <= _119_;
always @(posedge \add_20ns_20s_20_2_1_U15.top_add_20ns_20s_20_2_1_Adder_11_U.clk )
\add_20ns_20s_20_2_1_U15.top_add_20ns_20s_20_2_1_Adder_11_U.carry_s1  <= _118_;
assign _117_ = \add_20ns_20s_20_2_1_U15.top_add_20ns_20s_20_2_1_Adder_11_U.ce  ? \add_20ns_20s_20_2_1_U15.top_add_20ns_20s_20_2_1_Adder_11_U.b [19:10] : \add_20ns_20s_20_2_1_U15.top_add_20ns_20s_20_2_1_Adder_11_U.bin_s1 ;
assign _116_ = \add_20ns_20s_20_2_1_U15.top_add_20ns_20s_20_2_1_Adder_11_U.ce  ? \add_20ns_20s_20_2_1_U15.top_add_20ns_20s_20_2_1_Adder_11_U.a [19:10] : \add_20ns_20s_20_2_1_U15.top_add_20ns_20s_20_2_1_Adder_11_U.ain_s1 ;
assign _118_ = \add_20ns_20s_20_2_1_U15.top_add_20ns_20s_20_2_1_Adder_11_U.ce  ? \add_20ns_20s_20_2_1_U15.top_add_20ns_20s_20_2_1_Adder_11_U.facout_s1  : \add_20ns_20s_20_2_1_U15.top_add_20ns_20s_20_2_1_Adder_11_U.carry_s1 ;
assign _119_ = \add_20ns_20s_20_2_1_U15.top_add_20ns_20s_20_2_1_Adder_11_U.ce  ? \add_20ns_20s_20_2_1_U15.top_add_20ns_20s_20_2_1_Adder_11_U.fas_s1  : \add_20ns_20s_20_2_1_U15.top_add_20ns_20s_20_2_1_Adder_11_U.sum_s1 ;
assign _120_ = \add_20ns_20s_20_2_1_U15.top_add_20ns_20s_20_2_1_Adder_11_U.u1.a  + \add_20ns_20s_20_2_1_U15.top_add_20ns_20s_20_2_1_Adder_11_U.u1.b ;
assign { \add_20ns_20s_20_2_1_U15.top_add_20ns_20s_20_2_1_Adder_11_U.u1.cout , \add_20ns_20s_20_2_1_U15.top_add_20ns_20s_20_2_1_Adder_11_U.u1.s  } = _120_ + \add_20ns_20s_20_2_1_U15.top_add_20ns_20s_20_2_1_Adder_11_U.u1.cin ;
assign _121_ = \add_20ns_20s_20_2_1_U15.top_add_20ns_20s_20_2_1_Adder_11_U.u2.a  + \add_20ns_20s_20_2_1_U15.top_add_20ns_20s_20_2_1_Adder_11_U.u2.b ;
assign { \add_20ns_20s_20_2_1_U15.top_add_20ns_20s_20_2_1_Adder_11_U.u2.cout , \add_20ns_20s_20_2_1_U15.top_add_20ns_20s_20_2_1_Adder_11_U.u2.s  } = _121_ + \add_20ns_20s_20_2_1_U15.top_add_20ns_20s_20_2_1_Adder_11_U.u2.cin ;
always @(posedge \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_6_U.clk )
\add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_6_U.bin_s1  <= _123_;
always @(posedge \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_6_U.clk )
\add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_6_U.ain_s1  <= _122_;
always @(posedge \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_6_U.clk )
\add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_6_U.sum_s1  <= _125_;
always @(posedge \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_6_U.clk )
\add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_6_U.carry_s1  <= _124_;
assign _123_ = \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_6_U.ce  ? \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_6_U.b [1] : \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_6_U.bin_s1 ;
assign _122_ = \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_6_U.ce  ? \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_6_U.a [1] : \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_6_U.ain_s1 ;
assign _124_ = \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_6_U.ce  ? \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_6_U.facout_s1  : \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_6_U.carry_s1 ;
assign _125_ = \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_6_U.ce  ? \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_6_U.fas_s1  : \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_6_U.sum_s1 ;
assign _126_ = \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_6_U.u1.a  + \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_6_U.u1.b ;
assign { \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_6_U.u1.cout , \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_6_U.u1.s  } = _126_ + \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_6_U.u1.cin ;
assign _127_ = \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_6_U.u2.a  + \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_6_U.u2.b ;
assign { \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_6_U.u2.cout , \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_6_U.u2.s  } = _127_ + \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_6_U.u2.cin ;
always @(posedge \add_2ns_2ns_2_2_1_U18.top_add_2ns_2ns_2_2_1_Adder_6_U.clk )
\add_2ns_2ns_2_2_1_U18.top_add_2ns_2ns_2_2_1_Adder_6_U.bin_s1  <= _129_;
always @(posedge \add_2ns_2ns_2_2_1_U18.top_add_2ns_2ns_2_2_1_Adder_6_U.clk )
\add_2ns_2ns_2_2_1_U18.top_add_2ns_2ns_2_2_1_Adder_6_U.ain_s1  <= _128_;
always @(posedge \add_2ns_2ns_2_2_1_U18.top_add_2ns_2ns_2_2_1_Adder_6_U.clk )
\add_2ns_2ns_2_2_1_U18.top_add_2ns_2ns_2_2_1_Adder_6_U.sum_s1  <= _131_;
always @(posedge \add_2ns_2ns_2_2_1_U18.top_add_2ns_2ns_2_2_1_Adder_6_U.clk )
\add_2ns_2ns_2_2_1_U18.top_add_2ns_2ns_2_2_1_Adder_6_U.carry_s1  <= _130_;
assign _129_ = \add_2ns_2ns_2_2_1_U18.top_add_2ns_2ns_2_2_1_Adder_6_U.ce  ? \add_2ns_2ns_2_2_1_U18.top_add_2ns_2ns_2_2_1_Adder_6_U.b [1] : \add_2ns_2ns_2_2_1_U18.top_add_2ns_2ns_2_2_1_Adder_6_U.bin_s1 ;
assign _128_ = \add_2ns_2ns_2_2_1_U18.top_add_2ns_2ns_2_2_1_Adder_6_U.ce  ? \add_2ns_2ns_2_2_1_U18.top_add_2ns_2ns_2_2_1_Adder_6_U.a [1] : \add_2ns_2ns_2_2_1_U18.top_add_2ns_2ns_2_2_1_Adder_6_U.ain_s1 ;
assign _130_ = \add_2ns_2ns_2_2_1_U18.top_add_2ns_2ns_2_2_1_Adder_6_U.ce  ? \add_2ns_2ns_2_2_1_U18.top_add_2ns_2ns_2_2_1_Adder_6_U.facout_s1  : \add_2ns_2ns_2_2_1_U18.top_add_2ns_2ns_2_2_1_Adder_6_U.carry_s1 ;
assign _131_ = \add_2ns_2ns_2_2_1_U18.top_add_2ns_2ns_2_2_1_Adder_6_U.ce  ? \add_2ns_2ns_2_2_1_U18.top_add_2ns_2ns_2_2_1_Adder_6_U.fas_s1  : \add_2ns_2ns_2_2_1_U18.top_add_2ns_2ns_2_2_1_Adder_6_U.sum_s1 ;
assign _132_ = \add_2ns_2ns_2_2_1_U18.top_add_2ns_2ns_2_2_1_Adder_6_U.u1.a  + \add_2ns_2ns_2_2_1_U18.top_add_2ns_2ns_2_2_1_Adder_6_U.u1.b ;
assign { \add_2ns_2ns_2_2_1_U18.top_add_2ns_2ns_2_2_1_Adder_6_U.u1.cout , \add_2ns_2ns_2_2_1_U18.top_add_2ns_2ns_2_2_1_Adder_6_U.u1.s  } = _132_ + \add_2ns_2ns_2_2_1_U18.top_add_2ns_2ns_2_2_1_Adder_6_U.u1.cin ;
assign _133_ = \add_2ns_2ns_2_2_1_U18.top_add_2ns_2ns_2_2_1_Adder_6_U.u2.a  + \add_2ns_2ns_2_2_1_U18.top_add_2ns_2ns_2_2_1_Adder_6_U.u2.b ;
assign { \add_2ns_2ns_2_2_1_U18.top_add_2ns_2ns_2_2_1_Adder_6_U.u2.cout , \add_2ns_2ns_2_2_1_U18.top_add_2ns_2ns_2_2_1_Adder_6_U.u2.s  } = _133_ + \add_2ns_2ns_2_2_1_U18.top_add_2ns_2ns_2_2_1_Adder_6_U.u2.cin ;
always @(posedge \add_2ns_2s_2_2_1_U2.top_add_2ns_2s_2_2_1_Adder_0_U.clk )
\add_2ns_2s_2_2_1_U2.top_add_2ns_2s_2_2_1_Adder_0_U.bin_s1  <= _135_;
always @(posedge \add_2ns_2s_2_2_1_U2.top_add_2ns_2s_2_2_1_Adder_0_U.clk )
\add_2ns_2s_2_2_1_U2.top_add_2ns_2s_2_2_1_Adder_0_U.ain_s1  <= _134_;
always @(posedge \add_2ns_2s_2_2_1_U2.top_add_2ns_2s_2_2_1_Adder_0_U.clk )
\add_2ns_2s_2_2_1_U2.top_add_2ns_2s_2_2_1_Adder_0_U.sum_s1  <= _137_;
always @(posedge \add_2ns_2s_2_2_1_U2.top_add_2ns_2s_2_2_1_Adder_0_U.clk )
\add_2ns_2s_2_2_1_U2.top_add_2ns_2s_2_2_1_Adder_0_U.carry_s1  <= _136_;
assign _135_ = \add_2ns_2s_2_2_1_U2.top_add_2ns_2s_2_2_1_Adder_0_U.ce  ? \add_2ns_2s_2_2_1_U2.top_add_2ns_2s_2_2_1_Adder_0_U.b [1] : \add_2ns_2s_2_2_1_U2.top_add_2ns_2s_2_2_1_Adder_0_U.bin_s1 ;
assign _134_ = \add_2ns_2s_2_2_1_U2.top_add_2ns_2s_2_2_1_Adder_0_U.ce  ? \add_2ns_2s_2_2_1_U2.top_add_2ns_2s_2_2_1_Adder_0_U.a [1] : \add_2ns_2s_2_2_1_U2.top_add_2ns_2s_2_2_1_Adder_0_U.ain_s1 ;
assign _136_ = \add_2ns_2s_2_2_1_U2.top_add_2ns_2s_2_2_1_Adder_0_U.ce  ? \add_2ns_2s_2_2_1_U2.top_add_2ns_2s_2_2_1_Adder_0_U.facout_s1  : \add_2ns_2s_2_2_1_U2.top_add_2ns_2s_2_2_1_Adder_0_U.carry_s1 ;
assign _137_ = \add_2ns_2s_2_2_1_U2.top_add_2ns_2s_2_2_1_Adder_0_U.ce  ? \add_2ns_2s_2_2_1_U2.top_add_2ns_2s_2_2_1_Adder_0_U.fas_s1  : \add_2ns_2s_2_2_1_U2.top_add_2ns_2s_2_2_1_Adder_0_U.sum_s1 ;
assign _138_ = \add_2ns_2s_2_2_1_U2.top_add_2ns_2s_2_2_1_Adder_0_U.u1.a  + \add_2ns_2s_2_2_1_U2.top_add_2ns_2s_2_2_1_Adder_0_U.u1.b ;
assign { \add_2ns_2s_2_2_1_U2.top_add_2ns_2s_2_2_1_Adder_0_U.u1.cout , \add_2ns_2s_2_2_1_U2.top_add_2ns_2s_2_2_1_Adder_0_U.u1.s  } = _138_ + \add_2ns_2s_2_2_1_U2.top_add_2ns_2s_2_2_1_Adder_0_U.u1.cin ;
assign _139_ = \add_2ns_2s_2_2_1_U2.top_add_2ns_2s_2_2_1_Adder_0_U.u2.a  + \add_2ns_2s_2_2_1_U2.top_add_2ns_2s_2_2_1_Adder_0_U.u2.b ;
assign { \add_2ns_2s_2_2_1_U2.top_add_2ns_2s_2_2_1_Adder_0_U.u2.cout , \add_2ns_2s_2_2_1_U2.top_add_2ns_2s_2_2_1_Adder_0_U.u2.s  } = _139_ + \add_2ns_2s_2_2_1_U2.top_add_2ns_2s_2_2_1_Adder_0_U.u2.cin ;
always @(posedge \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.clk )
\add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.bin_s1  <= _141_;
always @(posedge \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.clk )
\add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.ain_s1  <= _140_;
always @(posedge \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.clk )
\add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.sum_s1  <= _143_;
always @(posedge \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.clk )
\add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.carry_s1  <= _142_;
assign _141_ = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.ce  ? \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.b [31:16] : \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.bin_s1 ;
assign _140_ = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.ce  ? \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.a [31:16] : \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.ain_s1 ;
assign _142_ = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.ce  ? \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.facout_s1  : \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.carry_s1 ;
assign _143_ = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.ce  ? \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.fas_s1  : \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.sum_s1 ;
assign _144_ = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.a  + \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.b ;
assign { \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.cout , \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.s  } = _144_ + \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.cin ;
assign _145_ = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.a  + \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.b ;
assign { \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.cout , \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.s  } = _145_ + \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.cin ;
always @(posedge \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.clk )
\add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.bin_s1  <= _147_;
always @(posedge \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.clk )
\add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.ain_s1  <= _146_;
always @(posedge \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.clk )
\add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.sum_s1  <= _149_;
always @(posedge \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.clk )
\add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.carry_s1  <= _148_;
assign _147_ = \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.ce  ? \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.b [31:16] : \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.bin_s1 ;
assign _146_ = \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.ce  ? \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.a [31:16] : \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.ain_s1 ;
assign _148_ = \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.ce  ? \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.facout_s1  : \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.carry_s1 ;
assign _149_ = \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.ce  ? \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.fas_s1  : \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.sum_s1 ;
assign _150_ = \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.a  + \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.b ;
assign { \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.cout , \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.s  } = _150_ + \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.cin ;
assign _151_ = \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.a  + \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.b ;
assign { \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.cout , \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.s  } = _151_ + \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.cin ;
always @(posedge \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.clk )
\add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.bin_s1  <= _153_;
always @(posedge \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.clk )
\add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.ain_s1  <= _152_;
always @(posedge \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.clk )
\add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.sum_s1  <= _155_;
always @(posedge \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.clk )
\add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.carry_s1  <= _154_;
assign _153_ = \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.ce  ? \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.b [31:16] : \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.bin_s1 ;
assign _152_ = \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.ce  ? \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.a [31:16] : \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.ain_s1 ;
assign _154_ = \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.ce  ? \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.facout_s1  : \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.carry_s1 ;
assign _155_ = \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.ce  ? \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.fas_s1  : \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.sum_s1 ;
assign _156_ = \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.a  + \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.b ;
assign { \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.cout , \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.s  } = _156_ + \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.cin ;
assign _157_ = \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.a  + \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.b ;
assign { \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.cout , \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.s  } = _157_ + \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.cin ;
always @(posedge \add_32ns_32ns_32_2_1_U26.top_add_32ns_32ns_32_2_1_Adder_15_U.clk )
\add_32ns_32ns_32_2_1_U26.top_add_32ns_32ns_32_2_1_Adder_15_U.bin_s1  <= _159_;
always @(posedge \add_32ns_32ns_32_2_1_U26.top_add_32ns_32ns_32_2_1_Adder_15_U.clk )
\add_32ns_32ns_32_2_1_U26.top_add_32ns_32ns_32_2_1_Adder_15_U.ain_s1  <= _158_;
always @(posedge \add_32ns_32ns_32_2_1_U26.top_add_32ns_32ns_32_2_1_Adder_15_U.clk )
\add_32ns_32ns_32_2_1_U26.top_add_32ns_32ns_32_2_1_Adder_15_U.sum_s1  <= _161_;
always @(posedge \add_32ns_32ns_32_2_1_U26.top_add_32ns_32ns_32_2_1_Adder_15_U.clk )
\add_32ns_32ns_32_2_1_U26.top_add_32ns_32ns_32_2_1_Adder_15_U.carry_s1  <= _160_;
assign _159_ = \add_32ns_32ns_32_2_1_U26.top_add_32ns_32ns_32_2_1_Adder_15_U.ce  ? \add_32ns_32ns_32_2_1_U26.top_add_32ns_32ns_32_2_1_Adder_15_U.b [31:16] : \add_32ns_32ns_32_2_1_U26.top_add_32ns_32ns_32_2_1_Adder_15_U.bin_s1 ;
assign _158_ = \add_32ns_32ns_32_2_1_U26.top_add_32ns_32ns_32_2_1_Adder_15_U.ce  ? \add_32ns_32ns_32_2_1_U26.top_add_32ns_32ns_32_2_1_Adder_15_U.a [31:16] : \add_32ns_32ns_32_2_1_U26.top_add_32ns_32ns_32_2_1_Adder_15_U.ain_s1 ;
assign _160_ = \add_32ns_32ns_32_2_1_U26.top_add_32ns_32ns_32_2_1_Adder_15_U.ce  ? \add_32ns_32ns_32_2_1_U26.top_add_32ns_32ns_32_2_1_Adder_15_U.facout_s1  : \add_32ns_32ns_32_2_1_U26.top_add_32ns_32ns_32_2_1_Adder_15_U.carry_s1 ;
assign _161_ = \add_32ns_32ns_32_2_1_U26.top_add_32ns_32ns_32_2_1_Adder_15_U.ce  ? \add_32ns_32ns_32_2_1_U26.top_add_32ns_32ns_32_2_1_Adder_15_U.fas_s1  : \add_32ns_32ns_32_2_1_U26.top_add_32ns_32ns_32_2_1_Adder_15_U.sum_s1 ;
assign _162_ = \add_32ns_32ns_32_2_1_U26.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.a  + \add_32ns_32ns_32_2_1_U26.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.b ;
assign { \add_32ns_32ns_32_2_1_U26.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.cout , \add_32ns_32ns_32_2_1_U26.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.s  } = _162_ + \add_32ns_32ns_32_2_1_U26.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.cin ;
assign _163_ = \add_32ns_32ns_32_2_1_U26.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.a  + \add_32ns_32ns_32_2_1_U26.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.b ;
assign { \add_32ns_32ns_32_2_1_U26.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.cout , \add_32ns_32ns_32_2_1_U26.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.s  } = _163_ + \add_32ns_32ns_32_2_1_U26.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.cin ;
always @(posedge \add_35s_35s_35_2_1_U24.top_add_35s_35s_35_2_1_Adder_17_U.clk )
\add_35s_35s_35_2_1_U24.top_add_35s_35s_35_2_1_Adder_17_U.bin_s1  <= _165_;
always @(posedge \add_35s_35s_35_2_1_U24.top_add_35s_35s_35_2_1_Adder_17_U.clk )
\add_35s_35s_35_2_1_U24.top_add_35s_35s_35_2_1_Adder_17_U.ain_s1  <= _164_;
always @(posedge \add_35s_35s_35_2_1_U24.top_add_35s_35s_35_2_1_Adder_17_U.clk )
\add_35s_35s_35_2_1_U24.top_add_35s_35s_35_2_1_Adder_17_U.sum_s1  <= _167_;
always @(posedge \add_35s_35s_35_2_1_U24.top_add_35s_35s_35_2_1_Adder_17_U.clk )
\add_35s_35s_35_2_1_U24.top_add_35s_35s_35_2_1_Adder_17_U.carry_s1  <= _166_;
assign _165_ = \add_35s_35s_35_2_1_U24.top_add_35s_35s_35_2_1_Adder_17_U.ce  ? \add_35s_35s_35_2_1_U24.top_add_35s_35s_35_2_1_Adder_17_U.b [34:17] : \add_35s_35s_35_2_1_U24.top_add_35s_35s_35_2_1_Adder_17_U.bin_s1 ;
assign _164_ = \add_35s_35s_35_2_1_U24.top_add_35s_35s_35_2_1_Adder_17_U.ce  ? \add_35s_35s_35_2_1_U24.top_add_35s_35s_35_2_1_Adder_17_U.a [34:17] : \add_35s_35s_35_2_1_U24.top_add_35s_35s_35_2_1_Adder_17_U.ain_s1 ;
assign _166_ = \add_35s_35s_35_2_1_U24.top_add_35s_35s_35_2_1_Adder_17_U.ce  ? \add_35s_35s_35_2_1_U24.top_add_35s_35s_35_2_1_Adder_17_U.facout_s1  : \add_35s_35s_35_2_1_U24.top_add_35s_35s_35_2_1_Adder_17_U.carry_s1 ;
assign _167_ = \add_35s_35s_35_2_1_U24.top_add_35s_35s_35_2_1_Adder_17_U.ce  ? \add_35s_35s_35_2_1_U24.top_add_35s_35s_35_2_1_Adder_17_U.fas_s1  : \add_35s_35s_35_2_1_U24.top_add_35s_35s_35_2_1_Adder_17_U.sum_s1 ;
assign _168_ = \add_35s_35s_35_2_1_U24.top_add_35s_35s_35_2_1_Adder_17_U.u1.a  + \add_35s_35s_35_2_1_U24.top_add_35s_35s_35_2_1_Adder_17_U.u1.b ;
assign { \add_35s_35s_35_2_1_U24.top_add_35s_35s_35_2_1_Adder_17_U.u1.cout , \add_35s_35s_35_2_1_U24.top_add_35s_35s_35_2_1_Adder_17_U.u1.s  } = _168_ + \add_35s_35s_35_2_1_U24.top_add_35s_35s_35_2_1_Adder_17_U.u1.cin ;
assign _169_ = \add_35s_35s_35_2_1_U24.top_add_35s_35s_35_2_1_Adder_17_U.u2.a  + \add_35s_35s_35_2_1_U24.top_add_35s_35s_35_2_1_Adder_17_U.u2.b ;
assign { \add_35s_35s_35_2_1_U24.top_add_35s_35s_35_2_1_Adder_17_U.u2.cout , \add_35s_35s_35_2_1_U24.top_add_35s_35s_35_2_1_Adder_17_U.u2.s  } = _169_ + \add_35s_35s_35_2_1_U24.top_add_35s_35s_35_2_1_Adder_17_U.u2.cin ;
always @(posedge \add_37s_37s_37_2_1_U20.top_add_37s_37s_37_2_1_Adder_14_U.clk )
\add_37s_37s_37_2_1_U20.top_add_37s_37s_37_2_1_Adder_14_U.bin_s1  <= _171_;
always @(posedge \add_37s_37s_37_2_1_U20.top_add_37s_37s_37_2_1_Adder_14_U.clk )
\add_37s_37s_37_2_1_U20.top_add_37s_37s_37_2_1_Adder_14_U.ain_s1  <= _170_;
always @(posedge \add_37s_37s_37_2_1_U20.top_add_37s_37s_37_2_1_Adder_14_U.clk )
\add_37s_37s_37_2_1_U20.top_add_37s_37s_37_2_1_Adder_14_U.sum_s1  <= _173_;
always @(posedge \add_37s_37s_37_2_1_U20.top_add_37s_37s_37_2_1_Adder_14_U.clk )
\add_37s_37s_37_2_1_U20.top_add_37s_37s_37_2_1_Adder_14_U.carry_s1  <= _172_;
assign _171_ = \add_37s_37s_37_2_1_U20.top_add_37s_37s_37_2_1_Adder_14_U.ce  ? \add_37s_37s_37_2_1_U20.top_add_37s_37s_37_2_1_Adder_14_U.b [36:18] : \add_37s_37s_37_2_1_U20.top_add_37s_37s_37_2_1_Adder_14_U.bin_s1 ;
assign _170_ = \add_37s_37s_37_2_1_U20.top_add_37s_37s_37_2_1_Adder_14_U.ce  ? \add_37s_37s_37_2_1_U20.top_add_37s_37s_37_2_1_Adder_14_U.a [36:18] : \add_37s_37s_37_2_1_U20.top_add_37s_37s_37_2_1_Adder_14_U.ain_s1 ;
assign _172_ = \add_37s_37s_37_2_1_U20.top_add_37s_37s_37_2_1_Adder_14_U.ce  ? \add_37s_37s_37_2_1_U20.top_add_37s_37s_37_2_1_Adder_14_U.facout_s1  : \add_37s_37s_37_2_1_U20.top_add_37s_37s_37_2_1_Adder_14_U.carry_s1 ;
assign _173_ = \add_37s_37s_37_2_1_U20.top_add_37s_37s_37_2_1_Adder_14_U.ce  ? \add_37s_37s_37_2_1_U20.top_add_37s_37s_37_2_1_Adder_14_U.fas_s1  : \add_37s_37s_37_2_1_U20.top_add_37s_37s_37_2_1_Adder_14_U.sum_s1 ;
assign _174_ = \add_37s_37s_37_2_1_U20.top_add_37s_37s_37_2_1_Adder_14_U.u1.a  + \add_37s_37s_37_2_1_U20.top_add_37s_37s_37_2_1_Adder_14_U.u1.b ;
assign { \add_37s_37s_37_2_1_U20.top_add_37s_37s_37_2_1_Adder_14_U.u1.cout , \add_37s_37s_37_2_1_U20.top_add_37s_37s_37_2_1_Adder_14_U.u1.s  } = _174_ + \add_37s_37s_37_2_1_U20.top_add_37s_37s_37_2_1_Adder_14_U.u1.cin ;
assign _175_ = \add_37s_37s_37_2_1_U20.top_add_37s_37s_37_2_1_Adder_14_U.u2.a  + \add_37s_37s_37_2_1_U20.top_add_37s_37s_37_2_1_Adder_14_U.u2.b ;
assign { \add_37s_37s_37_2_1_U20.top_add_37s_37s_37_2_1_Adder_14_U.u2.cout , \add_37s_37s_37_2_1_U20.top_add_37s_37s_37_2_1_Adder_14_U.u2.s  } = _175_ + \add_37s_37s_37_2_1_U20.top_add_37s_37s_37_2_1_Adder_14_U.u2.cin ;
always @(posedge \add_3s_3s_3_2_1_U4.top_add_3s_3s_3_2_1_Adder_2_U.clk )
\add_3s_3s_3_2_1_U4.top_add_3s_3s_3_2_1_Adder_2_U.bin_s1  <= _177_;
always @(posedge \add_3s_3s_3_2_1_U4.top_add_3s_3s_3_2_1_Adder_2_U.clk )
\add_3s_3s_3_2_1_U4.top_add_3s_3s_3_2_1_Adder_2_U.ain_s1  <= _176_;
always @(posedge \add_3s_3s_3_2_1_U4.top_add_3s_3s_3_2_1_Adder_2_U.clk )
\add_3s_3s_3_2_1_U4.top_add_3s_3s_3_2_1_Adder_2_U.sum_s1  <= _179_;
always @(posedge \add_3s_3s_3_2_1_U4.top_add_3s_3s_3_2_1_Adder_2_U.clk )
\add_3s_3s_3_2_1_U4.top_add_3s_3s_3_2_1_Adder_2_U.carry_s1  <= _178_;
assign _177_ = \add_3s_3s_3_2_1_U4.top_add_3s_3s_3_2_1_Adder_2_U.ce  ? \add_3s_3s_3_2_1_U4.top_add_3s_3s_3_2_1_Adder_2_U.b [2:1] : \add_3s_3s_3_2_1_U4.top_add_3s_3s_3_2_1_Adder_2_U.bin_s1 ;
assign _176_ = \add_3s_3s_3_2_1_U4.top_add_3s_3s_3_2_1_Adder_2_U.ce  ? \add_3s_3s_3_2_1_U4.top_add_3s_3s_3_2_1_Adder_2_U.a [2:1] : \add_3s_3s_3_2_1_U4.top_add_3s_3s_3_2_1_Adder_2_U.ain_s1 ;
assign _178_ = \add_3s_3s_3_2_1_U4.top_add_3s_3s_3_2_1_Adder_2_U.ce  ? \add_3s_3s_3_2_1_U4.top_add_3s_3s_3_2_1_Adder_2_U.facout_s1  : \add_3s_3s_3_2_1_U4.top_add_3s_3s_3_2_1_Adder_2_U.carry_s1 ;
assign _179_ = \add_3s_3s_3_2_1_U4.top_add_3s_3s_3_2_1_Adder_2_U.ce  ? \add_3s_3s_3_2_1_U4.top_add_3s_3s_3_2_1_Adder_2_U.fas_s1  : \add_3s_3s_3_2_1_U4.top_add_3s_3s_3_2_1_Adder_2_U.sum_s1 ;
assign _180_ = \add_3s_3s_3_2_1_U4.top_add_3s_3s_3_2_1_Adder_2_U.u1.a  + \add_3s_3s_3_2_1_U4.top_add_3s_3s_3_2_1_Adder_2_U.u1.b ;
assign { \add_3s_3s_3_2_1_U4.top_add_3s_3s_3_2_1_Adder_2_U.u1.cout , \add_3s_3s_3_2_1_U4.top_add_3s_3s_3_2_1_Adder_2_U.u1.s  } = _180_ + \add_3s_3s_3_2_1_U4.top_add_3s_3s_3_2_1_Adder_2_U.u1.cin ;
assign _181_ = \add_3s_3s_3_2_1_U4.top_add_3s_3s_3_2_1_Adder_2_U.u2.a  + \add_3s_3s_3_2_1_U4.top_add_3s_3s_3_2_1_Adder_2_U.u2.b ;
assign { \add_3s_3s_3_2_1_U4.top_add_3s_3s_3_2_1_Adder_2_U.u2.cout , \add_3s_3s_3_2_1_U4.top_add_3s_3s_3_2_1_Adder_2_U.u2.s  } = _181_ + \add_3s_3s_3_2_1_U4.top_add_3s_3s_3_2_1_Adder_2_U.u2.cin ;
always @(posedge \add_57s_57s_57_2_1_U22.top_add_57s_57s_57_2_1_Adder_16_U.clk )
\add_57s_57s_57_2_1_U22.top_add_57s_57s_57_2_1_Adder_16_U.bin_s1  <= _183_;
always @(posedge \add_57s_57s_57_2_1_U22.top_add_57s_57s_57_2_1_Adder_16_U.clk )
\add_57s_57s_57_2_1_U22.top_add_57s_57s_57_2_1_Adder_16_U.ain_s1  <= _182_;
always @(posedge \add_57s_57s_57_2_1_U22.top_add_57s_57s_57_2_1_Adder_16_U.clk )
\add_57s_57s_57_2_1_U22.top_add_57s_57s_57_2_1_Adder_16_U.sum_s1  <= _185_;
always @(posedge \add_57s_57s_57_2_1_U22.top_add_57s_57s_57_2_1_Adder_16_U.clk )
\add_57s_57s_57_2_1_U22.top_add_57s_57s_57_2_1_Adder_16_U.carry_s1  <= _184_;
assign _183_ = \add_57s_57s_57_2_1_U22.top_add_57s_57s_57_2_1_Adder_16_U.ce  ? \add_57s_57s_57_2_1_U22.top_add_57s_57s_57_2_1_Adder_16_U.b [56:28] : \add_57s_57s_57_2_1_U22.top_add_57s_57s_57_2_1_Adder_16_U.bin_s1 ;
assign _182_ = \add_57s_57s_57_2_1_U22.top_add_57s_57s_57_2_1_Adder_16_U.ce  ? \add_57s_57s_57_2_1_U22.top_add_57s_57s_57_2_1_Adder_16_U.a [56:28] : \add_57s_57s_57_2_1_U22.top_add_57s_57s_57_2_1_Adder_16_U.ain_s1 ;
assign _184_ = \add_57s_57s_57_2_1_U22.top_add_57s_57s_57_2_1_Adder_16_U.ce  ? \add_57s_57s_57_2_1_U22.top_add_57s_57s_57_2_1_Adder_16_U.facout_s1  : \add_57s_57s_57_2_1_U22.top_add_57s_57s_57_2_1_Adder_16_U.carry_s1 ;
assign _185_ = \add_57s_57s_57_2_1_U22.top_add_57s_57s_57_2_1_Adder_16_U.ce  ? \add_57s_57s_57_2_1_U22.top_add_57s_57s_57_2_1_Adder_16_U.fas_s1  : \add_57s_57s_57_2_1_U22.top_add_57s_57s_57_2_1_Adder_16_U.sum_s1 ;
assign _186_ = \add_57s_57s_57_2_1_U22.top_add_57s_57s_57_2_1_Adder_16_U.u1.a  + \add_57s_57s_57_2_1_U22.top_add_57s_57s_57_2_1_Adder_16_U.u1.b ;
assign { \add_57s_57s_57_2_1_U22.top_add_57s_57s_57_2_1_Adder_16_U.u1.cout , \add_57s_57s_57_2_1_U22.top_add_57s_57s_57_2_1_Adder_16_U.u1.s  } = _186_ + \add_57s_57s_57_2_1_U22.top_add_57s_57s_57_2_1_Adder_16_U.u1.cin ;
assign _187_ = \add_57s_57s_57_2_1_U22.top_add_57s_57s_57_2_1_Adder_16_U.u2.a  + \add_57s_57s_57_2_1_U22.top_add_57s_57s_57_2_1_Adder_16_U.u2.b ;
assign { \add_57s_57s_57_2_1_U22.top_add_57s_57s_57_2_1_Adder_16_U.u2.cout , \add_57s_57s_57_2_1_U22.top_add_57s_57s_57_2_1_Adder_16_U.u2.s  } = _187_ + \add_57s_57s_57_2_1_U22.top_add_57s_57s_57_2_1_Adder_16_U.u2.cin ;
always @(posedge \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_8_U.clk )
\add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_8_U.ain_s1  <= _188_;
always @(posedge \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_8_U.clk )
\add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_8_U.sum_s1  <= _191_;
always @(posedge \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_8_U.clk )
\add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_8_U.carry_s1  <= _190_;
always @(posedge \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_8_U.clk )
\add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_8_U.bin_s1  <= _189_;
assign _189_ = \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_8_U.ce  ? \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_8_U.b [5:3] : \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_8_U.bin_s1 ;
assign _188_ = \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_8_U.ce  ? \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_8_U.a [5:3] : \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_8_U.ain_s1 ;
assign _190_ = \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_8_U.ce  ? \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_8_U.facout_s1  : \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_8_U.carry_s1 ;
assign _191_ = \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_8_U.ce  ? \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_8_U.fas_s1  : \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_8_U.sum_s1 ;
assign _192_ = \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_8_U.u1.a  + \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_8_U.u1.b ;
assign { \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_8_U.u1.cout , \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_8_U.u1.s  } = _192_ + \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_8_U.u1.cin ;
assign _193_ = \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_8_U.u2.a  + \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_8_U.u2.b ;
assign { \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_8_U.u2.cout , \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_8_U.u2.s  } = _193_ + \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_8_U.u2.cin ;
always @(posedge \add_7ns_7ns_7_2_1_U3.top_add_7ns_7ns_7_2_1_Adder_1_U.clk )
\add_7ns_7ns_7_2_1_U3.top_add_7ns_7ns_7_2_1_Adder_1_U.bin_s1  <= _195_;
always @(posedge \add_7ns_7ns_7_2_1_U3.top_add_7ns_7ns_7_2_1_Adder_1_U.clk )
\add_7ns_7ns_7_2_1_U3.top_add_7ns_7ns_7_2_1_Adder_1_U.ain_s1  <= _194_;
always @(posedge \add_7ns_7ns_7_2_1_U3.top_add_7ns_7ns_7_2_1_Adder_1_U.clk )
\add_7ns_7ns_7_2_1_U3.top_add_7ns_7ns_7_2_1_Adder_1_U.sum_s1  <= _197_;
always @(posedge \add_7ns_7ns_7_2_1_U3.top_add_7ns_7ns_7_2_1_Adder_1_U.clk )
\add_7ns_7ns_7_2_1_U3.top_add_7ns_7ns_7_2_1_Adder_1_U.carry_s1  <= _196_;
assign _195_ = \add_7ns_7ns_7_2_1_U3.top_add_7ns_7ns_7_2_1_Adder_1_U.ce  ? \add_7ns_7ns_7_2_1_U3.top_add_7ns_7ns_7_2_1_Adder_1_U.b [6:3] : \add_7ns_7ns_7_2_1_U3.top_add_7ns_7ns_7_2_1_Adder_1_U.bin_s1 ;
assign _194_ = \add_7ns_7ns_7_2_1_U3.top_add_7ns_7ns_7_2_1_Adder_1_U.ce  ? \add_7ns_7ns_7_2_1_U3.top_add_7ns_7ns_7_2_1_Adder_1_U.a [6:3] : \add_7ns_7ns_7_2_1_U3.top_add_7ns_7ns_7_2_1_Adder_1_U.ain_s1 ;
assign _196_ = \add_7ns_7ns_7_2_1_U3.top_add_7ns_7ns_7_2_1_Adder_1_U.ce  ? \add_7ns_7ns_7_2_1_U3.top_add_7ns_7ns_7_2_1_Adder_1_U.facout_s1  : \add_7ns_7ns_7_2_1_U3.top_add_7ns_7ns_7_2_1_Adder_1_U.carry_s1 ;
assign _197_ = \add_7ns_7ns_7_2_1_U3.top_add_7ns_7ns_7_2_1_Adder_1_U.ce  ? \add_7ns_7ns_7_2_1_U3.top_add_7ns_7ns_7_2_1_Adder_1_U.fas_s1  : \add_7ns_7ns_7_2_1_U3.top_add_7ns_7ns_7_2_1_Adder_1_U.sum_s1 ;
assign _198_ = \add_7ns_7ns_7_2_1_U3.top_add_7ns_7ns_7_2_1_Adder_1_U.u1.a  + \add_7ns_7ns_7_2_1_U3.top_add_7ns_7ns_7_2_1_Adder_1_U.u1.b ;
assign { \add_7ns_7ns_7_2_1_U3.top_add_7ns_7ns_7_2_1_Adder_1_U.u1.cout , \add_7ns_7ns_7_2_1_U3.top_add_7ns_7ns_7_2_1_Adder_1_U.u1.s  } = _198_ + \add_7ns_7ns_7_2_1_U3.top_add_7ns_7ns_7_2_1_Adder_1_U.u1.cin ;
assign _199_ = \add_7ns_7ns_7_2_1_U3.top_add_7ns_7ns_7_2_1_Adder_1_U.u2.a  + \add_7ns_7ns_7_2_1_U3.top_add_7ns_7ns_7_2_1_Adder_1_U.u2.b ;
assign { \add_7ns_7ns_7_2_1_U3.top_add_7ns_7ns_7_2_1_Adder_1_U.u2.cout , \add_7ns_7ns_7_2_1_U3.top_add_7ns_7ns_7_2_1_Adder_1_U.u2.s  } = _199_ + \add_7ns_7ns_7_2_1_U3.top_add_7ns_7ns_7_2_1_Adder_1_U.u2.cin ;
always @(posedge \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_9_U.clk )
\add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_9_U.bin_s1  <= _201_;
always @(posedge \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_9_U.clk )
\add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_9_U.ain_s1  <= _200_;
always @(posedge \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_9_U.clk )
\add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_9_U.sum_s1  <= _203_;
always @(posedge \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_9_U.clk )
\add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_9_U.carry_s1  <= _202_;
assign _201_ = \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_9_U.ce  ? \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_9_U.b [6:3] : \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_9_U.bin_s1 ;
assign _200_ = \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_9_U.ce  ? \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_9_U.a [6:3] : \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_9_U.ain_s1 ;
assign _202_ = \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_9_U.ce  ? \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_9_U.facout_s1  : \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_9_U.carry_s1 ;
assign _203_ = \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_9_U.ce  ? \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_9_U.fas_s1  : \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_9_U.sum_s1 ;
assign _204_ = \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_9_U.u1.a  + \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_9_U.u1.b ;
assign { \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_9_U.u1.cout , \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_9_U.u1.s  } = _204_ + \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_9_U.u1.cin ;
assign _205_ = \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_9_U.u2.a  + \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_9_U.u2.b ;
assign { \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_9_U.u2.cout , \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_9_U.u2.s  } = _205_ + \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_9_U.u2.cin ;
always @(posedge \add_9ns_9s_9_2_1_U11.top_add_9ns_9s_9_2_1_Adder_7_U.clk )
\add_9ns_9s_9_2_1_U11.top_add_9ns_9s_9_2_1_Adder_7_U.bin_s1  <= _207_;
always @(posedge \add_9ns_9s_9_2_1_U11.top_add_9ns_9s_9_2_1_Adder_7_U.clk )
\add_9ns_9s_9_2_1_U11.top_add_9ns_9s_9_2_1_Adder_7_U.ain_s1  <= _206_;
always @(posedge \add_9ns_9s_9_2_1_U11.top_add_9ns_9s_9_2_1_Adder_7_U.clk )
\add_9ns_9s_9_2_1_U11.top_add_9ns_9s_9_2_1_Adder_7_U.sum_s1  <= _209_;
always @(posedge \add_9ns_9s_9_2_1_U11.top_add_9ns_9s_9_2_1_Adder_7_U.clk )
\add_9ns_9s_9_2_1_U11.top_add_9ns_9s_9_2_1_Adder_7_U.carry_s1  <= _208_;
assign _207_ = \add_9ns_9s_9_2_1_U11.top_add_9ns_9s_9_2_1_Adder_7_U.ce  ? \add_9ns_9s_9_2_1_U11.top_add_9ns_9s_9_2_1_Adder_7_U.b [8:4] : \add_9ns_9s_9_2_1_U11.top_add_9ns_9s_9_2_1_Adder_7_U.bin_s1 ;
assign _206_ = \add_9ns_9s_9_2_1_U11.top_add_9ns_9s_9_2_1_Adder_7_U.ce  ? \add_9ns_9s_9_2_1_U11.top_add_9ns_9s_9_2_1_Adder_7_U.a [8:4] : \add_9ns_9s_9_2_1_U11.top_add_9ns_9s_9_2_1_Adder_7_U.ain_s1 ;
assign _208_ = \add_9ns_9s_9_2_1_U11.top_add_9ns_9s_9_2_1_Adder_7_U.ce  ? \add_9ns_9s_9_2_1_U11.top_add_9ns_9s_9_2_1_Adder_7_U.facout_s1  : \add_9ns_9s_9_2_1_U11.top_add_9ns_9s_9_2_1_Adder_7_U.carry_s1 ;
assign _209_ = \add_9ns_9s_9_2_1_U11.top_add_9ns_9s_9_2_1_Adder_7_U.ce  ? \add_9ns_9s_9_2_1_U11.top_add_9ns_9s_9_2_1_Adder_7_U.fas_s1  : \add_9ns_9s_9_2_1_U11.top_add_9ns_9s_9_2_1_Adder_7_U.sum_s1 ;
assign _210_ = \add_9ns_9s_9_2_1_U11.top_add_9ns_9s_9_2_1_Adder_7_U.u1.a  + \add_9ns_9s_9_2_1_U11.top_add_9ns_9s_9_2_1_Adder_7_U.u1.b ;
assign { \add_9ns_9s_9_2_1_U11.top_add_9ns_9s_9_2_1_Adder_7_U.u1.cout , \add_9ns_9s_9_2_1_U11.top_add_9ns_9s_9_2_1_Adder_7_U.u1.s  } = _210_ + \add_9ns_9s_9_2_1_U11.top_add_9ns_9s_9_2_1_Adder_7_U.u1.cin ;
assign _211_ = \add_9ns_9s_9_2_1_U11.top_add_9ns_9s_9_2_1_Adder_7_U.u2.a  + \add_9ns_9s_9_2_1_U11.top_add_9ns_9s_9_2_1_Adder_7_U.u2.b ;
assign { \add_9ns_9s_9_2_1_U11.top_add_9ns_9s_9_2_1_Adder_7_U.u2.cout , \add_9ns_9s_9_2_1_U11.top_add_9ns_9s_9_2_1_Adder_7_U.u2.s  } = _211_ + \add_9ns_9s_9_2_1_U11.top_add_9ns_9s_9_2_1_Adder_7_U.u2.cin ;
always @(posedge \ashr_32s_16ns_32_7_1_U8.clk )
\ashr_32s_16ns_32_7_1_U8.dout_array[5]  <= _223_;
always @(posedge \ashr_32s_16ns_32_7_1_U8.clk )
\ashr_32s_16ns_32_7_1_U8.din1_cast_array[5]  <= _217_;
always @(posedge \ashr_32s_16ns_32_7_1_U8.clk )
\ashr_32s_16ns_32_7_1_U8.dout_array[4]  <= _222_;
always @(posedge \ashr_32s_16ns_32_7_1_U8.clk )
\ashr_32s_16ns_32_7_1_U8.din1_cast_array[4]  <= _216_;
always @(posedge \ashr_32s_16ns_32_7_1_U8.clk )
\ashr_32s_16ns_32_7_1_U8.dout_array[3]  <= _221_;
always @(posedge \ashr_32s_16ns_32_7_1_U8.clk )
\ashr_32s_16ns_32_7_1_U8.din1_cast_array[3]  <= _215_;
always @(posedge \ashr_32s_16ns_32_7_1_U8.clk )
\ashr_32s_16ns_32_7_1_U8.dout_array[2]  <= _220_;
always @(posedge \ashr_32s_16ns_32_7_1_U8.clk )
\ashr_32s_16ns_32_7_1_U8.din1_cast_array[2]  <= _214_;
always @(posedge \ashr_32s_16ns_32_7_1_U8.clk )
\ashr_32s_16ns_32_7_1_U8.dout_array[1]  <= _219_;
always @(posedge \ashr_32s_16ns_32_7_1_U8.clk )
\ashr_32s_16ns_32_7_1_U8.din1_cast_array[1]  <= _213_;
always @(posedge \ashr_32s_16ns_32_7_1_U8.clk )
\ashr_32s_16ns_32_7_1_U8.dout_array[0]  <= _218_;
always @(posedge \ashr_32s_16ns_32_7_1_U8.clk )
\ashr_32s_16ns_32_7_1_U8.din1_cast_array[0]  <= _212_;
assign _224_ = \ashr_32s_16ns_32_7_1_U8.ce  ? \ashr_32s_16ns_32_7_1_U8.din1_cast_array[4]  : \ashr_32s_16ns_32_7_1_U8.din1_cast_array[5] ;
assign _217_ = \ashr_32s_16ns_32_7_1_U8.reset  ? 16'h0000 : _224_;
assign _225_ = \ashr_32s_16ns_32_7_1_U8.ce  ? _240_ : \ashr_32s_16ns_32_7_1_U8.dout_array[5] ;
assign _223_ = \ashr_32s_16ns_32_7_1_U8.reset  ? 32'd0 : _225_;
assign _226_ = \ashr_32s_16ns_32_7_1_U8.ce  ? \ashr_32s_16ns_32_7_1_U8.din1_cast_array[3]  : \ashr_32s_16ns_32_7_1_U8.din1_cast_array[4] ;
assign _216_ = \ashr_32s_16ns_32_7_1_U8.reset  ? 16'h0000 : _226_;
assign _227_ = \ashr_32s_16ns_32_7_1_U8.ce  ? _239_ : \ashr_32s_16ns_32_7_1_U8.dout_array[4] ;
assign _222_ = \ashr_32s_16ns_32_7_1_U8.reset  ? 32'd0 : _227_;
assign _228_ = \ashr_32s_16ns_32_7_1_U8.ce  ? \ashr_32s_16ns_32_7_1_U8.din1_cast_array[2]  : \ashr_32s_16ns_32_7_1_U8.din1_cast_array[3] ;
assign _215_ = \ashr_32s_16ns_32_7_1_U8.reset  ? 16'h0000 : _228_;
assign _229_ = \ashr_32s_16ns_32_7_1_U8.ce  ? _238_ : \ashr_32s_16ns_32_7_1_U8.dout_array[3] ;
assign _221_ = \ashr_32s_16ns_32_7_1_U8.reset  ? 32'd0 : _229_;
assign _230_ = \ashr_32s_16ns_32_7_1_U8.ce  ? \ashr_32s_16ns_32_7_1_U8.din1_cast_array[1]  : \ashr_32s_16ns_32_7_1_U8.din1_cast_array[2] ;
assign _214_ = \ashr_32s_16ns_32_7_1_U8.reset  ? 16'h0000 : _230_;
assign _231_ = \ashr_32s_16ns_32_7_1_U8.ce  ? _237_ : \ashr_32s_16ns_32_7_1_U8.dout_array[2] ;
assign _220_ = \ashr_32s_16ns_32_7_1_U8.reset  ? 32'd0 : _231_;
assign _232_ = \ashr_32s_16ns_32_7_1_U8.ce  ? \ashr_32s_16ns_32_7_1_U8.din1_cast_array[0]  : \ashr_32s_16ns_32_7_1_U8.din1_cast_array[1] ;
assign _213_ = \ashr_32s_16ns_32_7_1_U8.reset  ? 16'h0000 : _232_;
assign _233_ = \ashr_32s_16ns_32_7_1_U8.ce  ? _236_ : \ashr_32s_16ns_32_7_1_U8.dout_array[1] ;
assign _219_ = \ashr_32s_16ns_32_7_1_U8.reset  ? 32'd0 : _233_;
assign _234_ = \ashr_32s_16ns_32_7_1_U8.ce  ? \ashr_32s_16ns_32_7_1_U8.din1 [15:0] : \ashr_32s_16ns_32_7_1_U8.din1_cast_array[0] ;
assign _212_ = \ashr_32s_16ns_32_7_1_U8.reset  ? 16'h0000 : _234_;
assign _235_ = \ashr_32s_16ns_32_7_1_U8.ce  ? \ashr_32s_16ns_32_7_1_U8.din0  : \ashr_32s_16ns_32_7_1_U8.dout_array[0] ;
assign _218_ = \ashr_32s_16ns_32_7_1_U8.reset  ? 32'd0 : _235_;
assign _236_ = $signed(\ashr_32s_16ns_32_7_1_U8.dout_array[0] ) >>> { \ashr_32s_16ns_32_7_1_U8.din1_cast_array[0] [15], 15'h0000 };
assign _237_ = $signed(\ashr_32s_16ns_32_7_1_U8.dout_array[1] ) >>> { \ashr_32s_16ns_32_7_1_U8.din1_cast_array[1] [14:12], 12'h000 };
assign _238_ = $signed(\ashr_32s_16ns_32_7_1_U8.dout_array[2] ) >>> { \ashr_32s_16ns_32_7_1_U8.din1_cast_array[2] [11:9], 9'h000 };
assign _239_ = $signed(\ashr_32s_16ns_32_7_1_U8.dout_array[3] ) >>> { \ashr_32s_16ns_32_7_1_U8.din1_cast_array[3] [8:6], 6'h00 };
assign _240_ = $signed(\ashr_32s_16ns_32_7_1_U8.dout_array[4] ) >>> { \ashr_32s_16ns_32_7_1_U8.din1_cast_array[4] [5:3], 3'h0 };
assign \ashr_32s_16ns_32_7_1_U8.dout  = $signed(\ashr_32s_16ns_32_7_1_U8.dout_array[5] ) >>> \ashr_32s_16ns_32_7_1_U8.din1_cast_array[5] [2:0];
assign \mul_8s_2s_10_7_1_U1.top_mul_8s_2s_10_7_1_Mul_DSP_0_U.tmp_product  = $signed(\mul_8s_2s_10_7_1_U1.top_mul_8s_2s_10_7_1_Mul_DSP_0_U.a_reg0 ) * $signed(\mul_8s_2s_10_7_1_U1.top_mul_8s_2s_10_7_1_Mul_DSP_0_U.b_reg0 );
always @(posedge \mul_8s_2s_10_7_1_U1.top_mul_8s_2s_10_7_1_Mul_DSP_0_U.clk )
\mul_8s_2s_10_7_1_U1.top_mul_8s_2s_10_7_1_Mul_DSP_0_U.a_reg0  <= _241_;
always @(posedge \mul_8s_2s_10_7_1_U1.top_mul_8s_2s_10_7_1_Mul_DSP_0_U.clk )
\mul_8s_2s_10_7_1_U1.top_mul_8s_2s_10_7_1_Mul_DSP_0_U.b_reg0  <= _242_;
always @(posedge \mul_8s_2s_10_7_1_U1.top_mul_8s_2s_10_7_1_Mul_DSP_0_U.clk )
\mul_8s_2s_10_7_1_U1.top_mul_8s_2s_10_7_1_Mul_DSP_0_U.buff0  <= _243_;
always @(posedge \mul_8s_2s_10_7_1_U1.top_mul_8s_2s_10_7_1_Mul_DSP_0_U.clk )
\mul_8s_2s_10_7_1_U1.top_mul_8s_2s_10_7_1_Mul_DSP_0_U.buff1  <= _244_;
always @(posedge \mul_8s_2s_10_7_1_U1.top_mul_8s_2s_10_7_1_Mul_DSP_0_U.clk )
\mul_8s_2s_10_7_1_U1.top_mul_8s_2s_10_7_1_Mul_DSP_0_U.buff2  <= _245_;
always @(posedge \mul_8s_2s_10_7_1_U1.top_mul_8s_2s_10_7_1_Mul_DSP_0_U.clk )
\mul_8s_2s_10_7_1_U1.top_mul_8s_2s_10_7_1_Mul_DSP_0_U.buff3  <= _246_;
always @(posedge \mul_8s_2s_10_7_1_U1.top_mul_8s_2s_10_7_1_Mul_DSP_0_U.clk )
\mul_8s_2s_10_7_1_U1.top_mul_8s_2s_10_7_1_Mul_DSP_0_U.buff4  <= _247_;
assign _247_ = \mul_8s_2s_10_7_1_U1.top_mul_8s_2s_10_7_1_Mul_DSP_0_U.ce  ? \mul_8s_2s_10_7_1_U1.top_mul_8s_2s_10_7_1_Mul_DSP_0_U.buff3  : \mul_8s_2s_10_7_1_U1.top_mul_8s_2s_10_7_1_Mul_DSP_0_U.buff4 ;
assign _246_ = \mul_8s_2s_10_7_1_U1.top_mul_8s_2s_10_7_1_Mul_DSP_0_U.ce  ? \mul_8s_2s_10_7_1_U1.top_mul_8s_2s_10_7_1_Mul_DSP_0_U.buff2  : \mul_8s_2s_10_7_1_U1.top_mul_8s_2s_10_7_1_Mul_DSP_0_U.buff3 ;
assign _245_ = \mul_8s_2s_10_7_1_U1.top_mul_8s_2s_10_7_1_Mul_DSP_0_U.ce  ? \mul_8s_2s_10_7_1_U1.top_mul_8s_2s_10_7_1_Mul_DSP_0_U.buff1  : \mul_8s_2s_10_7_1_U1.top_mul_8s_2s_10_7_1_Mul_DSP_0_U.buff2 ;
assign _244_ = \mul_8s_2s_10_7_1_U1.top_mul_8s_2s_10_7_1_Mul_DSP_0_U.ce  ? \mul_8s_2s_10_7_1_U1.top_mul_8s_2s_10_7_1_Mul_DSP_0_U.buff0  : \mul_8s_2s_10_7_1_U1.top_mul_8s_2s_10_7_1_Mul_DSP_0_U.buff1 ;
assign _243_ = \mul_8s_2s_10_7_1_U1.top_mul_8s_2s_10_7_1_Mul_DSP_0_U.ce  ? \mul_8s_2s_10_7_1_U1.top_mul_8s_2s_10_7_1_Mul_DSP_0_U.tmp_product  : \mul_8s_2s_10_7_1_U1.top_mul_8s_2s_10_7_1_Mul_DSP_0_U.buff0 ;
assign _242_ = \mul_8s_2s_10_7_1_U1.top_mul_8s_2s_10_7_1_Mul_DSP_0_U.ce  ? \mul_8s_2s_10_7_1_U1.top_mul_8s_2s_10_7_1_Mul_DSP_0_U.b  : \mul_8s_2s_10_7_1_U1.top_mul_8s_2s_10_7_1_Mul_DSP_0_U.b_reg0 ;
assign _241_ = \mul_8s_2s_10_7_1_U1.top_mul_8s_2s_10_7_1_Mul_DSP_0_U.ce  ? \mul_8s_2s_10_7_1_U1.top_mul_8s_2s_10_7_1_Mul_DSP_0_U.a  : \mul_8s_2s_10_7_1_U1.top_mul_8s_2s_10_7_1_Mul_DSP_0_U.a_reg0 ;
always @(posedge \shl_32s_16ns_32_7_1_U9.clk )
\shl_32s_16ns_32_7_1_U9.dout_array[5]  <= _259_;
always @(posedge \shl_32s_16ns_32_7_1_U9.clk )
\shl_32s_16ns_32_7_1_U9.din1_cast_array[5]  <= _253_;
always @(posedge \shl_32s_16ns_32_7_1_U9.clk )
\shl_32s_16ns_32_7_1_U9.dout_array[4]  <= _258_;
always @(posedge \shl_32s_16ns_32_7_1_U9.clk )
\shl_32s_16ns_32_7_1_U9.din1_cast_array[4]  <= _252_;
always @(posedge \shl_32s_16ns_32_7_1_U9.clk )
\shl_32s_16ns_32_7_1_U9.dout_array[3]  <= _257_;
always @(posedge \shl_32s_16ns_32_7_1_U9.clk )
\shl_32s_16ns_32_7_1_U9.din1_cast_array[3]  <= _251_;
always @(posedge \shl_32s_16ns_32_7_1_U9.clk )
\shl_32s_16ns_32_7_1_U9.dout_array[2]  <= _256_;
always @(posedge \shl_32s_16ns_32_7_1_U9.clk )
\shl_32s_16ns_32_7_1_U9.din1_cast_array[2]  <= _250_;
always @(posedge \shl_32s_16ns_32_7_1_U9.clk )
\shl_32s_16ns_32_7_1_U9.dout_array[1]  <= _255_;
always @(posedge \shl_32s_16ns_32_7_1_U9.clk )
\shl_32s_16ns_32_7_1_U9.din1_cast_array[1]  <= _249_;
always @(posedge \shl_32s_16ns_32_7_1_U9.clk )
\shl_32s_16ns_32_7_1_U9.dout_array[0]  <= _254_;
always @(posedge \shl_32s_16ns_32_7_1_U9.clk )
\shl_32s_16ns_32_7_1_U9.din1_cast_array[0]  <= _248_;
assign _260_ = \shl_32s_16ns_32_7_1_U9.ce  ? \shl_32s_16ns_32_7_1_U9.din1_cast_array[4]  : \shl_32s_16ns_32_7_1_U9.din1_cast_array[5] ;
assign _253_ = \shl_32s_16ns_32_7_1_U9.reset  ? 16'h0000 : _260_;
assign _261_ = \shl_32s_16ns_32_7_1_U9.ce  ? _276_ : \shl_32s_16ns_32_7_1_U9.dout_array[5] ;
assign _259_ = \shl_32s_16ns_32_7_1_U9.reset  ? 32'd0 : _261_;
assign _262_ = \shl_32s_16ns_32_7_1_U9.ce  ? \shl_32s_16ns_32_7_1_U9.din1_cast_array[3]  : \shl_32s_16ns_32_7_1_U9.din1_cast_array[4] ;
assign _252_ = \shl_32s_16ns_32_7_1_U9.reset  ? 16'h0000 : _262_;
assign _263_ = \shl_32s_16ns_32_7_1_U9.ce  ? _275_ : \shl_32s_16ns_32_7_1_U9.dout_array[4] ;
assign _258_ = \shl_32s_16ns_32_7_1_U9.reset  ? 32'd0 : _263_;
assign _264_ = \shl_32s_16ns_32_7_1_U9.ce  ? \shl_32s_16ns_32_7_1_U9.din1_cast_array[2]  : \shl_32s_16ns_32_7_1_U9.din1_cast_array[3] ;
assign _251_ = \shl_32s_16ns_32_7_1_U9.reset  ? 16'h0000 : _264_;
assign _265_ = \shl_32s_16ns_32_7_1_U9.ce  ? _274_ : \shl_32s_16ns_32_7_1_U9.dout_array[3] ;
assign _257_ = \shl_32s_16ns_32_7_1_U9.reset  ? 32'd0 : _265_;
assign _266_ = \shl_32s_16ns_32_7_1_U9.ce  ? \shl_32s_16ns_32_7_1_U9.din1_cast_array[1]  : \shl_32s_16ns_32_7_1_U9.din1_cast_array[2] ;
assign _250_ = \shl_32s_16ns_32_7_1_U9.reset  ? 16'h0000 : _266_;
assign _267_ = \shl_32s_16ns_32_7_1_U9.ce  ? _273_ : \shl_32s_16ns_32_7_1_U9.dout_array[2] ;
assign _256_ = \shl_32s_16ns_32_7_1_U9.reset  ? 32'd0 : _267_;
assign _268_ = \shl_32s_16ns_32_7_1_U9.ce  ? \shl_32s_16ns_32_7_1_U9.din1_cast_array[0]  : \shl_32s_16ns_32_7_1_U9.din1_cast_array[1] ;
assign _249_ = \shl_32s_16ns_32_7_1_U9.reset  ? 16'h0000 : _268_;
assign _269_ = \shl_32s_16ns_32_7_1_U9.ce  ? _272_ : \shl_32s_16ns_32_7_1_U9.dout_array[1] ;
assign _255_ = \shl_32s_16ns_32_7_1_U9.reset  ? 32'd0 : _269_;
assign _270_ = \shl_32s_16ns_32_7_1_U9.ce  ? \shl_32s_16ns_32_7_1_U9.din1 [15:0] : \shl_32s_16ns_32_7_1_U9.din1_cast_array[0] ;
assign _248_ = \shl_32s_16ns_32_7_1_U9.reset  ? 16'h0000 : _270_;
assign _271_ = \shl_32s_16ns_32_7_1_U9.ce  ? \shl_32s_16ns_32_7_1_U9.din0  : \shl_32s_16ns_32_7_1_U9.dout_array[0] ;
assign _254_ = \shl_32s_16ns_32_7_1_U9.reset  ? 32'd0 : _271_;
assign _272_ = \shl_32s_16ns_32_7_1_U9.dout_array[0]  << { \shl_32s_16ns_32_7_1_U9.din1_cast_array[0] [15], 15'h0000 };
assign _273_ = \shl_32s_16ns_32_7_1_U9.dout_array[1]  << { \shl_32s_16ns_32_7_1_U9.din1_cast_array[1] [14:12], 12'h000 };
assign _274_ = \shl_32s_16ns_32_7_1_U9.dout_array[2]  << { \shl_32s_16ns_32_7_1_U9.din1_cast_array[2] [11:9], 9'h000 };
assign _275_ = \shl_32s_16ns_32_7_1_U9.dout_array[3]  << { \shl_32s_16ns_32_7_1_U9.din1_cast_array[3] [8:6], 6'h00 };
assign _276_ = \shl_32s_16ns_32_7_1_U9.dout_array[4]  << { \shl_32s_16ns_32_7_1_U9.din1_cast_array[4] [5:3], 3'h0 };
assign \shl_32s_16ns_32_7_1_U9.dout  = \shl_32s_16ns_32_7_1_U9.dout_array[5]  << \shl_32s_16ns_32_7_1_U9.din1_cast_array[5] [2:0];
assign \sub_11s_11s_11_2_1_U5.top_sub_11s_11s_11_2_1_Adder_3_U.bin_s0  = ~ \sub_11s_11s_11_2_1_U5.top_sub_11s_11s_11_2_1_Adder_3_U.b ;
always @(posedge \sub_11s_11s_11_2_1_U5.top_sub_11s_11s_11_2_1_Adder_3_U.clk )
\sub_11s_11s_11_2_1_U5.top_sub_11s_11s_11_2_1_Adder_3_U.bin_s1  <= _278_;
always @(posedge \sub_11s_11s_11_2_1_U5.top_sub_11s_11s_11_2_1_Adder_3_U.clk )
\sub_11s_11s_11_2_1_U5.top_sub_11s_11s_11_2_1_Adder_3_U.ain_s1  <= _277_;
always @(posedge \sub_11s_11s_11_2_1_U5.top_sub_11s_11s_11_2_1_Adder_3_U.clk )
\sub_11s_11s_11_2_1_U5.top_sub_11s_11s_11_2_1_Adder_3_U.sum_s1  <= _280_;
always @(posedge \sub_11s_11s_11_2_1_U5.top_sub_11s_11s_11_2_1_Adder_3_U.clk )
\sub_11s_11s_11_2_1_U5.top_sub_11s_11s_11_2_1_Adder_3_U.carry_s1  <= _279_;
assign _278_ = \sub_11s_11s_11_2_1_U5.top_sub_11s_11s_11_2_1_Adder_3_U.ce  ? \sub_11s_11s_11_2_1_U5.top_sub_11s_11s_11_2_1_Adder_3_U.bin_s0 [10:5] : \sub_11s_11s_11_2_1_U5.top_sub_11s_11s_11_2_1_Adder_3_U.bin_s1 ;
assign _277_ = \sub_11s_11s_11_2_1_U5.top_sub_11s_11s_11_2_1_Adder_3_U.ce  ? \sub_11s_11s_11_2_1_U5.top_sub_11s_11s_11_2_1_Adder_3_U.a [10:5] : \sub_11s_11s_11_2_1_U5.top_sub_11s_11s_11_2_1_Adder_3_U.ain_s1 ;
assign _279_ = \sub_11s_11s_11_2_1_U5.top_sub_11s_11s_11_2_1_Adder_3_U.ce  ? \sub_11s_11s_11_2_1_U5.top_sub_11s_11s_11_2_1_Adder_3_U.facout_s1  : \sub_11s_11s_11_2_1_U5.top_sub_11s_11s_11_2_1_Adder_3_U.carry_s1 ;
assign _280_ = \sub_11s_11s_11_2_1_U5.top_sub_11s_11s_11_2_1_Adder_3_U.ce  ? \sub_11s_11s_11_2_1_U5.top_sub_11s_11s_11_2_1_Adder_3_U.fas_s1  : \sub_11s_11s_11_2_1_U5.top_sub_11s_11s_11_2_1_Adder_3_U.sum_s1 ;
assign _281_ = \sub_11s_11s_11_2_1_U5.top_sub_11s_11s_11_2_1_Adder_3_U.u1.a  + \sub_11s_11s_11_2_1_U5.top_sub_11s_11s_11_2_1_Adder_3_U.u1.b ;
assign { \sub_11s_11s_11_2_1_U5.top_sub_11s_11s_11_2_1_Adder_3_U.u1.cout , \sub_11s_11s_11_2_1_U5.top_sub_11s_11s_11_2_1_Adder_3_U.u1.s  } = _281_ + \sub_11s_11s_11_2_1_U5.top_sub_11s_11s_11_2_1_Adder_3_U.u1.cin ;
assign _282_ = \sub_11s_11s_11_2_1_U5.top_sub_11s_11s_11_2_1_Adder_3_U.u2.a  + \sub_11s_11s_11_2_1_U5.top_sub_11s_11s_11_2_1_Adder_3_U.u2.b ;
assign { \sub_11s_11s_11_2_1_U5.top_sub_11s_11s_11_2_1_Adder_3_U.u2.cout , \sub_11s_11s_11_2_1_U5.top_sub_11s_11s_11_2_1_Adder_3_U.u2.s  } = _282_ + \sub_11s_11s_11_2_1_U5.top_sub_11s_11s_11_2_1_Adder_3_U.u2.cin ;
assign \sub_8ns_8s_8_2_1_U6.top_sub_8ns_8s_8_2_1_Adder_4_U.bin_s0  = ~ \sub_8ns_8s_8_2_1_U6.top_sub_8ns_8s_8_2_1_Adder_4_U.b ;
always @(posedge \sub_8ns_8s_8_2_1_U6.top_sub_8ns_8s_8_2_1_Adder_4_U.clk )
\sub_8ns_8s_8_2_1_U6.top_sub_8ns_8s_8_2_1_Adder_4_U.bin_s1  <= _284_;
always @(posedge \sub_8ns_8s_8_2_1_U6.top_sub_8ns_8s_8_2_1_Adder_4_U.clk )
\sub_8ns_8s_8_2_1_U6.top_sub_8ns_8s_8_2_1_Adder_4_U.ain_s1  <= _283_;
always @(posedge \sub_8ns_8s_8_2_1_U6.top_sub_8ns_8s_8_2_1_Adder_4_U.clk )
\sub_8ns_8s_8_2_1_U6.top_sub_8ns_8s_8_2_1_Adder_4_U.sum_s1  <= _286_;
always @(posedge \sub_8ns_8s_8_2_1_U6.top_sub_8ns_8s_8_2_1_Adder_4_U.clk )
\sub_8ns_8s_8_2_1_U6.top_sub_8ns_8s_8_2_1_Adder_4_U.carry_s1  <= _285_;
assign _284_ = \sub_8ns_8s_8_2_1_U6.top_sub_8ns_8s_8_2_1_Adder_4_U.ce  ? \sub_8ns_8s_8_2_1_U6.top_sub_8ns_8s_8_2_1_Adder_4_U.bin_s0 [7:4] : \sub_8ns_8s_8_2_1_U6.top_sub_8ns_8s_8_2_1_Adder_4_U.bin_s1 ;
assign _283_ = \sub_8ns_8s_8_2_1_U6.top_sub_8ns_8s_8_2_1_Adder_4_U.ce  ? \sub_8ns_8s_8_2_1_U6.top_sub_8ns_8s_8_2_1_Adder_4_U.a [7:4] : \sub_8ns_8s_8_2_1_U6.top_sub_8ns_8s_8_2_1_Adder_4_U.ain_s1 ;
assign _285_ = \sub_8ns_8s_8_2_1_U6.top_sub_8ns_8s_8_2_1_Adder_4_U.ce  ? \sub_8ns_8s_8_2_1_U6.top_sub_8ns_8s_8_2_1_Adder_4_U.facout_s1  : \sub_8ns_8s_8_2_1_U6.top_sub_8ns_8s_8_2_1_Adder_4_U.carry_s1 ;
assign _286_ = \sub_8ns_8s_8_2_1_U6.top_sub_8ns_8s_8_2_1_Adder_4_U.ce  ? \sub_8ns_8s_8_2_1_U6.top_sub_8ns_8s_8_2_1_Adder_4_U.fas_s1  : \sub_8ns_8s_8_2_1_U6.top_sub_8ns_8s_8_2_1_Adder_4_U.sum_s1 ;
assign _287_ = \sub_8ns_8s_8_2_1_U6.top_sub_8ns_8s_8_2_1_Adder_4_U.u1.a  + \sub_8ns_8s_8_2_1_U6.top_sub_8ns_8s_8_2_1_Adder_4_U.u1.b ;
assign { \sub_8ns_8s_8_2_1_U6.top_sub_8ns_8s_8_2_1_Adder_4_U.u1.cout , \sub_8ns_8s_8_2_1_U6.top_sub_8ns_8s_8_2_1_Adder_4_U.u1.s  } = _287_ + \sub_8ns_8s_8_2_1_U6.top_sub_8ns_8s_8_2_1_Adder_4_U.u1.cin ;
assign _288_ = \sub_8ns_8s_8_2_1_U6.top_sub_8ns_8s_8_2_1_Adder_4_U.u2.a  + \sub_8ns_8s_8_2_1_U6.top_sub_8ns_8s_8_2_1_Adder_4_U.u2.b ;
assign { \sub_8ns_8s_8_2_1_U6.top_sub_8ns_8s_8_2_1_Adder_4_U.u2.cout , \sub_8ns_8s_8_2_1_U6.top_sub_8ns_8s_8_2_1_Adder_4_U.u2.s  } = _288_ + \sub_8ns_8s_8_2_1_U6.top_sub_8ns_8s_8_2_1_Adder_4_U.u2.cin ;
assign _289_ = | { tmp_5_reg_1279, 1'h0, p_Result_s_20_reg_1285 };
assign _290_ = p_Result_s_20_reg_1285 != 2'h3;
assign _291_ = | trunc_ln851_2_reg_1158;
assign _292_ = | trunc_ln851_4_reg_1342;
assign _293_ = | op_16[3:0];
assign _294_ = | op_17[23:0];
assign _295_ = | op_18[1:0];
assign op_8_V_fu_356_p2 = op_4[7:0] | { op_2_V_reg_1084[1], op_2_V_reg_1084[1], op_2_V_reg_1084[1], op_2_V_reg_1084[1], op_2_V_reg_1084[1], op_2_V_reg_1084[1], op_2_V_reg_1084 };
assign or_ln384_fu_713_p2 = underflow_fu_701_p2 | overflow_reg_1311;
assign or_ln786_fu_697_p2 = icmp_ln786_reg_1317 | icmp_ln786_1_reg_1301;
always @(posedge ap_clk)
trunc_ln769_reg_1258 <= _062_;
always @(posedge ap_clk)
trunc_ln546_reg_1253 <= _061_;
always @(posedge ap_clk)
sh_V_1_reg_1163 <= _058_;
always @(posedge ap_clk)
sext_ln850_reg_1372 <= _057_;
always @(posedge ap_clk)
select_ln353_reg_1456 <= _054_;
always @(posedge ap_clk)
select_ln353_1_reg_1493 <= _053_;
always @(posedge ap_clk)
ret_reg_1127 <= _052_;
always @(posedge ap_clk)
ret_V_5_reg_1243 <= _050_;
always @(posedge ap_clk)
ret_V_30_reg_1530 <= _048_;
always @(posedge ap_clk)
select_ln69_1_reg_1535 <= _055_;
always @(posedge ap_clk)
ret_V_26_reg_1384 <= _044_;
always @(posedge ap_clk)
select_ln69_reg_1389 <= _056_;
always @(posedge ap_clk)
ret_V_25_reg_1362 <= _043_;
always @(posedge ap_clk)
tmp_1_reg_1367 <= _059_;
always @(posedge ap_clk)
ret_V_29_reg_1513 <= _047_;
always @(posedge ap_clk)
ret_V_25_cast_reg_1518 <= _042_;
always @(posedge ap_clk)
ret_V_22_reg_1201 <= _039_;
always @(posedge ap_clk)
ret_V_28_reg_1476 <= _046_;
always @(posedge ap_clk)
ret_V_22_cast_reg_1481 <= _038_;
always @(posedge ap_clk)
ret_V_20_reg_1248 <= _036_;
always @(posedge ap_clk)
ret_V_19_reg_1231 <= _034_;
always @(posedge ap_clk)
ret_V_4_reg_1236 <= _049_;
always @(posedge ap_clk)
ret_V_27_reg_1439 <= _045_;
always @(posedge ap_clk)
ret_V_19_cast_reg_1444 <= _033_;
always @(posedge ap_clk)
ret_V_21_reg_1152 <= _037_;
always @(posedge ap_clk)
trunc_ln851_2_reg_1158 <= _063_;
always @(posedge ap_clk)
ret_V_23_reg_1168 <= _040_;
always @(posedge ap_clk)
ret_V_12_cast_reg_1173 <= _031_;
always @(posedge ap_clk)
ret_V_10_reg_1206 <= _030_;
always @(posedge ap_clk)
r_V_reg_1057 <= _028_;
always @(posedge ap_clk)
ret_V_reg_1062 <= _051_;
always @(posedge ap_clk)
trunc_ln851_reg_1069 <= _065_;
always @(posedge ap_clk)
r_reg_1268 <= _029_;
always @(posedge ap_clk)
p_Result_11_reg_1273 <= _026_;
always @(posedge ap_clk)
tmp_5_reg_1279 <= _060_;
always @(posedge ap_clk)
p_Result_s_20_reg_1285 <= _027_;
always @(posedge ap_clk)
ret_V_18_reg_1095 <= _032_;
always @(posedge ap_clk)
op_8_V_reg_1112 <= _023_;
always @(posedge ap_clk)
p_Result_10_reg_1117 <= _025_;
always @(posedge ap_clk)
op_2_V_reg_1084 <= _022_;
always @(posedge ap_clk)
ret_V_1_reg_1090 <= _035_;
always @(posedge ap_clk)
op_26_V_reg_1419 <= _021_;
always @(posedge ap_clk)
op_12_V_reg_1332 <= _019_;
always @(posedge ap_clk)
op_22_V_reg_1337 <= _020_;
always @(posedge ap_clk)
trunc_ln851_4_reg_1342 <= _064_;
always @(posedge ap_clk)
icmp_ln851_reg_1079 <= _018_;
always @(posedge ap_clk)
icmp_ln851_6_reg_1508 <= _017_;
always @(posedge ap_clk)
icmp_ln851_5_reg_1471 <= _016_;
always @(posedge ap_clk)
icmp_ln851_4_reg_1434 <= _015_;
always @(posedge ap_clk)
icmp_ln851_3_reg_1357 <= _014_;
always @(posedge ap_clk)
icmp_ln851_2_reg_1052 <= _013_;
always @(posedge ap_clk)
icmp_ln851_1_reg_1221 <= _012_;
always @(posedge ap_clk)
ret_V_24_reg_1226 <= _041_;
always @(posedge ap_clk)
icmp_ln850_reg_1180 <= _011_;
always @(posedge ap_clk)
overflow_reg_1311 <= _024_;
always @(posedge ap_clk)
icmp_ln786_reg_1317 <= _010_;
always @(posedge ap_clk)
icmp_ln785_reg_1296 <= _008_;
always @(posedge ap_clk)
icmp_ln786_1_reg_1301 <= _009_;
always @(posedge ap_clk)
add_ln69_reg_1306 <= _006_;
always @(posedge ap_clk)
add_ln69_2_reg_1404 <= _004_;
always @(posedge ap_clk)
add_ln69_3_reg_1409 <= _005_;
always @(posedge ap_clk)
add_ln691_reg_1379 <= _003_;
always @(posedge ap_clk)
add_ln691_3_reg_1525 <= _002_;
always @(posedge ap_clk)
add_ln691_2_reg_1488 <= _001_;
always @(posedge ap_clk)
add_ln691_1_reg_1451 <= _000_;
always @(posedge ap_clk)
ap_CS_fsm <= _007_;
assign _066_ = _077_ ? 2'h2 : 2'h1;
assign _296_ = ap_CS_fsm == 1'h1;
function [48:0] _823_;
input [48:0] a;
input [2400:0] b;
input [48:0] s;
case (s)
49'b0000000000000000000000000000000000000000000000001:
_823_ = b[48:0];
49'b0000000000000000000000000000000000000000000000010:
_823_ = b[97:49];
49'b0000000000000000000000000000000000000000000000100:
_823_ = b[146:98];
49'b0000000000000000000000000000000000000000000001000:
_823_ = b[195:147];
49'b0000000000000000000000000000000000000000000010000:
_823_ = b[244:196];
49'b0000000000000000000000000000000000000000000100000:
_823_ = b[293:245];
49'b0000000000000000000000000000000000000000001000000:
_823_ = b[342:294];
49'b0000000000000000000000000000000000000000010000000:
_823_ = b[391:343];
49'b0000000000000000000000000000000000000000100000000:
_823_ = b[440:392];
49'b0000000000000000000000000000000000000001000000000:
_823_ = b[489:441];
49'b0000000000000000000000000000000000000010000000000:
_823_ = b[538:490];
49'b0000000000000000000000000000000000000100000000000:
_823_ = b[587:539];
49'b0000000000000000000000000000000000001000000000000:
_823_ = b[636:588];
49'b0000000000000000000000000000000000010000000000000:
_823_ = b[685:637];
49'b0000000000000000000000000000000000100000000000000:
_823_ = b[734:686];
49'b0000000000000000000000000000000001000000000000000:
_823_ = b[783:735];
49'b0000000000000000000000000000000010000000000000000:
_823_ = b[832:784];
49'b0000000000000000000000000000000100000000000000000:
_823_ = b[881:833];
49'b0000000000000000000000000000001000000000000000000:
_823_ = b[930:882];
49'b0000000000000000000000000000010000000000000000000:
_823_ = b[979:931];
49'b0000000000000000000000000000100000000000000000000:
_823_ = b[1028:980];
49'b0000000000000000000000000001000000000000000000000:
_823_ = b[1077:1029];
49'b0000000000000000000000000010000000000000000000000:
_823_ = b[1126:1078];
49'b0000000000000000000000000100000000000000000000000:
_823_ = b[1175:1127];
49'b0000000000000000000000001000000000000000000000000:
_823_ = b[1224:1176];
49'b0000000000000000000000010000000000000000000000000:
_823_ = b[1273:1225];
49'b0000000000000000000000100000000000000000000000000:
_823_ = b[1322:1274];
49'b0000000000000000000001000000000000000000000000000:
_823_ = b[1371:1323];
49'b0000000000000000000010000000000000000000000000000:
_823_ = b[1420:1372];
49'b0000000000000000000100000000000000000000000000000:
_823_ = b[1469:1421];
49'b0000000000000000001000000000000000000000000000000:
_823_ = b[1518:1470];
49'b0000000000000000010000000000000000000000000000000:
_823_ = b[1567:1519];
49'b0000000000000000100000000000000000000000000000000:
_823_ = b[1616:1568];
49'b0000000000000001000000000000000000000000000000000:
_823_ = b[1665:1617];
49'b0000000000000010000000000000000000000000000000000:
_823_ = b[1714:1666];
49'b0000000000000100000000000000000000000000000000000:
_823_ = b[1763:1715];
49'b0000000000001000000000000000000000000000000000000:
_823_ = b[1812:1764];
49'b0000000000010000000000000000000000000000000000000:
_823_ = b[1861:1813];
49'b0000000000100000000000000000000000000000000000000:
_823_ = b[1910:1862];
49'b0000000001000000000000000000000000000000000000000:
_823_ = b[1959:1911];
49'b0000000010000000000000000000000000000000000000000:
_823_ = b[2008:1960];
49'b0000000100000000000000000000000000000000000000000:
_823_ = b[2057:2009];
49'b0000001000000000000000000000000000000000000000000:
_823_ = b[2106:2058];
49'b0000010000000000000000000000000000000000000000000:
_823_ = b[2155:2107];
49'b0000100000000000000000000000000000000000000000000:
_823_ = b[2204:2156];
49'b0001000000000000000000000000000000000000000000000:
_823_ = b[2253:2205];
49'b0010000000000000000000000000000000000000000000000:
_823_ = b[2302:2254];
49'b0100000000000000000000000000000000000000000000000:
_823_ = b[2351:2303];
49'b1000000000000000000000000000000000000000000000000:
_823_ = b[2400:2352];
49'b0000000000000000000000000000000000000000000000000:
_823_ = a;
default:
_823_ = 49'bx;
endcase
endfunction
assign ap_NS_fsm = _823_(49'hxxxxxxxxxxxxx, { 47'h000000000000, _066_, 2352'h000000000002000000000002000000000002000000000002000000000002000000000002000000000002000000000002000000000002000000000002000000000002000000000002000000000002000000000002000000000002000000000002000000000002000000000002000000000002000000000002000000000002000000000002000000000002000000000002000000000002000000000002000000000002000000000002000000000002000000000002000000000002000000000002000000000002000000000002000000000002000000000002000000000002000000000002000000000002000000000002000000000002000000000002000000000002000000000002000000000002000000000002000000000002000000000000000000000001 }, { _296_, _344_, _343_, _342_, _341_, _340_, _339_, _338_, _337_, _336_, _335_, _334_, _333_, _332_, _331_, _330_, _329_, _328_, _327_, _326_, _325_, _324_, _323_, _322_, _321_, _320_, _319_, _318_, _317_, _316_, _315_, _314_, _313_, _312_, _311_, _310_, _309_, _308_, _307_, _306_, _305_, _304_, _303_, _302_, _301_, _300_, _299_, _298_, _297_ });
assign _297_ = ap_CS_fsm == 49'h1000000000000;
assign _298_ = ap_CS_fsm == 48'h800000000000;
assign _299_ = ap_CS_fsm == 47'h400000000000;
assign _300_ = ap_CS_fsm == 46'h200000000000;
assign _301_ = ap_CS_fsm == 45'h100000000000;
assign _302_ = ap_CS_fsm == 44'h80000000000;
assign _303_ = ap_CS_fsm == 43'h40000000000;
assign _304_ = ap_CS_fsm == 42'h20000000000;
assign _305_ = ap_CS_fsm == 41'h10000000000;
assign _306_ = ap_CS_fsm == 40'h8000000000;
assign _307_ = ap_CS_fsm == 39'h4000000000;
assign _308_ = ap_CS_fsm == 38'h2000000000;
assign _309_ = ap_CS_fsm == 37'h1000000000;
assign _310_ = ap_CS_fsm == 36'h800000000;
assign _311_ = ap_CS_fsm == 35'h400000000;
assign _312_ = ap_CS_fsm == 34'h200000000;
assign _313_ = ap_CS_fsm == 33'h100000000;
assign _314_ = ap_CS_fsm == 32'd2147483648;
assign _315_ = ap_CS_fsm == 31'h40000000;
assign _316_ = ap_CS_fsm == 30'h20000000;
assign _317_ = ap_CS_fsm == 29'h10000000;
assign _318_ = ap_CS_fsm == 28'h8000000;
assign _319_ = ap_CS_fsm == 27'h4000000;
assign _320_ = ap_CS_fsm == 26'h2000000;
assign _321_ = ap_CS_fsm == 25'h1000000;
assign _322_ = ap_CS_fsm == 24'h800000;
assign _323_ = ap_CS_fsm == 23'h400000;
assign _324_ = ap_CS_fsm == 22'h200000;
assign _325_ = ap_CS_fsm == 21'h100000;
assign _326_ = ap_CS_fsm == 20'h80000;
assign _327_ = ap_CS_fsm == 19'h40000;
assign _328_ = ap_CS_fsm == 18'h20000;
assign _329_ = ap_CS_fsm == 17'h10000;
assign _330_ = ap_CS_fsm == 16'h8000;
assign _331_ = ap_CS_fsm == 15'h4000;
assign _332_ = ap_CS_fsm == 14'h2000;
assign _333_ = ap_CS_fsm == 13'h1000;
assign _334_ = ap_CS_fsm == 12'h800;
assign _335_ = ap_CS_fsm == 11'h400;
assign _336_ = ap_CS_fsm == 10'h200;
assign _337_ = ap_CS_fsm == 9'h100;
assign _338_ = ap_CS_fsm == 8'h80;
assign _339_ = ap_CS_fsm == 7'h40;
assign _340_ = ap_CS_fsm == 6'h20;
assign _341_ = ap_CS_fsm == 5'h10;
assign _342_ = ap_CS_fsm == 4'h8;
assign _343_ = ap_CS_fsm == 3'h4;
assign _344_ = ap_CS_fsm == 2'h2;
assign op_30_ap_vld = ap_CS_fsm[48] ? 1'h1 : 1'h0;
assign ap_idle = _076_ ? 1'h1 : 1'h0;
assign _062_ = _075_ ? grp_fu_461_p2[3:0] : trunc_ln769_reg_1258;
assign _061_ = _074_ ? grp_fu_448_p2[2:0] : trunc_ln546_reg_1253;
assign _058_ = _073_ ? grp_fu_393_p2 : sh_V_1_reg_1163;
assign _057_ = ap_CS_fsm[25] ? { tmp_1_reg_1367[17], tmp_1_reg_1367 } : sext_ln850_reg_1372;
assign _054_ = ap_CS_fsm[36] ? select_ln353_fu_880_p3 : select_ln353_reg_1456;
assign _053_ = ap_CS_fsm[41] ? select_ln353_1_fu_945_p3 : select_ln353_1_reg_1493;
assign _052_ = ap_CS_fsm[10] ? grp_fu_343_p2 : ret_reg_1127;
assign _050_ = _072_ ? grp_fu_558_p2 : ret_V_5_reg_1243;
assign _055_ = ap_CS_fsm[46] ? select_ln69_1_fu_1017_p3 : select_ln69_1_reg_1535;
assign _048_ = ap_CS_fsm[46] ? ret_V_30_fu_1010_p3 : ret_V_30_reg_1530;
assign _056_ = ap_CS_fsm[27] ? select_ln69_fu_789_p3 : select_ln69_reg_1389;
assign _044_ = ap_CS_fsm[27] ? ret_V_26_fu_782_p3 : ret_V_26_reg_1384;
assign _059_ = ap_CS_fsm[24] ? grp_fu_740_p2[19:2] : tmp_1_reg_1367;
assign _043_ = ap_CS_fsm[24] ? grp_fu_740_p2 : ret_V_25_reg_1362;
assign _042_ = ap_CS_fsm[43] ? grp_fu_967_p2[33:2] : ret_V_25_cast_reg_1518;
assign _047_ = ap_CS_fsm[43] ? grp_fu_967_p2 : ret_V_29_reg_1513;
assign _039_ = ap_CS_fsm[13] ? ret_V_22_fu_491_p2 : ret_V_22_reg_1201;
assign _038_ = ap_CS_fsm[38] ? grp_fu_902_p2[55:24] : ret_V_22_cast_reg_1481;
assign _046_ = ap_CS_fsm[38] ? grp_fu_902_p2 : ret_V_28_reg_1476;
assign _036_ = ap_CS_fsm[18] ? ret_V_20_fu_575_p3 : ret_V_20_reg_1248;
assign _049_ = ap_CS_fsm[15] ? grp_fu_513_p2[8:3] : ret_V_4_reg_1236;
assign _034_ = ap_CS_fsm[15] ? grp_fu_513_p2 : ret_V_19_reg_1231;
assign _033_ = ap_CS_fsm[33] ? grp_fu_837_p2[35:4] : ret_V_19_cast_reg_1444;
assign _045_ = ap_CS_fsm[33] ? grp_fu_837_p2 : ret_V_27_reg_1439;
assign _031_ = ap_CS_fsm[11] ? grp_fu_413_p2[4:3] : ret_V_12_cast_reg_1173;
assign _040_ = ap_CS_fsm[11] ? grp_fu_413_p2 : ret_V_23_reg_1168;
assign _063_ = ap_CS_fsm[11] ? grp_fu_387_p2[2:0] : trunc_ln851_2_reg_1158;
assign _037_ = ap_CS_fsm[11] ? grp_fu_387_p2 : ret_V_21_reg_1152;
assign _030_ = _071_ ? grp_fu_467_p2 : ret_V_10_reg_1206;
assign _065_ = ap_CS_fsm[6] ? grp_fu_269_p2[2:0] : trunc_ln851_reg_1069;
assign _051_ = ap_CS_fsm[6] ? grp_fu_269_p2[9:3] : ret_V_reg_1062;
assign _028_ = ap_CS_fsm[6] ? grp_fu_269_p2 : r_V_reg_1057;
assign _027_ = ap_CS_fsm[19] ? r_fu_596_p3[3:2] : p_Result_s_20_reg_1285;
assign _060_ = ap_CS_fsm[19] ? r_fu_596_p3[1] : tmp_5_reg_1279;
assign _026_ = ap_CS_fsm[19] ? r_fu_596_p3[3] : p_Result_11_reg_1273;
assign _029_ = ap_CS_fsm[19] ? r_fu_596_p3 : r_reg_1268;
assign _025_ = ap_CS_fsm[9] ? ret_V_18_fu_330_p3[6] : p_Result_10_reg_1117;
assign _023_ = ap_CS_fsm[9] ? op_8_V_fu_356_p2 : op_8_V_reg_1112;
assign _032_ = ap_CS_fsm[9] ? ret_V_18_fu_330_p3 : ret_V_18_reg_1095;
assign _035_ = ap_CS_fsm[8] ? grp_fu_313_p2 : ret_V_1_reg_1090;
assign _022_ = ap_CS_fsm[8] ? grp_fu_303_p2 : op_2_V_reg_1084;
assign _021_ = ap_CS_fsm[31] ? grp_fu_817_p2 : op_26_V_reg_1419;
assign _064_ = ap_CS_fsm[22] ? op_12_V_fu_718_p3[1:0] : trunc_ln851_4_reg_1342;
assign _020_ = ap_CS_fsm[22] ? grp_fu_686_p2 : op_22_V_reg_1337;
assign _019_ = ap_CS_fsm[22] ? op_12_V_fu_718_p3 : op_12_V_reg_1332;
assign _018_ = ap_CS_fsm[7] ? icmp_ln851_fu_308_p2 : icmp_ln851_reg_1079;
assign _017_ = ap_CS_fsm[42] ? icmp_ln851_6_fu_977_p2 : icmp_ln851_6_reg_1508;
assign _016_ = ap_CS_fsm[37] ? icmp_ln851_5_fu_912_p2 : icmp_ln851_5_reg_1471;
assign _015_ = ap_CS_fsm[32] ? icmp_ln851_4_fu_847_p2 : icmp_ln851_4_reg_1434;
assign _014_ = ap_CS_fsm[23] ? icmp_ln851_3_fu_746_p2 : icmp_ln851_3_reg_1357;
assign _013_ = ap_CS_fsm[0] ? icmp_ln851_2_fu_279_p2 : icmp_ln851_2_reg_1052;
assign _041_ = ap_CS_fsm[14] ? ret_V_24_fu_541_p3 : ret_V_24_reg_1226;
assign _012_ = ap_CS_fsm[14] ? icmp_ln851_1_fu_523_p2 : icmp_ln851_1_reg_1221;
assign _011_ = ap_CS_fsm[12] ? icmp_ln850_fu_433_p2 : icmp_ln850_reg_1180;
assign _010_ = ap_CS_fsm[21] ? icmp_ln786_fu_673_p2 : icmp_ln786_reg_1317;
assign _024_ = ap_CS_fsm[21] ? overflow_fu_668_p2 : overflow_reg_1311;
assign _006_ = ap_CS_fsm[20] ? grp_fu_631_p2 : add_ln69_reg_1306;
assign _009_ = ap_CS_fsm[20] ? icmp_ln786_1_fu_651_p2 : icmp_ln786_1_reg_1301;
assign _008_ = ap_CS_fsm[20] ? icmp_ln785_fu_645_p2 : icmp_ln785_reg_1296;
assign _005_ = ap_CS_fsm[29] ? grp_fu_809_p2 : add_ln69_3_reg_1409;
assign _004_ = ap_CS_fsm[29] ? grp_fu_804_p2 : add_ln69_2_reg_1404;
assign _003_ = _070_ ? grp_fu_764_p2 : add_ln691_reg_1379;
assign _002_ = _069_ ? grp_fu_993_p2 : add_ln691_3_reg_1525;
assign _001_ = _068_ ? grp_fu_928_p2 : add_ln691_2_reg_1488;
assign _000_ = _067_ ? grp_fu_863_p2 : add_ln691_1_reg_1451;
assign _007_ = ap_rst ? 49'h0000000000001 : ap_NS_fsm;
assign icmp_ln785_fu_645_p2 = _289_ ? 1'h1 : 1'h0;
assign icmp_ln786_1_fu_651_p2 = _290_ ? 1'h1 : 1'h0;
assign icmp_ln786_fu_673_p2 = _082_ ? 1'h1 : 1'h0;
assign icmp_ln850_fu_433_p2 = _291_ ? 1'h1 : 1'h0;
assign icmp_ln851_1_fu_523_p2 = _083_ ? 1'h1 : 1'h0;
assign icmp_ln851_2_fu_279_p2 = _084_ ? 1'h1 : 1'h0;
assign icmp_ln851_3_fu_746_p2 = _292_ ? 1'h1 : 1'h0;
assign icmp_ln851_4_fu_847_p2 = _293_ ? 1'h1 : 1'h0;
assign icmp_ln851_5_fu_912_p2 = _294_ ? 1'h1 : 1'h0;
assign icmp_ln851_6_fu_977_p2 = _295_ ? 1'h1 : 1'h0;
assign icmp_ln851_fu_308_p2 = _085_ ? 1'h1 : 1'h0;
assign op_12_V_fu_718_p3 = or_ln384_fu_713_p2 ? select_ln384_fu_706_p3 : { r_reg_1268[1:0], 2'h0 };
assign r_fu_596_p3 = p_Result_10_reg_1117 ? { trunc_ln546_reg_1253[2], trunc_ln546_reg_1253 } : trunc_ln769_reg_1258;
assign ret_V_18_fu_330_p3 = r_V_reg_1057[9] ? select_ln850_fu_325_p3 : ret_V_reg_1062;
assign ret_V_20_fu_575_p3 = ret_V_19_reg_1231[8] ? select_ln850_1_fu_570_p3 : ret_V_4_reg_1236;
assign ret_V_24_fu_541_p3 = ret_V_23_reg_1168[11] ? select_ln850_3_fu_536_p3 : ret_V_12_cast_reg_1173;
assign ret_V_26_fu_782_p3 = ret_V_25_reg_1362[19] ? select_ln850_4_fu_777_p3 : sext_ln850_reg_1372;
assign ret_V_30_fu_1010_p3 = ret_V_29_reg_1513[34] ? select_ln850_7_fu_1005_p3 : ret_V_25_cast_reg_1518;
assign select_ln353_1_fu_945_p3 = ret_V_28_reg_1476[56] ? select_ln850_8_fu_940_p3 : ret_V_22_cast_reg_1481;
assign select_ln353_fu_880_p3 = ret_V_27_reg_1439[36] ? select_ln850_6_fu_875_p3 : ret_V_19_cast_reg_1444;
assign select_ln384_fu_706_p3 = overflow_reg_1311 ? 4'h7 : 4'h8;
assign select_ln69_1_fu_1017_p3 = op_19 ? 32'd4294967295 : 32'd0;
assign select_ln69_fu_789_p3 = op_15 ? 2'h3 : 2'h0;
assign select_ln850_1_fu_570_p3 = icmp_ln851_1_reg_1221 ? ret_V_4_reg_1236 : ret_V_5_reg_1243;
assign select_ln850_3_fu_536_p3 = icmp_ln851_2_reg_1052 ? ret_V_12_cast_reg_1173 : ret_V_10_reg_1206;
assign select_ln850_4_fu_777_p3 = icmp_ln851_3_reg_1357 ? add_ln691_reg_1379 : sext_ln850_reg_1372;
assign select_ln850_6_fu_875_p3 = icmp_ln851_4_reg_1434 ? add_ln691_1_reg_1451 : ret_V_19_cast_reg_1444;
assign select_ln850_7_fu_1005_p3 = icmp_ln851_6_reg_1508 ? add_ln691_3_reg_1525 : ret_V_25_cast_reg_1518;
assign select_ln850_8_fu_940_p3 = icmp_ln851_5_reg_1471 ? add_ln691_2_reg_1488 : ret_V_22_cast_reg_1481;
assign select_ln850_fu_325_p3 = icmp_ln851_reg_1079 ? ret_V_reg_1062 : ret_V_1_reg_1090;
assign ret_V_22_fu_491_p2 = ret_V_21_reg_1152[3] ^ and_ln353_fu_486_p2;
assign and_ln_fu_656_p3 = { tmp_5_reg_1279, 3'h0 };
assign ap_CS_fsm_state1 = ap_CS_fsm[0];
assign ap_CS_fsm_state10 = ap_CS_fsm[9];
assign ap_CS_fsm_state11 = ap_CS_fsm[10];
assign ap_CS_fsm_state12 = ap_CS_fsm[11];
assign ap_CS_fsm_state13 = ap_CS_fsm[12];
assign ap_CS_fsm_state14 = ap_CS_fsm[13];
assign ap_CS_fsm_state15 = ap_CS_fsm[14];
assign ap_CS_fsm_state16 = ap_CS_fsm[15];
assign ap_CS_fsm_state17 = ap_CS_fsm[16];
assign ap_CS_fsm_state18 = ap_CS_fsm[17];
assign ap_CS_fsm_state19 = ap_CS_fsm[18];
assign ap_CS_fsm_state20 = ap_CS_fsm[19];
assign ap_CS_fsm_state21 = ap_CS_fsm[20];
assign ap_CS_fsm_state22 = ap_CS_fsm[21];
assign ap_CS_fsm_state23 = ap_CS_fsm[22];
assign ap_CS_fsm_state24 = ap_CS_fsm[23];
assign ap_CS_fsm_state25 = ap_CS_fsm[24];
assign ap_CS_fsm_state26 = ap_CS_fsm[25];
assign ap_CS_fsm_state27 = ap_CS_fsm[26];
assign ap_CS_fsm_state28 = ap_CS_fsm[27];
assign ap_CS_fsm_state29 = ap_CS_fsm[28];
assign ap_CS_fsm_state30 = ap_CS_fsm[29];
assign ap_CS_fsm_state31 = ap_CS_fsm[30];
assign ap_CS_fsm_state32 = ap_CS_fsm[31];
assign ap_CS_fsm_state33 = ap_CS_fsm[32];
assign ap_CS_fsm_state34 = ap_CS_fsm[33];
assign ap_CS_fsm_state35 = ap_CS_fsm[34];
assign ap_CS_fsm_state36 = ap_CS_fsm[35];
assign ap_CS_fsm_state37 = ap_CS_fsm[36];
assign ap_CS_fsm_state38 = ap_CS_fsm[37];
assign ap_CS_fsm_state39 = ap_CS_fsm[38];
assign ap_CS_fsm_state40 = ap_CS_fsm[39];
assign ap_CS_fsm_state41 = ap_CS_fsm[40];
assign ap_CS_fsm_state42 = ap_CS_fsm[41];
assign ap_CS_fsm_state43 = ap_CS_fsm[42];
assign ap_CS_fsm_state44 = ap_CS_fsm[43];
assign ap_CS_fsm_state45 = ap_CS_fsm[44];
assign ap_CS_fsm_state46 = ap_CS_fsm[45];
assign ap_CS_fsm_state47 = ap_CS_fsm[46];
assign ap_CS_fsm_state48 = ap_CS_fsm[47];
assign ap_CS_fsm_state49 = ap_CS_fsm[48];
assign ap_CS_fsm_state7 = ap_CS_fsm[6];
assign ap_CS_fsm_state8 = ap_CS_fsm[7];
assign ap_CS_fsm_state9 = ap_CS_fsm[8];
assign ap_done = op_30_ap_vld;
assign ap_ready = op_30_ap_vld;
assign grp_fu_303_p0 = op_0[1:0];
assign grp_fu_343_p0 = { op_2_V_reg_1084[1], op_2_V_reg_1084 };
assign grp_fu_343_p1 = { op_1[1], op_1 };
assign grp_fu_387_p0 = { op_3[7], op_3[7], op_3[7], op_3 };
assign grp_fu_387_p1 = { ret_V_18_reg_1095[6], ret_V_18_reg_1095, 3'h0 };
assign grp_fu_393_p1 = { ret_V_18_reg_1095[6], ret_V_18_reg_1095 };
assign grp_fu_413_p0 = { op_8_V_reg_1112[7], op_8_V_reg_1112, 3'h0 };
assign grp_fu_413_p1 = { op_3[7], op_3[7], op_3[7], op_3[7], op_3 };
assign grp_fu_448_p1 = { 16'h0000, sh_V_1_reg_1163[7], sh_V_1_reg_1163[7], sh_V_1_reg_1163[7], sh_V_1_reg_1163[7], sh_V_1_reg_1163[7], sh_V_1_reg_1163[7], sh_V_1_reg_1163[7], sh_V_1_reg_1163[7], sh_V_1_reg_1163 };
assign grp_fu_461_p1 = { 16'h0000, ret_V_18_reg_1095[6], ret_V_18_reg_1095[6], ret_V_18_reg_1095[6], ret_V_18_reg_1095[6], ret_V_18_reg_1095[6], ret_V_18_reg_1095[6], ret_V_18_reg_1095[6], ret_V_18_reg_1095[6], ret_V_18_reg_1095[6], ret_V_18_reg_1095 };
assign grp_fu_513_p0 = { 2'h0, op_7, 3'h0 };
assign grp_fu_513_p1 = { op_9[7], op_9 };
assign grp_fu_631_p0 = { ret_V_20_reg_1248[5], ret_V_20_reg_1248 };
assign grp_fu_631_p1 = { ret_V_24_reg_1226[1], ret_V_24_reg_1226[1], ret_V_24_reg_1226[1], ret_V_24_reg_1226[1], ret_V_24_reg_1226[1], ret_V_24_reg_1226 };
assign grp_fu_686_p0 = { add_ln69_reg_1306[6], add_ln69_reg_1306[6], add_ln69_reg_1306[6], add_ln69_reg_1306[6], add_ln69_reg_1306[6], add_ln69_reg_1306[6], add_ln69_reg_1306[6], add_ln69_reg_1306[6], add_ln69_reg_1306[6], add_ln69_reg_1306[6], add_ln69_reg_1306[6], add_ln69_reg_1306 };
assign grp_fu_686_p1 = { 2'h0, op_11 };
assign grp_fu_740_p0 = { op_22_V_reg_1337, 2'h0 };
assign grp_fu_740_p1 = { op_12_V_reg_1332[3], op_12_V_reg_1332[3], op_12_V_reg_1332[3], op_12_V_reg_1332[3], op_12_V_reg_1332[3], op_12_V_reg_1332[3], op_12_V_reg_1332[3], op_12_V_reg_1332[3], op_12_V_reg_1332[3], op_12_V_reg_1332[3], op_12_V_reg_1332[3], op_12_V_reg_1332[3], op_12_V_reg_1332[3], op_12_V_reg_1332[3], op_12_V_reg_1332[3], op_12_V_reg_1332[3], op_12_V_reg_1332 };
assign grp_fu_764_p0 = { tmp_1_reg_1367[17], tmp_1_reg_1367 };
assign grp_fu_804_p1 = { op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14 };
assign grp_fu_809_p1 = { 1'h0, ret_V_22_reg_1201 };
assign grp_fu_817_p0 = { add_ln69_3_reg_1409[1], add_ln69_3_reg_1409[1], add_ln69_3_reg_1409[1], add_ln69_3_reg_1409[1], add_ln69_3_reg_1409[1], add_ln69_3_reg_1409[1], add_ln69_3_reg_1409[1], add_ln69_3_reg_1409[1], add_ln69_3_reg_1409[1], add_ln69_3_reg_1409[1], add_ln69_3_reg_1409[1], add_ln69_3_reg_1409[1], add_ln69_3_reg_1409[1], add_ln69_3_reg_1409[1], add_ln69_3_reg_1409[1], add_ln69_3_reg_1409[1], add_ln69_3_reg_1409[1], add_ln69_3_reg_1409 };
assign grp_fu_837_p0 = { op_26_V_reg_1419[18], op_26_V_reg_1419[18], op_26_V_reg_1419[18], op_26_V_reg_1419[18], op_26_V_reg_1419[18], op_26_V_reg_1419[18], op_26_V_reg_1419[18], op_26_V_reg_1419[18], op_26_V_reg_1419[18], op_26_V_reg_1419[18], op_26_V_reg_1419[18], op_26_V_reg_1419[18], op_26_V_reg_1419[18], op_26_V_reg_1419[18], op_26_V_reg_1419, 4'h0 };
assign grp_fu_837_p1 = { op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16 };
assign grp_fu_902_p0 = { select_ln353_reg_1456[31], select_ln353_reg_1456, 24'h000000 };
assign grp_fu_902_p1 = { op_17[31], op_17[31], op_17[31], op_17[31], op_17[31], op_17[31], op_17[31], op_17[31], op_17[31], op_17[31], op_17[31], op_17[31], op_17[31], op_17[31], op_17[31], op_17[31], op_17[31], op_17[31], op_17[31], op_17[31], op_17[31], op_17[31], op_17[31], op_17[31], op_17[31], op_17 };
assign grp_fu_967_p0 = { select_ln353_1_reg_1493[31], select_ln353_1_reg_1493, 2'h0 };
assign grp_fu_967_p1 = { op_18[7], op_18[7], op_18[7], op_18[7], op_18[7], op_18[7], op_18[7], op_18[7], op_18[7], op_18[7], op_18[7], op_18[7], op_18[7], op_18[7], op_18[7], op_18[7], op_18[7], op_18[7], op_18[7], op_18[7], op_18[7], op_18[7], op_18[7], op_18[7], op_18[7], op_18[7], op_18[7], op_18 };
assign lhs_fu_497_p3 = { op_7, 3'h0 };
assign op_30 = grp_fu_1025_p2;
assign or_ln_fu_637_p4 = { tmp_5_reg_1279, 1'h0, p_Result_s_20_reg_1285 };
assign p_Result_1_fu_563_p3 = ret_V_19_reg_1231[8];
assign p_Result_2_fu_479_p3 = ret_V_21_reg_1152[10];
assign p_Result_5_fu_529_p3 = ret_V_23_reg_1168[11];
assign p_Result_6_fu_770_p3 = ret_V_25_reg_1362[19];
assign p_Result_7_fu_868_p3 = ret_V_27_reg_1439[36];
assign p_Result_8_fu_933_p3 = ret_V_28_reg_1476[56];
assign p_Result_9_fu_998_p3 = ret_V_29_reg_1513[34];
assign p_Result_s_fu_318_p3 = r_V_reg_1057[9];
assign p_Val2_5_fu_692_p2 = { r_reg_1268[1:0], 2'h0 };
assign rhs_2_fu_376_p3 = { ret_V_18_reg_1095, 3'h0 };
assign rhs_4_fu_402_p3 = { op_8_V_reg_1112, 3'h0 };
assign rhs_8_fu_891_p3 = { select_ln353_reg_1456, 24'h000000 };
assign rhs_9_fu_956_p3 = { select_ln353_1_reg_1493, 2'h0 };
assign sext_ln1193_fu_373_p0 = op_3;
assign sext_ln1349_fu_349_p1 = { op_2_V_reg_1084[1], op_2_V_reg_1084[1], op_2_V_reg_1084[1], op_2_V_reg_1084[1], op_2_V_reg_1084[1], op_2_V_reg_1084[1], op_2_V_reg_1084 };
assign sext_ln215_fu_337_p0 = op_1;
assign sext_ln546_1_fu_593_p1 = { trunc_ln546_reg_1253[2], trunc_ln546_reg_1253 };
assign sext_ln546_2_fu_454_p1 = { ret_V_18_reg_1095[6], ret_V_18_reg_1095[6], ret_V_18_reg_1095[6], ret_V_18_reg_1095[6], ret_V_18_reg_1095[6], ret_V_18_reg_1095[6], ret_V_18_reg_1095[6], ret_V_18_reg_1095[6], ret_V_18_reg_1095[6], ret_V_18_reg_1095 };
assign sext_ln546_fu_441_p1 = { sh_V_1_reg_1163[7], sh_V_1_reg_1163[7], sh_V_1_reg_1163[7], sh_V_1_reg_1163[7], sh_V_1_reg_1163[7], sh_V_1_reg_1163[7], sh_V_1_reg_1163[7], sh_V_1_reg_1163[7], sh_V_1_reg_1163 };
assign sext_ln703_1_fu_399_p0 = op_3;
assign sext_ln703_2_fu_822_p0 = op_16;
assign sext_ln703_3_fu_887_p0 = op_17;
assign sext_ln703_4_fu_952_p0 = op_18;
assign sext_ln703_fu_509_p0 = op_9;
assign sext_ln781_fu_438_p1 = { ret_reg_1127[2], ret_reg_1127[2], ret_reg_1127[2], ret_reg_1127[2], ret_reg_1127[2], ret_reg_1127[2], ret_reg_1127[2], ret_reg_1127[2], ret_reg_1127[2], ret_reg_1127[2], ret_reg_1127[2], ret_reg_1127[2], ret_reg_1127[2], ret_reg_1127[2], ret_reg_1127[2], ret_reg_1127[2], ret_reg_1127[2], ret_reg_1127[2], ret_reg_1127[2], ret_reg_1127[2], ret_reg_1127[2], ret_reg_1127[2], ret_reg_1127[2], ret_reg_1127[2], ret_reg_1127[2], ret_reg_1127[2], ret_reg_1127[2], ret_reg_1127[2], ret_reg_1127[2], ret_reg_1127 };
assign sext_ln850_fu_761_p1 = { tmp_1_reg_1367[17], tmp_1_reg_1367 };
assign tmp_8_fu_826_p3 = { op_26_V_reg_1419, 4'h0 };
assign tmp_fu_472_p3 = ret_V_21_reg_1152[3];
assign trunc_ln1349_fu_352_p1 = op_4[7:0];
assign trunc_ln546_fu_582_p1 = grp_fu_448_p2[2:0];
assign trunc_ln769_fu_586_p1 = grp_fu_461_p2[3:0];
assign trunc_ln851_1_fu_519_p0 = op_9;
assign trunc_ln851_1_fu_519_p1 = op_9[2:0];
assign trunc_ln851_2_fu_419_p1 = grp_fu_387_p2[2:0];
assign trunc_ln851_3_fu_275_p0 = op_3;
assign trunc_ln851_3_fu_275_p1 = op_3[2:0];
assign trunc_ln851_4_fu_726_p1 = op_12_V_fu_718_p3[1:0];
assign trunc_ln851_5_fu_843_p0 = op_16;
assign trunc_ln851_5_fu_843_p1 = op_16[3:0];
assign trunc_ln851_6_fu_908_p0 = op_17;
assign trunc_ln851_6_fu_908_p1 = op_17[23:0];
assign trunc_ln851_7_fu_973_p0 = op_18;
assign trunc_ln851_7_fu_973_p1 = op_18[1:0];
assign trunc_ln851_fu_295_p1 = grp_fu_269_p2[2:0];
assign \sub_8ns_8s_8_2_1_U6.top_sub_8ns_8s_8_2_1_Adder_4_U.ain_s0  = \sub_8ns_8s_8_2_1_U6.top_sub_8ns_8s_8_2_1_Adder_4_U.a ;
assign \sub_8ns_8s_8_2_1_U6.top_sub_8ns_8s_8_2_1_Adder_4_U.s  = { \sub_8ns_8s_8_2_1_U6.top_sub_8ns_8s_8_2_1_Adder_4_U.fas_s2 , \sub_8ns_8s_8_2_1_U6.top_sub_8ns_8s_8_2_1_Adder_4_U.sum_s1  };
assign \sub_8ns_8s_8_2_1_U6.top_sub_8ns_8s_8_2_1_Adder_4_U.u2.a  = \sub_8ns_8s_8_2_1_U6.top_sub_8ns_8s_8_2_1_Adder_4_U.ain_s1 ;
assign \sub_8ns_8s_8_2_1_U6.top_sub_8ns_8s_8_2_1_Adder_4_U.u2.b  = \sub_8ns_8s_8_2_1_U6.top_sub_8ns_8s_8_2_1_Adder_4_U.bin_s1 ;
assign \sub_8ns_8s_8_2_1_U6.top_sub_8ns_8s_8_2_1_Adder_4_U.u2.cin  = \sub_8ns_8s_8_2_1_U6.top_sub_8ns_8s_8_2_1_Adder_4_U.carry_s1 ;
assign \sub_8ns_8s_8_2_1_U6.top_sub_8ns_8s_8_2_1_Adder_4_U.facout_s2  = \sub_8ns_8s_8_2_1_U6.top_sub_8ns_8s_8_2_1_Adder_4_U.u2.cout ;
assign \sub_8ns_8s_8_2_1_U6.top_sub_8ns_8s_8_2_1_Adder_4_U.fas_s2  = \sub_8ns_8s_8_2_1_U6.top_sub_8ns_8s_8_2_1_Adder_4_U.u2.s ;
assign \sub_8ns_8s_8_2_1_U6.top_sub_8ns_8s_8_2_1_Adder_4_U.u1.a  = \sub_8ns_8s_8_2_1_U6.top_sub_8ns_8s_8_2_1_Adder_4_U.a [3:0];
assign \sub_8ns_8s_8_2_1_U6.top_sub_8ns_8s_8_2_1_Adder_4_U.u1.b  = \sub_8ns_8s_8_2_1_U6.top_sub_8ns_8s_8_2_1_Adder_4_U.bin_s0 [3:0];
assign \sub_8ns_8s_8_2_1_U6.top_sub_8ns_8s_8_2_1_Adder_4_U.u1.cin  = 1'h1;
assign \sub_8ns_8s_8_2_1_U6.top_sub_8ns_8s_8_2_1_Adder_4_U.facout_s1  = \sub_8ns_8s_8_2_1_U6.top_sub_8ns_8s_8_2_1_Adder_4_U.u1.cout ;
assign \sub_8ns_8s_8_2_1_U6.top_sub_8ns_8s_8_2_1_Adder_4_U.fas_s1  = \sub_8ns_8s_8_2_1_U6.top_sub_8ns_8s_8_2_1_Adder_4_U.u1.s ;
assign \sub_8ns_8s_8_2_1_U6.top_sub_8ns_8s_8_2_1_Adder_4_U.a  = \sub_8ns_8s_8_2_1_U6.din0 ;
assign \sub_8ns_8s_8_2_1_U6.top_sub_8ns_8s_8_2_1_Adder_4_U.b  = \sub_8ns_8s_8_2_1_U6.din1 ;
assign \sub_8ns_8s_8_2_1_U6.top_sub_8ns_8s_8_2_1_Adder_4_U.ce  = \sub_8ns_8s_8_2_1_U6.ce ;
assign \sub_8ns_8s_8_2_1_U6.top_sub_8ns_8s_8_2_1_Adder_4_U.clk  = \sub_8ns_8s_8_2_1_U6.clk ;
assign \sub_8ns_8s_8_2_1_U6.top_sub_8ns_8s_8_2_1_Adder_4_U.reset  = \sub_8ns_8s_8_2_1_U6.reset ;
assign \sub_8ns_8s_8_2_1_U6.dout  = \sub_8ns_8s_8_2_1_U6.top_sub_8ns_8s_8_2_1_Adder_4_U.s ;
assign \sub_8ns_8s_8_2_1_U6.ce  = 1'h1;
assign \sub_8ns_8s_8_2_1_U6.clk  = ap_clk;
assign \sub_8ns_8s_8_2_1_U6.din0  = 8'h00;
assign \sub_8ns_8s_8_2_1_U6.din1  = { ret_V_18_reg_1095[6], ret_V_18_reg_1095 };
assign grp_fu_393_p2 = \sub_8ns_8s_8_2_1_U6.dout ;
assign \sub_8ns_8s_8_2_1_U6.reset  = ap_rst;
assign \sub_11s_11s_11_2_1_U5.top_sub_11s_11s_11_2_1_Adder_3_U.ain_s0  = \sub_11s_11s_11_2_1_U5.top_sub_11s_11s_11_2_1_Adder_3_U.a ;
assign \sub_11s_11s_11_2_1_U5.top_sub_11s_11s_11_2_1_Adder_3_U.s  = { \sub_11s_11s_11_2_1_U5.top_sub_11s_11s_11_2_1_Adder_3_U.fas_s2 , \sub_11s_11s_11_2_1_U5.top_sub_11s_11s_11_2_1_Adder_3_U.sum_s1  };
assign \sub_11s_11s_11_2_1_U5.top_sub_11s_11s_11_2_1_Adder_3_U.u2.a  = \sub_11s_11s_11_2_1_U5.top_sub_11s_11s_11_2_1_Adder_3_U.ain_s1 ;
assign \sub_11s_11s_11_2_1_U5.top_sub_11s_11s_11_2_1_Adder_3_U.u2.b  = \sub_11s_11s_11_2_1_U5.top_sub_11s_11s_11_2_1_Adder_3_U.bin_s1 ;
assign \sub_11s_11s_11_2_1_U5.top_sub_11s_11s_11_2_1_Adder_3_U.u2.cin  = \sub_11s_11s_11_2_1_U5.top_sub_11s_11s_11_2_1_Adder_3_U.carry_s1 ;
assign \sub_11s_11s_11_2_1_U5.top_sub_11s_11s_11_2_1_Adder_3_U.facout_s2  = \sub_11s_11s_11_2_1_U5.top_sub_11s_11s_11_2_1_Adder_3_U.u2.cout ;
assign \sub_11s_11s_11_2_1_U5.top_sub_11s_11s_11_2_1_Adder_3_U.fas_s2  = \sub_11s_11s_11_2_1_U5.top_sub_11s_11s_11_2_1_Adder_3_U.u2.s ;
assign \sub_11s_11s_11_2_1_U5.top_sub_11s_11s_11_2_1_Adder_3_U.u1.a  = \sub_11s_11s_11_2_1_U5.top_sub_11s_11s_11_2_1_Adder_3_U.a [4:0];
assign \sub_11s_11s_11_2_1_U5.top_sub_11s_11s_11_2_1_Adder_3_U.u1.b  = \sub_11s_11s_11_2_1_U5.top_sub_11s_11s_11_2_1_Adder_3_U.bin_s0 [4:0];
assign \sub_11s_11s_11_2_1_U5.top_sub_11s_11s_11_2_1_Adder_3_U.u1.cin  = 1'h1;
assign \sub_11s_11s_11_2_1_U5.top_sub_11s_11s_11_2_1_Adder_3_U.facout_s1  = \sub_11s_11s_11_2_1_U5.top_sub_11s_11s_11_2_1_Adder_3_U.u1.cout ;
assign \sub_11s_11s_11_2_1_U5.top_sub_11s_11s_11_2_1_Adder_3_U.fas_s1  = \sub_11s_11s_11_2_1_U5.top_sub_11s_11s_11_2_1_Adder_3_U.u1.s ;
assign \sub_11s_11s_11_2_1_U5.top_sub_11s_11s_11_2_1_Adder_3_U.a  = \sub_11s_11s_11_2_1_U5.din0 ;
assign \sub_11s_11s_11_2_1_U5.top_sub_11s_11s_11_2_1_Adder_3_U.b  = \sub_11s_11s_11_2_1_U5.din1 ;
assign \sub_11s_11s_11_2_1_U5.top_sub_11s_11s_11_2_1_Adder_3_U.ce  = \sub_11s_11s_11_2_1_U5.ce ;
assign \sub_11s_11s_11_2_1_U5.top_sub_11s_11s_11_2_1_Adder_3_U.clk  = \sub_11s_11s_11_2_1_U5.clk ;
assign \sub_11s_11s_11_2_1_U5.top_sub_11s_11s_11_2_1_Adder_3_U.reset  = \sub_11s_11s_11_2_1_U5.reset ;
assign \sub_11s_11s_11_2_1_U5.dout  = \sub_11s_11s_11_2_1_U5.top_sub_11s_11s_11_2_1_Adder_3_U.s ;
assign \sub_11s_11s_11_2_1_U5.ce  = 1'h1;
assign \sub_11s_11s_11_2_1_U5.clk  = ap_clk;
assign \sub_11s_11s_11_2_1_U5.din0  = { op_3[7], op_3[7], op_3[7], op_3 };
assign \sub_11s_11s_11_2_1_U5.din1  = { ret_V_18_reg_1095[6], ret_V_18_reg_1095, 3'h0 };
assign grp_fu_387_p2 = \sub_11s_11s_11_2_1_U5.dout ;
assign \sub_11s_11s_11_2_1_U5.reset  = ap_rst;
assign \shl_32s_16ns_32_7_1_U9.din1_cast  = \shl_32s_16ns_32_7_1_U9.din1 [15:0];
assign \shl_32s_16ns_32_7_1_U9.din1_mask  = 16'h0007;
assign \shl_32s_16ns_32_7_1_U9.ce  = 1'h1;
assign \shl_32s_16ns_32_7_1_U9.clk  = ap_clk;
assign \shl_32s_16ns_32_7_1_U9.din0  = { ret_reg_1127[2], ret_reg_1127[2], ret_reg_1127[2], ret_reg_1127[2], ret_reg_1127[2], ret_reg_1127[2], ret_reg_1127[2], ret_reg_1127[2], ret_reg_1127[2], ret_reg_1127[2], ret_reg_1127[2], ret_reg_1127[2], ret_reg_1127[2], ret_reg_1127[2], ret_reg_1127[2], ret_reg_1127[2], ret_reg_1127[2], ret_reg_1127[2], ret_reg_1127[2], ret_reg_1127[2], ret_reg_1127[2], ret_reg_1127[2], ret_reg_1127[2], ret_reg_1127[2], ret_reg_1127[2], ret_reg_1127[2], ret_reg_1127[2], ret_reg_1127[2], ret_reg_1127[2], ret_reg_1127 };
assign \shl_32s_16ns_32_7_1_U9.din1  = { 16'h0000, ret_V_18_reg_1095[6], ret_V_18_reg_1095[6], ret_V_18_reg_1095[6], ret_V_18_reg_1095[6], ret_V_18_reg_1095[6], ret_V_18_reg_1095[6], ret_V_18_reg_1095[6], ret_V_18_reg_1095[6], ret_V_18_reg_1095[6], ret_V_18_reg_1095 };
assign grp_fu_461_p2 = \shl_32s_16ns_32_7_1_U9.dout ;
assign \shl_32s_16ns_32_7_1_U9.reset  = ap_rst;
assign \mul_8s_2s_10_7_1_U1.top_mul_8s_2s_10_7_1_Mul_DSP_0_U.p  = \mul_8s_2s_10_7_1_U1.top_mul_8s_2s_10_7_1_Mul_DSP_0_U.buff4 ;
assign \mul_8s_2s_10_7_1_U1.top_mul_8s_2s_10_7_1_Mul_DSP_0_U.a  = \mul_8s_2s_10_7_1_U1.din0 ;
assign \mul_8s_2s_10_7_1_U1.top_mul_8s_2s_10_7_1_Mul_DSP_0_U.b  = \mul_8s_2s_10_7_1_U1.din1 ;
assign \mul_8s_2s_10_7_1_U1.top_mul_8s_2s_10_7_1_Mul_DSP_0_U.ce  = \mul_8s_2s_10_7_1_U1.ce ;
assign \mul_8s_2s_10_7_1_U1.top_mul_8s_2s_10_7_1_Mul_DSP_0_U.clk  = \mul_8s_2s_10_7_1_U1.clk ;
assign \mul_8s_2s_10_7_1_U1.dout  = \mul_8s_2s_10_7_1_U1.top_mul_8s_2s_10_7_1_Mul_DSP_0_U.p ;
assign \mul_8s_2s_10_7_1_U1.ce  = 1'h1;
assign \mul_8s_2s_10_7_1_U1.clk  = ap_clk;
assign \mul_8s_2s_10_7_1_U1.din0  = op_3;
assign \mul_8s_2s_10_7_1_U1.din1  = op_1;
assign grp_fu_269_p2 = \mul_8s_2s_10_7_1_U1.dout ;
assign \mul_8s_2s_10_7_1_U1.reset  = ap_rst;
assign \ashr_32s_16ns_32_7_1_U8.din1_cast  = \ashr_32s_16ns_32_7_1_U8.din1 [15:0];
assign \ashr_32s_16ns_32_7_1_U8.din1_mask  = 16'h0007;
assign \ashr_32s_16ns_32_7_1_U8.ce  = 1'h1;
assign \ashr_32s_16ns_32_7_1_U8.clk  = ap_clk;
assign \ashr_32s_16ns_32_7_1_U8.din0  = { ret_reg_1127[2], ret_reg_1127[2], ret_reg_1127[2], ret_reg_1127[2], ret_reg_1127[2], ret_reg_1127[2], ret_reg_1127[2], ret_reg_1127[2], ret_reg_1127[2], ret_reg_1127[2], ret_reg_1127[2], ret_reg_1127[2], ret_reg_1127[2], ret_reg_1127[2], ret_reg_1127[2], ret_reg_1127[2], ret_reg_1127[2], ret_reg_1127[2], ret_reg_1127[2], ret_reg_1127[2], ret_reg_1127[2], ret_reg_1127[2], ret_reg_1127[2], ret_reg_1127[2], ret_reg_1127[2], ret_reg_1127[2], ret_reg_1127[2], ret_reg_1127[2], ret_reg_1127[2], ret_reg_1127 };
assign \ashr_32s_16ns_32_7_1_U8.din1  = { 16'h0000, sh_V_1_reg_1163[7], sh_V_1_reg_1163[7], sh_V_1_reg_1163[7], sh_V_1_reg_1163[7], sh_V_1_reg_1163[7], sh_V_1_reg_1163[7], sh_V_1_reg_1163[7], sh_V_1_reg_1163[7], sh_V_1_reg_1163 };
assign grp_fu_448_p2 = \ashr_32s_16ns_32_7_1_U8.dout ;
assign \ashr_32s_16ns_32_7_1_U8.reset  = ap_rst;
assign \add_9ns_9s_9_2_1_U11.top_add_9ns_9s_9_2_1_Adder_7_U.ain_s0  = \add_9ns_9s_9_2_1_U11.top_add_9ns_9s_9_2_1_Adder_7_U.a ;
assign \add_9ns_9s_9_2_1_U11.top_add_9ns_9s_9_2_1_Adder_7_U.bin_s0  = \add_9ns_9s_9_2_1_U11.top_add_9ns_9s_9_2_1_Adder_7_U.b ;
assign \add_9ns_9s_9_2_1_U11.top_add_9ns_9s_9_2_1_Adder_7_U.s  = { \add_9ns_9s_9_2_1_U11.top_add_9ns_9s_9_2_1_Adder_7_U.fas_s2 , \add_9ns_9s_9_2_1_U11.top_add_9ns_9s_9_2_1_Adder_7_U.sum_s1  };
assign \add_9ns_9s_9_2_1_U11.top_add_9ns_9s_9_2_1_Adder_7_U.u2.a  = \add_9ns_9s_9_2_1_U11.top_add_9ns_9s_9_2_1_Adder_7_U.ain_s1 ;
assign \add_9ns_9s_9_2_1_U11.top_add_9ns_9s_9_2_1_Adder_7_U.u2.b  = \add_9ns_9s_9_2_1_U11.top_add_9ns_9s_9_2_1_Adder_7_U.bin_s1 ;
assign \add_9ns_9s_9_2_1_U11.top_add_9ns_9s_9_2_1_Adder_7_U.u2.cin  = \add_9ns_9s_9_2_1_U11.top_add_9ns_9s_9_2_1_Adder_7_U.carry_s1 ;
assign \add_9ns_9s_9_2_1_U11.top_add_9ns_9s_9_2_1_Adder_7_U.facout_s2  = \add_9ns_9s_9_2_1_U11.top_add_9ns_9s_9_2_1_Adder_7_U.u2.cout ;
assign \add_9ns_9s_9_2_1_U11.top_add_9ns_9s_9_2_1_Adder_7_U.fas_s2  = \add_9ns_9s_9_2_1_U11.top_add_9ns_9s_9_2_1_Adder_7_U.u2.s ;
assign \add_9ns_9s_9_2_1_U11.top_add_9ns_9s_9_2_1_Adder_7_U.u1.a  = \add_9ns_9s_9_2_1_U11.top_add_9ns_9s_9_2_1_Adder_7_U.a [3:0];
assign \add_9ns_9s_9_2_1_U11.top_add_9ns_9s_9_2_1_Adder_7_U.u1.b  = \add_9ns_9s_9_2_1_U11.top_add_9ns_9s_9_2_1_Adder_7_U.b [3:0];
assign \add_9ns_9s_9_2_1_U11.top_add_9ns_9s_9_2_1_Adder_7_U.u1.cin  = 1'h0;
assign \add_9ns_9s_9_2_1_U11.top_add_9ns_9s_9_2_1_Adder_7_U.facout_s1  = \add_9ns_9s_9_2_1_U11.top_add_9ns_9s_9_2_1_Adder_7_U.u1.cout ;
assign \add_9ns_9s_9_2_1_U11.top_add_9ns_9s_9_2_1_Adder_7_U.fas_s1  = \add_9ns_9s_9_2_1_U11.top_add_9ns_9s_9_2_1_Adder_7_U.u1.s ;
assign \add_9ns_9s_9_2_1_U11.top_add_9ns_9s_9_2_1_Adder_7_U.a  = \add_9ns_9s_9_2_1_U11.din0 ;
assign \add_9ns_9s_9_2_1_U11.top_add_9ns_9s_9_2_1_Adder_7_U.b  = \add_9ns_9s_9_2_1_U11.din1 ;
assign \add_9ns_9s_9_2_1_U11.top_add_9ns_9s_9_2_1_Adder_7_U.ce  = \add_9ns_9s_9_2_1_U11.ce ;
assign \add_9ns_9s_9_2_1_U11.top_add_9ns_9s_9_2_1_Adder_7_U.clk  = \add_9ns_9s_9_2_1_U11.clk ;
assign \add_9ns_9s_9_2_1_U11.top_add_9ns_9s_9_2_1_Adder_7_U.reset  = \add_9ns_9s_9_2_1_U11.reset ;
assign \add_9ns_9s_9_2_1_U11.dout  = \add_9ns_9s_9_2_1_U11.top_add_9ns_9s_9_2_1_Adder_7_U.s ;
assign \add_9ns_9s_9_2_1_U11.ce  = 1'h1;
assign \add_9ns_9s_9_2_1_U11.clk  = ap_clk;
assign \add_9ns_9s_9_2_1_U11.din0  = { 2'h0, op_7, 3'h0 };
assign \add_9ns_9s_9_2_1_U11.din1  = { op_9[7], op_9 };
assign grp_fu_513_p2 = \add_9ns_9s_9_2_1_U11.dout ;
assign \add_9ns_9s_9_2_1_U11.reset  = ap_rst;
assign \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_9_U.ain_s0  = \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_9_U.a ;
assign \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_9_U.bin_s0  = \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_9_U.b ;
assign \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_9_U.s  = { \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_9_U.fas_s2 , \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_9_U.sum_s1  };
assign \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_9_U.u2.a  = \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_9_U.ain_s1 ;
assign \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_9_U.u2.b  = \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_9_U.bin_s1 ;
assign \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_9_U.u2.cin  = \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_9_U.carry_s1 ;
assign \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_9_U.facout_s2  = \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_9_U.u2.cout ;
assign \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_9_U.fas_s2  = \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_9_U.u2.s ;
assign \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_9_U.u1.a  = \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_9_U.a [2:0];
assign \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_9_U.u1.b  = \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_9_U.b [2:0];
assign \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_9_U.u1.cin  = 1'h0;
assign \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_9_U.facout_s1  = \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_9_U.u1.cout ;
assign \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_9_U.fas_s1  = \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_9_U.u1.s ;
assign \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_9_U.a  = \add_7s_7s_7_2_1_U13.din0 ;
assign \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_9_U.b  = \add_7s_7s_7_2_1_U13.din1 ;
assign \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_9_U.ce  = \add_7s_7s_7_2_1_U13.ce ;
assign \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_9_U.clk  = \add_7s_7s_7_2_1_U13.clk ;
assign \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_9_U.reset  = \add_7s_7s_7_2_1_U13.reset ;
assign \add_7s_7s_7_2_1_U13.dout  = \add_7s_7s_7_2_1_U13.top_add_7s_7s_7_2_1_Adder_9_U.s ;
assign \add_7s_7s_7_2_1_U13.ce  = 1'h1;
assign \add_7s_7s_7_2_1_U13.clk  = ap_clk;
assign \add_7s_7s_7_2_1_U13.din0  = { ret_V_20_reg_1248[5], ret_V_20_reg_1248 };
assign \add_7s_7s_7_2_1_U13.din1  = { ret_V_24_reg_1226[1], ret_V_24_reg_1226[1], ret_V_24_reg_1226[1], ret_V_24_reg_1226[1], ret_V_24_reg_1226[1], ret_V_24_reg_1226 };
assign grp_fu_631_p2 = \add_7s_7s_7_2_1_U13.dout ;
assign \add_7s_7s_7_2_1_U13.reset  = ap_rst;
assign \add_7ns_7ns_7_2_1_U3.top_add_7ns_7ns_7_2_1_Adder_1_U.ain_s0  = \add_7ns_7ns_7_2_1_U3.top_add_7ns_7ns_7_2_1_Adder_1_U.a ;
assign \add_7ns_7ns_7_2_1_U3.top_add_7ns_7ns_7_2_1_Adder_1_U.bin_s0  = \add_7ns_7ns_7_2_1_U3.top_add_7ns_7ns_7_2_1_Adder_1_U.b ;
assign \add_7ns_7ns_7_2_1_U3.top_add_7ns_7ns_7_2_1_Adder_1_U.s  = { \add_7ns_7ns_7_2_1_U3.top_add_7ns_7ns_7_2_1_Adder_1_U.fas_s2 , \add_7ns_7ns_7_2_1_U3.top_add_7ns_7ns_7_2_1_Adder_1_U.sum_s1  };
assign \add_7ns_7ns_7_2_1_U3.top_add_7ns_7ns_7_2_1_Adder_1_U.u2.a  = \add_7ns_7ns_7_2_1_U3.top_add_7ns_7ns_7_2_1_Adder_1_U.ain_s1 ;
assign \add_7ns_7ns_7_2_1_U3.top_add_7ns_7ns_7_2_1_Adder_1_U.u2.b  = \add_7ns_7ns_7_2_1_U3.top_add_7ns_7ns_7_2_1_Adder_1_U.bin_s1 ;
assign \add_7ns_7ns_7_2_1_U3.top_add_7ns_7ns_7_2_1_Adder_1_U.u2.cin  = \add_7ns_7ns_7_2_1_U3.top_add_7ns_7ns_7_2_1_Adder_1_U.carry_s1 ;
assign \add_7ns_7ns_7_2_1_U3.top_add_7ns_7ns_7_2_1_Adder_1_U.facout_s2  = \add_7ns_7ns_7_2_1_U3.top_add_7ns_7ns_7_2_1_Adder_1_U.u2.cout ;
assign \add_7ns_7ns_7_2_1_U3.top_add_7ns_7ns_7_2_1_Adder_1_U.fas_s2  = \add_7ns_7ns_7_2_1_U3.top_add_7ns_7ns_7_2_1_Adder_1_U.u2.s ;
assign \add_7ns_7ns_7_2_1_U3.top_add_7ns_7ns_7_2_1_Adder_1_U.u1.a  = \add_7ns_7ns_7_2_1_U3.top_add_7ns_7ns_7_2_1_Adder_1_U.a [2:0];
assign \add_7ns_7ns_7_2_1_U3.top_add_7ns_7ns_7_2_1_Adder_1_U.u1.b  = \add_7ns_7ns_7_2_1_U3.top_add_7ns_7ns_7_2_1_Adder_1_U.b [2:0];
assign \add_7ns_7ns_7_2_1_U3.top_add_7ns_7ns_7_2_1_Adder_1_U.u1.cin  = 1'h0;
assign \add_7ns_7ns_7_2_1_U3.top_add_7ns_7ns_7_2_1_Adder_1_U.facout_s1  = \add_7ns_7ns_7_2_1_U3.top_add_7ns_7ns_7_2_1_Adder_1_U.u1.cout ;
assign \add_7ns_7ns_7_2_1_U3.top_add_7ns_7ns_7_2_1_Adder_1_U.fas_s1  = \add_7ns_7ns_7_2_1_U3.top_add_7ns_7ns_7_2_1_Adder_1_U.u1.s ;
assign \add_7ns_7ns_7_2_1_U3.top_add_7ns_7ns_7_2_1_Adder_1_U.a  = \add_7ns_7ns_7_2_1_U3.din0 ;
assign \add_7ns_7ns_7_2_1_U3.top_add_7ns_7ns_7_2_1_Adder_1_U.b  = \add_7ns_7ns_7_2_1_U3.din1 ;
assign \add_7ns_7ns_7_2_1_U3.top_add_7ns_7ns_7_2_1_Adder_1_U.ce  = \add_7ns_7ns_7_2_1_U3.ce ;
assign \add_7ns_7ns_7_2_1_U3.top_add_7ns_7ns_7_2_1_Adder_1_U.clk  = \add_7ns_7ns_7_2_1_U3.clk ;
assign \add_7ns_7ns_7_2_1_U3.top_add_7ns_7ns_7_2_1_Adder_1_U.reset  = \add_7ns_7ns_7_2_1_U3.reset ;
assign \add_7ns_7ns_7_2_1_U3.dout  = \add_7ns_7ns_7_2_1_U3.top_add_7ns_7ns_7_2_1_Adder_1_U.s ;
assign \add_7ns_7ns_7_2_1_U3.ce  = 1'h1;
assign \add_7ns_7ns_7_2_1_U3.clk  = ap_clk;
assign \add_7ns_7ns_7_2_1_U3.din0  = ret_V_reg_1062;
assign \add_7ns_7ns_7_2_1_U3.din1  = 7'h01;
assign grp_fu_313_p2 = \add_7ns_7ns_7_2_1_U3.dout ;
assign \add_7ns_7ns_7_2_1_U3.reset  = ap_rst;
assign \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_8_U.ain_s0  = \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_8_U.a ;
assign \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_8_U.bin_s0  = \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_8_U.b ;
assign \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_8_U.s  = { \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_8_U.fas_s2 , \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_8_U.sum_s1  };
assign \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_8_U.u2.a  = \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_8_U.ain_s1 ;
assign \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_8_U.u2.b  = \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_8_U.bin_s1 ;
assign \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_8_U.u2.cin  = \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_8_U.carry_s1 ;
assign \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_8_U.facout_s2  = \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_8_U.u2.cout ;
assign \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_8_U.fas_s2  = \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_8_U.u2.s ;
assign \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_8_U.u1.a  = \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_8_U.a [2:0];
assign \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_8_U.u1.b  = \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_8_U.b [2:0];
assign \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_8_U.u1.cin  = 1'h0;
assign \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_8_U.facout_s1  = \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_8_U.u1.cout ;
assign \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_8_U.fas_s1  = \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_8_U.u1.s ;
assign \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_8_U.a  = \add_6ns_6ns_6_2_1_U12.din0 ;
assign \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_8_U.b  = \add_6ns_6ns_6_2_1_U12.din1 ;
assign \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_8_U.ce  = \add_6ns_6ns_6_2_1_U12.ce ;
assign \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_8_U.clk  = \add_6ns_6ns_6_2_1_U12.clk ;
assign \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_8_U.reset  = \add_6ns_6ns_6_2_1_U12.reset ;
assign \add_6ns_6ns_6_2_1_U12.dout  = \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_8_U.s ;
assign \add_6ns_6ns_6_2_1_U12.ce  = 1'h1;
assign \add_6ns_6ns_6_2_1_U12.clk  = ap_clk;
assign \add_6ns_6ns_6_2_1_U12.din0  = ret_V_4_reg_1236;
assign \add_6ns_6ns_6_2_1_U12.din1  = 6'h01;
assign grp_fu_558_p2 = \add_6ns_6ns_6_2_1_U12.dout ;
assign \add_6ns_6ns_6_2_1_U12.reset  = ap_rst;
assign \add_57s_57s_57_2_1_U22.top_add_57s_57s_57_2_1_Adder_16_U.ain_s0  = \add_57s_57s_57_2_1_U22.top_add_57s_57s_57_2_1_Adder_16_U.a ;
assign \add_57s_57s_57_2_1_U22.top_add_57s_57s_57_2_1_Adder_16_U.bin_s0  = \add_57s_57s_57_2_1_U22.top_add_57s_57s_57_2_1_Adder_16_U.b ;
assign \add_57s_57s_57_2_1_U22.top_add_57s_57s_57_2_1_Adder_16_U.s  = { \add_57s_57s_57_2_1_U22.top_add_57s_57s_57_2_1_Adder_16_U.fas_s2 , \add_57s_57s_57_2_1_U22.top_add_57s_57s_57_2_1_Adder_16_U.sum_s1  };
assign \add_57s_57s_57_2_1_U22.top_add_57s_57s_57_2_1_Adder_16_U.u2.a  = \add_57s_57s_57_2_1_U22.top_add_57s_57s_57_2_1_Adder_16_U.ain_s1 ;
assign \add_57s_57s_57_2_1_U22.top_add_57s_57s_57_2_1_Adder_16_U.u2.b  = \add_57s_57s_57_2_1_U22.top_add_57s_57s_57_2_1_Adder_16_U.bin_s1 ;
assign \add_57s_57s_57_2_1_U22.top_add_57s_57s_57_2_1_Adder_16_U.u2.cin  = \add_57s_57s_57_2_1_U22.top_add_57s_57s_57_2_1_Adder_16_U.carry_s1 ;
assign \add_57s_57s_57_2_1_U22.top_add_57s_57s_57_2_1_Adder_16_U.facout_s2  = \add_57s_57s_57_2_1_U22.top_add_57s_57s_57_2_1_Adder_16_U.u2.cout ;
assign \add_57s_57s_57_2_1_U22.top_add_57s_57s_57_2_1_Adder_16_U.fas_s2  = \add_57s_57s_57_2_1_U22.top_add_57s_57s_57_2_1_Adder_16_U.u2.s ;
assign \add_57s_57s_57_2_1_U22.top_add_57s_57s_57_2_1_Adder_16_U.u1.a  = \add_57s_57s_57_2_1_U22.top_add_57s_57s_57_2_1_Adder_16_U.a [27:0];
assign \add_57s_57s_57_2_1_U22.top_add_57s_57s_57_2_1_Adder_16_U.u1.b  = \add_57s_57s_57_2_1_U22.top_add_57s_57s_57_2_1_Adder_16_U.b [27:0];
assign \add_57s_57s_57_2_1_U22.top_add_57s_57s_57_2_1_Adder_16_U.u1.cin  = 1'h0;
assign \add_57s_57s_57_2_1_U22.top_add_57s_57s_57_2_1_Adder_16_U.facout_s1  = \add_57s_57s_57_2_1_U22.top_add_57s_57s_57_2_1_Adder_16_U.u1.cout ;
assign \add_57s_57s_57_2_1_U22.top_add_57s_57s_57_2_1_Adder_16_U.fas_s1  = \add_57s_57s_57_2_1_U22.top_add_57s_57s_57_2_1_Adder_16_U.u1.s ;
assign \add_57s_57s_57_2_1_U22.top_add_57s_57s_57_2_1_Adder_16_U.a  = \add_57s_57s_57_2_1_U22.din0 ;
assign \add_57s_57s_57_2_1_U22.top_add_57s_57s_57_2_1_Adder_16_U.b  = \add_57s_57s_57_2_1_U22.din1 ;
assign \add_57s_57s_57_2_1_U22.top_add_57s_57s_57_2_1_Adder_16_U.ce  = \add_57s_57s_57_2_1_U22.ce ;
assign \add_57s_57s_57_2_1_U22.top_add_57s_57s_57_2_1_Adder_16_U.clk  = \add_57s_57s_57_2_1_U22.clk ;
assign \add_57s_57s_57_2_1_U22.top_add_57s_57s_57_2_1_Adder_16_U.reset  = \add_57s_57s_57_2_1_U22.reset ;
assign \add_57s_57s_57_2_1_U22.dout  = \add_57s_57s_57_2_1_U22.top_add_57s_57s_57_2_1_Adder_16_U.s ;
assign \add_57s_57s_57_2_1_U22.ce  = 1'h1;
assign \add_57s_57s_57_2_1_U22.clk  = ap_clk;
assign \add_57s_57s_57_2_1_U22.din0  = { select_ln353_reg_1456[31], select_ln353_reg_1456, 24'h000000 };
assign \add_57s_57s_57_2_1_U22.din1  = { op_17[31], op_17[31], op_17[31], op_17[31], op_17[31], op_17[31], op_17[31], op_17[31], op_17[31], op_17[31], op_17[31], op_17[31], op_17[31], op_17[31], op_17[31], op_17[31], op_17[31], op_17[31], op_17[31], op_17[31], op_17[31], op_17[31], op_17[31], op_17[31], op_17[31], op_17 };
assign grp_fu_902_p2 = \add_57s_57s_57_2_1_U22.dout ;
assign \add_57s_57s_57_2_1_U22.reset  = ap_rst;
assign \add_3s_3s_3_2_1_U4.top_add_3s_3s_3_2_1_Adder_2_U.ain_s0  = \add_3s_3s_3_2_1_U4.top_add_3s_3s_3_2_1_Adder_2_U.a ;
assign \add_3s_3s_3_2_1_U4.top_add_3s_3s_3_2_1_Adder_2_U.bin_s0  = \add_3s_3s_3_2_1_U4.top_add_3s_3s_3_2_1_Adder_2_U.b ;
assign \add_3s_3s_3_2_1_U4.top_add_3s_3s_3_2_1_Adder_2_U.s  = { \add_3s_3s_3_2_1_U4.top_add_3s_3s_3_2_1_Adder_2_U.fas_s2 , \add_3s_3s_3_2_1_U4.top_add_3s_3s_3_2_1_Adder_2_U.sum_s1  };
assign \add_3s_3s_3_2_1_U4.top_add_3s_3s_3_2_1_Adder_2_U.u2.a  = \add_3s_3s_3_2_1_U4.top_add_3s_3s_3_2_1_Adder_2_U.ain_s1 ;
assign \add_3s_3s_3_2_1_U4.top_add_3s_3s_3_2_1_Adder_2_U.u2.b  = \add_3s_3s_3_2_1_U4.top_add_3s_3s_3_2_1_Adder_2_U.bin_s1 ;
assign \add_3s_3s_3_2_1_U4.top_add_3s_3s_3_2_1_Adder_2_U.u2.cin  = \add_3s_3s_3_2_1_U4.top_add_3s_3s_3_2_1_Adder_2_U.carry_s1 ;
assign \add_3s_3s_3_2_1_U4.top_add_3s_3s_3_2_1_Adder_2_U.facout_s2  = \add_3s_3s_3_2_1_U4.top_add_3s_3s_3_2_1_Adder_2_U.u2.cout ;
assign \add_3s_3s_3_2_1_U4.top_add_3s_3s_3_2_1_Adder_2_U.fas_s2  = \add_3s_3s_3_2_1_U4.top_add_3s_3s_3_2_1_Adder_2_U.u2.s ;
assign \add_3s_3s_3_2_1_U4.top_add_3s_3s_3_2_1_Adder_2_U.u1.a  = \add_3s_3s_3_2_1_U4.top_add_3s_3s_3_2_1_Adder_2_U.a [0];
assign \add_3s_3s_3_2_1_U4.top_add_3s_3s_3_2_1_Adder_2_U.u1.b  = \add_3s_3s_3_2_1_U4.top_add_3s_3s_3_2_1_Adder_2_U.b [0];
assign \add_3s_3s_3_2_1_U4.top_add_3s_3s_3_2_1_Adder_2_U.u1.cin  = 1'h0;
assign \add_3s_3s_3_2_1_U4.top_add_3s_3s_3_2_1_Adder_2_U.facout_s1  = \add_3s_3s_3_2_1_U4.top_add_3s_3s_3_2_1_Adder_2_U.u1.cout ;
assign \add_3s_3s_3_2_1_U4.top_add_3s_3s_3_2_1_Adder_2_U.fas_s1  = \add_3s_3s_3_2_1_U4.top_add_3s_3s_3_2_1_Adder_2_U.u1.s ;
assign \add_3s_3s_3_2_1_U4.top_add_3s_3s_3_2_1_Adder_2_U.a  = \add_3s_3s_3_2_1_U4.din0 ;
assign \add_3s_3s_3_2_1_U4.top_add_3s_3s_3_2_1_Adder_2_U.b  = \add_3s_3s_3_2_1_U4.din1 ;
assign \add_3s_3s_3_2_1_U4.top_add_3s_3s_3_2_1_Adder_2_U.ce  = \add_3s_3s_3_2_1_U4.ce ;
assign \add_3s_3s_3_2_1_U4.top_add_3s_3s_3_2_1_Adder_2_U.clk  = \add_3s_3s_3_2_1_U4.clk ;
assign \add_3s_3s_3_2_1_U4.top_add_3s_3s_3_2_1_Adder_2_U.reset  = \add_3s_3s_3_2_1_U4.reset ;
assign \add_3s_3s_3_2_1_U4.dout  = \add_3s_3s_3_2_1_U4.top_add_3s_3s_3_2_1_Adder_2_U.s ;
assign \add_3s_3s_3_2_1_U4.ce  = 1'h1;
assign \add_3s_3s_3_2_1_U4.clk  = ap_clk;
assign \add_3s_3s_3_2_1_U4.din0  = { op_2_V_reg_1084[1], op_2_V_reg_1084 };
assign \add_3s_3s_3_2_1_U4.din1  = { op_1[1], op_1 };
assign grp_fu_343_p2 = \add_3s_3s_3_2_1_U4.dout ;
assign \add_3s_3s_3_2_1_U4.reset  = ap_rst;
assign \add_37s_37s_37_2_1_U20.top_add_37s_37s_37_2_1_Adder_14_U.ain_s0  = \add_37s_37s_37_2_1_U20.top_add_37s_37s_37_2_1_Adder_14_U.a ;
assign \add_37s_37s_37_2_1_U20.top_add_37s_37s_37_2_1_Adder_14_U.bin_s0  = \add_37s_37s_37_2_1_U20.top_add_37s_37s_37_2_1_Adder_14_U.b ;
assign \add_37s_37s_37_2_1_U20.top_add_37s_37s_37_2_1_Adder_14_U.s  = { \add_37s_37s_37_2_1_U20.top_add_37s_37s_37_2_1_Adder_14_U.fas_s2 , \add_37s_37s_37_2_1_U20.top_add_37s_37s_37_2_1_Adder_14_U.sum_s1  };
assign \add_37s_37s_37_2_1_U20.top_add_37s_37s_37_2_1_Adder_14_U.u2.a  = \add_37s_37s_37_2_1_U20.top_add_37s_37s_37_2_1_Adder_14_U.ain_s1 ;
assign \add_37s_37s_37_2_1_U20.top_add_37s_37s_37_2_1_Adder_14_U.u2.b  = \add_37s_37s_37_2_1_U20.top_add_37s_37s_37_2_1_Adder_14_U.bin_s1 ;
assign \add_37s_37s_37_2_1_U20.top_add_37s_37s_37_2_1_Adder_14_U.u2.cin  = \add_37s_37s_37_2_1_U20.top_add_37s_37s_37_2_1_Adder_14_U.carry_s1 ;
assign \add_37s_37s_37_2_1_U20.top_add_37s_37s_37_2_1_Adder_14_U.facout_s2  = \add_37s_37s_37_2_1_U20.top_add_37s_37s_37_2_1_Adder_14_U.u2.cout ;
assign \add_37s_37s_37_2_1_U20.top_add_37s_37s_37_2_1_Adder_14_U.fas_s2  = \add_37s_37s_37_2_1_U20.top_add_37s_37s_37_2_1_Adder_14_U.u2.s ;
assign \add_37s_37s_37_2_1_U20.top_add_37s_37s_37_2_1_Adder_14_U.u1.a  = \add_37s_37s_37_2_1_U20.top_add_37s_37s_37_2_1_Adder_14_U.a [17:0];
assign \add_37s_37s_37_2_1_U20.top_add_37s_37s_37_2_1_Adder_14_U.u1.b  = \add_37s_37s_37_2_1_U20.top_add_37s_37s_37_2_1_Adder_14_U.b [17:0];
assign \add_37s_37s_37_2_1_U20.top_add_37s_37s_37_2_1_Adder_14_U.u1.cin  = 1'h0;
assign \add_37s_37s_37_2_1_U20.top_add_37s_37s_37_2_1_Adder_14_U.facout_s1  = \add_37s_37s_37_2_1_U20.top_add_37s_37s_37_2_1_Adder_14_U.u1.cout ;
assign \add_37s_37s_37_2_1_U20.top_add_37s_37s_37_2_1_Adder_14_U.fas_s1  = \add_37s_37s_37_2_1_U20.top_add_37s_37s_37_2_1_Adder_14_U.u1.s ;
assign \add_37s_37s_37_2_1_U20.top_add_37s_37s_37_2_1_Adder_14_U.a  = \add_37s_37s_37_2_1_U20.din0 ;
assign \add_37s_37s_37_2_1_U20.top_add_37s_37s_37_2_1_Adder_14_U.b  = \add_37s_37s_37_2_1_U20.din1 ;
assign \add_37s_37s_37_2_1_U20.top_add_37s_37s_37_2_1_Adder_14_U.ce  = \add_37s_37s_37_2_1_U20.ce ;
assign \add_37s_37s_37_2_1_U20.top_add_37s_37s_37_2_1_Adder_14_U.clk  = \add_37s_37s_37_2_1_U20.clk ;
assign \add_37s_37s_37_2_1_U20.top_add_37s_37s_37_2_1_Adder_14_U.reset  = \add_37s_37s_37_2_1_U20.reset ;
assign \add_37s_37s_37_2_1_U20.dout  = \add_37s_37s_37_2_1_U20.top_add_37s_37s_37_2_1_Adder_14_U.s ;
assign \add_37s_37s_37_2_1_U20.ce  = 1'h1;
assign \add_37s_37s_37_2_1_U20.clk  = ap_clk;
assign \add_37s_37s_37_2_1_U20.din0  = { op_26_V_reg_1419[18], op_26_V_reg_1419[18], op_26_V_reg_1419[18], op_26_V_reg_1419[18], op_26_V_reg_1419[18], op_26_V_reg_1419[18], op_26_V_reg_1419[18], op_26_V_reg_1419[18], op_26_V_reg_1419[18], op_26_V_reg_1419[18], op_26_V_reg_1419[18], op_26_V_reg_1419[18], op_26_V_reg_1419[18], op_26_V_reg_1419[18], op_26_V_reg_1419, 4'h0 };
assign \add_37s_37s_37_2_1_U20.din1  = { op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16 };
assign grp_fu_837_p2 = \add_37s_37s_37_2_1_U20.dout ;
assign \add_37s_37s_37_2_1_U20.reset  = ap_rst;
assign \add_35s_35s_35_2_1_U24.top_add_35s_35s_35_2_1_Adder_17_U.ain_s0  = \add_35s_35s_35_2_1_U24.top_add_35s_35s_35_2_1_Adder_17_U.a ;
assign \add_35s_35s_35_2_1_U24.top_add_35s_35s_35_2_1_Adder_17_U.bin_s0  = \add_35s_35s_35_2_1_U24.top_add_35s_35s_35_2_1_Adder_17_U.b ;
assign \add_35s_35s_35_2_1_U24.top_add_35s_35s_35_2_1_Adder_17_U.s  = { \add_35s_35s_35_2_1_U24.top_add_35s_35s_35_2_1_Adder_17_U.fas_s2 , \add_35s_35s_35_2_1_U24.top_add_35s_35s_35_2_1_Adder_17_U.sum_s1  };
assign \add_35s_35s_35_2_1_U24.top_add_35s_35s_35_2_1_Adder_17_U.u2.a  = \add_35s_35s_35_2_1_U24.top_add_35s_35s_35_2_1_Adder_17_U.ain_s1 ;
assign \add_35s_35s_35_2_1_U24.top_add_35s_35s_35_2_1_Adder_17_U.u2.b  = \add_35s_35s_35_2_1_U24.top_add_35s_35s_35_2_1_Adder_17_U.bin_s1 ;
assign \add_35s_35s_35_2_1_U24.top_add_35s_35s_35_2_1_Adder_17_U.u2.cin  = \add_35s_35s_35_2_1_U24.top_add_35s_35s_35_2_1_Adder_17_U.carry_s1 ;
assign \add_35s_35s_35_2_1_U24.top_add_35s_35s_35_2_1_Adder_17_U.facout_s2  = \add_35s_35s_35_2_1_U24.top_add_35s_35s_35_2_1_Adder_17_U.u2.cout ;
assign \add_35s_35s_35_2_1_U24.top_add_35s_35s_35_2_1_Adder_17_U.fas_s2  = \add_35s_35s_35_2_1_U24.top_add_35s_35s_35_2_1_Adder_17_U.u2.s ;
assign \add_35s_35s_35_2_1_U24.top_add_35s_35s_35_2_1_Adder_17_U.u1.a  = \add_35s_35s_35_2_1_U24.top_add_35s_35s_35_2_1_Adder_17_U.a [16:0];
assign \add_35s_35s_35_2_1_U24.top_add_35s_35s_35_2_1_Adder_17_U.u1.b  = \add_35s_35s_35_2_1_U24.top_add_35s_35s_35_2_1_Adder_17_U.b [16:0];
assign \add_35s_35s_35_2_1_U24.top_add_35s_35s_35_2_1_Adder_17_U.u1.cin  = 1'h0;
assign \add_35s_35s_35_2_1_U24.top_add_35s_35s_35_2_1_Adder_17_U.facout_s1  = \add_35s_35s_35_2_1_U24.top_add_35s_35s_35_2_1_Adder_17_U.u1.cout ;
assign \add_35s_35s_35_2_1_U24.top_add_35s_35s_35_2_1_Adder_17_U.fas_s1  = \add_35s_35s_35_2_1_U24.top_add_35s_35s_35_2_1_Adder_17_U.u1.s ;
assign \add_35s_35s_35_2_1_U24.top_add_35s_35s_35_2_1_Adder_17_U.a  = \add_35s_35s_35_2_1_U24.din0 ;
assign \add_35s_35s_35_2_1_U24.top_add_35s_35s_35_2_1_Adder_17_U.b  = \add_35s_35s_35_2_1_U24.din1 ;
assign \add_35s_35s_35_2_1_U24.top_add_35s_35s_35_2_1_Adder_17_U.ce  = \add_35s_35s_35_2_1_U24.ce ;
assign \add_35s_35s_35_2_1_U24.top_add_35s_35s_35_2_1_Adder_17_U.clk  = \add_35s_35s_35_2_1_U24.clk ;
assign \add_35s_35s_35_2_1_U24.top_add_35s_35s_35_2_1_Adder_17_U.reset  = \add_35s_35s_35_2_1_U24.reset ;
assign \add_35s_35s_35_2_1_U24.dout  = \add_35s_35s_35_2_1_U24.top_add_35s_35s_35_2_1_Adder_17_U.s ;
assign \add_35s_35s_35_2_1_U24.ce  = 1'h1;
assign \add_35s_35s_35_2_1_U24.clk  = ap_clk;
assign \add_35s_35s_35_2_1_U24.din0  = { select_ln353_1_reg_1493[31], select_ln353_1_reg_1493, 2'h0 };
assign \add_35s_35s_35_2_1_U24.din1  = { op_18[7], op_18[7], op_18[7], op_18[7], op_18[7], op_18[7], op_18[7], op_18[7], op_18[7], op_18[7], op_18[7], op_18[7], op_18[7], op_18[7], op_18[7], op_18[7], op_18[7], op_18[7], op_18[7], op_18[7], op_18[7], op_18[7], op_18[7], op_18[7], op_18[7], op_18[7], op_18[7], op_18 };
assign grp_fu_967_p2 = \add_35s_35s_35_2_1_U24.dout ;
assign \add_35s_35s_35_2_1_U24.reset  = ap_rst;
assign \add_32ns_32ns_32_2_1_U26.top_add_32ns_32ns_32_2_1_Adder_15_U.ain_s0  = \add_32ns_32ns_32_2_1_U26.top_add_32ns_32ns_32_2_1_Adder_15_U.a ;
assign \add_32ns_32ns_32_2_1_U26.top_add_32ns_32ns_32_2_1_Adder_15_U.bin_s0  = \add_32ns_32ns_32_2_1_U26.top_add_32ns_32ns_32_2_1_Adder_15_U.b ;
assign \add_32ns_32ns_32_2_1_U26.top_add_32ns_32ns_32_2_1_Adder_15_U.s  = { \add_32ns_32ns_32_2_1_U26.top_add_32ns_32ns_32_2_1_Adder_15_U.fas_s2 , \add_32ns_32ns_32_2_1_U26.top_add_32ns_32ns_32_2_1_Adder_15_U.sum_s1  };
assign \add_32ns_32ns_32_2_1_U26.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.a  = \add_32ns_32ns_32_2_1_U26.top_add_32ns_32ns_32_2_1_Adder_15_U.ain_s1 ;
assign \add_32ns_32ns_32_2_1_U26.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.b  = \add_32ns_32ns_32_2_1_U26.top_add_32ns_32ns_32_2_1_Adder_15_U.bin_s1 ;
assign \add_32ns_32ns_32_2_1_U26.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.cin  = \add_32ns_32ns_32_2_1_U26.top_add_32ns_32ns_32_2_1_Adder_15_U.carry_s1 ;
assign \add_32ns_32ns_32_2_1_U26.top_add_32ns_32ns_32_2_1_Adder_15_U.facout_s2  = \add_32ns_32ns_32_2_1_U26.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.cout ;
assign \add_32ns_32ns_32_2_1_U26.top_add_32ns_32ns_32_2_1_Adder_15_U.fas_s2  = \add_32ns_32ns_32_2_1_U26.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.s ;
assign \add_32ns_32ns_32_2_1_U26.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.a  = \add_32ns_32ns_32_2_1_U26.top_add_32ns_32ns_32_2_1_Adder_15_U.a [15:0];
assign \add_32ns_32ns_32_2_1_U26.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.b  = \add_32ns_32ns_32_2_1_U26.top_add_32ns_32ns_32_2_1_Adder_15_U.b [15:0];
assign \add_32ns_32ns_32_2_1_U26.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.cin  = 1'h0;
assign \add_32ns_32ns_32_2_1_U26.top_add_32ns_32ns_32_2_1_Adder_15_U.facout_s1  = \add_32ns_32ns_32_2_1_U26.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.cout ;
assign \add_32ns_32ns_32_2_1_U26.top_add_32ns_32ns_32_2_1_Adder_15_U.fas_s1  = \add_32ns_32ns_32_2_1_U26.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.s ;
assign \add_32ns_32ns_32_2_1_U26.top_add_32ns_32ns_32_2_1_Adder_15_U.a  = \add_32ns_32ns_32_2_1_U26.din0 ;
assign \add_32ns_32ns_32_2_1_U26.top_add_32ns_32ns_32_2_1_Adder_15_U.b  = \add_32ns_32ns_32_2_1_U26.din1 ;
assign \add_32ns_32ns_32_2_1_U26.top_add_32ns_32ns_32_2_1_Adder_15_U.ce  = \add_32ns_32ns_32_2_1_U26.ce ;
assign \add_32ns_32ns_32_2_1_U26.top_add_32ns_32ns_32_2_1_Adder_15_U.clk  = \add_32ns_32ns_32_2_1_U26.clk ;
assign \add_32ns_32ns_32_2_1_U26.top_add_32ns_32ns_32_2_1_Adder_15_U.reset  = \add_32ns_32ns_32_2_1_U26.reset ;
assign \add_32ns_32ns_32_2_1_U26.dout  = \add_32ns_32ns_32_2_1_U26.top_add_32ns_32ns_32_2_1_Adder_15_U.s ;
assign \add_32ns_32ns_32_2_1_U26.ce  = 1'h1;
assign \add_32ns_32ns_32_2_1_U26.clk  = ap_clk;
assign \add_32ns_32ns_32_2_1_U26.din0  = ret_V_30_reg_1530;
assign \add_32ns_32ns_32_2_1_U26.din1  = select_ln69_1_reg_1535;
assign grp_fu_1025_p2 = \add_32ns_32ns_32_2_1_U26.dout ;
assign \add_32ns_32ns_32_2_1_U26.reset  = ap_rst;
assign \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.ain_s0  = \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.a ;
assign \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.bin_s0  = \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.b ;
assign \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.s  = { \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.fas_s2 , \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.sum_s1  };
assign \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.a  = \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.ain_s1 ;
assign \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.b  = \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.bin_s1 ;
assign \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.cin  = \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.carry_s1 ;
assign \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.facout_s2  = \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.cout ;
assign \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.fas_s2  = \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.s ;
assign \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.a  = \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.a [15:0];
assign \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.b  = \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.b [15:0];
assign \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.cin  = 1'h0;
assign \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.facout_s1  = \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.cout ;
assign \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.fas_s1  = \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.s ;
assign \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.a  = \add_32ns_32ns_32_2_1_U25.din0 ;
assign \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.b  = \add_32ns_32ns_32_2_1_U25.din1 ;
assign \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.ce  = \add_32ns_32ns_32_2_1_U25.ce ;
assign \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.clk  = \add_32ns_32ns_32_2_1_U25.clk ;
assign \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.reset  = \add_32ns_32ns_32_2_1_U25.reset ;
assign \add_32ns_32ns_32_2_1_U25.dout  = \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_15_U.s ;
assign \add_32ns_32ns_32_2_1_U25.ce  = 1'h1;
assign \add_32ns_32ns_32_2_1_U25.clk  = ap_clk;
assign \add_32ns_32ns_32_2_1_U25.din0  = ret_V_25_cast_reg_1518;
assign \add_32ns_32ns_32_2_1_U25.din1  = 32'd1;
assign grp_fu_993_p2 = \add_32ns_32ns_32_2_1_U25.dout ;
assign \add_32ns_32ns_32_2_1_U25.reset  = ap_rst;
assign \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.ain_s0  = \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.a ;
assign \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.bin_s0  = \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.b ;
assign \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.s  = { \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.fas_s2 , \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.sum_s1  };
assign \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.a  = \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.ain_s1 ;
assign \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.b  = \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.bin_s1 ;
assign \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.cin  = \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.carry_s1 ;
assign \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.facout_s2  = \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.cout ;
assign \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.fas_s2  = \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.s ;
assign \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.a  = \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.a [15:0];
assign \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.b  = \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.b [15:0];
assign \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.cin  = 1'h0;
assign \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.facout_s1  = \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.cout ;
assign \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.fas_s1  = \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.s ;
assign \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.a  = \add_32ns_32ns_32_2_1_U23.din0 ;
assign \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.b  = \add_32ns_32ns_32_2_1_U23.din1 ;
assign \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.ce  = \add_32ns_32ns_32_2_1_U23.ce ;
assign \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.clk  = \add_32ns_32ns_32_2_1_U23.clk ;
assign \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.reset  = \add_32ns_32ns_32_2_1_U23.reset ;
assign \add_32ns_32ns_32_2_1_U23.dout  = \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.s ;
assign \add_32ns_32ns_32_2_1_U23.ce  = 1'h1;
assign \add_32ns_32ns_32_2_1_U23.clk  = ap_clk;
assign \add_32ns_32ns_32_2_1_U23.din0  = ret_V_22_cast_reg_1481;
assign \add_32ns_32ns_32_2_1_U23.din1  = 32'd1;
assign grp_fu_928_p2 = \add_32ns_32ns_32_2_1_U23.dout ;
assign \add_32ns_32ns_32_2_1_U23.reset  = ap_rst;
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.ain_s0  = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.a ;
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.bin_s0  = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.b ;
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.s  = { \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.fas_s2 , \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.sum_s1  };
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.a  = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.ain_s1 ;
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.b  = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.bin_s1 ;
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.cin  = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.carry_s1 ;
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.facout_s2  = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.cout ;
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.fas_s2  = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.s ;
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.a  = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.a [15:0];
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.b  = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.b [15:0];
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.cin  = 1'h0;
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.facout_s1  = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.cout ;
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.fas_s1  = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.s ;
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.a  = \add_32ns_32ns_32_2_1_U21.din0 ;
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.b  = \add_32ns_32ns_32_2_1_U21.din1 ;
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.ce  = \add_32ns_32ns_32_2_1_U21.ce ;
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.clk  = \add_32ns_32ns_32_2_1_U21.clk ;
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.reset  = \add_32ns_32ns_32_2_1_U21.reset ;
assign \add_32ns_32ns_32_2_1_U21.dout  = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.s ;
assign \add_32ns_32ns_32_2_1_U21.ce  = 1'h1;
assign \add_32ns_32ns_32_2_1_U21.clk  = ap_clk;
assign \add_32ns_32ns_32_2_1_U21.din0  = ret_V_19_cast_reg_1444;
assign \add_32ns_32ns_32_2_1_U21.din1  = 32'd1;
assign grp_fu_863_p2 = \add_32ns_32ns_32_2_1_U21.dout ;
assign \add_32ns_32ns_32_2_1_U21.reset  = ap_rst;
assign \add_2ns_2s_2_2_1_U2.top_add_2ns_2s_2_2_1_Adder_0_U.ain_s0  = \add_2ns_2s_2_2_1_U2.top_add_2ns_2s_2_2_1_Adder_0_U.a ;
assign \add_2ns_2s_2_2_1_U2.top_add_2ns_2s_2_2_1_Adder_0_U.bin_s0  = \add_2ns_2s_2_2_1_U2.top_add_2ns_2s_2_2_1_Adder_0_U.b ;
assign \add_2ns_2s_2_2_1_U2.top_add_2ns_2s_2_2_1_Adder_0_U.s  = { \add_2ns_2s_2_2_1_U2.top_add_2ns_2s_2_2_1_Adder_0_U.fas_s2 , \add_2ns_2s_2_2_1_U2.top_add_2ns_2s_2_2_1_Adder_0_U.sum_s1  };
assign \add_2ns_2s_2_2_1_U2.top_add_2ns_2s_2_2_1_Adder_0_U.u2.a  = \add_2ns_2s_2_2_1_U2.top_add_2ns_2s_2_2_1_Adder_0_U.ain_s1 ;
assign \add_2ns_2s_2_2_1_U2.top_add_2ns_2s_2_2_1_Adder_0_U.u2.b  = \add_2ns_2s_2_2_1_U2.top_add_2ns_2s_2_2_1_Adder_0_U.bin_s1 ;
assign \add_2ns_2s_2_2_1_U2.top_add_2ns_2s_2_2_1_Adder_0_U.u2.cin  = \add_2ns_2s_2_2_1_U2.top_add_2ns_2s_2_2_1_Adder_0_U.carry_s1 ;
assign \add_2ns_2s_2_2_1_U2.top_add_2ns_2s_2_2_1_Adder_0_U.facout_s2  = \add_2ns_2s_2_2_1_U2.top_add_2ns_2s_2_2_1_Adder_0_U.u2.cout ;
assign \add_2ns_2s_2_2_1_U2.top_add_2ns_2s_2_2_1_Adder_0_U.fas_s2  = \add_2ns_2s_2_2_1_U2.top_add_2ns_2s_2_2_1_Adder_0_U.u2.s ;
assign \add_2ns_2s_2_2_1_U2.top_add_2ns_2s_2_2_1_Adder_0_U.u1.a  = \add_2ns_2s_2_2_1_U2.top_add_2ns_2s_2_2_1_Adder_0_U.a [0];
assign \add_2ns_2s_2_2_1_U2.top_add_2ns_2s_2_2_1_Adder_0_U.u1.b  = \add_2ns_2s_2_2_1_U2.top_add_2ns_2s_2_2_1_Adder_0_U.b [0];
assign \add_2ns_2s_2_2_1_U2.top_add_2ns_2s_2_2_1_Adder_0_U.u1.cin  = 1'h0;
assign \add_2ns_2s_2_2_1_U2.top_add_2ns_2s_2_2_1_Adder_0_U.facout_s1  = \add_2ns_2s_2_2_1_U2.top_add_2ns_2s_2_2_1_Adder_0_U.u1.cout ;
assign \add_2ns_2s_2_2_1_U2.top_add_2ns_2s_2_2_1_Adder_0_U.fas_s1  = \add_2ns_2s_2_2_1_U2.top_add_2ns_2s_2_2_1_Adder_0_U.u1.s ;
assign \add_2ns_2s_2_2_1_U2.top_add_2ns_2s_2_2_1_Adder_0_U.a  = \add_2ns_2s_2_2_1_U2.din0 ;
assign \add_2ns_2s_2_2_1_U2.top_add_2ns_2s_2_2_1_Adder_0_U.b  = \add_2ns_2s_2_2_1_U2.din1 ;
assign \add_2ns_2s_2_2_1_U2.top_add_2ns_2s_2_2_1_Adder_0_U.ce  = \add_2ns_2s_2_2_1_U2.ce ;
assign \add_2ns_2s_2_2_1_U2.top_add_2ns_2s_2_2_1_Adder_0_U.clk  = \add_2ns_2s_2_2_1_U2.clk ;
assign \add_2ns_2s_2_2_1_U2.top_add_2ns_2s_2_2_1_Adder_0_U.reset  = \add_2ns_2s_2_2_1_U2.reset ;
assign \add_2ns_2s_2_2_1_U2.dout  = \add_2ns_2s_2_2_1_U2.top_add_2ns_2s_2_2_1_Adder_0_U.s ;
assign \add_2ns_2s_2_2_1_U2.ce  = 1'h1;
assign \add_2ns_2s_2_2_1_U2.clk  = ap_clk;
assign \add_2ns_2s_2_2_1_U2.din0  = op_0[1:0];
assign \add_2ns_2s_2_2_1_U2.din1  = op_1;
assign grp_fu_303_p2 = \add_2ns_2s_2_2_1_U2.dout ;
assign \add_2ns_2s_2_2_1_U2.reset  = ap_rst;
assign \add_2ns_2ns_2_2_1_U18.top_add_2ns_2ns_2_2_1_Adder_6_U.ain_s0  = \add_2ns_2ns_2_2_1_U18.top_add_2ns_2ns_2_2_1_Adder_6_U.a ;
assign \add_2ns_2ns_2_2_1_U18.top_add_2ns_2ns_2_2_1_Adder_6_U.bin_s0  = \add_2ns_2ns_2_2_1_U18.top_add_2ns_2ns_2_2_1_Adder_6_U.b ;
assign \add_2ns_2ns_2_2_1_U18.top_add_2ns_2ns_2_2_1_Adder_6_U.s  = { \add_2ns_2ns_2_2_1_U18.top_add_2ns_2ns_2_2_1_Adder_6_U.fas_s2 , \add_2ns_2ns_2_2_1_U18.top_add_2ns_2ns_2_2_1_Adder_6_U.sum_s1  };
assign \add_2ns_2ns_2_2_1_U18.top_add_2ns_2ns_2_2_1_Adder_6_U.u2.a  = \add_2ns_2ns_2_2_1_U18.top_add_2ns_2ns_2_2_1_Adder_6_U.ain_s1 ;
assign \add_2ns_2ns_2_2_1_U18.top_add_2ns_2ns_2_2_1_Adder_6_U.u2.b  = \add_2ns_2ns_2_2_1_U18.top_add_2ns_2ns_2_2_1_Adder_6_U.bin_s1 ;
assign \add_2ns_2ns_2_2_1_U18.top_add_2ns_2ns_2_2_1_Adder_6_U.u2.cin  = \add_2ns_2ns_2_2_1_U18.top_add_2ns_2ns_2_2_1_Adder_6_U.carry_s1 ;
assign \add_2ns_2ns_2_2_1_U18.top_add_2ns_2ns_2_2_1_Adder_6_U.facout_s2  = \add_2ns_2ns_2_2_1_U18.top_add_2ns_2ns_2_2_1_Adder_6_U.u2.cout ;
assign \add_2ns_2ns_2_2_1_U18.top_add_2ns_2ns_2_2_1_Adder_6_U.fas_s2  = \add_2ns_2ns_2_2_1_U18.top_add_2ns_2ns_2_2_1_Adder_6_U.u2.s ;
assign \add_2ns_2ns_2_2_1_U18.top_add_2ns_2ns_2_2_1_Adder_6_U.u1.a  = \add_2ns_2ns_2_2_1_U18.top_add_2ns_2ns_2_2_1_Adder_6_U.a [0];
assign \add_2ns_2ns_2_2_1_U18.top_add_2ns_2ns_2_2_1_Adder_6_U.u1.b  = \add_2ns_2ns_2_2_1_U18.top_add_2ns_2ns_2_2_1_Adder_6_U.b [0];
assign \add_2ns_2ns_2_2_1_U18.top_add_2ns_2ns_2_2_1_Adder_6_U.u1.cin  = 1'h0;
assign \add_2ns_2ns_2_2_1_U18.top_add_2ns_2ns_2_2_1_Adder_6_U.facout_s1  = \add_2ns_2ns_2_2_1_U18.top_add_2ns_2ns_2_2_1_Adder_6_U.u1.cout ;
assign \add_2ns_2ns_2_2_1_U18.top_add_2ns_2ns_2_2_1_Adder_6_U.fas_s1  = \add_2ns_2ns_2_2_1_U18.top_add_2ns_2ns_2_2_1_Adder_6_U.u1.s ;
assign \add_2ns_2ns_2_2_1_U18.top_add_2ns_2ns_2_2_1_Adder_6_U.a  = \add_2ns_2ns_2_2_1_U18.din0 ;
assign \add_2ns_2ns_2_2_1_U18.top_add_2ns_2ns_2_2_1_Adder_6_U.b  = \add_2ns_2ns_2_2_1_U18.din1 ;
assign \add_2ns_2ns_2_2_1_U18.top_add_2ns_2ns_2_2_1_Adder_6_U.ce  = \add_2ns_2ns_2_2_1_U18.ce ;
assign \add_2ns_2ns_2_2_1_U18.top_add_2ns_2ns_2_2_1_Adder_6_U.clk  = \add_2ns_2ns_2_2_1_U18.clk ;
assign \add_2ns_2ns_2_2_1_U18.top_add_2ns_2ns_2_2_1_Adder_6_U.reset  = \add_2ns_2ns_2_2_1_U18.reset ;
assign \add_2ns_2ns_2_2_1_U18.dout  = \add_2ns_2ns_2_2_1_U18.top_add_2ns_2ns_2_2_1_Adder_6_U.s ;
assign \add_2ns_2ns_2_2_1_U18.ce  = 1'h1;
assign \add_2ns_2ns_2_2_1_U18.clk  = ap_clk;
assign \add_2ns_2ns_2_2_1_U18.din0  = select_ln69_reg_1389;
assign \add_2ns_2ns_2_2_1_U18.din1  = { 1'h0, ret_V_22_reg_1201 };
assign grp_fu_809_p2 = \add_2ns_2ns_2_2_1_U18.dout ;
assign \add_2ns_2ns_2_2_1_U18.reset  = ap_rst;
assign \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_6_U.ain_s0  = \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_6_U.a ;
assign \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_6_U.bin_s0  = \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_6_U.b ;
assign \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_6_U.s  = { \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_6_U.fas_s2 , \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_6_U.sum_s1  };
assign \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_6_U.u2.a  = \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_6_U.ain_s1 ;
assign \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_6_U.u2.b  = \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_6_U.bin_s1 ;
assign \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_6_U.u2.cin  = \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_6_U.carry_s1 ;
assign \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_6_U.facout_s2  = \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_6_U.u2.cout ;
assign \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_6_U.fas_s2  = \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_6_U.u2.s ;
assign \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_6_U.u1.a  = \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_6_U.a [0];
assign \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_6_U.u1.b  = \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_6_U.b [0];
assign \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_6_U.u1.cin  = 1'h0;
assign \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_6_U.facout_s1  = \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_6_U.u1.cout ;
assign \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_6_U.fas_s1  = \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_6_U.u1.s ;
assign \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_6_U.a  = \add_2ns_2ns_2_2_1_U10.din0 ;
assign \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_6_U.b  = \add_2ns_2ns_2_2_1_U10.din1 ;
assign \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_6_U.ce  = \add_2ns_2ns_2_2_1_U10.ce ;
assign \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_6_U.clk  = \add_2ns_2ns_2_2_1_U10.clk ;
assign \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_6_U.reset  = \add_2ns_2ns_2_2_1_U10.reset ;
assign \add_2ns_2ns_2_2_1_U10.dout  = \add_2ns_2ns_2_2_1_U10.top_add_2ns_2ns_2_2_1_Adder_6_U.s ;
assign \add_2ns_2ns_2_2_1_U10.ce  = 1'h1;
assign \add_2ns_2ns_2_2_1_U10.clk  = ap_clk;
assign \add_2ns_2ns_2_2_1_U10.din0  = ret_V_12_cast_reg_1173;
assign \add_2ns_2ns_2_2_1_U10.din1  = 2'h1;
assign grp_fu_467_p2 = \add_2ns_2ns_2_2_1_U10.dout ;
assign \add_2ns_2ns_2_2_1_U10.reset  = ap_rst;
assign \add_20ns_20s_20_2_1_U15.top_add_20ns_20s_20_2_1_Adder_11_U.ain_s0  = \add_20ns_20s_20_2_1_U15.top_add_20ns_20s_20_2_1_Adder_11_U.a ;
assign \add_20ns_20s_20_2_1_U15.top_add_20ns_20s_20_2_1_Adder_11_U.bin_s0  = \add_20ns_20s_20_2_1_U15.top_add_20ns_20s_20_2_1_Adder_11_U.b ;
assign \add_20ns_20s_20_2_1_U15.top_add_20ns_20s_20_2_1_Adder_11_U.s  = { \add_20ns_20s_20_2_1_U15.top_add_20ns_20s_20_2_1_Adder_11_U.fas_s2 , \add_20ns_20s_20_2_1_U15.top_add_20ns_20s_20_2_1_Adder_11_U.sum_s1  };
assign \add_20ns_20s_20_2_1_U15.top_add_20ns_20s_20_2_1_Adder_11_U.u2.a  = \add_20ns_20s_20_2_1_U15.top_add_20ns_20s_20_2_1_Adder_11_U.ain_s1 ;
assign \add_20ns_20s_20_2_1_U15.top_add_20ns_20s_20_2_1_Adder_11_U.u2.b  = \add_20ns_20s_20_2_1_U15.top_add_20ns_20s_20_2_1_Adder_11_U.bin_s1 ;
assign \add_20ns_20s_20_2_1_U15.top_add_20ns_20s_20_2_1_Adder_11_U.u2.cin  = \add_20ns_20s_20_2_1_U15.top_add_20ns_20s_20_2_1_Adder_11_U.carry_s1 ;
assign \add_20ns_20s_20_2_1_U15.top_add_20ns_20s_20_2_1_Adder_11_U.facout_s2  = \add_20ns_20s_20_2_1_U15.top_add_20ns_20s_20_2_1_Adder_11_U.u2.cout ;
assign \add_20ns_20s_20_2_1_U15.top_add_20ns_20s_20_2_1_Adder_11_U.fas_s2  = \add_20ns_20s_20_2_1_U15.top_add_20ns_20s_20_2_1_Adder_11_U.u2.s ;
assign \add_20ns_20s_20_2_1_U15.top_add_20ns_20s_20_2_1_Adder_11_U.u1.a  = \add_20ns_20s_20_2_1_U15.top_add_20ns_20s_20_2_1_Adder_11_U.a [9:0];
assign \add_20ns_20s_20_2_1_U15.top_add_20ns_20s_20_2_1_Adder_11_U.u1.b  = \add_20ns_20s_20_2_1_U15.top_add_20ns_20s_20_2_1_Adder_11_U.b [9:0];
assign \add_20ns_20s_20_2_1_U15.top_add_20ns_20s_20_2_1_Adder_11_U.u1.cin  = 1'h0;
assign \add_20ns_20s_20_2_1_U15.top_add_20ns_20s_20_2_1_Adder_11_U.facout_s1  = \add_20ns_20s_20_2_1_U15.top_add_20ns_20s_20_2_1_Adder_11_U.u1.cout ;
assign \add_20ns_20s_20_2_1_U15.top_add_20ns_20s_20_2_1_Adder_11_U.fas_s1  = \add_20ns_20s_20_2_1_U15.top_add_20ns_20s_20_2_1_Adder_11_U.u1.s ;
assign \add_20ns_20s_20_2_1_U15.top_add_20ns_20s_20_2_1_Adder_11_U.a  = \add_20ns_20s_20_2_1_U15.din0 ;
assign \add_20ns_20s_20_2_1_U15.top_add_20ns_20s_20_2_1_Adder_11_U.b  = \add_20ns_20s_20_2_1_U15.din1 ;
assign \add_20ns_20s_20_2_1_U15.top_add_20ns_20s_20_2_1_Adder_11_U.ce  = \add_20ns_20s_20_2_1_U15.ce ;
assign \add_20ns_20s_20_2_1_U15.top_add_20ns_20s_20_2_1_Adder_11_U.clk  = \add_20ns_20s_20_2_1_U15.clk ;
assign \add_20ns_20s_20_2_1_U15.top_add_20ns_20s_20_2_1_Adder_11_U.reset  = \add_20ns_20s_20_2_1_U15.reset ;
assign \add_20ns_20s_20_2_1_U15.dout  = \add_20ns_20s_20_2_1_U15.top_add_20ns_20s_20_2_1_Adder_11_U.s ;
assign \add_20ns_20s_20_2_1_U15.ce  = 1'h1;
assign \add_20ns_20s_20_2_1_U15.clk  = ap_clk;
assign \add_20ns_20s_20_2_1_U15.din0  = { op_22_V_reg_1337, 2'h0 };
assign \add_20ns_20s_20_2_1_U15.din1  = { op_12_V_reg_1332[3], op_12_V_reg_1332[3], op_12_V_reg_1332[3], op_12_V_reg_1332[3], op_12_V_reg_1332[3], op_12_V_reg_1332[3], op_12_V_reg_1332[3], op_12_V_reg_1332[3], op_12_V_reg_1332[3], op_12_V_reg_1332[3], op_12_V_reg_1332[3], op_12_V_reg_1332[3], op_12_V_reg_1332[3], op_12_V_reg_1332[3], op_12_V_reg_1332[3], op_12_V_reg_1332[3], op_12_V_reg_1332 };
assign grp_fu_740_p2 = \add_20ns_20s_20_2_1_U15.dout ;
assign \add_20ns_20s_20_2_1_U15.reset  = ap_rst;
assign \add_19s_19ns_19_2_1_U19.top_add_19s_19ns_19_2_1_Adder_12_U.ain_s0  = \add_19s_19ns_19_2_1_U19.top_add_19s_19ns_19_2_1_Adder_12_U.a ;
assign \add_19s_19ns_19_2_1_U19.top_add_19s_19ns_19_2_1_Adder_12_U.bin_s0  = \add_19s_19ns_19_2_1_U19.top_add_19s_19ns_19_2_1_Adder_12_U.b ;
assign \add_19s_19ns_19_2_1_U19.top_add_19s_19ns_19_2_1_Adder_12_U.s  = { \add_19s_19ns_19_2_1_U19.top_add_19s_19ns_19_2_1_Adder_12_U.fas_s2 , \add_19s_19ns_19_2_1_U19.top_add_19s_19ns_19_2_1_Adder_12_U.sum_s1  };
assign \add_19s_19ns_19_2_1_U19.top_add_19s_19ns_19_2_1_Adder_12_U.u2.a  = \add_19s_19ns_19_2_1_U19.top_add_19s_19ns_19_2_1_Adder_12_U.ain_s1 ;
assign \add_19s_19ns_19_2_1_U19.top_add_19s_19ns_19_2_1_Adder_12_U.u2.b  = \add_19s_19ns_19_2_1_U19.top_add_19s_19ns_19_2_1_Adder_12_U.bin_s1 ;
assign \add_19s_19ns_19_2_1_U19.top_add_19s_19ns_19_2_1_Adder_12_U.u2.cin  = \add_19s_19ns_19_2_1_U19.top_add_19s_19ns_19_2_1_Adder_12_U.carry_s1 ;
assign \add_19s_19ns_19_2_1_U19.top_add_19s_19ns_19_2_1_Adder_12_U.facout_s2  = \add_19s_19ns_19_2_1_U19.top_add_19s_19ns_19_2_1_Adder_12_U.u2.cout ;
assign \add_19s_19ns_19_2_1_U19.top_add_19s_19ns_19_2_1_Adder_12_U.fas_s2  = \add_19s_19ns_19_2_1_U19.top_add_19s_19ns_19_2_1_Adder_12_U.u2.s ;
assign \add_19s_19ns_19_2_1_U19.top_add_19s_19ns_19_2_1_Adder_12_U.u1.a  = \add_19s_19ns_19_2_1_U19.top_add_19s_19ns_19_2_1_Adder_12_U.a [8:0];
assign \add_19s_19ns_19_2_1_U19.top_add_19s_19ns_19_2_1_Adder_12_U.u1.b  = \add_19s_19ns_19_2_1_U19.top_add_19s_19ns_19_2_1_Adder_12_U.b [8:0];
assign \add_19s_19ns_19_2_1_U19.top_add_19s_19ns_19_2_1_Adder_12_U.u1.cin  = 1'h0;
assign \add_19s_19ns_19_2_1_U19.top_add_19s_19ns_19_2_1_Adder_12_U.facout_s1  = \add_19s_19ns_19_2_1_U19.top_add_19s_19ns_19_2_1_Adder_12_U.u1.cout ;
assign \add_19s_19ns_19_2_1_U19.top_add_19s_19ns_19_2_1_Adder_12_U.fas_s1  = \add_19s_19ns_19_2_1_U19.top_add_19s_19ns_19_2_1_Adder_12_U.u1.s ;
assign \add_19s_19ns_19_2_1_U19.top_add_19s_19ns_19_2_1_Adder_12_U.a  = \add_19s_19ns_19_2_1_U19.din0 ;
assign \add_19s_19ns_19_2_1_U19.top_add_19s_19ns_19_2_1_Adder_12_U.b  = \add_19s_19ns_19_2_1_U19.din1 ;
assign \add_19s_19ns_19_2_1_U19.top_add_19s_19ns_19_2_1_Adder_12_U.ce  = \add_19s_19ns_19_2_1_U19.ce ;
assign \add_19s_19ns_19_2_1_U19.top_add_19s_19ns_19_2_1_Adder_12_U.clk  = \add_19s_19ns_19_2_1_U19.clk ;
assign \add_19s_19ns_19_2_1_U19.top_add_19s_19ns_19_2_1_Adder_12_U.reset  = \add_19s_19ns_19_2_1_U19.reset ;
assign \add_19s_19ns_19_2_1_U19.dout  = \add_19s_19ns_19_2_1_U19.top_add_19s_19ns_19_2_1_Adder_12_U.s ;
assign \add_19s_19ns_19_2_1_U19.ce  = 1'h1;
assign \add_19s_19ns_19_2_1_U19.clk  = ap_clk;
assign \add_19s_19ns_19_2_1_U19.din0  = { add_ln69_3_reg_1409[1], add_ln69_3_reg_1409[1], add_ln69_3_reg_1409[1], add_ln69_3_reg_1409[1], add_ln69_3_reg_1409[1], add_ln69_3_reg_1409[1], add_ln69_3_reg_1409[1], add_ln69_3_reg_1409[1], add_ln69_3_reg_1409[1], add_ln69_3_reg_1409[1], add_ln69_3_reg_1409[1], add_ln69_3_reg_1409[1], add_ln69_3_reg_1409[1], add_ln69_3_reg_1409[1], add_ln69_3_reg_1409[1], add_ln69_3_reg_1409[1], add_ln69_3_reg_1409[1], add_ln69_3_reg_1409 };
assign \add_19s_19ns_19_2_1_U19.din1  = add_ln69_2_reg_1404;
assign grp_fu_817_p2 = \add_19s_19ns_19_2_1_U19.dout ;
assign \add_19s_19ns_19_2_1_U19.reset  = ap_rst;
assign \add_19s_19ns_19_2_1_U16.top_add_19s_19ns_19_2_1_Adder_12_U.ain_s0  = \add_19s_19ns_19_2_1_U16.top_add_19s_19ns_19_2_1_Adder_12_U.a ;
assign \add_19s_19ns_19_2_1_U16.top_add_19s_19ns_19_2_1_Adder_12_U.bin_s0  = \add_19s_19ns_19_2_1_U16.top_add_19s_19ns_19_2_1_Adder_12_U.b ;
assign \add_19s_19ns_19_2_1_U16.top_add_19s_19ns_19_2_1_Adder_12_U.s  = { \add_19s_19ns_19_2_1_U16.top_add_19s_19ns_19_2_1_Adder_12_U.fas_s2 , \add_19s_19ns_19_2_1_U16.top_add_19s_19ns_19_2_1_Adder_12_U.sum_s1  };
assign \add_19s_19ns_19_2_1_U16.top_add_19s_19ns_19_2_1_Adder_12_U.u2.a  = \add_19s_19ns_19_2_1_U16.top_add_19s_19ns_19_2_1_Adder_12_U.ain_s1 ;
assign \add_19s_19ns_19_2_1_U16.top_add_19s_19ns_19_2_1_Adder_12_U.u2.b  = \add_19s_19ns_19_2_1_U16.top_add_19s_19ns_19_2_1_Adder_12_U.bin_s1 ;
assign \add_19s_19ns_19_2_1_U16.top_add_19s_19ns_19_2_1_Adder_12_U.u2.cin  = \add_19s_19ns_19_2_1_U16.top_add_19s_19ns_19_2_1_Adder_12_U.carry_s1 ;
assign \add_19s_19ns_19_2_1_U16.top_add_19s_19ns_19_2_1_Adder_12_U.facout_s2  = \add_19s_19ns_19_2_1_U16.top_add_19s_19ns_19_2_1_Adder_12_U.u2.cout ;
assign \add_19s_19ns_19_2_1_U16.top_add_19s_19ns_19_2_1_Adder_12_U.fas_s2  = \add_19s_19ns_19_2_1_U16.top_add_19s_19ns_19_2_1_Adder_12_U.u2.s ;
assign \add_19s_19ns_19_2_1_U16.top_add_19s_19ns_19_2_1_Adder_12_U.u1.a  = \add_19s_19ns_19_2_1_U16.top_add_19s_19ns_19_2_1_Adder_12_U.a [8:0];
assign \add_19s_19ns_19_2_1_U16.top_add_19s_19ns_19_2_1_Adder_12_U.u1.b  = \add_19s_19ns_19_2_1_U16.top_add_19s_19ns_19_2_1_Adder_12_U.b [8:0];
assign \add_19s_19ns_19_2_1_U16.top_add_19s_19ns_19_2_1_Adder_12_U.u1.cin  = 1'h0;
assign \add_19s_19ns_19_2_1_U16.top_add_19s_19ns_19_2_1_Adder_12_U.facout_s1  = \add_19s_19ns_19_2_1_U16.top_add_19s_19ns_19_2_1_Adder_12_U.u1.cout ;
assign \add_19s_19ns_19_2_1_U16.top_add_19s_19ns_19_2_1_Adder_12_U.fas_s1  = \add_19s_19ns_19_2_1_U16.top_add_19s_19ns_19_2_1_Adder_12_U.u1.s ;
assign \add_19s_19ns_19_2_1_U16.top_add_19s_19ns_19_2_1_Adder_12_U.a  = \add_19s_19ns_19_2_1_U16.din0 ;
assign \add_19s_19ns_19_2_1_U16.top_add_19s_19ns_19_2_1_Adder_12_U.b  = \add_19s_19ns_19_2_1_U16.din1 ;
assign \add_19s_19ns_19_2_1_U16.top_add_19s_19ns_19_2_1_Adder_12_U.ce  = \add_19s_19ns_19_2_1_U16.ce ;
assign \add_19s_19ns_19_2_1_U16.top_add_19s_19ns_19_2_1_Adder_12_U.clk  = \add_19s_19ns_19_2_1_U16.clk ;
assign \add_19s_19ns_19_2_1_U16.top_add_19s_19ns_19_2_1_Adder_12_U.reset  = \add_19s_19ns_19_2_1_U16.reset ;
assign \add_19s_19ns_19_2_1_U16.dout  = \add_19s_19ns_19_2_1_U16.top_add_19s_19ns_19_2_1_Adder_12_U.s ;
assign \add_19s_19ns_19_2_1_U16.ce  = 1'h1;
assign \add_19s_19ns_19_2_1_U16.clk  = ap_clk;
assign \add_19s_19ns_19_2_1_U16.din0  = { tmp_1_reg_1367[17], tmp_1_reg_1367 };
assign \add_19s_19ns_19_2_1_U16.din1  = 19'h00001;
assign grp_fu_764_p2 = \add_19s_19ns_19_2_1_U16.dout ;
assign \add_19s_19ns_19_2_1_U16.reset  = ap_rst;
assign \add_19ns_19s_19_2_1_U17.top_add_19ns_19s_19_2_1_Adder_13_U.ain_s0  = \add_19ns_19s_19_2_1_U17.top_add_19ns_19s_19_2_1_Adder_13_U.a ;
assign \add_19ns_19s_19_2_1_U17.top_add_19ns_19s_19_2_1_Adder_13_U.bin_s0  = \add_19ns_19s_19_2_1_U17.top_add_19ns_19s_19_2_1_Adder_13_U.b ;
assign \add_19ns_19s_19_2_1_U17.top_add_19ns_19s_19_2_1_Adder_13_U.s  = { \add_19ns_19s_19_2_1_U17.top_add_19ns_19s_19_2_1_Adder_13_U.fas_s2 , \add_19ns_19s_19_2_1_U17.top_add_19ns_19s_19_2_1_Adder_13_U.sum_s1  };
assign \add_19ns_19s_19_2_1_U17.top_add_19ns_19s_19_2_1_Adder_13_U.u2.a  = \add_19ns_19s_19_2_1_U17.top_add_19ns_19s_19_2_1_Adder_13_U.ain_s1 ;
assign \add_19ns_19s_19_2_1_U17.top_add_19ns_19s_19_2_1_Adder_13_U.u2.b  = \add_19ns_19s_19_2_1_U17.top_add_19ns_19s_19_2_1_Adder_13_U.bin_s1 ;
assign \add_19ns_19s_19_2_1_U17.top_add_19ns_19s_19_2_1_Adder_13_U.u2.cin  = \add_19ns_19s_19_2_1_U17.top_add_19ns_19s_19_2_1_Adder_13_U.carry_s1 ;
assign \add_19ns_19s_19_2_1_U17.top_add_19ns_19s_19_2_1_Adder_13_U.facout_s2  = \add_19ns_19s_19_2_1_U17.top_add_19ns_19s_19_2_1_Adder_13_U.u2.cout ;
assign \add_19ns_19s_19_2_1_U17.top_add_19ns_19s_19_2_1_Adder_13_U.fas_s2  = \add_19ns_19s_19_2_1_U17.top_add_19ns_19s_19_2_1_Adder_13_U.u2.s ;
assign \add_19ns_19s_19_2_1_U17.top_add_19ns_19s_19_2_1_Adder_13_U.u1.a  = \add_19ns_19s_19_2_1_U17.top_add_19ns_19s_19_2_1_Adder_13_U.a [8:0];
assign \add_19ns_19s_19_2_1_U17.top_add_19ns_19s_19_2_1_Adder_13_U.u1.b  = \add_19ns_19s_19_2_1_U17.top_add_19ns_19s_19_2_1_Adder_13_U.b [8:0];
assign \add_19ns_19s_19_2_1_U17.top_add_19ns_19s_19_2_1_Adder_13_U.u1.cin  = 1'h0;
assign \add_19ns_19s_19_2_1_U17.top_add_19ns_19s_19_2_1_Adder_13_U.facout_s1  = \add_19ns_19s_19_2_1_U17.top_add_19ns_19s_19_2_1_Adder_13_U.u1.cout ;
assign \add_19ns_19s_19_2_1_U17.top_add_19ns_19s_19_2_1_Adder_13_U.fas_s1  = \add_19ns_19s_19_2_1_U17.top_add_19ns_19s_19_2_1_Adder_13_U.u1.s ;
assign \add_19ns_19s_19_2_1_U17.top_add_19ns_19s_19_2_1_Adder_13_U.a  = \add_19ns_19s_19_2_1_U17.din0 ;
assign \add_19ns_19s_19_2_1_U17.top_add_19ns_19s_19_2_1_Adder_13_U.b  = \add_19ns_19s_19_2_1_U17.din1 ;
assign \add_19ns_19s_19_2_1_U17.top_add_19ns_19s_19_2_1_Adder_13_U.ce  = \add_19ns_19s_19_2_1_U17.ce ;
assign \add_19ns_19s_19_2_1_U17.top_add_19ns_19s_19_2_1_Adder_13_U.clk  = \add_19ns_19s_19_2_1_U17.clk ;
assign \add_19ns_19s_19_2_1_U17.top_add_19ns_19s_19_2_1_Adder_13_U.reset  = \add_19ns_19s_19_2_1_U17.reset ;
assign \add_19ns_19s_19_2_1_U17.dout  = \add_19ns_19s_19_2_1_U17.top_add_19ns_19s_19_2_1_Adder_13_U.s ;
assign \add_19ns_19s_19_2_1_U17.ce  = 1'h1;
assign \add_19ns_19s_19_2_1_U17.clk  = ap_clk;
assign \add_19ns_19s_19_2_1_U17.din0  = ret_V_26_reg_1384;
assign \add_19ns_19s_19_2_1_U17.din1  = { op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14[3], op_14 };
assign grp_fu_804_p2 = \add_19ns_19s_19_2_1_U17.dout ;
assign \add_19ns_19s_19_2_1_U17.reset  = ap_rst;
assign \add_18s_18ns_18_2_1_U14.top_add_18s_18ns_18_2_1_Adder_10_U.ain_s0  = \add_18s_18ns_18_2_1_U14.top_add_18s_18ns_18_2_1_Adder_10_U.a ;
assign \add_18s_18ns_18_2_1_U14.top_add_18s_18ns_18_2_1_Adder_10_U.bin_s0  = \add_18s_18ns_18_2_1_U14.top_add_18s_18ns_18_2_1_Adder_10_U.b ;
assign \add_18s_18ns_18_2_1_U14.top_add_18s_18ns_18_2_1_Adder_10_U.s  = { \add_18s_18ns_18_2_1_U14.top_add_18s_18ns_18_2_1_Adder_10_U.fas_s2 , \add_18s_18ns_18_2_1_U14.top_add_18s_18ns_18_2_1_Adder_10_U.sum_s1  };
assign \add_18s_18ns_18_2_1_U14.top_add_18s_18ns_18_2_1_Adder_10_U.u2.a  = \add_18s_18ns_18_2_1_U14.top_add_18s_18ns_18_2_1_Adder_10_U.ain_s1 ;
assign \add_18s_18ns_18_2_1_U14.top_add_18s_18ns_18_2_1_Adder_10_U.u2.b  = \add_18s_18ns_18_2_1_U14.top_add_18s_18ns_18_2_1_Adder_10_U.bin_s1 ;
assign \add_18s_18ns_18_2_1_U14.top_add_18s_18ns_18_2_1_Adder_10_U.u2.cin  = \add_18s_18ns_18_2_1_U14.top_add_18s_18ns_18_2_1_Adder_10_U.carry_s1 ;
assign \add_18s_18ns_18_2_1_U14.top_add_18s_18ns_18_2_1_Adder_10_U.facout_s2  = \add_18s_18ns_18_2_1_U14.top_add_18s_18ns_18_2_1_Adder_10_U.u2.cout ;
assign \add_18s_18ns_18_2_1_U14.top_add_18s_18ns_18_2_1_Adder_10_U.fas_s2  = \add_18s_18ns_18_2_1_U14.top_add_18s_18ns_18_2_1_Adder_10_U.u2.s ;
assign \add_18s_18ns_18_2_1_U14.top_add_18s_18ns_18_2_1_Adder_10_U.u1.a  = \add_18s_18ns_18_2_1_U14.top_add_18s_18ns_18_2_1_Adder_10_U.a [8:0];
assign \add_18s_18ns_18_2_1_U14.top_add_18s_18ns_18_2_1_Adder_10_U.u1.b  = \add_18s_18ns_18_2_1_U14.top_add_18s_18ns_18_2_1_Adder_10_U.b [8:0];
assign \add_18s_18ns_18_2_1_U14.top_add_18s_18ns_18_2_1_Adder_10_U.u1.cin  = 1'h0;
assign \add_18s_18ns_18_2_1_U14.top_add_18s_18ns_18_2_1_Adder_10_U.facout_s1  = \add_18s_18ns_18_2_1_U14.top_add_18s_18ns_18_2_1_Adder_10_U.u1.cout ;
assign \add_18s_18ns_18_2_1_U14.top_add_18s_18ns_18_2_1_Adder_10_U.fas_s1  = \add_18s_18ns_18_2_1_U14.top_add_18s_18ns_18_2_1_Adder_10_U.u1.s ;
assign \add_18s_18ns_18_2_1_U14.top_add_18s_18ns_18_2_1_Adder_10_U.a  = \add_18s_18ns_18_2_1_U14.din0 ;
assign \add_18s_18ns_18_2_1_U14.top_add_18s_18ns_18_2_1_Adder_10_U.b  = \add_18s_18ns_18_2_1_U14.din1 ;
assign \add_18s_18ns_18_2_1_U14.top_add_18s_18ns_18_2_1_Adder_10_U.ce  = \add_18s_18ns_18_2_1_U14.ce ;
assign \add_18s_18ns_18_2_1_U14.top_add_18s_18ns_18_2_1_Adder_10_U.clk  = \add_18s_18ns_18_2_1_U14.clk ;
assign \add_18s_18ns_18_2_1_U14.top_add_18s_18ns_18_2_1_Adder_10_U.reset  = \add_18s_18ns_18_2_1_U14.reset ;
assign \add_18s_18ns_18_2_1_U14.dout  = \add_18s_18ns_18_2_1_U14.top_add_18s_18ns_18_2_1_Adder_10_U.s ;
assign \add_18s_18ns_18_2_1_U14.ce  = 1'h1;
assign \add_18s_18ns_18_2_1_U14.clk  = ap_clk;
assign \add_18s_18ns_18_2_1_U14.din0  = { add_ln69_reg_1306[6], add_ln69_reg_1306[6], add_ln69_reg_1306[6], add_ln69_reg_1306[6], add_ln69_reg_1306[6], add_ln69_reg_1306[6], add_ln69_reg_1306[6], add_ln69_reg_1306[6], add_ln69_reg_1306[6], add_ln69_reg_1306[6], add_ln69_reg_1306[6], add_ln69_reg_1306 };
assign \add_18s_18ns_18_2_1_U14.din1  = { 2'h0, op_11 };
assign grp_fu_686_p2 = \add_18s_18ns_18_2_1_U14.dout ;
assign \add_18s_18ns_18_2_1_U14.reset  = ap_rst;
assign \add_12s_12s_12_2_1_U7.top_add_12s_12s_12_2_1_Adder_5_U.ain_s0  = \add_12s_12s_12_2_1_U7.top_add_12s_12s_12_2_1_Adder_5_U.a ;
assign \add_12s_12s_12_2_1_U7.top_add_12s_12s_12_2_1_Adder_5_U.bin_s0  = \add_12s_12s_12_2_1_U7.top_add_12s_12s_12_2_1_Adder_5_U.b ;
assign \add_12s_12s_12_2_1_U7.top_add_12s_12s_12_2_1_Adder_5_U.s  = { \add_12s_12s_12_2_1_U7.top_add_12s_12s_12_2_1_Adder_5_U.fas_s2 , \add_12s_12s_12_2_1_U7.top_add_12s_12s_12_2_1_Adder_5_U.sum_s1  };
assign \add_12s_12s_12_2_1_U7.top_add_12s_12s_12_2_1_Adder_5_U.u2.a  = \add_12s_12s_12_2_1_U7.top_add_12s_12s_12_2_1_Adder_5_U.ain_s1 ;
assign \add_12s_12s_12_2_1_U7.top_add_12s_12s_12_2_1_Adder_5_U.u2.b  = \add_12s_12s_12_2_1_U7.top_add_12s_12s_12_2_1_Adder_5_U.bin_s1 ;
assign \add_12s_12s_12_2_1_U7.top_add_12s_12s_12_2_1_Adder_5_U.u2.cin  = \add_12s_12s_12_2_1_U7.top_add_12s_12s_12_2_1_Adder_5_U.carry_s1 ;
assign \add_12s_12s_12_2_1_U7.top_add_12s_12s_12_2_1_Adder_5_U.facout_s2  = \add_12s_12s_12_2_1_U7.top_add_12s_12s_12_2_1_Adder_5_U.u2.cout ;
assign \add_12s_12s_12_2_1_U7.top_add_12s_12s_12_2_1_Adder_5_U.fas_s2  = \add_12s_12s_12_2_1_U7.top_add_12s_12s_12_2_1_Adder_5_U.u2.s ;
assign \add_12s_12s_12_2_1_U7.top_add_12s_12s_12_2_1_Adder_5_U.u1.a  = \add_12s_12s_12_2_1_U7.top_add_12s_12s_12_2_1_Adder_5_U.a [5:0];
assign \add_12s_12s_12_2_1_U7.top_add_12s_12s_12_2_1_Adder_5_U.u1.b  = \add_12s_12s_12_2_1_U7.top_add_12s_12s_12_2_1_Adder_5_U.b [5:0];
assign \add_12s_12s_12_2_1_U7.top_add_12s_12s_12_2_1_Adder_5_U.u1.cin  = 1'h0;
assign \add_12s_12s_12_2_1_U7.top_add_12s_12s_12_2_1_Adder_5_U.facout_s1  = \add_12s_12s_12_2_1_U7.top_add_12s_12s_12_2_1_Adder_5_U.u1.cout ;
assign \add_12s_12s_12_2_1_U7.top_add_12s_12s_12_2_1_Adder_5_U.fas_s1  = \add_12s_12s_12_2_1_U7.top_add_12s_12s_12_2_1_Adder_5_U.u1.s ;
assign \add_12s_12s_12_2_1_U7.top_add_12s_12s_12_2_1_Adder_5_U.a  = \add_12s_12s_12_2_1_U7.din0 ;
assign \add_12s_12s_12_2_1_U7.top_add_12s_12s_12_2_1_Adder_5_U.b  = \add_12s_12s_12_2_1_U7.din1 ;
assign \add_12s_12s_12_2_1_U7.top_add_12s_12s_12_2_1_Adder_5_U.ce  = \add_12s_12s_12_2_1_U7.ce ;
assign \add_12s_12s_12_2_1_U7.top_add_12s_12s_12_2_1_Adder_5_U.clk  = \add_12s_12s_12_2_1_U7.clk ;
assign \add_12s_12s_12_2_1_U7.top_add_12s_12s_12_2_1_Adder_5_U.reset  = \add_12s_12s_12_2_1_U7.reset ;
assign \add_12s_12s_12_2_1_U7.dout  = \add_12s_12s_12_2_1_U7.top_add_12s_12s_12_2_1_Adder_5_U.s ;
assign \add_12s_12s_12_2_1_U7.ce  = 1'h1;
assign \add_12s_12s_12_2_1_U7.clk  = ap_clk;
assign \add_12s_12s_12_2_1_U7.din0  = { op_8_V_reg_1112[7], op_8_V_reg_1112, 3'h0 };
assign \add_12s_12s_12_2_1_U7.din1  = { op_3[7], op_3[7], op_3[7], op_3[7], op_3 };
assign grp_fu_413_p2 = \add_12s_12s_12_2_1_U7.dout ;
assign \add_12s_12s_12_2_1_U7.reset  = ap_rst;
endmodule


// Product machine:
module top_A_times_top_B (ap_start, op_0, op_1, op_11, op_14, op_15, op_16, op_17, op_18, op_19, op_3, op_4, op_7, op_9, ap_clk, unsafe_signal);
input ap_start;
input [3:0] op_0;
input [1:0] op_1;
input [15:0] op_11;
input [3:0] op_14;
input op_15;
input [7:0] op_16;
input [31:0] op_17;
input [7:0] op_18;
input op_19;
input [7:0] op_3;
input [15:0] op_4;
input [3:0] op_7;
input [7:0] op_9;
input ap_clk;
output unsafe_signal;
reg _setup;
initial _setup = 1'b0;
always @ (posedge ap_clk) _setup <= 1'b1;
reg ap_start_internal;
always @ (posedge ap_clk) if (!_setup) ap_start_internal <= ap_start;
reg [3:0] op_0_internal;
always @ (posedge ap_clk) if (!_setup) op_0_internal <= op_0;
reg [1:0] op_1_internal;
always @ (posedge ap_clk) if (!_setup) op_1_internal <= op_1;
reg [15:0] op_11_internal;
always @ (posedge ap_clk) if (!_setup) op_11_internal <= op_11;
reg [3:0] op_14_internal;
always @ (posedge ap_clk) if (!_setup) op_14_internal <= op_14;
reg op_15_internal;
always @ (posedge ap_clk) if (!_setup) op_15_internal <= op_15;
reg [7:0] op_16_internal;
always @ (posedge ap_clk) if (!_setup) op_16_internal <= op_16;
reg [31:0] op_17_internal;
always @ (posedge ap_clk) if (!_setup) op_17_internal <= op_17;
reg [7:0] op_18_internal;
always @ (posedge ap_clk) if (!_setup) op_18_internal <= op_18;
reg op_19_internal;
always @ (posedge ap_clk) if (!_setup) op_19_internal <= op_19;
reg [7:0] op_3_internal;
always @ (posedge ap_clk) if (!_setup) op_3_internal <= op_3;
reg [15:0] op_4_internal;
always @ (posedge ap_clk) if (!_setup) op_4_internal <= op_4;
reg [3:0] op_7_internal;
always @ (posedge ap_clk) if (!_setup) op_7_internal <= op_7;
reg [7:0] op_9_internal;
always @ (posedge ap_clk) if (!_setup) op_9_internal <= op_9;
wire ap_done_A;
wire ap_done_B;
wire ap_done_eq;
assign ap_done_eq = ap_done_A == ap_done_B;
wire ap_idle_A;
wire ap_idle_B;
wire ap_idle_eq;
assign ap_idle_eq = ap_idle_A == ap_idle_B;
wire ap_ready_A;
wire ap_ready_B;
wire ap_ready_eq;
assign ap_ready_eq = ap_ready_A == ap_ready_B;
wire [31:0] op_30_A;
wire [31:0] op_30_B;
wire op_30_eq;
assign op_30_eq = op_30_A == op_30_B;
wire op_30_ap_vld_A;
wire op_30_ap_vld_B;
wire clk_enable_A;
wire clk_enable_B;
assign clk_enable_A = _setup & (~op_30_ap_vld_A | op_30_ap_vld_B);
assign clk_enable_B = _setup;
wire divergent;
assign divergent = ~(ap_done_eq & ap_idle_eq & ap_ready_eq & op_30_eq);
assign unsafe_signal = op_30_ap_vld_A & op_30_ap_vld_B & divergent;
top_A instance_A (
    .ap_clk(ap_clk),
    .clk_enable(clk_enable_A),
    .ap_start(ap_start_internal),
    .op_0(op_0_internal),
    .op_1(op_1_internal),
    .op_11(op_11_internal),
    .op_14(op_14_internal),
    .op_15(op_15_internal),
    .op_16(op_16_internal),
    .op_17(op_17_internal),
    .op_18(op_18_internal),
    .op_19(op_19_internal),
    .op_3(op_3_internal),
    .op_4(op_4_internal),
    .op_7(op_7_internal),
    .op_9(op_9_internal),
    .ap_done(ap_done_A),
    .ap_idle(ap_idle_A),
    .ap_ready(ap_ready_A),
    .op_30(op_30_A),
    .op_30_ap_vld(op_30_ap_vld_A)
);
top_B instance_B (
    .ap_clk(ap_clk),
    .clk_enable(clk_enable_B),
    .ap_start(ap_start_internal),
    .op_0(op_0_internal),
    .op_1(op_1_internal),
    .op_11(op_11_internal),
    .op_14(op_14_internal),
    .op_15(op_15_internal),
    .op_16(op_16_internal),
    .op_17(op_17_internal),
    .op_18(op_18_internal),
    .op_19(op_19_internal),
    .op_3(op_3_internal),
    .op_4(op_4_internal),
    .op_7(op_7_internal),
    .op_9(op_9_internal),
    .ap_done(ap_done_B),
    .ap_idle(ap_idle_B),
    .ap_ready(ap_ready_B),
    .op_30(op_30_B),
    .op_30_ap_vld(op_30_ap_vld_B)
);
endmodule
