// Processed by function `construct_kairos` in `verilog_tricks.py`.
// Machine A:
// Processed by function `add_clk_enable_signal` in `verilog_tricks.py`.
// Processed by function `remove_reset_signal` in `verilog_tricks.py`.
module top_A (
  ap_clk,
  ap_start,
  ap_done,
  ap_idle,
  ap_ready,
  op_0,
  op_1,
  op_2,
  op_4,
  op_5,
  op_6,
  op_8,
  op_9,
  op_10,
  op_12,
  op_13,
  op_14,
  op_15,
  op_16,
  op_17,
  op_18,
  op_32,
  op_32_ap_vld,
clk_enable
);
input clk_enable;


input ap_clk;
wire ap_rst;
assign ap_rst = op_32_ap_vld;
input ap_start;
input op_0;
input [3:0] op_1;
input [7:0] op_10;
input [3:0] op_12;
input [7:0] op_13;
input [1:0] op_14;
input [7:0] op_15;
input [7:0] op_16;
input [3:0] op_17;
input [1:0] op_18;
input [3:0] op_2;
input [15:0] op_4;
input [7:0] op_5;
input [15:0] op_6;
input [3:0] op_8;
input [3:0] op_9;
output ap_done;
output ap_idle;
output ap_ready;
output [31:0] op_32;
output op_32_ap_vld;


reg Range1_all_zeros_reg_1354;
reg [4:0] \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_10_U.ain_s1 ;
reg [4:0] \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_10_U.bin_s1 ;
reg \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_10_U.carry_s1 ;
reg [4:0] \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_10_U.sum_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_4_U.ain_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_4_U.bin_s1 ;
reg \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_4_U.carry_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_4_U.sum_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_4_U.ain_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_4_U.bin_s1 ;
reg \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_4_U.carry_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_4_U.sum_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_4_U.ain_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_4_U.bin_s1 ;
reg \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_4_U.carry_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_4_U.sum_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.ain_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.bin_s1 ;
reg \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.carry_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.sum_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.ain_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.bin_s1 ;
reg \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.carry_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.sum_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_4_U.ain_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_4_U.bin_s1 ;
reg \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_4_U.carry_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_4_U.sum_s1 ;
reg [15:0] \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_5_U.ain_s1 ;
reg [15:0] \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_5_U.bin_s1 ;
reg \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_5_U.carry_s1 ;
reg [15:0] \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_5_U.sum_s1 ;
reg [15:0] \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_5_U.ain_s1 ;
reg [15:0] \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_5_U.bin_s1 ;
reg \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_5_U.carry_s1 ;
reg [15:0] \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_5_U.sum_s1 ;
reg [15:0] \add_32ns_32s_32_2_1_U6.top_add_32ns_32s_32_2_1_Adder_5_U.ain_s1 ;
reg [15:0] \add_32ns_32s_32_2_1_U6.top_add_32ns_32s_32_2_1_Adder_5_U.bin_s1 ;
reg \add_32ns_32s_32_2_1_U6.top_add_32ns_32s_32_2_1_Adder_5_U.carry_s1 ;
reg [15:0] \add_32ns_32s_32_2_1_U6.top_add_32ns_32s_32_2_1_Adder_5_U.sum_s1 ;
reg [15:0] \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_11_U.ain_s1 ;
reg [15:0] \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_11_U.bin_s1 ;
reg \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_11_U.carry_s1 ;
reg [15:0] \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_11_U.sum_s1 ;
reg [16:0] \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_13_U.ain_s1 ;
reg [16:0] \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_13_U.bin_s1 ;
reg \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_13_U.carry_s1 ;
reg [16:0] \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_13_U.sum_s1 ;
reg [16:0] \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_13_U.ain_s1 ;
reg [16:0] \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_13_U.bin_s1 ;
reg \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_13_U.carry_s1 ;
reg [16:0] \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_13_U.sum_s1 ;
reg [17:0] \add_36s_36s_36_2_1_U11.top_add_36s_36s_36_2_1_Adder_6_U.ain_s1 ;
reg [17:0] \add_36s_36s_36_2_1_U11.top_add_36s_36s_36_2_1_Adder_6_U.bin_s1 ;
reg \add_36s_36s_36_2_1_U11.top_add_36s_36s_36_2_1_Adder_6_U.carry_s1 ;
reg [17:0] \add_36s_36s_36_2_1_U11.top_add_36s_36s_36_2_1_Adder_6_U.sum_s1 ;
reg [17:0] \add_36s_36s_36_2_1_U7.top_add_36s_36s_36_2_1_Adder_6_U.ain_s1 ;
reg [17:0] \add_36s_36s_36_2_1_U7.top_add_36s_36s_36_2_1_Adder_6_U.bin_s1 ;
reg \add_36s_36s_36_2_1_U7.top_add_36s_36s_36_2_1_Adder_6_U.carry_s1 ;
reg [17:0] \add_36s_36s_36_2_1_U7.top_add_36s_36s_36_2_1_Adder_6_U.sum_s1 ;
reg [21:0] \add_44s_44s_44_2_1_U4.top_add_44s_44s_44_2_1_Adder_3_U.ain_s1 ;
reg [21:0] \add_44s_44s_44_2_1_U4.top_add_44s_44s_44_2_1_Adder_3_U.bin_s1 ;
reg \add_44s_44s_44_2_1_U4.top_add_44s_44s_44_2_1_Adder_3_U.carry_s1 ;
reg [21:0] \add_44s_44s_44_2_1_U4.top_add_44s_44s_44_2_1_Adder_3_U.sum_s1 ;
reg [1:0] \add_4ns_4ns_4_2_1_U19.top_add_4ns_4ns_4_2_1_Adder_12_U.ain_s1 ;
reg [1:0] \add_4ns_4ns_4_2_1_U19.top_add_4ns_4ns_4_2_1_Adder_12_U.bin_s1 ;
reg \add_4ns_4ns_4_2_1_U19.top_add_4ns_4ns_4_2_1_Adder_12_U.carry_s1 ;
reg [1:0] \add_4ns_4ns_4_2_1_U19.top_add_4ns_4ns_4_2_1_Adder_12_U.sum_s1 ;
reg [2:0] \add_5s_5ns_5_2_1_U1.top_add_5s_5ns_5_2_1_Adder_0_U.ain_s1 ;
reg [2:0] \add_5s_5ns_5_2_1_U1.top_add_5s_5ns_5_2_1_Adder_0_U.bin_s1 ;
reg \add_5s_5ns_5_2_1_U1.top_add_5s_5ns_5_2_1_Adder_0_U.carry_s1 ;
reg [1:0] \add_5s_5ns_5_2_1_U1.top_add_5s_5ns_5_2_1_Adder_0_U.sum_s1 ;
reg [3:0] \add_7s_7ns_7_2_1_U3.top_add_7s_7ns_7_2_1_Adder_2_U.ain_s1 ;
reg [3:0] \add_7s_7ns_7_2_1_U3.top_add_7s_7ns_7_2_1_Adder_2_U.bin_s1 ;
reg \add_7s_7ns_7_2_1_U3.top_add_7s_7ns_7_2_1_Adder_2_U.carry_s1 ;
reg [2:0] \add_7s_7ns_7_2_1_U3.top_add_7s_7ns_7_2_1_Adder_2_U.sum_s1 ;
reg [3:0] \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_8_U.ain_s1 ;
reg [3:0] \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_8_U.bin_s1 ;
reg \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_8_U.carry_s1 ;
reg [3:0] \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_8_U.sum_s1 ;
reg [3:0] \add_8s_8s_8_2_1_U15.top_add_8s_8s_8_2_1_Adder_9_U.ain_s1 ;
reg [3:0] \add_8s_8s_8_2_1_U15.top_add_8s_8s_8_2_1_Adder_9_U.bin_s1 ;
reg \add_8s_8s_8_2_1_U15.top_add_8s_8s_8_2_1_Adder_9_U.carry_s1 ;
reg [3:0] \add_8s_8s_8_2_1_U15.top_add_8s_8s_8_2_1_Adder_9_U.sum_s1 ;
reg [4:0] \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_1_U.ain_s1 ;
reg [4:0] \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_1_U.bin_s1 ;
reg \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_1_U.carry_s1 ;
reg [3:0] \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_1_U.sum_s1 ;
reg [4:0] \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_1_U.ain_s1 ;
reg [4:0] \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_1_U.bin_s1 ;
reg \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_1_U.carry_s1 ;
reg [3:0] \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_1_U.sum_s1 ;
reg [7:0] add_ln1192_1_reg_1246;
reg [31:0] add_ln691_1_reg_1060;
reg [31:0] add_ln691_2_reg_1107;
reg [31:0] add_ln691_3_reg_1189;
reg [31:0] add_ln691_4_reg_1373;
reg [31:0] add_ln691_5_reg_1431;
reg [6:0] add_ln691_reg_1023;
reg [9:0] add_ln69_reg_1276;
reg and_ln412_reg_1281;
reg and_ln786_reg_1367;
reg [42:0] ap_CS_fsm = 43'h00000000001;
reg carry_1_reg_1348;
reg deleted_zeros_reg_1361;
reg icmp_ln410_reg_1179;
reg icmp_ln851_1_reg_1043;
reg icmp_ln851_2_reg_1090;
reg icmp_ln851_3_reg_1147;
reg icmp_ln851_reg_1001;
reg [7:0] op_11_V_reg_1194;
reg [3:0] op_19_V_reg_1398;
reg [31:0] op_23_V_reg_1075;
reg [31:0] op_25_V_reg_1122;
reg [31:0] op_29_V_reg_1296;
reg or_ln340_reg_1378;
reg p_Result_11_reg_1251;
reg p_Result_13_reg_1265;
reg p_Result_14_reg_1312;
reg [3:0] p_Val2_4_reg_1260;
reg [3:0] p_Val2_5_reg_1306;
reg r_reg_1226;
reg [31:0] ret_V_14_cast_reg_1172;
reg [8:0] ret_V_15_reg_1006;
reg [43:0] ret_V_17_reg_1048;
reg [31:0] ret_V_18_reg_1065;
reg [35:0] ret_V_20_reg_1095;
reg [31:0] ret_V_21_cast_reg_1341;
reg [31:0] ret_V_21_reg_1112;
reg [35:0] ret_V_22_reg_1167;
reg [31:0] ret_V_23_reg_1206;
reg [31:0] ret_V_24_cast_reg_1424;
reg [31:0] ret_V_24_reg_1271;
reg [33:0] ret_V_25_reg_1336;
reg [31:0] ret_V_26_reg_1383;
reg [31:0] ret_V_27_reg_1404;
reg [33:0] ret_V_28_reg_1419;
reg [31:0] ret_V_4_cast_reg_1053;
reg [31:0] ret_V_8_cast_reg_1100;
reg [4:0] ret_reg_986;
reg [4:0] select_ln215_reg_976;
reg [3:0] select_ln340_reg_1388;
reg [6:0] select_ln353_reg_1028;
reg [6:0] sext_ln850_reg_1016;
reg [8:0] \sub_17s_17ns_17_2_1_U10.top_sub_17s_17ns_17_2_1_Adder_7_U.ain_s1 ;
reg [8:0] \sub_17s_17ns_17_2_1_U10.top_sub_17s_17ns_17_2_1_Adder_7_U.bin_s1 ;
reg \sub_17s_17ns_17_2_1_U10.top_sub_17s_17ns_17_2_1_Adder_7_U.carry_s1 ;
reg [7:0] \sub_17s_17ns_17_2_1_U10.top_sub_17s_17ns_17_2_1_Adder_7_U.sum_s1 ;
reg [5:0] tmp_1_reg_1011;
reg tmp_reg_1157;
reg trunc_ln410_reg_1162;
reg [2:0] trunc_ln718_reg_1201;
reg [7:0] trunc_ln_reg_1152;
reg xor_ln416_reg_1330;
wire _000_;
wire [7:0] _001_;
wire [31:0] _002_;
wire [31:0] _003_;
wire [31:0] _004_;
wire [31:0] _005_;
wire [31:0] _006_;
wire [6:0] _007_;
wire [9:0] _008_;
wire _009_;
wire _010_;
wire [42:0] _011_;
wire _012_;
wire _013_;
wire _014_;
wire _015_;
wire _016_;
wire _017_;
wire _018_;
wire [7:0] _019_;
wire [3:0] _020_;
wire [31:0] _021_;
wire [31:0] _022_;
wire [31:0] _023_;
wire _024_;
wire _025_;
wire _026_;
wire _027_;
wire [3:0] _028_;
wire [3:0] _029_;
wire _030_;
wire [31:0] _031_;
wire [8:0] _032_;
wire [43:0] _033_;
wire [31:0] _034_;
wire [35:0] _035_;
wire [31:0] _036_;
wire [31:0] _037_;
wire [35:0] _038_;
wire [31:0] _039_;
wire [31:0] _040_;
wire [31:0] _041_;
wire [33:0] _042_;
wire [31:0] _043_;
wire [31:0] _044_;
wire [33:0] _045_;
wire [31:0] _046_;
wire [31:0] _047_;
wire [4:0] _048_;
wire [4:0] _049_;
wire [3:0] _050_;
wire [6:0] _051_;
wire [6:0] _052_;
wire [5:0] _053_;
wire _054_;
wire _055_;
wire [2:0] _056_;
wire [7:0] _057_;
wire _058_;
wire [1:0] _059_;
wire _060_;
wire _061_;
wire _062_;
wire _063_;
wire _064_;
wire _065_;
wire _066_;
wire _067_;
wire [4:0] _068_;
wire [4:0] _069_;
wire _070_;
wire [4:0] _071_;
wire [5:0] _072_;
wire [5:0] _073_;
wire [15:0] _074_;
wire [15:0] _075_;
wire _076_;
wire [15:0] _077_;
wire [16:0] _078_;
wire [16:0] _079_;
wire [15:0] _080_;
wire [15:0] _081_;
wire _082_;
wire [15:0] _083_;
wire [16:0] _084_;
wire [16:0] _085_;
wire [15:0] _086_;
wire [15:0] _087_;
wire _088_;
wire [15:0] _089_;
wire [16:0] _090_;
wire [16:0] _091_;
wire [15:0] _092_;
wire [15:0] _093_;
wire _094_;
wire [15:0] _095_;
wire [16:0] _096_;
wire [16:0] _097_;
wire [15:0] _098_;
wire [15:0] _099_;
wire _100_;
wire [15:0] _101_;
wire [16:0] _102_;
wire [16:0] _103_;
wire [15:0] _104_;
wire [15:0] _105_;
wire _106_;
wire [15:0] _107_;
wire [16:0] _108_;
wire [16:0] _109_;
wire [15:0] _110_;
wire [15:0] _111_;
wire _112_;
wire [15:0] _113_;
wire [16:0] _114_;
wire [16:0] _115_;
wire [15:0] _116_;
wire [15:0] _117_;
wire _118_;
wire [15:0] _119_;
wire [16:0] _120_;
wire [16:0] _121_;
wire [15:0] _122_;
wire [15:0] _123_;
wire _124_;
wire [15:0] _125_;
wire [16:0] _126_;
wire [16:0] _127_;
wire [15:0] _128_;
wire [15:0] _129_;
wire _130_;
wire [15:0] _131_;
wire [16:0] _132_;
wire [16:0] _133_;
wire [16:0] _134_;
wire [16:0] _135_;
wire _136_;
wire [16:0] _137_;
wire [17:0] _138_;
wire [17:0] _139_;
wire [16:0] _140_;
wire [16:0] _141_;
wire _142_;
wire [16:0] _143_;
wire [17:0] _144_;
wire [17:0] _145_;
wire [17:0] _146_;
wire [17:0] _147_;
wire _148_;
wire [17:0] _149_;
wire [18:0] _150_;
wire [18:0] _151_;
wire [17:0] _152_;
wire [17:0] _153_;
wire _154_;
wire [17:0] _155_;
wire [18:0] _156_;
wire [18:0] _157_;
wire [21:0] _158_;
wire [21:0] _159_;
wire _160_;
wire [21:0] _161_;
wire [22:0] _162_;
wire [22:0] _163_;
wire [1:0] _164_;
wire [1:0] _165_;
wire _166_;
wire [1:0] _167_;
wire [2:0] _168_;
wire [2:0] _169_;
wire [2:0] _170_;
wire [2:0] _171_;
wire _172_;
wire [1:0] _173_;
wire [2:0] _174_;
wire [3:0] _175_;
wire [3:0] _176_;
wire [3:0] _177_;
wire _178_;
wire [2:0] _179_;
wire [3:0] _180_;
wire [4:0] _181_;
wire [3:0] _182_;
wire [3:0] _183_;
wire _184_;
wire [3:0] _185_;
wire [4:0] _186_;
wire [4:0] _187_;
wire [3:0] _188_;
wire [3:0] _189_;
wire _190_;
wire [3:0] _191_;
wire [4:0] _192_;
wire [4:0] _193_;
wire [4:0] _194_;
wire [4:0] _195_;
wire _196_;
wire [3:0] _197_;
wire [4:0] _198_;
wire [5:0] _199_;
wire [4:0] _200_;
wire [4:0] _201_;
wire _202_;
wire [3:0] _203_;
wire [4:0] _204_;
wire [5:0] _205_;
wire [8:0] _206_;
wire [8:0] _207_;
wire _208_;
wire [7:0] _209_;
wire [8:0] _210_;
wire [9:0] _211_;
wire _212_;
wire _213_;
wire _214_;
wire _215_;
wire _216_;
wire _217_;
wire _218_;
wire _219_;
wire _220_;
wire _221_;
wire _222_;
wire _223_;
wire _224_;
wire _225_;
wire _226_;
wire _227_;
wire _228_;
wire _229_;
wire _230_;
wire _231_;
wire _232_;
wire _233_;
wire _234_;
wire _235_;
wire _236_;
wire _237_;
wire _238_;
wire _239_;
wire _240_;
wire _241_;
wire _242_;
wire _243_;
wire _244_;
wire _245_;
wire _246_;
wire _247_;
wire _248_;
wire _249_;
wire _250_;
wire _251_;
wire _252_;
wire _253_;
wire _254_;
wire _255_;
wire _256_;
wire _257_;
wire _258_;
wire _259_;
wire Range1_all_zeros_fu_793_p2;
wire \add_10s_10ns_10_2_1_U17.ce ;
wire \add_10s_10ns_10_2_1_U17.clk ;
wire [9:0] \add_10s_10ns_10_2_1_U17.din0 ;
wire [9:0] \add_10s_10ns_10_2_1_U17.din1 ;
wire [9:0] \add_10s_10ns_10_2_1_U17.dout ;
wire \add_10s_10ns_10_2_1_U17.reset ;
wire [9:0] \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_10_U.a ;
wire [9:0] \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_10_U.ain_s0 ;
wire [9:0] \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_10_U.b ;
wire [9:0] \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_10_U.bin_s0 ;
wire \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_10_U.ce ;
wire \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_10_U.clk ;
wire \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_10_U.facout_s1 ;
wire \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_10_U.facout_s2 ;
wire [4:0] \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_10_U.fas_s1 ;
wire [4:0] \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_10_U.fas_s2 ;
wire \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_10_U.reset ;
wire [9:0] \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_10_U.s ;
wire [4:0] \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_10_U.u1.a ;
wire [4:0] \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_10_U.u1.b ;
wire \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_10_U.u1.cin ;
wire \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_10_U.u1.cout ;
wire [4:0] \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_10_U.u1.s ;
wire [4:0] \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_10_U.u2.a ;
wire [4:0] \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_10_U.u2.b ;
wire \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_10_U.u2.cin ;
wire \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_10_U.u2.cout ;
wire [4:0] \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_10_U.u2.s ;
wire \add_32ns_32ns_32_2_1_U12.ce ;
wire \add_32ns_32ns_32_2_1_U12.clk ;
wire [31:0] \add_32ns_32ns_32_2_1_U12.din0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U12.din1 ;
wire [31:0] \add_32ns_32ns_32_2_1_U12.dout ;
wire \add_32ns_32ns_32_2_1_U12.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_4_U.a ;
wire [31:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_4_U.ain_s0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_4_U.b ;
wire [31:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_4_U.bin_s0 ;
wire \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_4_U.ce ;
wire \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_4_U.clk ;
wire \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_4_U.facout_s1 ;
wire \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_4_U.facout_s2 ;
wire [15:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_4_U.fas_s1 ;
wire [15:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_4_U.fas_s2 ;
wire \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_4_U.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_4_U.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.b ;
wire \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.cin ;
wire \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.b ;
wire \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.cin ;
wire \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.s ;
wire \add_32ns_32ns_32_2_1_U21.ce ;
wire \add_32ns_32ns_32_2_1_U21.clk ;
wire [31:0] \add_32ns_32ns_32_2_1_U21.din0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U21.din1 ;
wire [31:0] \add_32ns_32ns_32_2_1_U21.dout ;
wire \add_32ns_32ns_32_2_1_U21.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_4_U.a ;
wire [31:0] \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_4_U.ain_s0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_4_U.b ;
wire [31:0] \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_4_U.bin_s0 ;
wire \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_4_U.ce ;
wire \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_4_U.clk ;
wire \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_4_U.facout_s1 ;
wire \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_4_U.facout_s2 ;
wire [15:0] \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_4_U.fas_s1 ;
wire [15:0] \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_4_U.fas_s2 ;
wire \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_4_U.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_4_U.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.b ;
wire \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.cin ;
wire \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.b ;
wire \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.cin ;
wire \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.s ;
wire \add_32ns_32ns_32_2_1_U24.ce ;
wire \add_32ns_32ns_32_2_1_U24.clk ;
wire [31:0] \add_32ns_32ns_32_2_1_U24.din0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U24.din1 ;
wire [31:0] \add_32ns_32ns_32_2_1_U24.dout ;
wire \add_32ns_32ns_32_2_1_U24.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_4_U.a ;
wire [31:0] \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_4_U.ain_s0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_4_U.b ;
wire [31:0] \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_4_U.bin_s0 ;
wire \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_4_U.ce ;
wire \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_4_U.clk ;
wire \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_4_U.facout_s1 ;
wire \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_4_U.facout_s2 ;
wire [15:0] \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_4_U.fas_s1 ;
wire [15:0] \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_4_U.fas_s2 ;
wire \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_4_U.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_4_U.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.b ;
wire \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.cin ;
wire \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.b ;
wire \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.cin ;
wire \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.s ;
wire \add_32ns_32ns_32_2_1_U5.ce ;
wire \add_32ns_32ns_32_2_1_U5.clk ;
wire [31:0] \add_32ns_32ns_32_2_1_U5.din0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U5.din1 ;
wire [31:0] \add_32ns_32ns_32_2_1_U5.dout ;
wire \add_32ns_32ns_32_2_1_U5.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.a ;
wire [31:0] \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.ain_s0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.b ;
wire [31:0] \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.bin_s0 ;
wire \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.ce ;
wire \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.clk ;
wire \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.facout_s1 ;
wire \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.facout_s2 ;
wire [15:0] \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.fas_s1 ;
wire [15:0] \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.fas_s2 ;
wire \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.b ;
wire \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.cin ;
wire \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.b ;
wire \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.cin ;
wire \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.s ;
wire \add_32ns_32ns_32_2_1_U8.ce ;
wire \add_32ns_32ns_32_2_1_U8.clk ;
wire [31:0] \add_32ns_32ns_32_2_1_U8.din0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U8.din1 ;
wire [31:0] \add_32ns_32ns_32_2_1_U8.dout ;
wire \add_32ns_32ns_32_2_1_U8.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.a ;
wire [31:0] \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.ain_s0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.b ;
wire [31:0] \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.bin_s0 ;
wire \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.ce ;
wire \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.clk ;
wire \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.facout_s1 ;
wire \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.facout_s2 ;
wire [15:0] \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.fas_s1 ;
wire [15:0] \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.fas_s2 ;
wire \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.b ;
wire \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.cin ;
wire \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.b ;
wire \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.cin ;
wire \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.s ;
wire \add_32ns_32ns_32_2_1_U9.ce ;
wire \add_32ns_32ns_32_2_1_U9.clk ;
wire [31:0] \add_32ns_32ns_32_2_1_U9.din0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U9.din1 ;
wire [31:0] \add_32ns_32ns_32_2_1_U9.dout ;
wire \add_32ns_32ns_32_2_1_U9.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_4_U.a ;
wire [31:0] \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_4_U.ain_s0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_4_U.b ;
wire [31:0] \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_4_U.bin_s0 ;
wire \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_4_U.ce ;
wire \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_4_U.clk ;
wire \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_4_U.facout_s1 ;
wire \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_4_U.facout_s2 ;
wire [15:0] \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_4_U.fas_s1 ;
wire [15:0] \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_4_U.fas_s2 ;
wire \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_4_U.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_4_U.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.b ;
wire \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.cin ;
wire \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.b ;
wire \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.cin ;
wire \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.s ;
wire \add_32ns_32s_32_2_1_U16.ce ;
wire \add_32ns_32s_32_2_1_U16.clk ;
wire [31:0] \add_32ns_32s_32_2_1_U16.din0 ;
wire [31:0] \add_32ns_32s_32_2_1_U16.din1 ;
wire [31:0] \add_32ns_32s_32_2_1_U16.dout ;
wire \add_32ns_32s_32_2_1_U16.reset ;
wire [31:0] \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_5_U.a ;
wire [31:0] \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_5_U.ain_s0 ;
wire [31:0] \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_5_U.b ;
wire [31:0] \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_5_U.bin_s0 ;
wire \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_5_U.ce ;
wire \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_5_U.clk ;
wire \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_5_U.facout_s1 ;
wire \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_5_U.facout_s2 ;
wire [15:0] \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_5_U.fas_s1 ;
wire [15:0] \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_5_U.fas_s2 ;
wire \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_5_U.reset ;
wire [31:0] \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_5_U.s ;
wire [15:0] \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_5_U.u1.a ;
wire [15:0] \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_5_U.u1.b ;
wire \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_5_U.u1.cin ;
wire \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_5_U.u1.cout ;
wire [15:0] \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_5_U.u1.s ;
wire [15:0] \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_5_U.u2.a ;
wire [15:0] \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_5_U.u2.b ;
wire \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_5_U.u2.cin ;
wire \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_5_U.u2.cout ;
wire [15:0] \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_5_U.u2.s ;
wire \add_32ns_32s_32_2_1_U22.ce ;
wire \add_32ns_32s_32_2_1_U22.clk ;
wire [31:0] \add_32ns_32s_32_2_1_U22.din0 ;
wire [31:0] \add_32ns_32s_32_2_1_U22.din1 ;
wire [31:0] \add_32ns_32s_32_2_1_U22.dout ;
wire \add_32ns_32s_32_2_1_U22.reset ;
wire [31:0] \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_5_U.a ;
wire [31:0] \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_5_U.ain_s0 ;
wire [31:0] \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_5_U.b ;
wire [31:0] \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_5_U.bin_s0 ;
wire \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_5_U.ce ;
wire \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_5_U.clk ;
wire \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_5_U.facout_s1 ;
wire \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_5_U.facout_s2 ;
wire [15:0] \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_5_U.fas_s1 ;
wire [15:0] \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_5_U.fas_s2 ;
wire \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_5_U.reset ;
wire [31:0] \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_5_U.s ;
wire [15:0] \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_5_U.u1.a ;
wire [15:0] \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_5_U.u1.b ;
wire \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_5_U.u1.cin ;
wire \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_5_U.u1.cout ;
wire [15:0] \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_5_U.u1.s ;
wire [15:0] \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_5_U.u2.a ;
wire [15:0] \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_5_U.u2.b ;
wire \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_5_U.u2.cin ;
wire \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_5_U.u2.cout ;
wire [15:0] \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_5_U.u2.s ;
wire \add_32ns_32s_32_2_1_U6.ce ;
wire \add_32ns_32s_32_2_1_U6.clk ;
wire [31:0] \add_32ns_32s_32_2_1_U6.din0 ;
wire [31:0] \add_32ns_32s_32_2_1_U6.din1 ;
wire [31:0] \add_32ns_32s_32_2_1_U6.dout ;
wire \add_32ns_32s_32_2_1_U6.reset ;
wire [31:0] \add_32ns_32s_32_2_1_U6.top_add_32ns_32s_32_2_1_Adder_5_U.a ;
wire [31:0] \add_32ns_32s_32_2_1_U6.top_add_32ns_32s_32_2_1_Adder_5_U.ain_s0 ;
wire [31:0] \add_32ns_32s_32_2_1_U6.top_add_32ns_32s_32_2_1_Adder_5_U.b ;
wire [31:0] \add_32ns_32s_32_2_1_U6.top_add_32ns_32s_32_2_1_Adder_5_U.bin_s0 ;
wire \add_32ns_32s_32_2_1_U6.top_add_32ns_32s_32_2_1_Adder_5_U.ce ;
wire \add_32ns_32s_32_2_1_U6.top_add_32ns_32s_32_2_1_Adder_5_U.clk ;
wire \add_32ns_32s_32_2_1_U6.top_add_32ns_32s_32_2_1_Adder_5_U.facout_s1 ;
wire \add_32ns_32s_32_2_1_U6.top_add_32ns_32s_32_2_1_Adder_5_U.facout_s2 ;
wire [15:0] \add_32ns_32s_32_2_1_U6.top_add_32ns_32s_32_2_1_Adder_5_U.fas_s1 ;
wire [15:0] \add_32ns_32s_32_2_1_U6.top_add_32ns_32s_32_2_1_Adder_5_U.fas_s2 ;
wire \add_32ns_32s_32_2_1_U6.top_add_32ns_32s_32_2_1_Adder_5_U.reset ;
wire [31:0] \add_32ns_32s_32_2_1_U6.top_add_32ns_32s_32_2_1_Adder_5_U.s ;
wire [15:0] \add_32ns_32s_32_2_1_U6.top_add_32ns_32s_32_2_1_Adder_5_U.u1.a ;
wire [15:0] \add_32ns_32s_32_2_1_U6.top_add_32ns_32s_32_2_1_Adder_5_U.u1.b ;
wire \add_32ns_32s_32_2_1_U6.top_add_32ns_32s_32_2_1_Adder_5_U.u1.cin ;
wire \add_32ns_32s_32_2_1_U6.top_add_32ns_32s_32_2_1_Adder_5_U.u1.cout ;
wire [15:0] \add_32ns_32s_32_2_1_U6.top_add_32ns_32s_32_2_1_Adder_5_U.u1.s ;
wire [15:0] \add_32ns_32s_32_2_1_U6.top_add_32ns_32s_32_2_1_Adder_5_U.u2.a ;
wire [15:0] \add_32ns_32s_32_2_1_U6.top_add_32ns_32s_32_2_1_Adder_5_U.u2.b ;
wire \add_32ns_32s_32_2_1_U6.top_add_32ns_32s_32_2_1_Adder_5_U.u2.cin ;
wire \add_32ns_32s_32_2_1_U6.top_add_32ns_32s_32_2_1_Adder_5_U.u2.cout ;
wire [15:0] \add_32ns_32s_32_2_1_U6.top_add_32ns_32s_32_2_1_Adder_5_U.u2.s ;
wire \add_32s_32ns_32_2_1_U18.ce ;
wire \add_32s_32ns_32_2_1_U18.clk ;
wire [31:0] \add_32s_32ns_32_2_1_U18.din0 ;
wire [31:0] \add_32s_32ns_32_2_1_U18.din1 ;
wire [31:0] \add_32s_32ns_32_2_1_U18.dout ;
wire \add_32s_32ns_32_2_1_U18.reset ;
wire [31:0] \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_11_U.a ;
wire [31:0] \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_11_U.ain_s0 ;
wire [31:0] \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_11_U.b ;
wire [31:0] \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_11_U.bin_s0 ;
wire \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_11_U.ce ;
wire \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_11_U.clk ;
wire \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_11_U.facout_s1 ;
wire \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_11_U.facout_s2 ;
wire [15:0] \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_11_U.fas_s1 ;
wire [15:0] \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_11_U.fas_s2 ;
wire \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_11_U.reset ;
wire [31:0] \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_11_U.s ;
wire [15:0] \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_11_U.u1.a ;
wire [15:0] \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_11_U.u1.b ;
wire \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_11_U.u1.cin ;
wire \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_11_U.u1.cout ;
wire [15:0] \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_11_U.u1.s ;
wire [15:0] \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_11_U.u2.a ;
wire [15:0] \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_11_U.u2.b ;
wire \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_11_U.u2.cin ;
wire \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_11_U.u2.cout ;
wire [15:0] \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_11_U.u2.s ;
wire \add_34s_34s_34_2_1_U20.ce ;
wire \add_34s_34s_34_2_1_U20.clk ;
wire [33:0] \add_34s_34s_34_2_1_U20.din0 ;
wire [33:0] \add_34s_34s_34_2_1_U20.din1 ;
wire [33:0] \add_34s_34s_34_2_1_U20.dout ;
wire \add_34s_34s_34_2_1_U20.reset ;
wire [33:0] \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_13_U.a ;
wire [33:0] \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_13_U.ain_s0 ;
wire [33:0] \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_13_U.b ;
wire [33:0] \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_13_U.bin_s0 ;
wire \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_13_U.ce ;
wire \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_13_U.clk ;
wire \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_13_U.facout_s1 ;
wire \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_13_U.facout_s2 ;
wire [16:0] \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_13_U.fas_s1 ;
wire [16:0] \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_13_U.fas_s2 ;
wire \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_13_U.reset ;
wire [33:0] \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_13_U.s ;
wire [16:0] \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_13_U.u1.a ;
wire [16:0] \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_13_U.u1.b ;
wire \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_13_U.u1.cin ;
wire \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_13_U.u1.cout ;
wire [16:0] \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_13_U.u1.s ;
wire [16:0] \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_13_U.u2.a ;
wire [16:0] \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_13_U.u2.b ;
wire \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_13_U.u2.cin ;
wire \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_13_U.u2.cout ;
wire [16:0] \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_13_U.u2.s ;
wire \add_34s_34s_34_2_1_U23.ce ;
wire \add_34s_34s_34_2_1_U23.clk ;
wire [33:0] \add_34s_34s_34_2_1_U23.din0 ;
wire [33:0] \add_34s_34s_34_2_1_U23.din1 ;
wire [33:0] \add_34s_34s_34_2_1_U23.dout ;
wire \add_34s_34s_34_2_1_U23.reset ;
wire [33:0] \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_13_U.a ;
wire [33:0] \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_13_U.ain_s0 ;
wire [33:0] \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_13_U.b ;
wire [33:0] \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_13_U.bin_s0 ;
wire \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_13_U.ce ;
wire \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_13_U.clk ;
wire \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_13_U.facout_s1 ;
wire \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_13_U.facout_s2 ;
wire [16:0] \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_13_U.fas_s1 ;
wire [16:0] \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_13_U.fas_s2 ;
wire \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_13_U.reset ;
wire [33:0] \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_13_U.s ;
wire [16:0] \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_13_U.u1.a ;
wire [16:0] \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_13_U.u1.b ;
wire \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_13_U.u1.cin ;
wire \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_13_U.u1.cout ;
wire [16:0] \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_13_U.u1.s ;
wire [16:0] \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_13_U.u2.a ;
wire [16:0] \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_13_U.u2.b ;
wire \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_13_U.u2.cin ;
wire \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_13_U.u2.cout ;
wire [16:0] \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_13_U.u2.s ;
wire \add_36s_36s_36_2_1_U11.ce ;
wire \add_36s_36s_36_2_1_U11.clk ;
wire [35:0] \add_36s_36s_36_2_1_U11.din0 ;
wire [35:0] \add_36s_36s_36_2_1_U11.din1 ;
wire [35:0] \add_36s_36s_36_2_1_U11.dout ;
wire \add_36s_36s_36_2_1_U11.reset ;
wire [35:0] \add_36s_36s_36_2_1_U11.top_add_36s_36s_36_2_1_Adder_6_U.a ;
wire [35:0] \add_36s_36s_36_2_1_U11.top_add_36s_36s_36_2_1_Adder_6_U.ain_s0 ;
wire [35:0] \add_36s_36s_36_2_1_U11.top_add_36s_36s_36_2_1_Adder_6_U.b ;
wire [35:0] \add_36s_36s_36_2_1_U11.top_add_36s_36s_36_2_1_Adder_6_U.bin_s0 ;
wire \add_36s_36s_36_2_1_U11.top_add_36s_36s_36_2_1_Adder_6_U.ce ;
wire \add_36s_36s_36_2_1_U11.top_add_36s_36s_36_2_1_Adder_6_U.clk ;
wire \add_36s_36s_36_2_1_U11.top_add_36s_36s_36_2_1_Adder_6_U.facout_s1 ;
wire \add_36s_36s_36_2_1_U11.top_add_36s_36s_36_2_1_Adder_6_U.facout_s2 ;
wire [17:0] \add_36s_36s_36_2_1_U11.top_add_36s_36s_36_2_1_Adder_6_U.fas_s1 ;
wire [17:0] \add_36s_36s_36_2_1_U11.top_add_36s_36s_36_2_1_Adder_6_U.fas_s2 ;
wire \add_36s_36s_36_2_1_U11.top_add_36s_36s_36_2_1_Adder_6_U.reset ;
wire [35:0] \add_36s_36s_36_2_1_U11.top_add_36s_36s_36_2_1_Adder_6_U.s ;
wire [17:0] \add_36s_36s_36_2_1_U11.top_add_36s_36s_36_2_1_Adder_6_U.u1.a ;
wire [17:0] \add_36s_36s_36_2_1_U11.top_add_36s_36s_36_2_1_Adder_6_U.u1.b ;
wire \add_36s_36s_36_2_1_U11.top_add_36s_36s_36_2_1_Adder_6_U.u1.cin ;
wire \add_36s_36s_36_2_1_U11.top_add_36s_36s_36_2_1_Adder_6_U.u1.cout ;
wire [17:0] \add_36s_36s_36_2_1_U11.top_add_36s_36s_36_2_1_Adder_6_U.u1.s ;
wire [17:0] \add_36s_36s_36_2_1_U11.top_add_36s_36s_36_2_1_Adder_6_U.u2.a ;
wire [17:0] \add_36s_36s_36_2_1_U11.top_add_36s_36s_36_2_1_Adder_6_U.u2.b ;
wire \add_36s_36s_36_2_1_U11.top_add_36s_36s_36_2_1_Adder_6_U.u2.cin ;
wire \add_36s_36s_36_2_1_U11.top_add_36s_36s_36_2_1_Adder_6_U.u2.cout ;
wire [17:0] \add_36s_36s_36_2_1_U11.top_add_36s_36s_36_2_1_Adder_6_U.u2.s ;
wire \add_36s_36s_36_2_1_U7.ce ;
wire \add_36s_36s_36_2_1_U7.clk ;
wire [35:0] \add_36s_36s_36_2_1_U7.din0 ;
wire [35:0] \add_36s_36s_36_2_1_U7.din1 ;
wire [35:0] \add_36s_36s_36_2_1_U7.dout ;
wire \add_36s_36s_36_2_1_U7.reset ;
wire [35:0] \add_36s_36s_36_2_1_U7.top_add_36s_36s_36_2_1_Adder_6_U.a ;
wire [35:0] \add_36s_36s_36_2_1_U7.top_add_36s_36s_36_2_1_Adder_6_U.ain_s0 ;
wire [35:0] \add_36s_36s_36_2_1_U7.top_add_36s_36s_36_2_1_Adder_6_U.b ;
wire [35:0] \add_36s_36s_36_2_1_U7.top_add_36s_36s_36_2_1_Adder_6_U.bin_s0 ;
wire \add_36s_36s_36_2_1_U7.top_add_36s_36s_36_2_1_Adder_6_U.ce ;
wire \add_36s_36s_36_2_1_U7.top_add_36s_36s_36_2_1_Adder_6_U.clk ;
wire \add_36s_36s_36_2_1_U7.top_add_36s_36s_36_2_1_Adder_6_U.facout_s1 ;
wire \add_36s_36s_36_2_1_U7.top_add_36s_36s_36_2_1_Adder_6_U.facout_s2 ;
wire [17:0] \add_36s_36s_36_2_1_U7.top_add_36s_36s_36_2_1_Adder_6_U.fas_s1 ;
wire [17:0] \add_36s_36s_36_2_1_U7.top_add_36s_36s_36_2_1_Adder_6_U.fas_s2 ;
wire \add_36s_36s_36_2_1_U7.top_add_36s_36s_36_2_1_Adder_6_U.reset ;
wire [35:0] \add_36s_36s_36_2_1_U7.top_add_36s_36s_36_2_1_Adder_6_U.s ;
wire [17:0] \add_36s_36s_36_2_1_U7.top_add_36s_36s_36_2_1_Adder_6_U.u1.a ;
wire [17:0] \add_36s_36s_36_2_1_U7.top_add_36s_36s_36_2_1_Adder_6_U.u1.b ;
wire \add_36s_36s_36_2_1_U7.top_add_36s_36s_36_2_1_Adder_6_U.u1.cin ;
wire \add_36s_36s_36_2_1_U7.top_add_36s_36s_36_2_1_Adder_6_U.u1.cout ;
wire [17:0] \add_36s_36s_36_2_1_U7.top_add_36s_36s_36_2_1_Adder_6_U.u1.s ;
wire [17:0] \add_36s_36s_36_2_1_U7.top_add_36s_36s_36_2_1_Adder_6_U.u2.a ;
wire [17:0] \add_36s_36s_36_2_1_U7.top_add_36s_36s_36_2_1_Adder_6_U.u2.b ;
wire \add_36s_36s_36_2_1_U7.top_add_36s_36s_36_2_1_Adder_6_U.u2.cin ;
wire \add_36s_36s_36_2_1_U7.top_add_36s_36s_36_2_1_Adder_6_U.u2.cout ;
wire [17:0] \add_36s_36s_36_2_1_U7.top_add_36s_36s_36_2_1_Adder_6_U.u2.s ;
wire \add_44s_44s_44_2_1_U4.ce ;
wire \add_44s_44s_44_2_1_U4.clk ;
wire [43:0] \add_44s_44s_44_2_1_U4.din0 ;
wire [43:0] \add_44s_44s_44_2_1_U4.din1 ;
wire [43:0] \add_44s_44s_44_2_1_U4.dout ;
wire \add_44s_44s_44_2_1_U4.reset ;
wire [43:0] \add_44s_44s_44_2_1_U4.top_add_44s_44s_44_2_1_Adder_3_U.a ;
wire [43:0] \add_44s_44s_44_2_1_U4.top_add_44s_44s_44_2_1_Adder_3_U.ain_s0 ;
wire [43:0] \add_44s_44s_44_2_1_U4.top_add_44s_44s_44_2_1_Adder_3_U.b ;
wire [43:0] \add_44s_44s_44_2_1_U4.top_add_44s_44s_44_2_1_Adder_3_U.bin_s0 ;
wire \add_44s_44s_44_2_1_U4.top_add_44s_44s_44_2_1_Adder_3_U.ce ;
wire \add_44s_44s_44_2_1_U4.top_add_44s_44s_44_2_1_Adder_3_U.clk ;
wire \add_44s_44s_44_2_1_U4.top_add_44s_44s_44_2_1_Adder_3_U.facout_s1 ;
wire \add_44s_44s_44_2_1_U4.top_add_44s_44s_44_2_1_Adder_3_U.facout_s2 ;
wire [21:0] \add_44s_44s_44_2_1_U4.top_add_44s_44s_44_2_1_Adder_3_U.fas_s1 ;
wire [21:0] \add_44s_44s_44_2_1_U4.top_add_44s_44s_44_2_1_Adder_3_U.fas_s2 ;
wire \add_44s_44s_44_2_1_U4.top_add_44s_44s_44_2_1_Adder_3_U.reset ;
wire [43:0] \add_44s_44s_44_2_1_U4.top_add_44s_44s_44_2_1_Adder_3_U.s ;
wire [21:0] \add_44s_44s_44_2_1_U4.top_add_44s_44s_44_2_1_Adder_3_U.u1.a ;
wire [21:0] \add_44s_44s_44_2_1_U4.top_add_44s_44s_44_2_1_Adder_3_U.u1.b ;
wire \add_44s_44s_44_2_1_U4.top_add_44s_44s_44_2_1_Adder_3_U.u1.cin ;
wire \add_44s_44s_44_2_1_U4.top_add_44s_44s_44_2_1_Adder_3_U.u1.cout ;
wire [21:0] \add_44s_44s_44_2_1_U4.top_add_44s_44s_44_2_1_Adder_3_U.u1.s ;
wire [21:0] \add_44s_44s_44_2_1_U4.top_add_44s_44s_44_2_1_Adder_3_U.u2.a ;
wire [21:0] \add_44s_44s_44_2_1_U4.top_add_44s_44s_44_2_1_Adder_3_U.u2.b ;
wire \add_44s_44s_44_2_1_U4.top_add_44s_44s_44_2_1_Adder_3_U.u2.cin ;
wire \add_44s_44s_44_2_1_U4.top_add_44s_44s_44_2_1_Adder_3_U.u2.cout ;
wire [21:0] \add_44s_44s_44_2_1_U4.top_add_44s_44s_44_2_1_Adder_3_U.u2.s ;
wire \add_4ns_4ns_4_2_1_U19.ce ;
wire \add_4ns_4ns_4_2_1_U19.clk ;
wire [3:0] \add_4ns_4ns_4_2_1_U19.din0 ;
wire [3:0] \add_4ns_4ns_4_2_1_U19.din1 ;
wire [3:0] \add_4ns_4ns_4_2_1_U19.dout ;
wire \add_4ns_4ns_4_2_1_U19.reset ;
wire [3:0] \add_4ns_4ns_4_2_1_U19.top_add_4ns_4ns_4_2_1_Adder_12_U.a ;
wire [3:0] \add_4ns_4ns_4_2_1_U19.top_add_4ns_4ns_4_2_1_Adder_12_U.ain_s0 ;
wire [3:0] \add_4ns_4ns_4_2_1_U19.top_add_4ns_4ns_4_2_1_Adder_12_U.b ;
wire [3:0] \add_4ns_4ns_4_2_1_U19.top_add_4ns_4ns_4_2_1_Adder_12_U.bin_s0 ;
wire \add_4ns_4ns_4_2_1_U19.top_add_4ns_4ns_4_2_1_Adder_12_U.ce ;
wire \add_4ns_4ns_4_2_1_U19.top_add_4ns_4ns_4_2_1_Adder_12_U.clk ;
wire \add_4ns_4ns_4_2_1_U19.top_add_4ns_4ns_4_2_1_Adder_12_U.facout_s1 ;
wire \add_4ns_4ns_4_2_1_U19.top_add_4ns_4ns_4_2_1_Adder_12_U.facout_s2 ;
wire [1:0] \add_4ns_4ns_4_2_1_U19.top_add_4ns_4ns_4_2_1_Adder_12_U.fas_s1 ;
wire [1:0] \add_4ns_4ns_4_2_1_U19.top_add_4ns_4ns_4_2_1_Adder_12_U.fas_s2 ;
wire \add_4ns_4ns_4_2_1_U19.top_add_4ns_4ns_4_2_1_Adder_12_U.reset ;
wire [3:0] \add_4ns_4ns_4_2_1_U19.top_add_4ns_4ns_4_2_1_Adder_12_U.s ;
wire [1:0] \add_4ns_4ns_4_2_1_U19.top_add_4ns_4ns_4_2_1_Adder_12_U.u1.a ;
wire [1:0] \add_4ns_4ns_4_2_1_U19.top_add_4ns_4ns_4_2_1_Adder_12_U.u1.b ;
wire \add_4ns_4ns_4_2_1_U19.top_add_4ns_4ns_4_2_1_Adder_12_U.u1.cin ;
wire \add_4ns_4ns_4_2_1_U19.top_add_4ns_4ns_4_2_1_Adder_12_U.u1.cout ;
wire [1:0] \add_4ns_4ns_4_2_1_U19.top_add_4ns_4ns_4_2_1_Adder_12_U.u1.s ;
wire [1:0] \add_4ns_4ns_4_2_1_U19.top_add_4ns_4ns_4_2_1_Adder_12_U.u2.a ;
wire [1:0] \add_4ns_4ns_4_2_1_U19.top_add_4ns_4ns_4_2_1_Adder_12_U.u2.b ;
wire \add_4ns_4ns_4_2_1_U19.top_add_4ns_4ns_4_2_1_Adder_12_U.u2.cin ;
wire \add_4ns_4ns_4_2_1_U19.top_add_4ns_4ns_4_2_1_Adder_12_U.u2.cout ;
wire [1:0] \add_4ns_4ns_4_2_1_U19.top_add_4ns_4ns_4_2_1_Adder_12_U.u2.s ;
wire \add_5s_5ns_5_2_1_U1.ce ;
wire \add_5s_5ns_5_2_1_U1.clk ;
wire [4:0] \add_5s_5ns_5_2_1_U1.din0 ;
wire [4:0] \add_5s_5ns_5_2_1_U1.din1 ;
wire [4:0] \add_5s_5ns_5_2_1_U1.dout ;
wire \add_5s_5ns_5_2_1_U1.reset ;
wire [4:0] \add_5s_5ns_5_2_1_U1.top_add_5s_5ns_5_2_1_Adder_0_U.a ;
wire [4:0] \add_5s_5ns_5_2_1_U1.top_add_5s_5ns_5_2_1_Adder_0_U.ain_s0 ;
wire [4:0] \add_5s_5ns_5_2_1_U1.top_add_5s_5ns_5_2_1_Adder_0_U.b ;
wire [4:0] \add_5s_5ns_5_2_1_U1.top_add_5s_5ns_5_2_1_Adder_0_U.bin_s0 ;
wire \add_5s_5ns_5_2_1_U1.top_add_5s_5ns_5_2_1_Adder_0_U.ce ;
wire \add_5s_5ns_5_2_1_U1.top_add_5s_5ns_5_2_1_Adder_0_U.clk ;
wire \add_5s_5ns_5_2_1_U1.top_add_5s_5ns_5_2_1_Adder_0_U.facout_s1 ;
wire \add_5s_5ns_5_2_1_U1.top_add_5s_5ns_5_2_1_Adder_0_U.facout_s2 ;
wire [1:0] \add_5s_5ns_5_2_1_U1.top_add_5s_5ns_5_2_1_Adder_0_U.fas_s1 ;
wire [2:0] \add_5s_5ns_5_2_1_U1.top_add_5s_5ns_5_2_1_Adder_0_U.fas_s2 ;
wire \add_5s_5ns_5_2_1_U1.top_add_5s_5ns_5_2_1_Adder_0_U.reset ;
wire [4:0] \add_5s_5ns_5_2_1_U1.top_add_5s_5ns_5_2_1_Adder_0_U.s ;
wire [1:0] \add_5s_5ns_5_2_1_U1.top_add_5s_5ns_5_2_1_Adder_0_U.u1.a ;
wire [1:0] \add_5s_5ns_5_2_1_U1.top_add_5s_5ns_5_2_1_Adder_0_U.u1.b ;
wire \add_5s_5ns_5_2_1_U1.top_add_5s_5ns_5_2_1_Adder_0_U.u1.cin ;
wire \add_5s_5ns_5_2_1_U1.top_add_5s_5ns_5_2_1_Adder_0_U.u1.cout ;
wire [1:0] \add_5s_5ns_5_2_1_U1.top_add_5s_5ns_5_2_1_Adder_0_U.u1.s ;
wire [2:0] \add_5s_5ns_5_2_1_U1.top_add_5s_5ns_5_2_1_Adder_0_U.u2.a ;
wire [2:0] \add_5s_5ns_5_2_1_U1.top_add_5s_5ns_5_2_1_Adder_0_U.u2.b ;
wire \add_5s_5ns_5_2_1_U1.top_add_5s_5ns_5_2_1_Adder_0_U.u2.cin ;
wire \add_5s_5ns_5_2_1_U1.top_add_5s_5ns_5_2_1_Adder_0_U.u2.cout ;
wire [2:0] \add_5s_5ns_5_2_1_U1.top_add_5s_5ns_5_2_1_Adder_0_U.u2.s ;
wire \add_7s_7ns_7_2_1_U3.ce ;
wire \add_7s_7ns_7_2_1_U3.clk ;
wire [6:0] \add_7s_7ns_7_2_1_U3.din0 ;
wire [6:0] \add_7s_7ns_7_2_1_U3.din1 ;
wire [6:0] \add_7s_7ns_7_2_1_U3.dout ;
wire \add_7s_7ns_7_2_1_U3.reset ;
wire [6:0] \add_7s_7ns_7_2_1_U3.top_add_7s_7ns_7_2_1_Adder_2_U.a ;
wire [6:0] \add_7s_7ns_7_2_1_U3.top_add_7s_7ns_7_2_1_Adder_2_U.ain_s0 ;
wire [6:0] \add_7s_7ns_7_2_1_U3.top_add_7s_7ns_7_2_1_Adder_2_U.b ;
wire [6:0] \add_7s_7ns_7_2_1_U3.top_add_7s_7ns_7_2_1_Adder_2_U.bin_s0 ;
wire \add_7s_7ns_7_2_1_U3.top_add_7s_7ns_7_2_1_Adder_2_U.ce ;
wire \add_7s_7ns_7_2_1_U3.top_add_7s_7ns_7_2_1_Adder_2_U.clk ;
wire \add_7s_7ns_7_2_1_U3.top_add_7s_7ns_7_2_1_Adder_2_U.facout_s1 ;
wire \add_7s_7ns_7_2_1_U3.top_add_7s_7ns_7_2_1_Adder_2_U.facout_s2 ;
wire [2:0] \add_7s_7ns_7_2_1_U3.top_add_7s_7ns_7_2_1_Adder_2_U.fas_s1 ;
wire [3:0] \add_7s_7ns_7_2_1_U3.top_add_7s_7ns_7_2_1_Adder_2_U.fas_s2 ;
wire \add_7s_7ns_7_2_1_U3.top_add_7s_7ns_7_2_1_Adder_2_U.reset ;
wire [6:0] \add_7s_7ns_7_2_1_U3.top_add_7s_7ns_7_2_1_Adder_2_U.s ;
wire [2:0] \add_7s_7ns_7_2_1_U3.top_add_7s_7ns_7_2_1_Adder_2_U.u1.a ;
wire [2:0] \add_7s_7ns_7_2_1_U3.top_add_7s_7ns_7_2_1_Adder_2_U.u1.b ;
wire \add_7s_7ns_7_2_1_U3.top_add_7s_7ns_7_2_1_Adder_2_U.u1.cin ;
wire \add_7s_7ns_7_2_1_U3.top_add_7s_7ns_7_2_1_Adder_2_U.u1.cout ;
wire [2:0] \add_7s_7ns_7_2_1_U3.top_add_7s_7ns_7_2_1_Adder_2_U.u1.s ;
wire [3:0] \add_7s_7ns_7_2_1_U3.top_add_7s_7ns_7_2_1_Adder_2_U.u2.a ;
wire [3:0] \add_7s_7ns_7_2_1_U3.top_add_7s_7ns_7_2_1_Adder_2_U.u2.b ;
wire \add_7s_7ns_7_2_1_U3.top_add_7s_7ns_7_2_1_Adder_2_U.u2.cin ;
wire \add_7s_7ns_7_2_1_U3.top_add_7s_7ns_7_2_1_Adder_2_U.u2.cout ;
wire [3:0] \add_7s_7ns_7_2_1_U3.top_add_7s_7ns_7_2_1_Adder_2_U.u2.s ;
wire \add_8ns_8ns_8_2_1_U13.ce ;
wire \add_8ns_8ns_8_2_1_U13.clk ;
wire [7:0] \add_8ns_8ns_8_2_1_U13.din0 ;
wire [7:0] \add_8ns_8ns_8_2_1_U13.din1 ;
wire [7:0] \add_8ns_8ns_8_2_1_U13.dout ;
wire \add_8ns_8ns_8_2_1_U13.reset ;
wire [7:0] \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_8_U.a ;
wire [7:0] \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_8_U.ain_s0 ;
wire [7:0] \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_8_U.b ;
wire [7:0] \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_8_U.bin_s0 ;
wire \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_8_U.ce ;
wire \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_8_U.clk ;
wire \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_8_U.facout_s1 ;
wire \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_8_U.facout_s2 ;
wire [3:0] \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_8_U.fas_s1 ;
wire [3:0] \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_8_U.fas_s2 ;
wire \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_8_U.reset ;
wire [7:0] \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_8_U.s ;
wire [3:0] \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_8_U.u1.a ;
wire [3:0] \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_8_U.u1.b ;
wire \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_8_U.u1.cin ;
wire \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_8_U.u1.cout ;
wire [3:0] \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_8_U.u1.s ;
wire [3:0] \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_8_U.u2.a ;
wire [3:0] \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_8_U.u2.b ;
wire \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_8_U.u2.cin ;
wire \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_8_U.u2.cout ;
wire [3:0] \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_8_U.u2.s ;
wire \add_8s_8s_8_2_1_U15.ce ;
wire \add_8s_8s_8_2_1_U15.clk ;
wire [7:0] \add_8s_8s_8_2_1_U15.din0 ;
wire [7:0] \add_8s_8s_8_2_1_U15.din1 ;
wire [7:0] \add_8s_8s_8_2_1_U15.dout ;
wire \add_8s_8s_8_2_1_U15.reset ;
wire [7:0] \add_8s_8s_8_2_1_U15.top_add_8s_8s_8_2_1_Adder_9_U.a ;
wire [7:0] \add_8s_8s_8_2_1_U15.top_add_8s_8s_8_2_1_Adder_9_U.ain_s0 ;
wire [7:0] \add_8s_8s_8_2_1_U15.top_add_8s_8s_8_2_1_Adder_9_U.b ;
wire [7:0] \add_8s_8s_8_2_1_U15.top_add_8s_8s_8_2_1_Adder_9_U.bin_s0 ;
wire \add_8s_8s_8_2_1_U15.top_add_8s_8s_8_2_1_Adder_9_U.ce ;
wire \add_8s_8s_8_2_1_U15.top_add_8s_8s_8_2_1_Adder_9_U.clk ;
wire \add_8s_8s_8_2_1_U15.top_add_8s_8s_8_2_1_Adder_9_U.facout_s1 ;
wire \add_8s_8s_8_2_1_U15.top_add_8s_8s_8_2_1_Adder_9_U.facout_s2 ;
wire [3:0] \add_8s_8s_8_2_1_U15.top_add_8s_8s_8_2_1_Adder_9_U.fas_s1 ;
wire [3:0] \add_8s_8s_8_2_1_U15.top_add_8s_8s_8_2_1_Adder_9_U.fas_s2 ;
wire \add_8s_8s_8_2_1_U15.top_add_8s_8s_8_2_1_Adder_9_U.reset ;
wire [7:0] \add_8s_8s_8_2_1_U15.top_add_8s_8s_8_2_1_Adder_9_U.s ;
wire [3:0] \add_8s_8s_8_2_1_U15.top_add_8s_8s_8_2_1_Adder_9_U.u1.a ;
wire [3:0] \add_8s_8s_8_2_1_U15.top_add_8s_8s_8_2_1_Adder_9_U.u1.b ;
wire \add_8s_8s_8_2_1_U15.top_add_8s_8s_8_2_1_Adder_9_U.u1.cin ;
wire \add_8s_8s_8_2_1_U15.top_add_8s_8s_8_2_1_Adder_9_U.u1.cout ;
wire [3:0] \add_8s_8s_8_2_1_U15.top_add_8s_8s_8_2_1_Adder_9_U.u1.s ;
wire [3:0] \add_8s_8s_8_2_1_U15.top_add_8s_8s_8_2_1_Adder_9_U.u2.a ;
wire [3:0] \add_8s_8s_8_2_1_U15.top_add_8s_8s_8_2_1_Adder_9_U.u2.b ;
wire \add_8s_8s_8_2_1_U15.top_add_8s_8s_8_2_1_Adder_9_U.u2.cin ;
wire \add_8s_8s_8_2_1_U15.top_add_8s_8s_8_2_1_Adder_9_U.u2.cout ;
wire [3:0] \add_8s_8s_8_2_1_U15.top_add_8s_8s_8_2_1_Adder_9_U.u2.s ;
wire \add_9s_9s_9_2_1_U14.ce ;
wire \add_9s_9s_9_2_1_U14.clk ;
wire [8:0] \add_9s_9s_9_2_1_U14.din0 ;
wire [8:0] \add_9s_9s_9_2_1_U14.din1 ;
wire [8:0] \add_9s_9s_9_2_1_U14.dout ;
wire \add_9s_9s_9_2_1_U14.reset ;
wire [8:0] \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_1_U.a ;
wire [8:0] \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_1_U.ain_s0 ;
wire [8:0] \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_1_U.b ;
wire [8:0] \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_1_U.bin_s0 ;
wire \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_1_U.ce ;
wire \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_1_U.clk ;
wire \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_1_U.facout_s1 ;
wire \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_1_U.facout_s2 ;
wire [3:0] \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_1_U.fas_s1 ;
wire [4:0] \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_1_U.fas_s2 ;
wire \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_1_U.reset ;
wire [8:0] \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_1_U.s ;
wire [3:0] \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_1_U.u1.a ;
wire [3:0] \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_1_U.u1.b ;
wire \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_1_U.u1.cin ;
wire \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_1_U.u1.cout ;
wire [3:0] \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_1_U.u1.s ;
wire [4:0] \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_1_U.u2.a ;
wire [4:0] \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_1_U.u2.b ;
wire \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_1_U.u2.cin ;
wire \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_1_U.u2.cout ;
wire [4:0] \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_1_U.u2.s ;
wire \add_9s_9s_9_2_1_U2.ce ;
wire \add_9s_9s_9_2_1_U2.clk ;
wire [8:0] \add_9s_9s_9_2_1_U2.din0 ;
wire [8:0] \add_9s_9s_9_2_1_U2.din1 ;
wire [8:0] \add_9s_9s_9_2_1_U2.dout ;
wire \add_9s_9s_9_2_1_U2.reset ;
wire [8:0] \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_1_U.a ;
wire [8:0] \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_1_U.ain_s0 ;
wire [8:0] \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_1_U.b ;
wire [8:0] \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_1_U.bin_s0 ;
wire \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_1_U.ce ;
wire \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_1_U.clk ;
wire \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_1_U.facout_s1 ;
wire \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_1_U.facout_s2 ;
wire [3:0] \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_1_U.fas_s1 ;
wire [4:0] \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_1_U.fas_s2 ;
wire \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_1_U.reset ;
wire [8:0] \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_1_U.s ;
wire [3:0] \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_1_U.u1.a ;
wire [3:0] \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_1_U.u1.b ;
wire \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_1_U.u1.cin ;
wire \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_1_U.u1.cout ;
wire [3:0] \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_1_U.u1.s ;
wire [4:0] \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_1_U.u2.a ;
wire [4:0] \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_1_U.u2.b ;
wire \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_1_U.u2.cin ;
wire \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_1_U.u2.cout ;
wire [4:0] \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_1_U.u2.s ;
wire and_ln412_fu_723_p2;
wire and_ln785_1_fu_906_p2;
wire and_ln785_fu_897_p2;
wire and_ln786_fu_813_p2;
wire [16:0] and_ln_fu_570_p4;
wire ap_CS_fsm_state1;
wire ap_CS_fsm_state10;
wire ap_CS_fsm_state11;
wire ap_CS_fsm_state12;
wire ap_CS_fsm_state13;
wire ap_CS_fsm_state14;
wire ap_CS_fsm_state15;
wire ap_CS_fsm_state16;
wire ap_CS_fsm_state17;
wire ap_CS_fsm_state18;
wire ap_CS_fsm_state19;
wire ap_CS_fsm_state2;
wire ap_CS_fsm_state20;
wire ap_CS_fsm_state21;
wire ap_CS_fsm_state22;
wire ap_CS_fsm_state23;
wire ap_CS_fsm_state24;
wire ap_CS_fsm_state25;
wire ap_CS_fsm_state26;
wire ap_CS_fsm_state27;
wire ap_CS_fsm_state28;
wire ap_CS_fsm_state29;
wire ap_CS_fsm_state3;
wire ap_CS_fsm_state30;
wire ap_CS_fsm_state31;
wire ap_CS_fsm_state32;
wire ap_CS_fsm_state33;
wire ap_CS_fsm_state34;
wire ap_CS_fsm_state35;
wire ap_CS_fsm_state36;
wire ap_CS_fsm_state37;
wire ap_CS_fsm_state38;
wire ap_CS_fsm_state39;
wire ap_CS_fsm_state4;
wire ap_CS_fsm_state40;
wire ap_CS_fsm_state41;
wire ap_CS_fsm_state42;
wire ap_CS_fsm_state43;
wire ap_CS_fsm_state5;
wire ap_CS_fsm_state6;
wire ap_CS_fsm_state7;
wire ap_CS_fsm_state8;
wire ap_CS_fsm_state9;
wire [42:0] ap_NS_fsm;
wire ap_clk;
wire ap_done;
wire ap_idle;
wire ap_ready;
wire ap_rst;
wire ap_start;
wire carry_1_fu_789_p2;
wire deleted_ones_fu_808_p3;
wire deleted_zeros_fu_803_p3;
wire [4:0] grp_fu_263_p0;
wire [4:0] grp_fu_263_p2;
wire [8:0] grp_fu_283_p0;
wire [8:0] grp_fu_283_p1;
wire [8:0] grp_fu_283_p2;
wire [6:0] grp_fu_312_p0;
wire [6:0] grp_fu_312_p2;
wire [43:0] grp_fu_352_p0;
wire [43:0] grp_fu_352_p1;
wire [43:0] grp_fu_352_p2;
wire [31:0] grp_fu_378_p2;
wire [31:0] grp_fu_406_p1;
wire [31:0] grp_fu_406_p2;
wire [35:0] grp_fu_426_p0;
wire [35:0] grp_fu_426_p1;
wire [35:0] grp_fu_426_p2;
wire [31:0] grp_fu_452_p2;
wire [31:0] grp_fu_480_p1;
wire [31:0] grp_fu_480_p2;
wire [16:0] grp_fu_501_p0;
wire [16:0] grp_fu_501_p1;
wire [16:0] grp_fu_501_p2;
wire [35:0] grp_fu_522_p0;
wire [35:0] grp_fu_522_p1;
wire [35:0] grp_fu_522_p2;
wire [31:0] grp_fu_584_p2;
wire [7:0] grp_fu_592_p1;
wire [7:0] grp_fu_592_p2;
wire [8:0] grp_fu_639_p0;
wire [8:0] grp_fu_639_p1;
wire [8:0] grp_fu_639_p2;
wire [7:0] grp_fu_645_p0;
wire [7:0] grp_fu_645_p2;
wire [31:0] grp_fu_659_p1;
wire [31:0] grp_fu_659_p2;
wire [9:0] grp_fu_672_p0;
wire [9:0] grp_fu_672_p1;
wire [9:0] grp_fu_672_p2;
wire [31:0] grp_fu_732_p0;
wire [31:0] grp_fu_732_p2;
wire [3:0] grp_fu_740_p1;
wire [3:0] grp_fu_740_p2;
wire [33:0] grp_fu_768_p0;
wire [33:0] grp_fu_768_p1;
wire [33:0] grp_fu_768_p2;
wire [31:0] grp_fu_798_p2;
wire [31:0] grp_fu_892_p1;
wire [31:0] grp_fu_892_p2;
wire [33:0] grp_fu_931_p0;
wire [33:0] grp_fu_931_p1;
wire [33:0] grp_fu_931_p2;
wire [31:0] grp_fu_947_p2;
wire icmp_ln410_fu_578_p2;
wire icmp_ln851_1_fu_362_p2;
wire icmp_ln851_2_fu_436_p2;
wire icmp_ln851_3_fu_532_p2;
wire icmp_ln851_fu_293_p2;
wire neg_src_fu_871_p2;
wire op_0;
wire [3:0] op_1;
wire [7:0] op_10;
wire [3:0] op_12;
wire [7:0] op_13;
wire [1:0] op_14;
wire [7:0] op_15;
wire [7:0] op_16;
wire [3:0] op_17;
wire [1:0] op_18;
wire [3:0] op_19_V_fu_911_p3;
wire [3:0] op_2;
wire [31:0] op_32;
wire op_32_ap_vld;
wire [15:0] op_4;
wire [7:0] op_5;
wire [15:0] op_6;
wire [3:0] op_8;
wire [3:0] op_9;
wire or_ln340_1_fu_876_p2;
wire or_ln340_fu_833_p2;
wire or_ln412_fu_718_p2;
wire or_ln781_fu_866_p2;
wire or_ln785_1_fu_901_p2;
wire or_ln785_fu_823_p2;
wire overflow_fu_828_p2;
wire p_Result_10_fu_952_p3;
wire p_Result_12_fu_711_p3;
wire p_Result_1_fu_383_p3;
wire p_Result_5_fu_704_p3;
wire p_Result_7_fu_457_p3;
wire p_Result_8_fu_601_p3;
wire p_Result_9_fu_838_p3;
wire p_Result_s_fu_318_p3;
wire r_fu_650_p2;
wire [31:0] ret_V_18_fu_395_p3;
wire [31:0] ret_V_21_fu_469_p3;
wire [31:0] ret_V_23_fu_613_p3;
wire [31:0] ret_V_26_fu_854_p3;
wire [32:0] rhs_10_fu_757_p3;
wire [32:0] rhs_13_fu_920_p3;
wire [7:0] rhs_1_fu_272_p3;
wire [9:0] rhs_2_fu_489_p3;
wire [6:0] rhs_3_fu_623_p3;
wire [34:0] rhs_5_fu_415_p3;
wire [34:0] rhs_7_fu_511_p3;
wire [4:0] select_ln215_fu_251_p3;
wire [3:0] select_ln340_fu_881_p3;
wire [6:0] select_ln353_fu_330_p3;
wire [31:0] select_ln850_1_fu_390_p3;
wire [31:0] select_ln850_2_fu_464_p3;
wire [31:0] select_ln850_3_fu_608_p3;
wire [31:0] select_ln850_4_fu_848_p3;
wire [31:0] select_ln850_5_fu_962_p3;
wire [6:0] select_ln850_fu_325_p3;
wire [7:0] sext_ln1192_fu_268_p0;
wire [15:0] sext_ln703_1_fu_337_p0;
wire [3:0] sext_ln703_3_fu_411_p0;
wire [3:0] sext_ln703_4_fu_507_p0;
wire [3:0] sext_ln703_5_fu_753_p0;
wire [6:0] sext_ln850_fu_309_p1;
wire \sub_17s_17ns_17_2_1_U10.ce ;
wire \sub_17s_17ns_17_2_1_U10.clk ;
wire [16:0] \sub_17s_17ns_17_2_1_U10.din0 ;
wire [16:0] \sub_17s_17ns_17_2_1_U10.din1 ;
wire [16:0] \sub_17s_17ns_17_2_1_U10.dout ;
wire \sub_17s_17ns_17_2_1_U10.reset ;
wire [16:0] \sub_17s_17ns_17_2_1_U10.top_sub_17s_17ns_17_2_1_Adder_7_U.a ;
wire [16:0] \sub_17s_17ns_17_2_1_U10.top_sub_17s_17ns_17_2_1_Adder_7_U.ain_s0 ;
wire [16:0] \sub_17s_17ns_17_2_1_U10.top_sub_17s_17ns_17_2_1_Adder_7_U.b ;
wire [16:0] \sub_17s_17ns_17_2_1_U10.top_sub_17s_17ns_17_2_1_Adder_7_U.bin_s0 ;
wire \sub_17s_17ns_17_2_1_U10.top_sub_17s_17ns_17_2_1_Adder_7_U.ce ;
wire \sub_17s_17ns_17_2_1_U10.top_sub_17s_17ns_17_2_1_Adder_7_U.clk ;
wire \sub_17s_17ns_17_2_1_U10.top_sub_17s_17ns_17_2_1_Adder_7_U.facout_s1 ;
wire \sub_17s_17ns_17_2_1_U10.top_sub_17s_17ns_17_2_1_Adder_7_U.facout_s2 ;
wire [7:0] \sub_17s_17ns_17_2_1_U10.top_sub_17s_17ns_17_2_1_Adder_7_U.fas_s1 ;
wire [8:0] \sub_17s_17ns_17_2_1_U10.top_sub_17s_17ns_17_2_1_Adder_7_U.fas_s2 ;
wire \sub_17s_17ns_17_2_1_U10.top_sub_17s_17ns_17_2_1_Adder_7_U.reset ;
wire [16:0] \sub_17s_17ns_17_2_1_U10.top_sub_17s_17ns_17_2_1_Adder_7_U.s ;
wire [7:0] \sub_17s_17ns_17_2_1_U10.top_sub_17s_17ns_17_2_1_Adder_7_U.u1.a ;
wire [7:0] \sub_17s_17ns_17_2_1_U10.top_sub_17s_17ns_17_2_1_Adder_7_U.u1.b ;
wire \sub_17s_17ns_17_2_1_U10.top_sub_17s_17ns_17_2_1_Adder_7_U.u1.cin ;
wire \sub_17s_17ns_17_2_1_U10.top_sub_17s_17ns_17_2_1_Adder_7_U.u1.cout ;
wire [7:0] \sub_17s_17ns_17_2_1_U10.top_sub_17s_17ns_17_2_1_Adder_7_U.u1.s ;
wire [8:0] \sub_17s_17ns_17_2_1_U10.top_sub_17s_17ns_17_2_1_Adder_7_U.u2.a ;
wire [8:0] \sub_17s_17ns_17_2_1_U10.top_sub_17s_17ns_17_2_1_Adder_7_U.u2.b ;
wire \sub_17s_17ns_17_2_1_U10.top_sub_17s_17ns_17_2_1_Adder_7_U.u2.cin ;
wire \sub_17s_17ns_17_2_1_U10.top_sub_17s_17ns_17_2_1_Adder_7_U.u2.cout ;
wire [8:0] \sub_17s_17ns_17_2_1_U10.top_sub_17s_17ns_17_2_1_Adder_7_U.u2.s ;
wire [17:0] tmp_2_fu_341_p3;
wire trunc_ln410_fu_556_p1;
wire [2:0] trunc_ln718_fu_597_p1;
wire [15:0] trunc_ln851_1_fu_358_p0;
wire [10:0] trunc_ln851_1_fu_358_p1;
wire [3:0] trunc_ln851_2_fu_432_p0;
wire [2:0] trunc_ln851_2_fu_432_p1;
wire [3:0] trunc_ln851_3_fu_528_p0;
wire [2:0] trunc_ln851_3_fu_528_p1;
wire [3:0] trunc_ln851_4_fu_845_p0;
wire trunc_ln851_4_fu_845_p1;
wire trunc_ln851_5_fu_959_p1;
wire [7:0] trunc_ln851_fu_289_p0;
wire [2:0] trunc_ln851_fu_289_p1;
wire xor_ln416_fu_774_p2;
wire xor_ln781_fu_861_p2;
wire xor_ln785_fu_818_p2;


assign _060_ = ap_CS_fsm[11] & icmp_ln851_1_reg_1043;
assign _061_ = icmp_ln851_2_reg_1090 & ap_CS_fsm[18];
assign _062_ = icmp_ln851_3_reg_1147 & ap_CS_fsm[25];
assign _063_ = ap_CS_fsm[6] & icmp_ln851_reg_1001;
assign _064_ = _066_ & ap_CS_fsm[0];
assign _065_ = ap_start & ap_CS_fsm[0];
assign and_ln412_fu_723_p2 = op_11_V_reg_1194[3] & or_ln412_fu_718_p2;
assign and_ln785_1_fu_906_p2 = or_ln785_1_fu_901_p2 & and_ln786_reg_1367;
assign and_ln785_fu_897_p2 = xor_ln416_reg_1330 & deleted_zeros_reg_1361;
assign and_ln786_fu_813_p2 = p_Result_14_reg_1312 & deleted_ones_fu_808_p3;
assign carry_1_fu_789_p2 = xor_ln416_reg_1330 & p_Result_13_reg_1265;
assign neg_src_fu_871_p2 = p_Result_11_reg_1251 & or_ln781_fu_866_p2;
assign overflow_fu_828_p2 = or_ln785_fu_823_p2 & Range1_all_zeros_reg_1354;
assign Range1_all_zeros_fu_793_p2 = ~ p_Result_11_reg_1251;
assign xor_ln781_fu_861_p2 = ~ p_Result_13_reg_1265;
assign xor_ln785_fu_818_p2 = ~ deleted_zeros_reg_1361;
assign xor_ln416_fu_774_p2 = ~ p_Result_14_reg_1312;
assign _066_ = ~ ap_start;
assign _067_ = { tmp_reg_1157, trunc_ln410_reg_1162 } == 1'h1;
always @(posedge \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_10_U.clk )
\add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_10_U.bin_s1  <= _069_;
always @(posedge \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_10_U.clk )
\add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_10_U.ain_s1  <= _068_;
always @(posedge \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_10_U.clk )
\add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_10_U.sum_s1  <= _071_;
always @(posedge \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_10_U.clk )
\add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_10_U.carry_s1  <= _070_;
assign _069_ = \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_10_U.ce  ? \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_10_U.b [9:5] : \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_10_U.bin_s1 ;
assign _068_ = \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_10_U.ce  ? \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_10_U.a [9:5] : \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_10_U.ain_s1 ;
assign _070_ = \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_10_U.ce  ? \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_10_U.facout_s1  : \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_10_U.carry_s1 ;
assign _071_ = \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_10_U.ce  ? \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_10_U.fas_s1  : \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_10_U.sum_s1 ;
assign _072_ = \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_10_U.u1.a  + \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_10_U.u1.b ;
assign { \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_10_U.u1.cout , \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_10_U.u1.s  } = _072_ + \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_10_U.u1.cin ;
assign _073_ = \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_10_U.u2.a  + \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_10_U.u2.b ;
assign { \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_10_U.u2.cout , \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_10_U.u2.s  } = _073_ + \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_10_U.u2.cin ;
always @(posedge \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_4_U.clk )
\add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_4_U.bin_s1  <= _075_;
always @(posedge \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_4_U.clk )
\add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_4_U.ain_s1  <= _074_;
always @(posedge \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_4_U.clk )
\add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_4_U.sum_s1  <= _077_;
always @(posedge \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_4_U.clk )
\add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_4_U.carry_s1  <= _076_;
assign _075_ = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_4_U.ce  ? \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_4_U.b [31:16] : \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_4_U.bin_s1 ;
assign _074_ = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_4_U.ce  ? \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_4_U.a [31:16] : \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_4_U.ain_s1 ;
assign _076_ = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_4_U.ce  ? \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_4_U.facout_s1  : \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_4_U.carry_s1 ;
assign _077_ = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_4_U.ce  ? \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_4_U.fas_s1  : \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_4_U.sum_s1 ;
assign _078_ = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.a  + \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.b ;
assign { \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.cout , \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.s  } = _078_ + \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.cin ;
assign _079_ = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.a  + \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.b ;
assign { \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.cout , \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.s  } = _079_ + \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.cin ;
always @(posedge \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_4_U.clk )
\add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_4_U.bin_s1  <= _081_;
always @(posedge \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_4_U.clk )
\add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_4_U.ain_s1  <= _080_;
always @(posedge \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_4_U.clk )
\add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_4_U.sum_s1  <= _083_;
always @(posedge \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_4_U.clk )
\add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_4_U.carry_s1  <= _082_;
assign _081_ = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_4_U.ce  ? \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_4_U.b [31:16] : \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_4_U.bin_s1 ;
assign _080_ = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_4_U.ce  ? \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_4_U.a [31:16] : \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_4_U.ain_s1 ;
assign _082_ = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_4_U.ce  ? \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_4_U.facout_s1  : \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_4_U.carry_s1 ;
assign _083_ = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_4_U.ce  ? \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_4_U.fas_s1  : \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_4_U.sum_s1 ;
assign _084_ = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.a  + \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.b ;
assign { \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.cout , \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.s  } = _084_ + \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.cin ;
assign _085_ = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.a  + \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.b ;
assign { \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.cout , \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.s  } = _085_ + \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.cin ;
always @(posedge \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_4_U.clk )
\add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_4_U.bin_s1  <= _087_;
always @(posedge \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_4_U.clk )
\add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_4_U.ain_s1  <= _086_;
always @(posedge \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_4_U.clk )
\add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_4_U.sum_s1  <= _089_;
always @(posedge \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_4_U.clk )
\add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_4_U.carry_s1  <= _088_;
assign _087_ = \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_4_U.ce  ? \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_4_U.b [31:16] : \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_4_U.bin_s1 ;
assign _086_ = \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_4_U.ce  ? \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_4_U.a [31:16] : \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_4_U.ain_s1 ;
assign _088_ = \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_4_U.ce  ? \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_4_U.facout_s1  : \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_4_U.carry_s1 ;
assign _089_ = \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_4_U.ce  ? \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_4_U.fas_s1  : \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_4_U.sum_s1 ;
assign _090_ = \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.a  + \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.b ;
assign { \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.cout , \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.s  } = _090_ + \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.cin ;
assign _091_ = \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.a  + \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.b ;
assign { \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.cout , \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.s  } = _091_ + \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.cin ;
always @(posedge \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.clk )
\add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.bin_s1  <= _093_;
always @(posedge \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.clk )
\add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.ain_s1  <= _092_;
always @(posedge \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.clk )
\add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.sum_s1  <= _095_;
always @(posedge \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.clk )
\add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.carry_s1  <= _094_;
assign _093_ = \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.ce  ? \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.b [31:16] : \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.bin_s1 ;
assign _092_ = \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.ce  ? \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.a [31:16] : \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.ain_s1 ;
assign _094_ = \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.ce  ? \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.facout_s1  : \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.carry_s1 ;
assign _095_ = \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.ce  ? \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.fas_s1  : \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.sum_s1 ;
assign _096_ = \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.a  + \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.b ;
assign { \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.cout , \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.s  } = _096_ + \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.cin ;
assign _097_ = \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.a  + \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.b ;
assign { \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.cout , \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.s  } = _097_ + \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.cin ;
always @(posedge \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.clk )
\add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.bin_s1  <= _099_;
always @(posedge \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.clk )
\add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.ain_s1  <= _098_;
always @(posedge \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.clk )
\add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.sum_s1  <= _101_;
always @(posedge \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.clk )
\add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.carry_s1  <= _100_;
assign _099_ = \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.ce  ? \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.b [31:16] : \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.bin_s1 ;
assign _098_ = \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.ce  ? \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.a [31:16] : \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.ain_s1 ;
assign _100_ = \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.ce  ? \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.facout_s1  : \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.carry_s1 ;
assign _101_ = \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.ce  ? \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.fas_s1  : \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.sum_s1 ;
assign _102_ = \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.a  + \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.b ;
assign { \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.cout , \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.s  } = _102_ + \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.cin ;
assign _103_ = \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.a  + \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.b ;
assign { \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.cout , \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.s  } = _103_ + \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.cin ;
always @(posedge \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_4_U.clk )
\add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_4_U.bin_s1  <= _105_;
always @(posedge \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_4_U.clk )
\add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_4_U.ain_s1  <= _104_;
always @(posedge \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_4_U.clk )
\add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_4_U.sum_s1  <= _107_;
always @(posedge \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_4_U.clk )
\add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_4_U.carry_s1  <= _106_;
assign _105_ = \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_4_U.ce  ? \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_4_U.b [31:16] : \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_4_U.bin_s1 ;
assign _104_ = \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_4_U.ce  ? \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_4_U.a [31:16] : \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_4_U.ain_s1 ;
assign _106_ = \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_4_U.ce  ? \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_4_U.facout_s1  : \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_4_U.carry_s1 ;
assign _107_ = \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_4_U.ce  ? \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_4_U.fas_s1  : \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_4_U.sum_s1 ;
assign _108_ = \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.a  + \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.b ;
assign { \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.cout , \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.s  } = _108_ + \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.cin ;
assign _109_ = \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.a  + \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.b ;
assign { \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.cout , \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.s  } = _109_ + \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.cin ;
always @(posedge \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_5_U.clk )
\add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_5_U.bin_s1  <= _111_;
always @(posedge \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_5_U.clk )
\add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_5_U.ain_s1  <= _110_;
always @(posedge \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_5_U.clk )
\add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_5_U.sum_s1  <= _113_;
always @(posedge \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_5_U.clk )
\add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_5_U.carry_s1  <= _112_;
assign _111_ = \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_5_U.ce  ? \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_5_U.b [31:16] : \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_5_U.bin_s1 ;
assign _110_ = \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_5_U.ce  ? \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_5_U.a [31:16] : \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_5_U.ain_s1 ;
assign _112_ = \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_5_U.ce  ? \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_5_U.facout_s1  : \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_5_U.carry_s1 ;
assign _113_ = \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_5_U.ce  ? \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_5_U.fas_s1  : \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_5_U.sum_s1 ;
assign _114_ = \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_5_U.u1.a  + \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_5_U.u1.b ;
assign { \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_5_U.u1.cout , \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_5_U.u1.s  } = _114_ + \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_5_U.u1.cin ;
assign _115_ = \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_5_U.u2.a  + \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_5_U.u2.b ;
assign { \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_5_U.u2.cout , \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_5_U.u2.s  } = _115_ + \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_5_U.u2.cin ;
always @(posedge \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_5_U.clk )
\add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_5_U.bin_s1  <= _117_;
always @(posedge \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_5_U.clk )
\add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_5_U.ain_s1  <= _116_;
always @(posedge \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_5_U.clk )
\add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_5_U.sum_s1  <= _119_;
always @(posedge \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_5_U.clk )
\add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_5_U.carry_s1  <= _118_;
assign _117_ = \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_5_U.ce  ? \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_5_U.b [31:16] : \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_5_U.bin_s1 ;
assign _116_ = \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_5_U.ce  ? \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_5_U.a [31:16] : \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_5_U.ain_s1 ;
assign _118_ = \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_5_U.ce  ? \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_5_U.facout_s1  : \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_5_U.carry_s1 ;
assign _119_ = \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_5_U.ce  ? \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_5_U.fas_s1  : \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_5_U.sum_s1 ;
assign _120_ = \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_5_U.u1.a  + \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_5_U.u1.b ;
assign { \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_5_U.u1.cout , \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_5_U.u1.s  } = _120_ + \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_5_U.u1.cin ;
assign _121_ = \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_5_U.u2.a  + \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_5_U.u2.b ;
assign { \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_5_U.u2.cout , \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_5_U.u2.s  } = _121_ + \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_5_U.u2.cin ;
always @(posedge \add_32ns_32s_32_2_1_U6.top_add_32ns_32s_32_2_1_Adder_5_U.clk )
\add_32ns_32s_32_2_1_U6.top_add_32ns_32s_32_2_1_Adder_5_U.bin_s1  <= _123_;
always @(posedge \add_32ns_32s_32_2_1_U6.top_add_32ns_32s_32_2_1_Adder_5_U.clk )
\add_32ns_32s_32_2_1_U6.top_add_32ns_32s_32_2_1_Adder_5_U.ain_s1  <= _122_;
always @(posedge \add_32ns_32s_32_2_1_U6.top_add_32ns_32s_32_2_1_Adder_5_U.clk )
\add_32ns_32s_32_2_1_U6.top_add_32ns_32s_32_2_1_Adder_5_U.sum_s1  <= _125_;
always @(posedge \add_32ns_32s_32_2_1_U6.top_add_32ns_32s_32_2_1_Adder_5_U.clk )
\add_32ns_32s_32_2_1_U6.top_add_32ns_32s_32_2_1_Adder_5_U.carry_s1  <= _124_;
assign _123_ = \add_32ns_32s_32_2_1_U6.top_add_32ns_32s_32_2_1_Adder_5_U.ce  ? \add_32ns_32s_32_2_1_U6.top_add_32ns_32s_32_2_1_Adder_5_U.b [31:16] : \add_32ns_32s_32_2_1_U6.top_add_32ns_32s_32_2_1_Adder_5_U.bin_s1 ;
assign _122_ = \add_32ns_32s_32_2_1_U6.top_add_32ns_32s_32_2_1_Adder_5_U.ce  ? \add_32ns_32s_32_2_1_U6.top_add_32ns_32s_32_2_1_Adder_5_U.a [31:16] : \add_32ns_32s_32_2_1_U6.top_add_32ns_32s_32_2_1_Adder_5_U.ain_s1 ;
assign _124_ = \add_32ns_32s_32_2_1_U6.top_add_32ns_32s_32_2_1_Adder_5_U.ce  ? \add_32ns_32s_32_2_1_U6.top_add_32ns_32s_32_2_1_Adder_5_U.facout_s1  : \add_32ns_32s_32_2_1_U6.top_add_32ns_32s_32_2_1_Adder_5_U.carry_s1 ;
assign _125_ = \add_32ns_32s_32_2_1_U6.top_add_32ns_32s_32_2_1_Adder_5_U.ce  ? \add_32ns_32s_32_2_1_U6.top_add_32ns_32s_32_2_1_Adder_5_U.fas_s1  : \add_32ns_32s_32_2_1_U6.top_add_32ns_32s_32_2_1_Adder_5_U.sum_s1 ;
assign _126_ = \add_32ns_32s_32_2_1_U6.top_add_32ns_32s_32_2_1_Adder_5_U.u1.a  + \add_32ns_32s_32_2_1_U6.top_add_32ns_32s_32_2_1_Adder_5_U.u1.b ;
assign { \add_32ns_32s_32_2_1_U6.top_add_32ns_32s_32_2_1_Adder_5_U.u1.cout , \add_32ns_32s_32_2_1_U6.top_add_32ns_32s_32_2_1_Adder_5_U.u1.s  } = _126_ + \add_32ns_32s_32_2_1_U6.top_add_32ns_32s_32_2_1_Adder_5_U.u1.cin ;
assign _127_ = \add_32ns_32s_32_2_1_U6.top_add_32ns_32s_32_2_1_Adder_5_U.u2.a  + \add_32ns_32s_32_2_1_U6.top_add_32ns_32s_32_2_1_Adder_5_U.u2.b ;
assign { \add_32ns_32s_32_2_1_U6.top_add_32ns_32s_32_2_1_Adder_5_U.u2.cout , \add_32ns_32s_32_2_1_U6.top_add_32ns_32s_32_2_1_Adder_5_U.u2.s  } = _127_ + \add_32ns_32s_32_2_1_U6.top_add_32ns_32s_32_2_1_Adder_5_U.u2.cin ;
always @(posedge \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_11_U.clk )
\add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_11_U.bin_s1  <= _129_;
always @(posedge \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_11_U.clk )
\add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_11_U.ain_s1  <= _128_;
always @(posedge \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_11_U.clk )
\add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_11_U.sum_s1  <= _131_;
always @(posedge \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_11_U.clk )
\add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_11_U.carry_s1  <= _130_;
assign _129_ = \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_11_U.ce  ? \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_11_U.b [31:16] : \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_11_U.bin_s1 ;
assign _128_ = \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_11_U.ce  ? \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_11_U.a [31:16] : \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_11_U.ain_s1 ;
assign _130_ = \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_11_U.ce  ? \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_11_U.facout_s1  : \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_11_U.carry_s1 ;
assign _131_ = \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_11_U.ce  ? \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_11_U.fas_s1  : \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_11_U.sum_s1 ;
assign _132_ = \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_11_U.u1.a  + \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_11_U.u1.b ;
assign { \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_11_U.u1.cout , \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_11_U.u1.s  } = _132_ + \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_11_U.u1.cin ;
assign _133_ = \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_11_U.u2.a  + \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_11_U.u2.b ;
assign { \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_11_U.u2.cout , \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_11_U.u2.s  } = _133_ + \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_11_U.u2.cin ;
always @(posedge \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_13_U.clk )
\add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_13_U.bin_s1  <= _135_;
always @(posedge \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_13_U.clk )
\add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_13_U.ain_s1  <= _134_;
always @(posedge \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_13_U.clk )
\add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_13_U.sum_s1  <= _137_;
always @(posedge \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_13_U.clk )
\add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_13_U.carry_s1  <= _136_;
assign _135_ = \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_13_U.ce  ? \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_13_U.b [33:17] : \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_13_U.bin_s1 ;
assign _134_ = \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_13_U.ce  ? \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_13_U.a [33:17] : \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_13_U.ain_s1 ;
assign _136_ = \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_13_U.ce  ? \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_13_U.facout_s1  : \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_13_U.carry_s1 ;
assign _137_ = \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_13_U.ce  ? \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_13_U.fas_s1  : \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_13_U.sum_s1 ;
assign _138_ = \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_13_U.u1.a  + \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_13_U.u1.b ;
assign { \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_13_U.u1.cout , \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_13_U.u1.s  } = _138_ + \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_13_U.u1.cin ;
assign _139_ = \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_13_U.u2.a  + \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_13_U.u2.b ;
assign { \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_13_U.u2.cout , \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_13_U.u2.s  } = _139_ + \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_13_U.u2.cin ;
always @(posedge \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_13_U.clk )
\add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_13_U.bin_s1  <= _141_;
always @(posedge \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_13_U.clk )
\add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_13_U.ain_s1  <= _140_;
always @(posedge \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_13_U.clk )
\add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_13_U.sum_s1  <= _143_;
always @(posedge \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_13_U.clk )
\add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_13_U.carry_s1  <= _142_;
assign _141_ = \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_13_U.ce  ? \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_13_U.b [33:17] : \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_13_U.bin_s1 ;
assign _140_ = \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_13_U.ce  ? \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_13_U.a [33:17] : \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_13_U.ain_s1 ;
assign _142_ = \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_13_U.ce  ? \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_13_U.facout_s1  : \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_13_U.carry_s1 ;
assign _143_ = \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_13_U.ce  ? \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_13_U.fas_s1  : \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_13_U.sum_s1 ;
assign _144_ = \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_13_U.u1.a  + \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_13_U.u1.b ;
assign { \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_13_U.u1.cout , \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_13_U.u1.s  } = _144_ + \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_13_U.u1.cin ;
assign _145_ = \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_13_U.u2.a  + \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_13_U.u2.b ;
assign { \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_13_U.u2.cout , \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_13_U.u2.s  } = _145_ + \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_13_U.u2.cin ;
always @(posedge \add_36s_36s_36_2_1_U11.top_add_36s_36s_36_2_1_Adder_6_U.clk )
\add_36s_36s_36_2_1_U11.top_add_36s_36s_36_2_1_Adder_6_U.bin_s1  <= _147_;
always @(posedge \add_36s_36s_36_2_1_U11.top_add_36s_36s_36_2_1_Adder_6_U.clk )
\add_36s_36s_36_2_1_U11.top_add_36s_36s_36_2_1_Adder_6_U.ain_s1  <= _146_;
always @(posedge \add_36s_36s_36_2_1_U11.top_add_36s_36s_36_2_1_Adder_6_U.clk )
\add_36s_36s_36_2_1_U11.top_add_36s_36s_36_2_1_Adder_6_U.sum_s1  <= _149_;
always @(posedge \add_36s_36s_36_2_1_U11.top_add_36s_36s_36_2_1_Adder_6_U.clk )
\add_36s_36s_36_2_1_U11.top_add_36s_36s_36_2_1_Adder_6_U.carry_s1  <= _148_;
assign _147_ = \add_36s_36s_36_2_1_U11.top_add_36s_36s_36_2_1_Adder_6_U.ce  ? \add_36s_36s_36_2_1_U11.top_add_36s_36s_36_2_1_Adder_6_U.b [35:18] : \add_36s_36s_36_2_1_U11.top_add_36s_36s_36_2_1_Adder_6_U.bin_s1 ;
assign _146_ = \add_36s_36s_36_2_1_U11.top_add_36s_36s_36_2_1_Adder_6_U.ce  ? \add_36s_36s_36_2_1_U11.top_add_36s_36s_36_2_1_Adder_6_U.a [35:18] : \add_36s_36s_36_2_1_U11.top_add_36s_36s_36_2_1_Adder_6_U.ain_s1 ;
assign _148_ = \add_36s_36s_36_2_1_U11.top_add_36s_36s_36_2_1_Adder_6_U.ce  ? \add_36s_36s_36_2_1_U11.top_add_36s_36s_36_2_1_Adder_6_U.facout_s1  : \add_36s_36s_36_2_1_U11.top_add_36s_36s_36_2_1_Adder_6_U.carry_s1 ;
assign _149_ = \add_36s_36s_36_2_1_U11.top_add_36s_36s_36_2_1_Adder_6_U.ce  ? \add_36s_36s_36_2_1_U11.top_add_36s_36s_36_2_1_Adder_6_U.fas_s1  : \add_36s_36s_36_2_1_U11.top_add_36s_36s_36_2_1_Adder_6_U.sum_s1 ;
assign _150_ = \add_36s_36s_36_2_1_U11.top_add_36s_36s_36_2_1_Adder_6_U.u1.a  + \add_36s_36s_36_2_1_U11.top_add_36s_36s_36_2_1_Adder_6_U.u1.b ;
assign { \add_36s_36s_36_2_1_U11.top_add_36s_36s_36_2_1_Adder_6_U.u1.cout , \add_36s_36s_36_2_1_U11.top_add_36s_36s_36_2_1_Adder_6_U.u1.s  } = _150_ + \add_36s_36s_36_2_1_U11.top_add_36s_36s_36_2_1_Adder_6_U.u1.cin ;
assign _151_ = \add_36s_36s_36_2_1_U11.top_add_36s_36s_36_2_1_Adder_6_U.u2.a  + \add_36s_36s_36_2_1_U11.top_add_36s_36s_36_2_1_Adder_6_U.u2.b ;
assign { \add_36s_36s_36_2_1_U11.top_add_36s_36s_36_2_1_Adder_6_U.u2.cout , \add_36s_36s_36_2_1_U11.top_add_36s_36s_36_2_1_Adder_6_U.u2.s  } = _151_ + \add_36s_36s_36_2_1_U11.top_add_36s_36s_36_2_1_Adder_6_U.u2.cin ;
always @(posedge \add_36s_36s_36_2_1_U7.top_add_36s_36s_36_2_1_Adder_6_U.clk )
\add_36s_36s_36_2_1_U7.top_add_36s_36s_36_2_1_Adder_6_U.bin_s1  <= _153_;
always @(posedge \add_36s_36s_36_2_1_U7.top_add_36s_36s_36_2_1_Adder_6_U.clk )
\add_36s_36s_36_2_1_U7.top_add_36s_36s_36_2_1_Adder_6_U.ain_s1  <= _152_;
always @(posedge \add_36s_36s_36_2_1_U7.top_add_36s_36s_36_2_1_Adder_6_U.clk )
\add_36s_36s_36_2_1_U7.top_add_36s_36s_36_2_1_Adder_6_U.sum_s1  <= _155_;
always @(posedge \add_36s_36s_36_2_1_U7.top_add_36s_36s_36_2_1_Adder_6_U.clk )
\add_36s_36s_36_2_1_U7.top_add_36s_36s_36_2_1_Adder_6_U.carry_s1  <= _154_;
assign _153_ = \add_36s_36s_36_2_1_U7.top_add_36s_36s_36_2_1_Adder_6_U.ce  ? \add_36s_36s_36_2_1_U7.top_add_36s_36s_36_2_1_Adder_6_U.b [35:18] : \add_36s_36s_36_2_1_U7.top_add_36s_36s_36_2_1_Adder_6_U.bin_s1 ;
assign _152_ = \add_36s_36s_36_2_1_U7.top_add_36s_36s_36_2_1_Adder_6_U.ce  ? \add_36s_36s_36_2_1_U7.top_add_36s_36s_36_2_1_Adder_6_U.a [35:18] : \add_36s_36s_36_2_1_U7.top_add_36s_36s_36_2_1_Adder_6_U.ain_s1 ;
assign _154_ = \add_36s_36s_36_2_1_U7.top_add_36s_36s_36_2_1_Adder_6_U.ce  ? \add_36s_36s_36_2_1_U7.top_add_36s_36s_36_2_1_Adder_6_U.facout_s1  : \add_36s_36s_36_2_1_U7.top_add_36s_36s_36_2_1_Adder_6_U.carry_s1 ;
assign _155_ = \add_36s_36s_36_2_1_U7.top_add_36s_36s_36_2_1_Adder_6_U.ce  ? \add_36s_36s_36_2_1_U7.top_add_36s_36s_36_2_1_Adder_6_U.fas_s1  : \add_36s_36s_36_2_1_U7.top_add_36s_36s_36_2_1_Adder_6_U.sum_s1 ;
assign _156_ = \add_36s_36s_36_2_1_U7.top_add_36s_36s_36_2_1_Adder_6_U.u1.a  + \add_36s_36s_36_2_1_U7.top_add_36s_36s_36_2_1_Adder_6_U.u1.b ;
assign { \add_36s_36s_36_2_1_U7.top_add_36s_36s_36_2_1_Adder_6_U.u1.cout , \add_36s_36s_36_2_1_U7.top_add_36s_36s_36_2_1_Adder_6_U.u1.s  } = _156_ + \add_36s_36s_36_2_1_U7.top_add_36s_36s_36_2_1_Adder_6_U.u1.cin ;
assign _157_ = \add_36s_36s_36_2_1_U7.top_add_36s_36s_36_2_1_Adder_6_U.u2.a  + \add_36s_36s_36_2_1_U7.top_add_36s_36s_36_2_1_Adder_6_U.u2.b ;
assign { \add_36s_36s_36_2_1_U7.top_add_36s_36s_36_2_1_Adder_6_U.u2.cout , \add_36s_36s_36_2_1_U7.top_add_36s_36s_36_2_1_Adder_6_U.u2.s  } = _157_ + \add_36s_36s_36_2_1_U7.top_add_36s_36s_36_2_1_Adder_6_U.u2.cin ;
always @(posedge \add_44s_44s_44_2_1_U4.top_add_44s_44s_44_2_1_Adder_3_U.clk )
\add_44s_44s_44_2_1_U4.top_add_44s_44s_44_2_1_Adder_3_U.bin_s1  <= _159_;
always @(posedge \add_44s_44s_44_2_1_U4.top_add_44s_44s_44_2_1_Adder_3_U.clk )
\add_44s_44s_44_2_1_U4.top_add_44s_44s_44_2_1_Adder_3_U.ain_s1  <= _158_;
always @(posedge \add_44s_44s_44_2_1_U4.top_add_44s_44s_44_2_1_Adder_3_U.clk )
\add_44s_44s_44_2_1_U4.top_add_44s_44s_44_2_1_Adder_3_U.sum_s1  <= _161_;
always @(posedge \add_44s_44s_44_2_1_U4.top_add_44s_44s_44_2_1_Adder_3_U.clk )
\add_44s_44s_44_2_1_U4.top_add_44s_44s_44_2_1_Adder_3_U.carry_s1  <= _160_;
assign _159_ = \add_44s_44s_44_2_1_U4.top_add_44s_44s_44_2_1_Adder_3_U.ce  ? \add_44s_44s_44_2_1_U4.top_add_44s_44s_44_2_1_Adder_3_U.b [43:22] : \add_44s_44s_44_2_1_U4.top_add_44s_44s_44_2_1_Adder_3_U.bin_s1 ;
assign _158_ = \add_44s_44s_44_2_1_U4.top_add_44s_44s_44_2_1_Adder_3_U.ce  ? \add_44s_44s_44_2_1_U4.top_add_44s_44s_44_2_1_Adder_3_U.a [43:22] : \add_44s_44s_44_2_1_U4.top_add_44s_44s_44_2_1_Adder_3_U.ain_s1 ;
assign _160_ = \add_44s_44s_44_2_1_U4.top_add_44s_44s_44_2_1_Adder_3_U.ce  ? \add_44s_44s_44_2_1_U4.top_add_44s_44s_44_2_1_Adder_3_U.facout_s1  : \add_44s_44s_44_2_1_U4.top_add_44s_44s_44_2_1_Adder_3_U.carry_s1 ;
assign _161_ = \add_44s_44s_44_2_1_U4.top_add_44s_44s_44_2_1_Adder_3_U.ce  ? \add_44s_44s_44_2_1_U4.top_add_44s_44s_44_2_1_Adder_3_U.fas_s1  : \add_44s_44s_44_2_1_U4.top_add_44s_44s_44_2_1_Adder_3_U.sum_s1 ;
assign _162_ = \add_44s_44s_44_2_1_U4.top_add_44s_44s_44_2_1_Adder_3_U.u1.a  + \add_44s_44s_44_2_1_U4.top_add_44s_44s_44_2_1_Adder_3_U.u1.b ;
assign { \add_44s_44s_44_2_1_U4.top_add_44s_44s_44_2_1_Adder_3_U.u1.cout , \add_44s_44s_44_2_1_U4.top_add_44s_44s_44_2_1_Adder_3_U.u1.s  } = _162_ + \add_44s_44s_44_2_1_U4.top_add_44s_44s_44_2_1_Adder_3_U.u1.cin ;
assign _163_ = \add_44s_44s_44_2_1_U4.top_add_44s_44s_44_2_1_Adder_3_U.u2.a  + \add_44s_44s_44_2_1_U4.top_add_44s_44s_44_2_1_Adder_3_U.u2.b ;
assign { \add_44s_44s_44_2_1_U4.top_add_44s_44s_44_2_1_Adder_3_U.u2.cout , \add_44s_44s_44_2_1_U4.top_add_44s_44s_44_2_1_Adder_3_U.u2.s  } = _163_ + \add_44s_44s_44_2_1_U4.top_add_44s_44s_44_2_1_Adder_3_U.u2.cin ;
always @(posedge \add_4ns_4ns_4_2_1_U19.top_add_4ns_4ns_4_2_1_Adder_12_U.clk )
\add_4ns_4ns_4_2_1_U19.top_add_4ns_4ns_4_2_1_Adder_12_U.bin_s1  <= _165_;
always @(posedge \add_4ns_4ns_4_2_1_U19.top_add_4ns_4ns_4_2_1_Adder_12_U.clk )
\add_4ns_4ns_4_2_1_U19.top_add_4ns_4ns_4_2_1_Adder_12_U.ain_s1  <= _164_;
always @(posedge \add_4ns_4ns_4_2_1_U19.top_add_4ns_4ns_4_2_1_Adder_12_U.clk )
\add_4ns_4ns_4_2_1_U19.top_add_4ns_4ns_4_2_1_Adder_12_U.sum_s1  <= _167_;
always @(posedge \add_4ns_4ns_4_2_1_U19.top_add_4ns_4ns_4_2_1_Adder_12_U.clk )
\add_4ns_4ns_4_2_1_U19.top_add_4ns_4ns_4_2_1_Adder_12_U.carry_s1  <= _166_;
assign _165_ = \add_4ns_4ns_4_2_1_U19.top_add_4ns_4ns_4_2_1_Adder_12_U.ce  ? \add_4ns_4ns_4_2_1_U19.top_add_4ns_4ns_4_2_1_Adder_12_U.b [3:2] : \add_4ns_4ns_4_2_1_U19.top_add_4ns_4ns_4_2_1_Adder_12_U.bin_s1 ;
assign _164_ = \add_4ns_4ns_4_2_1_U19.top_add_4ns_4ns_4_2_1_Adder_12_U.ce  ? \add_4ns_4ns_4_2_1_U19.top_add_4ns_4ns_4_2_1_Adder_12_U.a [3:2] : \add_4ns_4ns_4_2_1_U19.top_add_4ns_4ns_4_2_1_Adder_12_U.ain_s1 ;
assign _166_ = \add_4ns_4ns_4_2_1_U19.top_add_4ns_4ns_4_2_1_Adder_12_U.ce  ? \add_4ns_4ns_4_2_1_U19.top_add_4ns_4ns_4_2_1_Adder_12_U.facout_s1  : \add_4ns_4ns_4_2_1_U19.top_add_4ns_4ns_4_2_1_Adder_12_U.carry_s1 ;
assign _167_ = \add_4ns_4ns_4_2_1_U19.top_add_4ns_4ns_4_2_1_Adder_12_U.ce  ? \add_4ns_4ns_4_2_1_U19.top_add_4ns_4ns_4_2_1_Adder_12_U.fas_s1  : \add_4ns_4ns_4_2_1_U19.top_add_4ns_4ns_4_2_1_Adder_12_U.sum_s1 ;
assign _168_ = \add_4ns_4ns_4_2_1_U19.top_add_4ns_4ns_4_2_1_Adder_12_U.u1.a  + \add_4ns_4ns_4_2_1_U19.top_add_4ns_4ns_4_2_1_Adder_12_U.u1.b ;
assign { \add_4ns_4ns_4_2_1_U19.top_add_4ns_4ns_4_2_1_Adder_12_U.u1.cout , \add_4ns_4ns_4_2_1_U19.top_add_4ns_4ns_4_2_1_Adder_12_U.u1.s  } = _168_ + \add_4ns_4ns_4_2_1_U19.top_add_4ns_4ns_4_2_1_Adder_12_U.u1.cin ;
assign _169_ = \add_4ns_4ns_4_2_1_U19.top_add_4ns_4ns_4_2_1_Adder_12_U.u2.a  + \add_4ns_4ns_4_2_1_U19.top_add_4ns_4ns_4_2_1_Adder_12_U.u2.b ;
assign { \add_4ns_4ns_4_2_1_U19.top_add_4ns_4ns_4_2_1_Adder_12_U.u2.cout , \add_4ns_4ns_4_2_1_U19.top_add_4ns_4ns_4_2_1_Adder_12_U.u2.s  } = _169_ + \add_4ns_4ns_4_2_1_U19.top_add_4ns_4ns_4_2_1_Adder_12_U.u2.cin ;
always @(posedge \add_5s_5ns_5_2_1_U1.top_add_5s_5ns_5_2_1_Adder_0_U.clk )
\add_5s_5ns_5_2_1_U1.top_add_5s_5ns_5_2_1_Adder_0_U.bin_s1  <= _171_;
always @(posedge \add_5s_5ns_5_2_1_U1.top_add_5s_5ns_5_2_1_Adder_0_U.clk )
\add_5s_5ns_5_2_1_U1.top_add_5s_5ns_5_2_1_Adder_0_U.ain_s1  <= _170_;
always @(posedge \add_5s_5ns_5_2_1_U1.top_add_5s_5ns_5_2_1_Adder_0_U.clk )
\add_5s_5ns_5_2_1_U1.top_add_5s_5ns_5_2_1_Adder_0_U.sum_s1  <= _173_;
always @(posedge \add_5s_5ns_5_2_1_U1.top_add_5s_5ns_5_2_1_Adder_0_U.clk )
\add_5s_5ns_5_2_1_U1.top_add_5s_5ns_5_2_1_Adder_0_U.carry_s1  <= _172_;
assign _171_ = \add_5s_5ns_5_2_1_U1.top_add_5s_5ns_5_2_1_Adder_0_U.ce  ? \add_5s_5ns_5_2_1_U1.top_add_5s_5ns_5_2_1_Adder_0_U.b [4:2] : \add_5s_5ns_5_2_1_U1.top_add_5s_5ns_5_2_1_Adder_0_U.bin_s1 ;
assign _170_ = \add_5s_5ns_5_2_1_U1.top_add_5s_5ns_5_2_1_Adder_0_U.ce  ? \add_5s_5ns_5_2_1_U1.top_add_5s_5ns_5_2_1_Adder_0_U.a [4:2] : \add_5s_5ns_5_2_1_U1.top_add_5s_5ns_5_2_1_Adder_0_U.ain_s1 ;
assign _172_ = \add_5s_5ns_5_2_1_U1.top_add_5s_5ns_5_2_1_Adder_0_U.ce  ? \add_5s_5ns_5_2_1_U1.top_add_5s_5ns_5_2_1_Adder_0_U.facout_s1  : \add_5s_5ns_5_2_1_U1.top_add_5s_5ns_5_2_1_Adder_0_U.carry_s1 ;
assign _173_ = \add_5s_5ns_5_2_1_U1.top_add_5s_5ns_5_2_1_Adder_0_U.ce  ? \add_5s_5ns_5_2_1_U1.top_add_5s_5ns_5_2_1_Adder_0_U.fas_s1  : \add_5s_5ns_5_2_1_U1.top_add_5s_5ns_5_2_1_Adder_0_U.sum_s1 ;
assign _174_ = \add_5s_5ns_5_2_1_U1.top_add_5s_5ns_5_2_1_Adder_0_U.u1.a  + \add_5s_5ns_5_2_1_U1.top_add_5s_5ns_5_2_1_Adder_0_U.u1.b ;
assign { \add_5s_5ns_5_2_1_U1.top_add_5s_5ns_5_2_1_Adder_0_U.u1.cout , \add_5s_5ns_5_2_1_U1.top_add_5s_5ns_5_2_1_Adder_0_U.u1.s  } = _174_ + \add_5s_5ns_5_2_1_U1.top_add_5s_5ns_5_2_1_Adder_0_U.u1.cin ;
assign _175_ = \add_5s_5ns_5_2_1_U1.top_add_5s_5ns_5_2_1_Adder_0_U.u2.a  + \add_5s_5ns_5_2_1_U1.top_add_5s_5ns_5_2_1_Adder_0_U.u2.b ;
assign { \add_5s_5ns_5_2_1_U1.top_add_5s_5ns_5_2_1_Adder_0_U.u2.cout , \add_5s_5ns_5_2_1_U1.top_add_5s_5ns_5_2_1_Adder_0_U.u2.s  } = _175_ + \add_5s_5ns_5_2_1_U1.top_add_5s_5ns_5_2_1_Adder_0_U.u2.cin ;
always @(posedge \add_7s_7ns_7_2_1_U3.top_add_7s_7ns_7_2_1_Adder_2_U.clk )
\add_7s_7ns_7_2_1_U3.top_add_7s_7ns_7_2_1_Adder_2_U.bin_s1  <= _177_;
always @(posedge \add_7s_7ns_7_2_1_U3.top_add_7s_7ns_7_2_1_Adder_2_U.clk )
\add_7s_7ns_7_2_1_U3.top_add_7s_7ns_7_2_1_Adder_2_U.ain_s1  <= _176_;
always @(posedge \add_7s_7ns_7_2_1_U3.top_add_7s_7ns_7_2_1_Adder_2_U.clk )
\add_7s_7ns_7_2_1_U3.top_add_7s_7ns_7_2_1_Adder_2_U.sum_s1  <= _179_;
always @(posedge \add_7s_7ns_7_2_1_U3.top_add_7s_7ns_7_2_1_Adder_2_U.clk )
\add_7s_7ns_7_2_1_U3.top_add_7s_7ns_7_2_1_Adder_2_U.carry_s1  <= _178_;
assign _177_ = \add_7s_7ns_7_2_1_U3.top_add_7s_7ns_7_2_1_Adder_2_U.ce  ? \add_7s_7ns_7_2_1_U3.top_add_7s_7ns_7_2_1_Adder_2_U.b [6:3] : \add_7s_7ns_7_2_1_U3.top_add_7s_7ns_7_2_1_Adder_2_U.bin_s1 ;
assign _176_ = \add_7s_7ns_7_2_1_U3.top_add_7s_7ns_7_2_1_Adder_2_U.ce  ? \add_7s_7ns_7_2_1_U3.top_add_7s_7ns_7_2_1_Adder_2_U.a [6:3] : \add_7s_7ns_7_2_1_U3.top_add_7s_7ns_7_2_1_Adder_2_U.ain_s1 ;
assign _178_ = \add_7s_7ns_7_2_1_U3.top_add_7s_7ns_7_2_1_Adder_2_U.ce  ? \add_7s_7ns_7_2_1_U3.top_add_7s_7ns_7_2_1_Adder_2_U.facout_s1  : \add_7s_7ns_7_2_1_U3.top_add_7s_7ns_7_2_1_Adder_2_U.carry_s1 ;
assign _179_ = \add_7s_7ns_7_2_1_U3.top_add_7s_7ns_7_2_1_Adder_2_U.ce  ? \add_7s_7ns_7_2_1_U3.top_add_7s_7ns_7_2_1_Adder_2_U.fas_s1  : \add_7s_7ns_7_2_1_U3.top_add_7s_7ns_7_2_1_Adder_2_U.sum_s1 ;
assign _180_ = \add_7s_7ns_7_2_1_U3.top_add_7s_7ns_7_2_1_Adder_2_U.u1.a  + \add_7s_7ns_7_2_1_U3.top_add_7s_7ns_7_2_1_Adder_2_U.u1.b ;
assign { \add_7s_7ns_7_2_1_U3.top_add_7s_7ns_7_2_1_Adder_2_U.u1.cout , \add_7s_7ns_7_2_1_U3.top_add_7s_7ns_7_2_1_Adder_2_U.u1.s  } = _180_ + \add_7s_7ns_7_2_1_U3.top_add_7s_7ns_7_2_1_Adder_2_U.u1.cin ;
assign _181_ = \add_7s_7ns_7_2_1_U3.top_add_7s_7ns_7_2_1_Adder_2_U.u2.a  + \add_7s_7ns_7_2_1_U3.top_add_7s_7ns_7_2_1_Adder_2_U.u2.b ;
assign { \add_7s_7ns_7_2_1_U3.top_add_7s_7ns_7_2_1_Adder_2_U.u2.cout , \add_7s_7ns_7_2_1_U3.top_add_7s_7ns_7_2_1_Adder_2_U.u2.s  } = _181_ + \add_7s_7ns_7_2_1_U3.top_add_7s_7ns_7_2_1_Adder_2_U.u2.cin ;
always @(posedge \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_8_U.clk )
\add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_8_U.bin_s1  <= _183_;
always @(posedge \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_8_U.clk )
\add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_8_U.ain_s1  <= _182_;
always @(posedge \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_8_U.clk )
\add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_8_U.sum_s1  <= _185_;
always @(posedge \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_8_U.clk )
\add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_8_U.carry_s1  <= _184_;
assign _183_ = \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_8_U.ce  ? \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_8_U.b [7:4] : \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_8_U.bin_s1 ;
assign _182_ = \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_8_U.ce  ? \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_8_U.a [7:4] : \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_8_U.ain_s1 ;
assign _184_ = \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_8_U.ce  ? \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_8_U.facout_s1  : \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_8_U.carry_s1 ;
assign _185_ = \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_8_U.ce  ? \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_8_U.fas_s1  : \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_8_U.sum_s1 ;
assign _186_ = \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_8_U.u1.a  + \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_8_U.u1.b ;
assign { \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_8_U.u1.cout , \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_8_U.u1.s  } = _186_ + \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_8_U.u1.cin ;
assign _187_ = \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_8_U.u2.a  + \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_8_U.u2.b ;
assign { \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_8_U.u2.cout , \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_8_U.u2.s  } = _187_ + \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_8_U.u2.cin ;
always @(posedge \add_8s_8s_8_2_1_U15.top_add_8s_8s_8_2_1_Adder_9_U.clk )
\add_8s_8s_8_2_1_U15.top_add_8s_8s_8_2_1_Adder_9_U.bin_s1  <= _189_;
always @(posedge \add_8s_8s_8_2_1_U15.top_add_8s_8s_8_2_1_Adder_9_U.clk )
\add_8s_8s_8_2_1_U15.top_add_8s_8s_8_2_1_Adder_9_U.ain_s1  <= _188_;
always @(posedge \add_8s_8s_8_2_1_U15.top_add_8s_8s_8_2_1_Adder_9_U.clk )
\add_8s_8s_8_2_1_U15.top_add_8s_8s_8_2_1_Adder_9_U.sum_s1  <= _191_;
always @(posedge \add_8s_8s_8_2_1_U15.top_add_8s_8s_8_2_1_Adder_9_U.clk )
\add_8s_8s_8_2_1_U15.top_add_8s_8s_8_2_1_Adder_9_U.carry_s1  <= _190_;
assign _189_ = \add_8s_8s_8_2_1_U15.top_add_8s_8s_8_2_1_Adder_9_U.ce  ? \add_8s_8s_8_2_1_U15.top_add_8s_8s_8_2_1_Adder_9_U.b [7:4] : \add_8s_8s_8_2_1_U15.top_add_8s_8s_8_2_1_Adder_9_U.bin_s1 ;
assign _188_ = \add_8s_8s_8_2_1_U15.top_add_8s_8s_8_2_1_Adder_9_U.ce  ? \add_8s_8s_8_2_1_U15.top_add_8s_8s_8_2_1_Adder_9_U.a [7:4] : \add_8s_8s_8_2_1_U15.top_add_8s_8s_8_2_1_Adder_9_U.ain_s1 ;
assign _190_ = \add_8s_8s_8_2_1_U15.top_add_8s_8s_8_2_1_Adder_9_U.ce  ? \add_8s_8s_8_2_1_U15.top_add_8s_8s_8_2_1_Adder_9_U.facout_s1  : \add_8s_8s_8_2_1_U15.top_add_8s_8s_8_2_1_Adder_9_U.carry_s1 ;
assign _191_ = \add_8s_8s_8_2_1_U15.top_add_8s_8s_8_2_1_Adder_9_U.ce  ? \add_8s_8s_8_2_1_U15.top_add_8s_8s_8_2_1_Adder_9_U.fas_s1  : \add_8s_8s_8_2_1_U15.top_add_8s_8s_8_2_1_Adder_9_U.sum_s1 ;
assign _192_ = \add_8s_8s_8_2_1_U15.top_add_8s_8s_8_2_1_Adder_9_U.u1.a  + \add_8s_8s_8_2_1_U15.top_add_8s_8s_8_2_1_Adder_9_U.u1.b ;
assign { \add_8s_8s_8_2_1_U15.top_add_8s_8s_8_2_1_Adder_9_U.u1.cout , \add_8s_8s_8_2_1_U15.top_add_8s_8s_8_2_1_Adder_9_U.u1.s  } = _192_ + \add_8s_8s_8_2_1_U15.top_add_8s_8s_8_2_1_Adder_9_U.u1.cin ;
assign _193_ = \add_8s_8s_8_2_1_U15.top_add_8s_8s_8_2_1_Adder_9_U.u2.a  + \add_8s_8s_8_2_1_U15.top_add_8s_8s_8_2_1_Adder_9_U.u2.b ;
assign { \add_8s_8s_8_2_1_U15.top_add_8s_8s_8_2_1_Adder_9_U.u2.cout , \add_8s_8s_8_2_1_U15.top_add_8s_8s_8_2_1_Adder_9_U.u2.s  } = _193_ + \add_8s_8s_8_2_1_U15.top_add_8s_8s_8_2_1_Adder_9_U.u2.cin ;
always @(posedge \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_1_U.clk )
\add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_1_U.bin_s1  <= _195_;
always @(posedge \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_1_U.clk )
\add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_1_U.ain_s1  <= _194_;
always @(posedge \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_1_U.clk )
\add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_1_U.sum_s1  <= _197_;
always @(posedge \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_1_U.clk )
\add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_1_U.carry_s1  <= _196_;
assign _195_ = \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_1_U.ce  ? \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_1_U.b [8:4] : \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_1_U.bin_s1 ;
assign _194_ = \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_1_U.ce  ? \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_1_U.a [8:4] : \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_1_U.ain_s1 ;
assign _196_ = \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_1_U.ce  ? \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_1_U.facout_s1  : \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_1_U.carry_s1 ;
assign _197_ = \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_1_U.ce  ? \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_1_U.fas_s1  : \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_1_U.sum_s1 ;
assign _198_ = \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_1_U.u1.a  + \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_1_U.u1.b ;
assign { \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_1_U.u1.cout , \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_1_U.u1.s  } = _198_ + \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_1_U.u1.cin ;
assign _199_ = \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_1_U.u2.a  + \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_1_U.u2.b ;
assign { \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_1_U.u2.cout , \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_1_U.u2.s  } = _199_ + \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_1_U.u2.cin ;
always @(posedge \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_1_U.clk )
\add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_1_U.bin_s1  <= _201_;
always @(posedge \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_1_U.clk )
\add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_1_U.ain_s1  <= _200_;
always @(posedge \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_1_U.clk )
\add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_1_U.sum_s1  <= _203_;
always @(posedge \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_1_U.clk )
\add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_1_U.carry_s1  <= _202_;
assign _201_ = \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_1_U.ce  ? \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_1_U.b [8:4] : \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_1_U.bin_s1 ;
assign _200_ = \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_1_U.ce  ? \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_1_U.a [8:4] : \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_1_U.ain_s1 ;
assign _202_ = \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_1_U.ce  ? \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_1_U.facout_s1  : \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_1_U.carry_s1 ;
assign _203_ = \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_1_U.ce  ? \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_1_U.fas_s1  : \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_1_U.sum_s1 ;
assign _204_ = \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_1_U.u1.a  + \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_1_U.u1.b ;
assign { \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_1_U.u1.cout , \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_1_U.u1.s  } = _204_ + \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_1_U.u1.cin ;
assign _205_ = \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_1_U.u2.a  + \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_1_U.u2.b ;
assign { \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_1_U.u2.cout , \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_1_U.u2.s  } = _205_ + \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_1_U.u2.cin ;
assign \sub_17s_17ns_17_2_1_U10.top_sub_17s_17ns_17_2_1_Adder_7_U.bin_s0  = ~ \sub_17s_17ns_17_2_1_U10.top_sub_17s_17ns_17_2_1_Adder_7_U.b ;
always @(posedge \sub_17s_17ns_17_2_1_U10.top_sub_17s_17ns_17_2_1_Adder_7_U.clk )
\sub_17s_17ns_17_2_1_U10.top_sub_17s_17ns_17_2_1_Adder_7_U.bin_s1  <= _207_;
always @(posedge \sub_17s_17ns_17_2_1_U10.top_sub_17s_17ns_17_2_1_Adder_7_U.clk )
\sub_17s_17ns_17_2_1_U10.top_sub_17s_17ns_17_2_1_Adder_7_U.ain_s1  <= _206_;
always @(posedge \sub_17s_17ns_17_2_1_U10.top_sub_17s_17ns_17_2_1_Adder_7_U.clk )
\sub_17s_17ns_17_2_1_U10.top_sub_17s_17ns_17_2_1_Adder_7_U.sum_s1  <= _209_;
always @(posedge \sub_17s_17ns_17_2_1_U10.top_sub_17s_17ns_17_2_1_Adder_7_U.clk )
\sub_17s_17ns_17_2_1_U10.top_sub_17s_17ns_17_2_1_Adder_7_U.carry_s1  <= _208_;
assign _207_ = \sub_17s_17ns_17_2_1_U10.top_sub_17s_17ns_17_2_1_Adder_7_U.ce  ? \sub_17s_17ns_17_2_1_U10.top_sub_17s_17ns_17_2_1_Adder_7_U.bin_s0 [16:8] : \sub_17s_17ns_17_2_1_U10.top_sub_17s_17ns_17_2_1_Adder_7_U.bin_s1 ;
assign _206_ = \sub_17s_17ns_17_2_1_U10.top_sub_17s_17ns_17_2_1_Adder_7_U.ce  ? \sub_17s_17ns_17_2_1_U10.top_sub_17s_17ns_17_2_1_Adder_7_U.a [16:8] : \sub_17s_17ns_17_2_1_U10.top_sub_17s_17ns_17_2_1_Adder_7_U.ain_s1 ;
assign _208_ = \sub_17s_17ns_17_2_1_U10.top_sub_17s_17ns_17_2_1_Adder_7_U.ce  ? \sub_17s_17ns_17_2_1_U10.top_sub_17s_17ns_17_2_1_Adder_7_U.facout_s1  : \sub_17s_17ns_17_2_1_U10.top_sub_17s_17ns_17_2_1_Adder_7_U.carry_s1 ;
assign _209_ = \sub_17s_17ns_17_2_1_U10.top_sub_17s_17ns_17_2_1_Adder_7_U.ce  ? \sub_17s_17ns_17_2_1_U10.top_sub_17s_17ns_17_2_1_Adder_7_U.fas_s1  : \sub_17s_17ns_17_2_1_U10.top_sub_17s_17ns_17_2_1_Adder_7_U.sum_s1 ;
assign _210_ = \sub_17s_17ns_17_2_1_U10.top_sub_17s_17ns_17_2_1_Adder_7_U.u1.a  + \sub_17s_17ns_17_2_1_U10.top_sub_17s_17ns_17_2_1_Adder_7_U.u1.b ;
assign { \sub_17s_17ns_17_2_1_U10.top_sub_17s_17ns_17_2_1_Adder_7_U.u1.cout , \sub_17s_17ns_17_2_1_U10.top_sub_17s_17ns_17_2_1_Adder_7_U.u1.s  } = _210_ + \sub_17s_17ns_17_2_1_U10.top_sub_17s_17ns_17_2_1_Adder_7_U.u1.cin ;
assign _211_ = \sub_17s_17ns_17_2_1_U10.top_sub_17s_17ns_17_2_1_Adder_7_U.u2.a  + \sub_17s_17ns_17_2_1_U10.top_sub_17s_17ns_17_2_1_Adder_7_U.u2.b ;
assign { \sub_17s_17ns_17_2_1_U10.top_sub_17s_17ns_17_2_1_Adder_7_U.u2.cout , \sub_17s_17ns_17_2_1_U10.top_sub_17s_17ns_17_2_1_Adder_7_U.u2.s  } = _211_ + \sub_17s_17ns_17_2_1_U10.top_sub_17s_17ns_17_2_1_Adder_7_U.u2.cin ;
assign _212_ = | op_6[10:0];
assign _213_ = | op_9[2:0];
assign _214_ = | op_12[2:0];
assign _215_ = | op_5[2:0];
assign _216_ = | trunc_ln718_reg_1201;
assign or_ln340_1_fu_876_p2 = or_ln340_reg_1378 | neg_src_fu_871_p2;
assign or_ln340_fu_833_p2 = overflow_fu_828_p2 | and_ln786_reg_1367;
assign or_ln412_fu_718_p2 = r_reg_1226 | add_ln1192_1_reg_1246[4];
assign or_ln781_fu_866_p2 = xor_ln781_fu_861_p2 | p_Result_14_reg_1312;
assign or_ln785_1_fu_901_p2 = p_Result_11_reg_1251 | and_ln785_fu_897_p2;
assign or_ln785_fu_823_p2 = xor_ln785_fu_818_p2 | p_Result_14_reg_1312;
always @(posedge ap_clk)
sext_ln850_reg_1016 <= _052_;
always @(posedge ap_clk)
select_ln353_reg_1028 <= _051_;
always @(posedge ap_clk)
select_ln340_reg_1388 <= _050_;
always @(posedge ap_clk)
select_ln215_reg_976 <= _049_;
always @(posedge ap_clk)
ret_reg_986 <= _048_;
always @(posedge ap_clk)
ret_V_28_reg_1419 <= _045_;
always @(posedge ap_clk)
ret_V_24_cast_reg_1424 <= _040_;
always @(posedge ap_clk)
ret_V_21_reg_1112 <= _037_;
always @(posedge ap_clk)
xor_ln416_reg_1330 <= _058_;
always @(posedge ap_clk)
ret_V_25_reg_1336 <= _042_;
always @(posedge ap_clk)
ret_V_21_cast_reg_1341 <= _036_;
always @(posedge ap_clk)
ret_V_20_reg_1095 <= _035_;
always @(posedge ap_clk)
ret_V_8_cast_reg_1100 <= _047_;
always @(posedge ap_clk)
ret_V_18_reg_1065 <= _034_;
always @(posedge ap_clk)
ret_V_17_reg_1048 <= _033_;
always @(posedge ap_clk)
ret_V_4_cast_reg_1053 <= _046_;
always @(posedge ap_clk)
ret_V_15_reg_1006 <= _032_;
always @(posedge ap_clk)
tmp_1_reg_1011 <= _053_;
always @(posedge ap_clk)
trunc_ln_reg_1152 <= _057_;
always @(posedge ap_clk)
tmp_reg_1157 <= _054_;
always @(posedge ap_clk)
trunc_ln410_reg_1162 <= _055_;
always @(posedge ap_clk)
ret_V_22_reg_1167 <= _038_;
always @(posedge ap_clk)
ret_V_14_cast_reg_1172 <= _031_;
always @(posedge ap_clk)
r_reg_1226 <= _030_;
always @(posedge ap_clk)
p_Val2_5_reg_1306 <= _029_;
always @(posedge ap_clk)
p_Result_14_reg_1312 <= _027_;
always @(posedge ap_clk)
or_ln340_reg_1378 <= _024_;
always @(posedge ap_clk)
ret_V_26_reg_1383 <= _043_;
always @(posedge ap_clk)
op_29_V_reg_1296 <= _023_;
always @(posedge ap_clk)
op_25_V_reg_1122 <= _022_;
always @(posedge ap_clk)
op_23_V_reg_1075 <= _021_;
always @(posedge ap_clk)
op_19_V_reg_1398 <= _020_;
always @(posedge ap_clk)
ret_V_27_reg_1404 <= _044_;
always @(posedge ap_clk)
op_11_V_reg_1194 <= _019_;
always @(posedge ap_clk)
trunc_ln718_reg_1201 <= _056_;
always @(posedge ap_clk)
ret_V_23_reg_1206 <= _039_;
always @(posedge ap_clk)
icmp_ln851_reg_1001 <= _018_;
always @(posedge ap_clk)
icmp_ln851_3_reg_1147 <= _017_;
always @(posedge ap_clk)
icmp_ln851_2_reg_1090 <= _016_;
always @(posedge ap_clk)
icmp_ln851_1_reg_1043 <= _015_;
always @(posedge ap_clk)
icmp_ln410_reg_1179 <= _014_;
always @(posedge ap_clk)
and_ln412_reg_1281 <= _009_;
always @(posedge ap_clk)
add_ln691_reg_1023 <= _007_;
always @(posedge ap_clk)
add_ln691_5_reg_1431 <= _006_;
always @(posedge ap_clk)
deleted_zeros_reg_1361 <= _013_;
always @(posedge ap_clk)
and_ln786_reg_1367 <= _010_;
always @(posedge ap_clk)
add_ln691_4_reg_1373 <= _005_;
always @(posedge ap_clk)
add_ln691_3_reg_1189 <= _004_;
always @(posedge ap_clk)
add_ln691_2_reg_1107 <= _003_;
always @(posedge ap_clk)
add_ln691_1_reg_1060 <= _002_;
always @(posedge ap_clk)
add_ln1192_1_reg_1246 <= _001_;
always @(posedge ap_clk)
p_Result_11_reg_1251 <= _025_;
always @(posedge ap_clk)
p_Val2_4_reg_1260 <= _028_;
always @(posedge ap_clk)
p_Result_13_reg_1265 <= _026_;
always @(posedge ap_clk)
ret_V_24_reg_1271 <= _041_;
always @(posedge ap_clk)
add_ln69_reg_1276 <= _008_;
always @(posedge ap_clk)
carry_1_reg_1348 <= _012_;
always @(posedge ap_clk)
Range1_all_zeros_reg_1354 <= _000_;
always @(posedge ap_clk)
ap_CS_fsm <= _011_;
assign _059_ = _065_ ? 2'h2 : 2'h1;
assign _217_ = ap_CS_fsm == 1'h1;
function [42:0] _640_;
input [42:0] a;
input [1848:0] b;
input [42:0] s;
case (s)
43'b0000000000000000000000000000000000000000001:
_640_ = b[42:0];
43'b0000000000000000000000000000000000000000010:
_640_ = b[85:43];
43'b0000000000000000000000000000000000000000100:
_640_ = b[128:86];
43'b0000000000000000000000000000000000000001000:
_640_ = b[171:129];
43'b0000000000000000000000000000000000000010000:
_640_ = b[214:172];
43'b0000000000000000000000000000000000000100000:
_640_ = b[257:215];
43'b0000000000000000000000000000000000001000000:
_640_ = b[300:258];
43'b0000000000000000000000000000000000010000000:
_640_ = b[343:301];
43'b0000000000000000000000000000000000100000000:
_640_ = b[386:344];
43'b0000000000000000000000000000000001000000000:
_640_ = b[429:387];
43'b0000000000000000000000000000000010000000000:
_640_ = b[472:430];
43'b0000000000000000000000000000000100000000000:
_640_ = b[515:473];
43'b0000000000000000000000000000001000000000000:
_640_ = b[558:516];
43'b0000000000000000000000000000010000000000000:
_640_ = b[601:559];
43'b0000000000000000000000000000100000000000000:
_640_ = b[644:602];
43'b0000000000000000000000000001000000000000000:
_640_ = b[687:645];
43'b0000000000000000000000000010000000000000000:
_640_ = b[730:688];
43'b0000000000000000000000000100000000000000000:
_640_ = b[773:731];
43'b0000000000000000000000001000000000000000000:
_640_ = b[816:774];
43'b0000000000000000000000010000000000000000000:
_640_ = b[859:817];
43'b0000000000000000000000100000000000000000000:
_640_ = b[902:860];
43'b0000000000000000000001000000000000000000000:
_640_ = b[945:903];
43'b0000000000000000000010000000000000000000000:
_640_ = b[988:946];
43'b0000000000000000000100000000000000000000000:
_640_ = b[1031:989];
43'b0000000000000000001000000000000000000000000:
_640_ = b[1074:1032];
43'b0000000000000000010000000000000000000000000:
_640_ = b[1117:1075];
43'b0000000000000000100000000000000000000000000:
_640_ = b[1160:1118];
43'b0000000000000001000000000000000000000000000:
_640_ = b[1203:1161];
43'b0000000000000010000000000000000000000000000:
_640_ = b[1246:1204];
43'b0000000000000100000000000000000000000000000:
_640_ = b[1289:1247];
43'b0000000000001000000000000000000000000000000:
_640_ = b[1332:1290];
43'b0000000000010000000000000000000000000000000:
_640_ = b[1375:1333];
43'b0000000000100000000000000000000000000000000:
_640_ = b[1418:1376];
43'b0000000001000000000000000000000000000000000:
_640_ = b[1461:1419];
43'b0000000010000000000000000000000000000000000:
_640_ = b[1504:1462];
43'b0000000100000000000000000000000000000000000:
_640_ = b[1547:1505];
43'b0000001000000000000000000000000000000000000:
_640_ = b[1590:1548];
43'b0000010000000000000000000000000000000000000:
_640_ = b[1633:1591];
43'b0000100000000000000000000000000000000000000:
_640_ = b[1676:1634];
43'b0001000000000000000000000000000000000000000:
_640_ = b[1719:1677];
43'b0010000000000000000000000000000000000000000:
_640_ = b[1762:1720];
43'b0100000000000000000000000000000000000000000:
_640_ = b[1805:1763];
43'b1000000000000000000000000000000000000000000:
_640_ = b[1848:1806];
43'b0000000000000000000000000000000000000000000:
_640_ = a;
default:
_640_ = 43'bx;
endcase
endfunction
assign ap_NS_fsm = _640_(43'hxxxxxxxxxxx, { 41'h00000000000, _059_, 1806'h00000000002000000000080000000002000000000080000000002000000000080000000002000000000080000000002000000000080000000002000000000080000000002000000000080000000002000000000080000000002000000000080000000002000000000080000000002000000000080000000002000000000080000000002000000000080000000002000000000080000000002000000000080000000002000000000080000000002000000000080000000002000000000080000000002000000000080000000002000000000080000000002000000000000000000001 }, { _217_, _259_, _258_, _257_, _256_, _255_, _254_, _253_, _252_, _251_, _250_, _249_, _248_, _247_, _246_, _245_, _244_, _243_, _242_, _241_, _240_, _239_, _238_, _237_, _236_, _235_, _234_, _233_, _232_, _231_, _230_, _229_, _228_, _227_, _226_, _225_, _224_, _223_, _222_, _221_, _220_, _219_, _218_ });
assign _218_ = ap_CS_fsm == 43'h40000000000;
assign _219_ = ap_CS_fsm == 42'h20000000000;
assign _220_ = ap_CS_fsm == 41'h10000000000;
assign _221_ = ap_CS_fsm == 40'h8000000000;
assign _222_ = ap_CS_fsm == 39'h4000000000;
assign _223_ = ap_CS_fsm == 38'h2000000000;
assign _224_ = ap_CS_fsm == 37'h1000000000;
assign _225_ = ap_CS_fsm == 36'h800000000;
assign _226_ = ap_CS_fsm == 35'h400000000;
assign _227_ = ap_CS_fsm == 34'h200000000;
assign _228_ = ap_CS_fsm == 33'h100000000;
assign _229_ = ap_CS_fsm == 32'd2147483648;
assign _230_ = ap_CS_fsm == 31'h40000000;
assign _231_ = ap_CS_fsm == 30'h20000000;
assign _232_ = ap_CS_fsm == 29'h10000000;
assign _233_ = ap_CS_fsm == 28'h8000000;
assign _234_ = ap_CS_fsm == 27'h4000000;
assign _235_ = ap_CS_fsm == 26'h2000000;
assign _236_ = ap_CS_fsm == 25'h1000000;
assign _237_ = ap_CS_fsm == 24'h800000;
assign _238_ = ap_CS_fsm == 23'h400000;
assign _239_ = ap_CS_fsm == 22'h200000;
assign _240_ = ap_CS_fsm == 21'h100000;
assign _241_ = ap_CS_fsm == 20'h80000;
assign _242_ = ap_CS_fsm == 19'h40000;
assign _243_ = ap_CS_fsm == 18'h20000;
assign _244_ = ap_CS_fsm == 17'h10000;
assign _245_ = ap_CS_fsm == 16'h8000;
assign _246_ = ap_CS_fsm == 15'h4000;
assign _247_ = ap_CS_fsm == 14'h2000;
assign _248_ = ap_CS_fsm == 13'h1000;
assign _249_ = ap_CS_fsm == 12'h800;
assign _250_ = ap_CS_fsm == 11'h400;
assign _251_ = ap_CS_fsm == 10'h200;
assign _252_ = ap_CS_fsm == 9'h100;
assign _253_ = ap_CS_fsm == 8'h80;
assign _254_ = ap_CS_fsm == 7'h40;
assign _255_ = ap_CS_fsm == 6'h20;
assign _256_ = ap_CS_fsm == 5'h10;
assign _257_ = ap_CS_fsm == 4'h8;
assign _258_ = ap_CS_fsm == 3'h4;
assign _259_ = ap_CS_fsm == 2'h2;
assign op_32_ap_vld = ap_CS_fsm[42] ? 1'h1 : 1'h0;
assign ap_idle = _064_ ? 1'h1 : 1'h0;
assign _052_ = ap_CS_fsm[5] ? { tmp_1_reg_1011[5], tmp_1_reg_1011 } : sext_ln850_reg_1016;
assign _051_ = ap_CS_fsm[7] ? select_ln353_fu_330_p3 : select_ln353_reg_1028;
assign _050_ = ap_CS_fsm[36] ? select_ln340_fu_881_p3 : select_ln340_reg_1388;
assign _049_ = ap_CS_fsm[0] ? select_ln215_fu_251_p3 : select_ln215_reg_976;
assign _048_ = ap_CS_fsm[2] ? grp_fu_263_p2 : ret_reg_986;
assign _040_ = ap_CS_fsm[39] ? grp_fu_931_p2[32:1] : ret_V_24_cast_reg_1424;
assign _045_ = ap_CS_fsm[39] ? grp_fu_931_p2 : ret_V_28_reg_1419;
assign _037_ = ap_CS_fsm[19] ? ret_V_21_fu_469_p3 : ret_V_21_reg_1112;
assign _036_ = ap_CS_fsm[32] ? grp_fu_768_p2[32:1] : ret_V_21_cast_reg_1341;
assign _042_ = ap_CS_fsm[32] ? grp_fu_768_p2 : ret_V_25_reg_1336;
assign _058_ = ap_CS_fsm[32] ? xor_ln416_fu_774_p2 : xor_ln416_reg_1330;
assign _047_ = ap_CS_fsm[16] ? grp_fu_426_p2[34:3] : ret_V_8_cast_reg_1100;
assign _035_ = ap_CS_fsm[16] ? grp_fu_426_p2 : ret_V_20_reg_1095;
assign _034_ = ap_CS_fsm[12] ? ret_V_18_fu_395_p3 : ret_V_18_reg_1065;
assign _046_ = ap_CS_fsm[9] ? grp_fu_352_p2[42:11] : ret_V_4_cast_reg_1053;
assign _033_ = ap_CS_fsm[9] ? grp_fu_352_p2 : ret_V_17_reg_1048;
assign _053_ = ap_CS_fsm[4] ? grp_fu_283_p2[8:3] : tmp_1_reg_1011;
assign _032_ = ap_CS_fsm[4] ? grp_fu_283_p2 : ret_V_15_reg_1006;
assign _031_ = ap_CS_fsm[23] ? grp_fu_522_p2[34:3] : ret_V_14_cast_reg_1172;
assign _038_ = ap_CS_fsm[23] ? grp_fu_522_p2 : ret_V_22_reg_1167;
assign _055_ = ap_CS_fsm[23] ? grp_fu_501_p2[0] : trunc_ln410_reg_1162;
assign _054_ = ap_CS_fsm[23] ? grp_fu_501_p2[16] : tmp_reg_1157;
assign _057_ = ap_CS_fsm[23] ? grp_fu_501_p2[8:1] : trunc_ln_reg_1152;
assign _030_ = ap_CS_fsm[27] ? r_fu_650_p2 : r_reg_1226;
assign _027_ = ap_CS_fsm[31] ? grp_fu_740_p2[3] : p_Result_14_reg_1312;
assign _029_ = ap_CS_fsm[31] ? grp_fu_740_p2 : p_Val2_5_reg_1306;
assign _043_ = ap_CS_fsm[35] ? ret_V_26_fu_854_p3 : ret_V_26_reg_1383;
assign _024_ = ap_CS_fsm[35] ? or_ln340_fu_833_p2 : or_ln340_reg_1378;
assign _023_ = ap_CS_fsm[30] ? grp_fu_732_p2 : op_29_V_reg_1296;
assign _022_ = ap_CS_fsm[21] ? grp_fu_480_p2 : op_25_V_reg_1122;
assign _021_ = ap_CS_fsm[14] ? grp_fu_406_p2 : op_23_V_reg_1075;
assign _044_ = ap_CS_fsm[37] ? grp_fu_892_p2 : ret_V_27_reg_1404;
assign _020_ = ap_CS_fsm[37] ? op_19_V_fu_911_p3 : op_19_V_reg_1398;
assign _039_ = ap_CS_fsm[26] ? ret_V_23_fu_613_p3 : ret_V_23_reg_1206;
assign _056_ = ap_CS_fsm[26] ? grp_fu_592_p2[2:0] : trunc_ln718_reg_1201;
assign _019_ = ap_CS_fsm[26] ? grp_fu_592_p2 : op_11_V_reg_1194;
assign _018_ = ap_CS_fsm[3] ? icmp_ln851_fu_293_p2 : icmp_ln851_reg_1001;
assign _017_ = ap_CS_fsm[22] ? icmp_ln851_3_fu_532_p2 : icmp_ln851_3_reg_1147;
assign _016_ = ap_CS_fsm[15] ? icmp_ln851_2_fu_436_p2 : icmp_ln851_2_reg_1090;
assign _015_ = ap_CS_fsm[8] ? icmp_ln851_1_fu_362_p2 : icmp_ln851_1_reg_1043;
assign _014_ = ap_CS_fsm[24] ? icmp_ln410_fu_578_p2 : icmp_ln410_reg_1179;
assign _009_ = ap_CS_fsm[29] ? and_ln412_fu_723_p2 : and_ln412_reg_1281;
assign _007_ = _063_ ? grp_fu_312_p2 : add_ln691_reg_1023;
assign _006_ = ap_CS_fsm[41] ? grp_fu_947_p2 : add_ln691_5_reg_1431;
assign _005_ = ap_CS_fsm[34] ? grp_fu_798_p2 : add_ln691_4_reg_1373;
assign _010_ = ap_CS_fsm[34] ? and_ln786_fu_813_p2 : and_ln786_reg_1367;
assign _013_ = ap_CS_fsm[34] ? deleted_zeros_fu_803_p3 : deleted_zeros_reg_1361;
assign _004_ = _062_ ? grp_fu_584_p2 : add_ln691_3_reg_1189;
assign _003_ = _061_ ? grp_fu_452_p2 : add_ln691_2_reg_1107;
assign _002_ = _060_ ? grp_fu_378_p2 : add_ln691_1_reg_1060;
assign _008_ = ap_CS_fsm[28] ? grp_fu_672_p2 : add_ln69_reg_1276;
assign _041_ = ap_CS_fsm[28] ? grp_fu_659_p2 : ret_V_24_reg_1271;
assign _026_ = ap_CS_fsm[28] ? grp_fu_645_p2[7] : p_Result_13_reg_1265;
assign _028_ = ap_CS_fsm[28] ? grp_fu_645_p2[7:4] : p_Val2_4_reg_1260;
assign _025_ = ap_CS_fsm[28] ? grp_fu_639_p2[8] : p_Result_11_reg_1251;
assign _001_ = ap_CS_fsm[28] ? grp_fu_645_p2 : add_ln1192_1_reg_1246;
assign _000_ = ap_CS_fsm[33] ? Range1_all_zeros_fu_793_p2 : Range1_all_zeros_reg_1354;
assign _012_ = ap_CS_fsm[33] ? carry_1_fu_789_p2 : carry_1_reg_1348;
assign _011_ = ap_rst ? 43'h00000000001 : ap_NS_fsm;
assign deleted_ones_fu_808_p3 = carry_1_reg_1348 ? Range1_all_zeros_reg_1354 : p_Result_11_reg_1251;
assign deleted_zeros_fu_803_p3 = carry_1_reg_1348 ? p_Result_11_reg_1251 : Range1_all_zeros_reg_1354;
assign icmp_ln410_fu_578_p2 = _067_ ? 1'h1 : 1'h0;
assign icmp_ln851_1_fu_362_p2 = _212_ ? 1'h1 : 1'h0;
assign icmp_ln851_2_fu_436_p2 = _213_ ? 1'h1 : 1'h0;
assign icmp_ln851_3_fu_532_p2 = _214_ ? 1'h1 : 1'h0;
assign icmp_ln851_fu_293_p2 = _215_ ? 1'h1 : 1'h0;
assign op_19_V_fu_911_p3 = and_ln785_1_fu_906_p2 ? p_Val2_5_reg_1306 : select_ln340_reg_1388;
assign op_32 = ret_V_28_reg_1419[33] ? select_ln850_5_fu_962_p3 : ret_V_24_cast_reg_1424;
assign r_fu_650_p2 = _216_ ? 1'h1 : 1'h0;
assign ret_V_18_fu_395_p3 = ret_V_17_reg_1048[43] ? select_ln850_1_fu_390_p3 : ret_V_4_cast_reg_1053;
assign ret_V_21_fu_469_p3 = ret_V_20_reg_1095[35] ? select_ln850_2_fu_464_p3 : ret_V_8_cast_reg_1100;
assign ret_V_23_fu_613_p3 = ret_V_22_reg_1167[35] ? select_ln850_3_fu_608_p3 : ret_V_14_cast_reg_1172;
assign ret_V_26_fu_854_p3 = ret_V_25_reg_1336[33] ? select_ln850_4_fu_848_p3 : ret_V_21_cast_reg_1341;
assign select_ln215_fu_251_p3 = op_0 ? 5'h1f : 5'h00;
assign select_ln340_fu_881_p3 = or_ln340_1_fu_876_p2 ? 4'h0 : p_Val2_5_reg_1306;
assign select_ln353_fu_330_p3 = ret_V_15_reg_1006[8] ? select_ln850_fu_325_p3 : sext_ln850_reg_1016;
assign select_ln850_1_fu_390_p3 = icmp_ln851_1_reg_1043 ? add_ln691_1_reg_1060 : ret_V_4_cast_reg_1053;
assign select_ln850_2_fu_464_p3 = icmp_ln851_2_reg_1090 ? add_ln691_2_reg_1107 : ret_V_8_cast_reg_1100;
assign select_ln850_3_fu_608_p3 = icmp_ln851_3_reg_1147 ? add_ln691_3_reg_1189 : ret_V_14_cast_reg_1172;
assign select_ln850_4_fu_848_p3 = op_17[0] ? add_ln691_4_reg_1373 : ret_V_21_cast_reg_1341;
assign select_ln850_5_fu_962_p3 = op_19_V_reg_1398[0] ? add_ln691_5_reg_1431 : ret_V_24_cast_reg_1424;
assign select_ln850_fu_325_p3 = icmp_ln851_reg_1001 ? add_ln691_reg_1023 : sext_ln850_reg_1016;
assign and_ln_fu_570_p4 = { tmp_reg_1157, 15'h0000, trunc_ln410_reg_1162 };
assign ap_CS_fsm_state1 = ap_CS_fsm[0];
assign ap_CS_fsm_state10 = ap_CS_fsm[9];
assign ap_CS_fsm_state11 = ap_CS_fsm[10];
assign ap_CS_fsm_state12 = ap_CS_fsm[11];
assign ap_CS_fsm_state13 = ap_CS_fsm[12];
assign ap_CS_fsm_state14 = ap_CS_fsm[13];
assign ap_CS_fsm_state15 = ap_CS_fsm[14];
assign ap_CS_fsm_state16 = ap_CS_fsm[15];
assign ap_CS_fsm_state17 = ap_CS_fsm[16];
assign ap_CS_fsm_state18 = ap_CS_fsm[17];
assign ap_CS_fsm_state19 = ap_CS_fsm[18];
assign ap_CS_fsm_state2 = ap_CS_fsm[1];
assign ap_CS_fsm_state20 = ap_CS_fsm[19];
assign ap_CS_fsm_state21 = ap_CS_fsm[20];
assign ap_CS_fsm_state22 = ap_CS_fsm[21];
assign ap_CS_fsm_state23 = ap_CS_fsm[22];
assign ap_CS_fsm_state24 = ap_CS_fsm[23];
assign ap_CS_fsm_state25 = ap_CS_fsm[24];
assign ap_CS_fsm_state26 = ap_CS_fsm[25];
assign ap_CS_fsm_state27 = ap_CS_fsm[26];
assign ap_CS_fsm_state28 = ap_CS_fsm[27];
assign ap_CS_fsm_state29 = ap_CS_fsm[28];
assign ap_CS_fsm_state3 = ap_CS_fsm[2];
assign ap_CS_fsm_state30 = ap_CS_fsm[29];
assign ap_CS_fsm_state31 = ap_CS_fsm[30];
assign ap_CS_fsm_state32 = ap_CS_fsm[31];
assign ap_CS_fsm_state33 = ap_CS_fsm[32];
assign ap_CS_fsm_state34 = ap_CS_fsm[33];
assign ap_CS_fsm_state35 = ap_CS_fsm[34];
assign ap_CS_fsm_state36 = ap_CS_fsm[35];
assign ap_CS_fsm_state37 = ap_CS_fsm[36];
assign ap_CS_fsm_state38 = ap_CS_fsm[37];
assign ap_CS_fsm_state39 = ap_CS_fsm[38];
assign ap_CS_fsm_state4 = ap_CS_fsm[3];
assign ap_CS_fsm_state40 = ap_CS_fsm[39];
assign ap_CS_fsm_state41 = ap_CS_fsm[40];
assign ap_CS_fsm_state42 = ap_CS_fsm[41];
assign ap_CS_fsm_state43 = ap_CS_fsm[42];
assign ap_CS_fsm_state5 = ap_CS_fsm[4];
assign ap_CS_fsm_state6 = ap_CS_fsm[5];
assign ap_CS_fsm_state7 = ap_CS_fsm[6];
assign ap_CS_fsm_state8 = ap_CS_fsm[7];
assign ap_CS_fsm_state9 = ap_CS_fsm[8];
assign ap_done = op_32_ap_vld;
assign ap_ready = op_32_ap_vld;
assign grp_fu_263_p0 = { op_2[3], op_2 };
assign grp_fu_283_p0 = { ret_reg_986[4], ret_reg_986, 3'h0 };
assign grp_fu_283_p1 = { op_5[7], op_5 };
assign grp_fu_312_p0 = { tmp_1_reg_1011[5], tmp_1_reg_1011 };
assign grp_fu_352_p0 = { select_ln353_reg_1028[6], select_ln353_reg_1028[6], select_ln353_reg_1028[6], select_ln353_reg_1028[6], select_ln353_reg_1028[6], select_ln353_reg_1028[6], select_ln353_reg_1028[6], select_ln353_reg_1028[6], select_ln353_reg_1028[6], select_ln353_reg_1028[6], select_ln353_reg_1028[6], select_ln353_reg_1028[6], select_ln353_reg_1028[6], select_ln353_reg_1028[6], select_ln353_reg_1028[6], select_ln353_reg_1028[6], select_ln353_reg_1028[6], select_ln353_reg_1028[6], select_ln353_reg_1028[6], select_ln353_reg_1028[6], select_ln353_reg_1028[6], select_ln353_reg_1028[6], select_ln353_reg_1028[6], select_ln353_reg_1028[6], select_ln353_reg_1028[6], select_ln353_reg_1028[6], select_ln353_reg_1028, 11'h000 };
assign grp_fu_352_p1 = { op_6[15], op_6[15], op_6[15], op_6[15], op_6[15], op_6[15], op_6[15], op_6[15], op_6[15], op_6[15], op_6[15], op_6[15], op_6[15], op_6[15], op_6[15], op_6[15], op_6[15], op_6[15], op_6[15], op_6[15], op_6[15], op_6[15], op_6[15], op_6[15], op_6[15], op_6[15], op_6[15], op_6[15], op_6 };
assign grp_fu_406_p1 = { op_8[3], op_8[3], op_8[3], op_8[3], op_8[3], op_8[3], op_8[3], op_8[3], op_8[3], op_8[3], op_8[3], op_8[3], op_8[3], op_8[3], op_8[3], op_8[3], op_8[3], op_8[3], op_8[3], op_8[3], op_8[3], op_8[3], op_8[3], op_8[3], op_8[3], op_8[3], op_8[3], op_8[3], op_8 };
assign grp_fu_426_p0 = { op_23_V_reg_1075[31], op_23_V_reg_1075, 3'h0 };
assign grp_fu_426_p1 = { op_9[3], op_9[3], op_9[3], op_9[3], op_9[3], op_9[3], op_9[3], op_9[3], op_9[3], op_9[3], op_9[3], op_9[3], op_9[3], op_9[3], op_9[3], op_9[3], op_9[3], op_9[3], op_9[3], op_9[3], op_9[3], op_9[3], op_9[3], op_9[3], op_9[3], op_9[3], op_9[3], op_9[3], op_9[3], op_9[3], op_9[3], op_9[3], op_9 };
assign grp_fu_480_p1 = { 24'h000000, op_10 };
assign grp_fu_501_p0 = { op_4[15], op_4 };
assign grp_fu_501_p1 = { 7'h00, op_1, 6'h00 };
assign grp_fu_522_p0 = { op_25_V_reg_1122[31], op_25_V_reg_1122, 3'h0 };
assign grp_fu_522_p1 = { op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12 };
assign grp_fu_592_p1 = { 7'h00, icmp_ln410_reg_1179 };
assign grp_fu_639_p0 = { op_14[1], op_14[1], op_14, 5'h00 };
assign grp_fu_639_p1 = { op_11_V_reg_1194[7], op_11_V_reg_1194 };
assign grp_fu_645_p0 = { op_14[1], op_14, 5'h00 };
assign grp_fu_659_p1 = { op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13 };
assign grp_fu_672_p0 = { op_16[7], op_16[7], op_16 };
assign grp_fu_672_p1 = { 2'h0, op_15 };
assign grp_fu_732_p0 = { add_ln69_reg_1276[9], add_ln69_reg_1276[9], add_ln69_reg_1276[9], add_ln69_reg_1276[9], add_ln69_reg_1276[9], add_ln69_reg_1276[9], add_ln69_reg_1276[9], add_ln69_reg_1276[9], add_ln69_reg_1276[9], add_ln69_reg_1276[9], add_ln69_reg_1276[9], add_ln69_reg_1276[9], add_ln69_reg_1276[9], add_ln69_reg_1276[9], add_ln69_reg_1276[9], add_ln69_reg_1276[9], add_ln69_reg_1276[9], add_ln69_reg_1276[9], add_ln69_reg_1276[9], add_ln69_reg_1276[9], add_ln69_reg_1276[9], add_ln69_reg_1276[9], add_ln69_reg_1276 };
assign grp_fu_740_p1 = { 3'h0, and_ln412_reg_1281 };
assign grp_fu_768_p0 = { op_29_V_reg_1296[31], op_29_V_reg_1296, 1'h0 };
assign grp_fu_768_p1 = { op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17 };
assign grp_fu_892_p1 = { op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18 };
assign grp_fu_931_p0 = { ret_V_27_reg_1404[31], ret_V_27_reg_1404, 1'h0 };
assign grp_fu_931_p1 = { op_19_V_reg_1398[3], op_19_V_reg_1398[3], op_19_V_reg_1398[3], op_19_V_reg_1398[3], op_19_V_reg_1398[3], op_19_V_reg_1398[3], op_19_V_reg_1398[3], op_19_V_reg_1398[3], op_19_V_reg_1398[3], op_19_V_reg_1398[3], op_19_V_reg_1398[3], op_19_V_reg_1398[3], op_19_V_reg_1398[3], op_19_V_reg_1398[3], op_19_V_reg_1398[3], op_19_V_reg_1398[3], op_19_V_reg_1398[3], op_19_V_reg_1398[3], op_19_V_reg_1398[3], op_19_V_reg_1398[3], op_19_V_reg_1398[3], op_19_V_reg_1398[3], op_19_V_reg_1398[3], op_19_V_reg_1398[3], op_19_V_reg_1398[3], op_19_V_reg_1398[3], op_19_V_reg_1398[3], op_19_V_reg_1398[3], op_19_V_reg_1398[3], op_19_V_reg_1398[3], op_19_V_reg_1398 };
assign p_Result_10_fu_952_p3 = ret_V_28_reg_1419[33];
assign p_Result_12_fu_711_p3 = op_11_V_reg_1194[3];
assign p_Result_1_fu_383_p3 = ret_V_17_reg_1048[43];
assign p_Result_5_fu_704_p3 = add_ln1192_1_reg_1246[4];
assign p_Result_7_fu_457_p3 = ret_V_20_reg_1095[35];
assign p_Result_8_fu_601_p3 = ret_V_22_reg_1167[35];
assign p_Result_9_fu_838_p3 = ret_V_25_reg_1336[33];
assign p_Result_s_fu_318_p3 = ret_V_15_reg_1006[8];
assign rhs_10_fu_757_p3 = { op_29_V_reg_1296, 1'h0 };
assign rhs_13_fu_920_p3 = { ret_V_27_reg_1404, 1'h0 };
assign rhs_1_fu_272_p3 = { ret_reg_986, 3'h0 };
assign rhs_2_fu_489_p3 = { op_1, 6'h00 };
assign rhs_3_fu_623_p3 = { op_14, 5'h00 };
assign rhs_5_fu_415_p3 = { op_23_V_reg_1075, 3'h0 };
assign rhs_7_fu_511_p3 = { op_25_V_reg_1122, 3'h0 };
assign sext_ln1192_fu_268_p0 = op_5;
assign sext_ln703_1_fu_337_p0 = op_6;
assign sext_ln703_3_fu_411_p0 = op_9;
assign sext_ln703_4_fu_507_p0 = op_12;
assign sext_ln703_5_fu_753_p0 = op_17;
assign sext_ln850_fu_309_p1 = { tmp_1_reg_1011[5], tmp_1_reg_1011 };
assign tmp_2_fu_341_p3 = { select_ln353_reg_1028, 11'h000 };
assign trunc_ln410_fu_556_p1 = grp_fu_501_p2[0];
assign trunc_ln718_fu_597_p1 = grp_fu_592_p2[2:0];
assign trunc_ln851_1_fu_358_p0 = op_6;
assign trunc_ln851_1_fu_358_p1 = op_6[10:0];
assign trunc_ln851_2_fu_432_p0 = op_9;
assign trunc_ln851_2_fu_432_p1 = op_9[2:0];
assign trunc_ln851_3_fu_528_p0 = op_12;
assign trunc_ln851_3_fu_528_p1 = op_12[2:0];
assign trunc_ln851_4_fu_845_p0 = op_17;
assign trunc_ln851_4_fu_845_p1 = op_17[0];
assign trunc_ln851_5_fu_959_p1 = op_19_V_reg_1398[0];
assign trunc_ln851_fu_289_p0 = op_5;
assign trunc_ln851_fu_289_p1 = op_5[2:0];
assign \sub_17s_17ns_17_2_1_U10.top_sub_17s_17ns_17_2_1_Adder_7_U.ain_s0  = \sub_17s_17ns_17_2_1_U10.top_sub_17s_17ns_17_2_1_Adder_7_U.a ;
assign \sub_17s_17ns_17_2_1_U10.top_sub_17s_17ns_17_2_1_Adder_7_U.s  = { \sub_17s_17ns_17_2_1_U10.top_sub_17s_17ns_17_2_1_Adder_7_U.fas_s2 , \sub_17s_17ns_17_2_1_U10.top_sub_17s_17ns_17_2_1_Adder_7_U.sum_s1  };
assign \sub_17s_17ns_17_2_1_U10.top_sub_17s_17ns_17_2_1_Adder_7_U.u2.a  = \sub_17s_17ns_17_2_1_U10.top_sub_17s_17ns_17_2_1_Adder_7_U.ain_s1 ;
assign \sub_17s_17ns_17_2_1_U10.top_sub_17s_17ns_17_2_1_Adder_7_U.u2.b  = \sub_17s_17ns_17_2_1_U10.top_sub_17s_17ns_17_2_1_Adder_7_U.bin_s1 ;
assign \sub_17s_17ns_17_2_1_U10.top_sub_17s_17ns_17_2_1_Adder_7_U.u2.cin  = \sub_17s_17ns_17_2_1_U10.top_sub_17s_17ns_17_2_1_Adder_7_U.carry_s1 ;
assign \sub_17s_17ns_17_2_1_U10.top_sub_17s_17ns_17_2_1_Adder_7_U.facout_s2  = \sub_17s_17ns_17_2_1_U10.top_sub_17s_17ns_17_2_1_Adder_7_U.u2.cout ;
assign \sub_17s_17ns_17_2_1_U10.top_sub_17s_17ns_17_2_1_Adder_7_U.fas_s2  = \sub_17s_17ns_17_2_1_U10.top_sub_17s_17ns_17_2_1_Adder_7_U.u2.s ;
assign \sub_17s_17ns_17_2_1_U10.top_sub_17s_17ns_17_2_1_Adder_7_U.u1.a  = \sub_17s_17ns_17_2_1_U10.top_sub_17s_17ns_17_2_1_Adder_7_U.a [7:0];
assign \sub_17s_17ns_17_2_1_U10.top_sub_17s_17ns_17_2_1_Adder_7_U.u1.b  = \sub_17s_17ns_17_2_1_U10.top_sub_17s_17ns_17_2_1_Adder_7_U.bin_s0 [7:0];
assign \sub_17s_17ns_17_2_1_U10.top_sub_17s_17ns_17_2_1_Adder_7_U.u1.cin  = 1'h1;
assign \sub_17s_17ns_17_2_1_U10.top_sub_17s_17ns_17_2_1_Adder_7_U.facout_s1  = \sub_17s_17ns_17_2_1_U10.top_sub_17s_17ns_17_2_1_Adder_7_U.u1.cout ;
assign \sub_17s_17ns_17_2_1_U10.top_sub_17s_17ns_17_2_1_Adder_7_U.fas_s1  = \sub_17s_17ns_17_2_1_U10.top_sub_17s_17ns_17_2_1_Adder_7_U.u1.s ;
assign \sub_17s_17ns_17_2_1_U10.top_sub_17s_17ns_17_2_1_Adder_7_U.a  = \sub_17s_17ns_17_2_1_U10.din0 ;
assign \sub_17s_17ns_17_2_1_U10.top_sub_17s_17ns_17_2_1_Adder_7_U.b  = \sub_17s_17ns_17_2_1_U10.din1 ;
assign \sub_17s_17ns_17_2_1_U10.top_sub_17s_17ns_17_2_1_Adder_7_U.ce  = \sub_17s_17ns_17_2_1_U10.ce ;
assign \sub_17s_17ns_17_2_1_U10.top_sub_17s_17ns_17_2_1_Adder_7_U.clk  = \sub_17s_17ns_17_2_1_U10.clk ;
assign \sub_17s_17ns_17_2_1_U10.top_sub_17s_17ns_17_2_1_Adder_7_U.reset  = \sub_17s_17ns_17_2_1_U10.reset ;
assign \sub_17s_17ns_17_2_1_U10.dout  = \sub_17s_17ns_17_2_1_U10.top_sub_17s_17ns_17_2_1_Adder_7_U.s ;
assign \sub_17s_17ns_17_2_1_U10.ce  = 1'h1;
assign \sub_17s_17ns_17_2_1_U10.clk  = ap_clk;
assign \sub_17s_17ns_17_2_1_U10.din0  = { op_4[15], op_4 };
assign \sub_17s_17ns_17_2_1_U10.din1  = { 7'h00, op_1, 6'h00 };
assign grp_fu_501_p2 = \sub_17s_17ns_17_2_1_U10.dout ;
assign \sub_17s_17ns_17_2_1_U10.reset  = ap_rst;
assign \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_1_U.ain_s0  = \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_1_U.a ;
assign \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_1_U.bin_s0  = \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_1_U.b ;
assign \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_1_U.s  = { \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_1_U.fas_s2 , \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_1_U.sum_s1  };
assign \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_1_U.u2.a  = \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_1_U.ain_s1 ;
assign \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_1_U.u2.b  = \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_1_U.bin_s1 ;
assign \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_1_U.u2.cin  = \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_1_U.carry_s1 ;
assign \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_1_U.facout_s2  = \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_1_U.u2.cout ;
assign \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_1_U.fas_s2  = \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_1_U.u2.s ;
assign \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_1_U.u1.a  = \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_1_U.a [3:0];
assign \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_1_U.u1.b  = \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_1_U.b [3:0];
assign \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_1_U.u1.cin  = 1'h0;
assign \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_1_U.facout_s1  = \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_1_U.u1.cout ;
assign \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_1_U.fas_s1  = \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_1_U.u1.s ;
assign \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_1_U.a  = \add_9s_9s_9_2_1_U2.din0 ;
assign \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_1_U.b  = \add_9s_9s_9_2_1_U2.din1 ;
assign \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_1_U.ce  = \add_9s_9s_9_2_1_U2.ce ;
assign \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_1_U.clk  = \add_9s_9s_9_2_1_U2.clk ;
assign \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_1_U.reset  = \add_9s_9s_9_2_1_U2.reset ;
assign \add_9s_9s_9_2_1_U2.dout  = \add_9s_9s_9_2_1_U2.top_add_9s_9s_9_2_1_Adder_1_U.s ;
assign \add_9s_9s_9_2_1_U2.ce  = 1'h1;
assign \add_9s_9s_9_2_1_U2.clk  = ap_clk;
assign \add_9s_9s_9_2_1_U2.din0  = { ret_reg_986[4], ret_reg_986, 3'h0 };
assign \add_9s_9s_9_2_1_U2.din1  = { op_5[7], op_5 };
assign grp_fu_283_p2 = \add_9s_9s_9_2_1_U2.dout ;
assign \add_9s_9s_9_2_1_U2.reset  = ap_rst;
assign \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_1_U.ain_s0  = \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_1_U.a ;
assign \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_1_U.bin_s0  = \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_1_U.b ;
assign \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_1_U.s  = { \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_1_U.fas_s2 , \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_1_U.sum_s1  };
assign \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_1_U.u2.a  = \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_1_U.ain_s1 ;
assign \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_1_U.u2.b  = \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_1_U.bin_s1 ;
assign \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_1_U.u2.cin  = \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_1_U.carry_s1 ;
assign \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_1_U.facout_s2  = \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_1_U.u2.cout ;
assign \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_1_U.fas_s2  = \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_1_U.u2.s ;
assign \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_1_U.u1.a  = \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_1_U.a [3:0];
assign \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_1_U.u1.b  = \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_1_U.b [3:0];
assign \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_1_U.u1.cin  = 1'h0;
assign \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_1_U.facout_s1  = \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_1_U.u1.cout ;
assign \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_1_U.fas_s1  = \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_1_U.u1.s ;
assign \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_1_U.a  = \add_9s_9s_9_2_1_U14.din0 ;
assign \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_1_U.b  = \add_9s_9s_9_2_1_U14.din1 ;
assign \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_1_U.ce  = \add_9s_9s_9_2_1_U14.ce ;
assign \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_1_U.clk  = \add_9s_9s_9_2_1_U14.clk ;
assign \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_1_U.reset  = \add_9s_9s_9_2_1_U14.reset ;
assign \add_9s_9s_9_2_1_U14.dout  = \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_1_U.s ;
assign \add_9s_9s_9_2_1_U14.ce  = 1'h1;
assign \add_9s_9s_9_2_1_U14.clk  = ap_clk;
assign \add_9s_9s_9_2_1_U14.din0  = { op_14[1], op_14[1], op_14, 5'h00 };
assign \add_9s_9s_9_2_1_U14.din1  = { op_11_V_reg_1194[7], op_11_V_reg_1194 };
assign grp_fu_639_p2 = \add_9s_9s_9_2_1_U14.dout ;
assign \add_9s_9s_9_2_1_U14.reset  = ap_rst;
assign \add_8s_8s_8_2_1_U15.top_add_8s_8s_8_2_1_Adder_9_U.ain_s0  = \add_8s_8s_8_2_1_U15.top_add_8s_8s_8_2_1_Adder_9_U.a ;
assign \add_8s_8s_8_2_1_U15.top_add_8s_8s_8_2_1_Adder_9_U.bin_s0  = \add_8s_8s_8_2_1_U15.top_add_8s_8s_8_2_1_Adder_9_U.b ;
assign \add_8s_8s_8_2_1_U15.top_add_8s_8s_8_2_1_Adder_9_U.s  = { \add_8s_8s_8_2_1_U15.top_add_8s_8s_8_2_1_Adder_9_U.fas_s2 , \add_8s_8s_8_2_1_U15.top_add_8s_8s_8_2_1_Adder_9_U.sum_s1  };
assign \add_8s_8s_8_2_1_U15.top_add_8s_8s_8_2_1_Adder_9_U.u2.a  = \add_8s_8s_8_2_1_U15.top_add_8s_8s_8_2_1_Adder_9_U.ain_s1 ;
assign \add_8s_8s_8_2_1_U15.top_add_8s_8s_8_2_1_Adder_9_U.u2.b  = \add_8s_8s_8_2_1_U15.top_add_8s_8s_8_2_1_Adder_9_U.bin_s1 ;
assign \add_8s_8s_8_2_1_U15.top_add_8s_8s_8_2_1_Adder_9_U.u2.cin  = \add_8s_8s_8_2_1_U15.top_add_8s_8s_8_2_1_Adder_9_U.carry_s1 ;
assign \add_8s_8s_8_2_1_U15.top_add_8s_8s_8_2_1_Adder_9_U.facout_s2  = \add_8s_8s_8_2_1_U15.top_add_8s_8s_8_2_1_Adder_9_U.u2.cout ;
assign \add_8s_8s_8_2_1_U15.top_add_8s_8s_8_2_1_Adder_9_U.fas_s2  = \add_8s_8s_8_2_1_U15.top_add_8s_8s_8_2_1_Adder_9_U.u2.s ;
assign \add_8s_8s_8_2_1_U15.top_add_8s_8s_8_2_1_Adder_9_U.u1.a  = \add_8s_8s_8_2_1_U15.top_add_8s_8s_8_2_1_Adder_9_U.a [3:0];
assign \add_8s_8s_8_2_1_U15.top_add_8s_8s_8_2_1_Adder_9_U.u1.b  = \add_8s_8s_8_2_1_U15.top_add_8s_8s_8_2_1_Adder_9_U.b [3:0];
assign \add_8s_8s_8_2_1_U15.top_add_8s_8s_8_2_1_Adder_9_U.u1.cin  = 1'h0;
assign \add_8s_8s_8_2_1_U15.top_add_8s_8s_8_2_1_Adder_9_U.facout_s1  = \add_8s_8s_8_2_1_U15.top_add_8s_8s_8_2_1_Adder_9_U.u1.cout ;
assign \add_8s_8s_8_2_1_U15.top_add_8s_8s_8_2_1_Adder_9_U.fas_s1  = \add_8s_8s_8_2_1_U15.top_add_8s_8s_8_2_1_Adder_9_U.u1.s ;
assign \add_8s_8s_8_2_1_U15.top_add_8s_8s_8_2_1_Adder_9_U.a  = \add_8s_8s_8_2_1_U15.din0 ;
assign \add_8s_8s_8_2_1_U15.top_add_8s_8s_8_2_1_Adder_9_U.b  = \add_8s_8s_8_2_1_U15.din1 ;
assign \add_8s_8s_8_2_1_U15.top_add_8s_8s_8_2_1_Adder_9_U.ce  = \add_8s_8s_8_2_1_U15.ce ;
assign \add_8s_8s_8_2_1_U15.top_add_8s_8s_8_2_1_Adder_9_U.clk  = \add_8s_8s_8_2_1_U15.clk ;
assign \add_8s_8s_8_2_1_U15.top_add_8s_8s_8_2_1_Adder_9_U.reset  = \add_8s_8s_8_2_1_U15.reset ;
assign \add_8s_8s_8_2_1_U15.dout  = \add_8s_8s_8_2_1_U15.top_add_8s_8s_8_2_1_Adder_9_U.s ;
assign \add_8s_8s_8_2_1_U15.ce  = 1'h1;
assign \add_8s_8s_8_2_1_U15.clk  = ap_clk;
assign \add_8s_8s_8_2_1_U15.din0  = { op_14[1], op_14, 5'h00 };
assign \add_8s_8s_8_2_1_U15.din1  = op_11_V_reg_1194;
assign grp_fu_645_p2 = \add_8s_8s_8_2_1_U15.dout ;
assign \add_8s_8s_8_2_1_U15.reset  = ap_rst;
assign \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_8_U.ain_s0  = \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_8_U.a ;
assign \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_8_U.bin_s0  = \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_8_U.b ;
assign \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_8_U.s  = { \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_8_U.fas_s2 , \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_8_U.sum_s1  };
assign \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_8_U.u2.a  = \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_8_U.ain_s1 ;
assign \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_8_U.u2.b  = \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_8_U.bin_s1 ;
assign \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_8_U.u2.cin  = \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_8_U.carry_s1 ;
assign \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_8_U.facout_s2  = \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_8_U.u2.cout ;
assign \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_8_U.fas_s2  = \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_8_U.u2.s ;
assign \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_8_U.u1.a  = \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_8_U.a [3:0];
assign \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_8_U.u1.b  = \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_8_U.b [3:0];
assign \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_8_U.u1.cin  = 1'h0;
assign \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_8_U.facout_s1  = \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_8_U.u1.cout ;
assign \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_8_U.fas_s1  = \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_8_U.u1.s ;
assign \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_8_U.a  = \add_8ns_8ns_8_2_1_U13.din0 ;
assign \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_8_U.b  = \add_8ns_8ns_8_2_1_U13.din1 ;
assign \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_8_U.ce  = \add_8ns_8ns_8_2_1_U13.ce ;
assign \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_8_U.clk  = \add_8ns_8ns_8_2_1_U13.clk ;
assign \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_8_U.reset  = \add_8ns_8ns_8_2_1_U13.reset ;
assign \add_8ns_8ns_8_2_1_U13.dout  = \add_8ns_8ns_8_2_1_U13.top_add_8ns_8ns_8_2_1_Adder_8_U.s ;
assign \add_8ns_8ns_8_2_1_U13.ce  = 1'h1;
assign \add_8ns_8ns_8_2_1_U13.clk  = ap_clk;
assign \add_8ns_8ns_8_2_1_U13.din0  = trunc_ln_reg_1152;
assign \add_8ns_8ns_8_2_1_U13.din1  = { 7'h00, icmp_ln410_reg_1179 };
assign grp_fu_592_p2 = \add_8ns_8ns_8_2_1_U13.dout ;
assign \add_8ns_8ns_8_2_1_U13.reset  = ap_rst;
assign \add_7s_7ns_7_2_1_U3.top_add_7s_7ns_7_2_1_Adder_2_U.ain_s0  = \add_7s_7ns_7_2_1_U3.top_add_7s_7ns_7_2_1_Adder_2_U.a ;
assign \add_7s_7ns_7_2_1_U3.top_add_7s_7ns_7_2_1_Adder_2_U.bin_s0  = \add_7s_7ns_7_2_1_U3.top_add_7s_7ns_7_2_1_Adder_2_U.b ;
assign \add_7s_7ns_7_2_1_U3.top_add_7s_7ns_7_2_1_Adder_2_U.s  = { \add_7s_7ns_7_2_1_U3.top_add_7s_7ns_7_2_1_Adder_2_U.fas_s2 , \add_7s_7ns_7_2_1_U3.top_add_7s_7ns_7_2_1_Adder_2_U.sum_s1  };
assign \add_7s_7ns_7_2_1_U3.top_add_7s_7ns_7_2_1_Adder_2_U.u2.a  = \add_7s_7ns_7_2_1_U3.top_add_7s_7ns_7_2_1_Adder_2_U.ain_s1 ;
assign \add_7s_7ns_7_2_1_U3.top_add_7s_7ns_7_2_1_Adder_2_U.u2.b  = \add_7s_7ns_7_2_1_U3.top_add_7s_7ns_7_2_1_Adder_2_U.bin_s1 ;
assign \add_7s_7ns_7_2_1_U3.top_add_7s_7ns_7_2_1_Adder_2_U.u2.cin  = \add_7s_7ns_7_2_1_U3.top_add_7s_7ns_7_2_1_Adder_2_U.carry_s1 ;
assign \add_7s_7ns_7_2_1_U3.top_add_7s_7ns_7_2_1_Adder_2_U.facout_s2  = \add_7s_7ns_7_2_1_U3.top_add_7s_7ns_7_2_1_Adder_2_U.u2.cout ;
assign \add_7s_7ns_7_2_1_U3.top_add_7s_7ns_7_2_1_Adder_2_U.fas_s2  = \add_7s_7ns_7_2_1_U3.top_add_7s_7ns_7_2_1_Adder_2_U.u2.s ;
assign \add_7s_7ns_7_2_1_U3.top_add_7s_7ns_7_2_1_Adder_2_U.u1.a  = \add_7s_7ns_7_2_1_U3.top_add_7s_7ns_7_2_1_Adder_2_U.a [2:0];
assign \add_7s_7ns_7_2_1_U3.top_add_7s_7ns_7_2_1_Adder_2_U.u1.b  = \add_7s_7ns_7_2_1_U3.top_add_7s_7ns_7_2_1_Adder_2_U.b [2:0];
assign \add_7s_7ns_7_2_1_U3.top_add_7s_7ns_7_2_1_Adder_2_U.u1.cin  = 1'h0;
assign \add_7s_7ns_7_2_1_U3.top_add_7s_7ns_7_2_1_Adder_2_U.facout_s1  = \add_7s_7ns_7_2_1_U3.top_add_7s_7ns_7_2_1_Adder_2_U.u1.cout ;
assign \add_7s_7ns_7_2_1_U3.top_add_7s_7ns_7_2_1_Adder_2_U.fas_s1  = \add_7s_7ns_7_2_1_U3.top_add_7s_7ns_7_2_1_Adder_2_U.u1.s ;
assign \add_7s_7ns_7_2_1_U3.top_add_7s_7ns_7_2_1_Adder_2_U.a  = \add_7s_7ns_7_2_1_U3.din0 ;
assign \add_7s_7ns_7_2_1_U3.top_add_7s_7ns_7_2_1_Adder_2_U.b  = \add_7s_7ns_7_2_1_U3.din1 ;
assign \add_7s_7ns_7_2_1_U3.top_add_7s_7ns_7_2_1_Adder_2_U.ce  = \add_7s_7ns_7_2_1_U3.ce ;
assign \add_7s_7ns_7_2_1_U3.top_add_7s_7ns_7_2_1_Adder_2_U.clk  = \add_7s_7ns_7_2_1_U3.clk ;
assign \add_7s_7ns_7_2_1_U3.top_add_7s_7ns_7_2_1_Adder_2_U.reset  = \add_7s_7ns_7_2_1_U3.reset ;
assign \add_7s_7ns_7_2_1_U3.dout  = \add_7s_7ns_7_2_1_U3.top_add_7s_7ns_7_2_1_Adder_2_U.s ;
assign \add_7s_7ns_7_2_1_U3.ce  = 1'h1;
assign \add_7s_7ns_7_2_1_U3.clk  = ap_clk;
assign \add_7s_7ns_7_2_1_U3.din0  = { tmp_1_reg_1011[5], tmp_1_reg_1011 };
assign \add_7s_7ns_7_2_1_U3.din1  = 7'h01;
assign grp_fu_312_p2 = \add_7s_7ns_7_2_1_U3.dout ;
assign \add_7s_7ns_7_2_1_U3.reset  = ap_rst;
assign \add_5s_5ns_5_2_1_U1.top_add_5s_5ns_5_2_1_Adder_0_U.ain_s0  = \add_5s_5ns_5_2_1_U1.top_add_5s_5ns_5_2_1_Adder_0_U.a ;
assign \add_5s_5ns_5_2_1_U1.top_add_5s_5ns_5_2_1_Adder_0_U.bin_s0  = \add_5s_5ns_5_2_1_U1.top_add_5s_5ns_5_2_1_Adder_0_U.b ;
assign \add_5s_5ns_5_2_1_U1.top_add_5s_5ns_5_2_1_Adder_0_U.s  = { \add_5s_5ns_5_2_1_U1.top_add_5s_5ns_5_2_1_Adder_0_U.fas_s2 , \add_5s_5ns_5_2_1_U1.top_add_5s_5ns_5_2_1_Adder_0_U.sum_s1  };
assign \add_5s_5ns_5_2_1_U1.top_add_5s_5ns_5_2_1_Adder_0_U.u2.a  = \add_5s_5ns_5_2_1_U1.top_add_5s_5ns_5_2_1_Adder_0_U.ain_s1 ;
assign \add_5s_5ns_5_2_1_U1.top_add_5s_5ns_5_2_1_Adder_0_U.u2.b  = \add_5s_5ns_5_2_1_U1.top_add_5s_5ns_5_2_1_Adder_0_U.bin_s1 ;
assign \add_5s_5ns_5_2_1_U1.top_add_5s_5ns_5_2_1_Adder_0_U.u2.cin  = \add_5s_5ns_5_2_1_U1.top_add_5s_5ns_5_2_1_Adder_0_U.carry_s1 ;
assign \add_5s_5ns_5_2_1_U1.top_add_5s_5ns_5_2_1_Adder_0_U.facout_s2  = \add_5s_5ns_5_2_1_U1.top_add_5s_5ns_5_2_1_Adder_0_U.u2.cout ;
assign \add_5s_5ns_5_2_1_U1.top_add_5s_5ns_5_2_1_Adder_0_U.fas_s2  = \add_5s_5ns_5_2_1_U1.top_add_5s_5ns_5_2_1_Adder_0_U.u2.s ;
assign \add_5s_5ns_5_2_1_U1.top_add_5s_5ns_5_2_1_Adder_0_U.u1.a  = \add_5s_5ns_5_2_1_U1.top_add_5s_5ns_5_2_1_Adder_0_U.a [1:0];
assign \add_5s_5ns_5_2_1_U1.top_add_5s_5ns_5_2_1_Adder_0_U.u1.b  = \add_5s_5ns_5_2_1_U1.top_add_5s_5ns_5_2_1_Adder_0_U.b [1:0];
assign \add_5s_5ns_5_2_1_U1.top_add_5s_5ns_5_2_1_Adder_0_U.u1.cin  = 1'h0;
assign \add_5s_5ns_5_2_1_U1.top_add_5s_5ns_5_2_1_Adder_0_U.facout_s1  = \add_5s_5ns_5_2_1_U1.top_add_5s_5ns_5_2_1_Adder_0_U.u1.cout ;
assign \add_5s_5ns_5_2_1_U1.top_add_5s_5ns_5_2_1_Adder_0_U.fas_s1  = \add_5s_5ns_5_2_1_U1.top_add_5s_5ns_5_2_1_Adder_0_U.u1.s ;
assign \add_5s_5ns_5_2_1_U1.top_add_5s_5ns_5_2_1_Adder_0_U.a  = \add_5s_5ns_5_2_1_U1.din0 ;
assign \add_5s_5ns_5_2_1_U1.top_add_5s_5ns_5_2_1_Adder_0_U.b  = \add_5s_5ns_5_2_1_U1.din1 ;
assign \add_5s_5ns_5_2_1_U1.top_add_5s_5ns_5_2_1_Adder_0_U.ce  = \add_5s_5ns_5_2_1_U1.ce ;
assign \add_5s_5ns_5_2_1_U1.top_add_5s_5ns_5_2_1_Adder_0_U.clk  = \add_5s_5ns_5_2_1_U1.clk ;
assign \add_5s_5ns_5_2_1_U1.top_add_5s_5ns_5_2_1_Adder_0_U.reset  = \add_5s_5ns_5_2_1_U1.reset ;
assign \add_5s_5ns_5_2_1_U1.dout  = \add_5s_5ns_5_2_1_U1.top_add_5s_5ns_5_2_1_Adder_0_U.s ;
assign \add_5s_5ns_5_2_1_U1.ce  = 1'h1;
assign \add_5s_5ns_5_2_1_U1.clk  = ap_clk;
assign \add_5s_5ns_5_2_1_U1.din0  = { op_2[3], op_2 };
assign \add_5s_5ns_5_2_1_U1.din1  = select_ln215_reg_976;
assign grp_fu_263_p2 = \add_5s_5ns_5_2_1_U1.dout ;
assign \add_5s_5ns_5_2_1_U1.reset  = ap_rst;
assign \add_4ns_4ns_4_2_1_U19.top_add_4ns_4ns_4_2_1_Adder_12_U.ain_s0  = \add_4ns_4ns_4_2_1_U19.top_add_4ns_4ns_4_2_1_Adder_12_U.a ;
assign \add_4ns_4ns_4_2_1_U19.top_add_4ns_4ns_4_2_1_Adder_12_U.bin_s0  = \add_4ns_4ns_4_2_1_U19.top_add_4ns_4ns_4_2_1_Adder_12_U.b ;
assign \add_4ns_4ns_4_2_1_U19.top_add_4ns_4ns_4_2_1_Adder_12_U.s  = { \add_4ns_4ns_4_2_1_U19.top_add_4ns_4ns_4_2_1_Adder_12_U.fas_s2 , \add_4ns_4ns_4_2_1_U19.top_add_4ns_4ns_4_2_1_Adder_12_U.sum_s1  };
assign \add_4ns_4ns_4_2_1_U19.top_add_4ns_4ns_4_2_1_Adder_12_U.u2.a  = \add_4ns_4ns_4_2_1_U19.top_add_4ns_4ns_4_2_1_Adder_12_U.ain_s1 ;
assign \add_4ns_4ns_4_2_1_U19.top_add_4ns_4ns_4_2_1_Adder_12_U.u2.b  = \add_4ns_4ns_4_2_1_U19.top_add_4ns_4ns_4_2_1_Adder_12_U.bin_s1 ;
assign \add_4ns_4ns_4_2_1_U19.top_add_4ns_4ns_4_2_1_Adder_12_U.u2.cin  = \add_4ns_4ns_4_2_1_U19.top_add_4ns_4ns_4_2_1_Adder_12_U.carry_s1 ;
assign \add_4ns_4ns_4_2_1_U19.top_add_4ns_4ns_4_2_1_Adder_12_U.facout_s2  = \add_4ns_4ns_4_2_1_U19.top_add_4ns_4ns_4_2_1_Adder_12_U.u2.cout ;
assign \add_4ns_4ns_4_2_1_U19.top_add_4ns_4ns_4_2_1_Adder_12_U.fas_s2  = \add_4ns_4ns_4_2_1_U19.top_add_4ns_4ns_4_2_1_Adder_12_U.u2.s ;
assign \add_4ns_4ns_4_2_1_U19.top_add_4ns_4ns_4_2_1_Adder_12_U.u1.a  = \add_4ns_4ns_4_2_1_U19.top_add_4ns_4ns_4_2_1_Adder_12_U.a [1:0];
assign \add_4ns_4ns_4_2_1_U19.top_add_4ns_4ns_4_2_1_Adder_12_U.u1.b  = \add_4ns_4ns_4_2_1_U19.top_add_4ns_4ns_4_2_1_Adder_12_U.b [1:0];
assign \add_4ns_4ns_4_2_1_U19.top_add_4ns_4ns_4_2_1_Adder_12_U.u1.cin  = 1'h0;
assign \add_4ns_4ns_4_2_1_U19.top_add_4ns_4ns_4_2_1_Adder_12_U.facout_s1  = \add_4ns_4ns_4_2_1_U19.top_add_4ns_4ns_4_2_1_Adder_12_U.u1.cout ;
assign \add_4ns_4ns_4_2_1_U19.top_add_4ns_4ns_4_2_1_Adder_12_U.fas_s1  = \add_4ns_4ns_4_2_1_U19.top_add_4ns_4ns_4_2_1_Adder_12_U.u1.s ;
assign \add_4ns_4ns_4_2_1_U19.top_add_4ns_4ns_4_2_1_Adder_12_U.a  = \add_4ns_4ns_4_2_1_U19.din0 ;
assign \add_4ns_4ns_4_2_1_U19.top_add_4ns_4ns_4_2_1_Adder_12_U.b  = \add_4ns_4ns_4_2_1_U19.din1 ;
assign \add_4ns_4ns_4_2_1_U19.top_add_4ns_4ns_4_2_1_Adder_12_U.ce  = \add_4ns_4ns_4_2_1_U19.ce ;
assign \add_4ns_4ns_4_2_1_U19.top_add_4ns_4ns_4_2_1_Adder_12_U.clk  = \add_4ns_4ns_4_2_1_U19.clk ;
assign \add_4ns_4ns_4_2_1_U19.top_add_4ns_4ns_4_2_1_Adder_12_U.reset  = \add_4ns_4ns_4_2_1_U19.reset ;
assign \add_4ns_4ns_4_2_1_U19.dout  = \add_4ns_4ns_4_2_1_U19.top_add_4ns_4ns_4_2_1_Adder_12_U.s ;
assign \add_4ns_4ns_4_2_1_U19.ce  = 1'h1;
assign \add_4ns_4ns_4_2_1_U19.clk  = ap_clk;
assign \add_4ns_4ns_4_2_1_U19.din0  = p_Val2_4_reg_1260;
assign \add_4ns_4ns_4_2_1_U19.din1  = { 3'h0, and_ln412_reg_1281 };
assign grp_fu_740_p2 = \add_4ns_4ns_4_2_1_U19.dout ;
assign \add_4ns_4ns_4_2_1_U19.reset  = ap_rst;
assign \add_44s_44s_44_2_1_U4.top_add_44s_44s_44_2_1_Adder_3_U.ain_s0  = \add_44s_44s_44_2_1_U4.top_add_44s_44s_44_2_1_Adder_3_U.a ;
assign \add_44s_44s_44_2_1_U4.top_add_44s_44s_44_2_1_Adder_3_U.bin_s0  = \add_44s_44s_44_2_1_U4.top_add_44s_44s_44_2_1_Adder_3_U.b ;
assign \add_44s_44s_44_2_1_U4.top_add_44s_44s_44_2_1_Adder_3_U.s  = { \add_44s_44s_44_2_1_U4.top_add_44s_44s_44_2_1_Adder_3_U.fas_s2 , \add_44s_44s_44_2_1_U4.top_add_44s_44s_44_2_1_Adder_3_U.sum_s1  };
assign \add_44s_44s_44_2_1_U4.top_add_44s_44s_44_2_1_Adder_3_U.u2.a  = \add_44s_44s_44_2_1_U4.top_add_44s_44s_44_2_1_Adder_3_U.ain_s1 ;
assign \add_44s_44s_44_2_1_U4.top_add_44s_44s_44_2_1_Adder_3_U.u2.b  = \add_44s_44s_44_2_1_U4.top_add_44s_44s_44_2_1_Adder_3_U.bin_s1 ;
assign \add_44s_44s_44_2_1_U4.top_add_44s_44s_44_2_1_Adder_3_U.u2.cin  = \add_44s_44s_44_2_1_U4.top_add_44s_44s_44_2_1_Adder_3_U.carry_s1 ;
assign \add_44s_44s_44_2_1_U4.top_add_44s_44s_44_2_1_Adder_3_U.facout_s2  = \add_44s_44s_44_2_1_U4.top_add_44s_44s_44_2_1_Adder_3_U.u2.cout ;
assign \add_44s_44s_44_2_1_U4.top_add_44s_44s_44_2_1_Adder_3_U.fas_s2  = \add_44s_44s_44_2_1_U4.top_add_44s_44s_44_2_1_Adder_3_U.u2.s ;
assign \add_44s_44s_44_2_1_U4.top_add_44s_44s_44_2_1_Adder_3_U.u1.a  = \add_44s_44s_44_2_1_U4.top_add_44s_44s_44_2_1_Adder_3_U.a [21:0];
assign \add_44s_44s_44_2_1_U4.top_add_44s_44s_44_2_1_Adder_3_U.u1.b  = \add_44s_44s_44_2_1_U4.top_add_44s_44s_44_2_1_Adder_3_U.b [21:0];
assign \add_44s_44s_44_2_1_U4.top_add_44s_44s_44_2_1_Adder_3_U.u1.cin  = 1'h0;
assign \add_44s_44s_44_2_1_U4.top_add_44s_44s_44_2_1_Adder_3_U.facout_s1  = \add_44s_44s_44_2_1_U4.top_add_44s_44s_44_2_1_Adder_3_U.u1.cout ;
assign \add_44s_44s_44_2_1_U4.top_add_44s_44s_44_2_1_Adder_3_U.fas_s1  = \add_44s_44s_44_2_1_U4.top_add_44s_44s_44_2_1_Adder_3_U.u1.s ;
assign \add_44s_44s_44_2_1_U4.top_add_44s_44s_44_2_1_Adder_3_U.a  = \add_44s_44s_44_2_1_U4.din0 ;
assign \add_44s_44s_44_2_1_U4.top_add_44s_44s_44_2_1_Adder_3_U.b  = \add_44s_44s_44_2_1_U4.din1 ;
assign \add_44s_44s_44_2_1_U4.top_add_44s_44s_44_2_1_Adder_3_U.ce  = \add_44s_44s_44_2_1_U4.ce ;
assign \add_44s_44s_44_2_1_U4.top_add_44s_44s_44_2_1_Adder_3_U.clk  = \add_44s_44s_44_2_1_U4.clk ;
assign \add_44s_44s_44_2_1_U4.top_add_44s_44s_44_2_1_Adder_3_U.reset  = \add_44s_44s_44_2_1_U4.reset ;
assign \add_44s_44s_44_2_1_U4.dout  = \add_44s_44s_44_2_1_U4.top_add_44s_44s_44_2_1_Adder_3_U.s ;
assign \add_44s_44s_44_2_1_U4.ce  = 1'h1;
assign \add_44s_44s_44_2_1_U4.clk  = ap_clk;
assign \add_44s_44s_44_2_1_U4.din0  = { select_ln353_reg_1028[6], select_ln353_reg_1028[6], select_ln353_reg_1028[6], select_ln353_reg_1028[6], select_ln353_reg_1028[6], select_ln353_reg_1028[6], select_ln353_reg_1028[6], select_ln353_reg_1028[6], select_ln353_reg_1028[6], select_ln353_reg_1028[6], select_ln353_reg_1028[6], select_ln353_reg_1028[6], select_ln353_reg_1028[6], select_ln353_reg_1028[6], select_ln353_reg_1028[6], select_ln353_reg_1028[6], select_ln353_reg_1028[6], select_ln353_reg_1028[6], select_ln353_reg_1028[6], select_ln353_reg_1028[6], select_ln353_reg_1028[6], select_ln353_reg_1028[6], select_ln353_reg_1028[6], select_ln353_reg_1028[6], select_ln353_reg_1028[6], select_ln353_reg_1028[6], select_ln353_reg_1028, 11'h000 };
assign \add_44s_44s_44_2_1_U4.din1  = { op_6[15], op_6[15], op_6[15], op_6[15], op_6[15], op_6[15], op_6[15], op_6[15], op_6[15], op_6[15], op_6[15], op_6[15], op_6[15], op_6[15], op_6[15], op_6[15], op_6[15], op_6[15], op_6[15], op_6[15], op_6[15], op_6[15], op_6[15], op_6[15], op_6[15], op_6[15], op_6[15], op_6[15], op_6 };
assign grp_fu_352_p2 = \add_44s_44s_44_2_1_U4.dout ;
assign \add_44s_44s_44_2_1_U4.reset  = ap_rst;
assign \add_36s_36s_36_2_1_U7.top_add_36s_36s_36_2_1_Adder_6_U.ain_s0  = \add_36s_36s_36_2_1_U7.top_add_36s_36s_36_2_1_Adder_6_U.a ;
assign \add_36s_36s_36_2_1_U7.top_add_36s_36s_36_2_1_Adder_6_U.bin_s0  = \add_36s_36s_36_2_1_U7.top_add_36s_36s_36_2_1_Adder_6_U.b ;
assign \add_36s_36s_36_2_1_U7.top_add_36s_36s_36_2_1_Adder_6_U.s  = { \add_36s_36s_36_2_1_U7.top_add_36s_36s_36_2_1_Adder_6_U.fas_s2 , \add_36s_36s_36_2_1_U7.top_add_36s_36s_36_2_1_Adder_6_U.sum_s1  };
assign \add_36s_36s_36_2_1_U7.top_add_36s_36s_36_2_1_Adder_6_U.u2.a  = \add_36s_36s_36_2_1_U7.top_add_36s_36s_36_2_1_Adder_6_U.ain_s1 ;
assign \add_36s_36s_36_2_1_U7.top_add_36s_36s_36_2_1_Adder_6_U.u2.b  = \add_36s_36s_36_2_1_U7.top_add_36s_36s_36_2_1_Adder_6_U.bin_s1 ;
assign \add_36s_36s_36_2_1_U7.top_add_36s_36s_36_2_1_Adder_6_U.u2.cin  = \add_36s_36s_36_2_1_U7.top_add_36s_36s_36_2_1_Adder_6_U.carry_s1 ;
assign \add_36s_36s_36_2_1_U7.top_add_36s_36s_36_2_1_Adder_6_U.facout_s2  = \add_36s_36s_36_2_1_U7.top_add_36s_36s_36_2_1_Adder_6_U.u2.cout ;
assign \add_36s_36s_36_2_1_U7.top_add_36s_36s_36_2_1_Adder_6_U.fas_s2  = \add_36s_36s_36_2_1_U7.top_add_36s_36s_36_2_1_Adder_6_U.u2.s ;
assign \add_36s_36s_36_2_1_U7.top_add_36s_36s_36_2_1_Adder_6_U.u1.a  = \add_36s_36s_36_2_1_U7.top_add_36s_36s_36_2_1_Adder_6_U.a [17:0];
assign \add_36s_36s_36_2_1_U7.top_add_36s_36s_36_2_1_Adder_6_U.u1.b  = \add_36s_36s_36_2_1_U7.top_add_36s_36s_36_2_1_Adder_6_U.b [17:0];
assign \add_36s_36s_36_2_1_U7.top_add_36s_36s_36_2_1_Adder_6_U.u1.cin  = 1'h0;
assign \add_36s_36s_36_2_1_U7.top_add_36s_36s_36_2_1_Adder_6_U.facout_s1  = \add_36s_36s_36_2_1_U7.top_add_36s_36s_36_2_1_Adder_6_U.u1.cout ;
assign \add_36s_36s_36_2_1_U7.top_add_36s_36s_36_2_1_Adder_6_U.fas_s1  = \add_36s_36s_36_2_1_U7.top_add_36s_36s_36_2_1_Adder_6_U.u1.s ;
assign \add_36s_36s_36_2_1_U7.top_add_36s_36s_36_2_1_Adder_6_U.a  = \add_36s_36s_36_2_1_U7.din0 ;
assign \add_36s_36s_36_2_1_U7.top_add_36s_36s_36_2_1_Adder_6_U.b  = \add_36s_36s_36_2_1_U7.din1 ;
assign \add_36s_36s_36_2_1_U7.top_add_36s_36s_36_2_1_Adder_6_U.ce  = \add_36s_36s_36_2_1_U7.ce ;
assign \add_36s_36s_36_2_1_U7.top_add_36s_36s_36_2_1_Adder_6_U.clk  = \add_36s_36s_36_2_1_U7.clk ;
assign \add_36s_36s_36_2_1_U7.top_add_36s_36s_36_2_1_Adder_6_U.reset  = \add_36s_36s_36_2_1_U7.reset ;
assign \add_36s_36s_36_2_1_U7.dout  = \add_36s_36s_36_2_1_U7.top_add_36s_36s_36_2_1_Adder_6_U.s ;
assign \add_36s_36s_36_2_1_U7.ce  = 1'h1;
assign \add_36s_36s_36_2_1_U7.clk  = ap_clk;
assign \add_36s_36s_36_2_1_U7.din0  = { op_23_V_reg_1075[31], op_23_V_reg_1075, 3'h0 };
assign \add_36s_36s_36_2_1_U7.din1  = { op_9[3], op_9[3], op_9[3], op_9[3], op_9[3], op_9[3], op_9[3], op_9[3], op_9[3], op_9[3], op_9[3], op_9[3], op_9[3], op_9[3], op_9[3], op_9[3], op_9[3], op_9[3], op_9[3], op_9[3], op_9[3], op_9[3], op_9[3], op_9[3], op_9[3], op_9[3], op_9[3], op_9[3], op_9[3], op_9[3], op_9[3], op_9[3], op_9 };
assign grp_fu_426_p2 = \add_36s_36s_36_2_1_U7.dout ;
assign \add_36s_36s_36_2_1_U7.reset  = ap_rst;
assign \add_36s_36s_36_2_1_U11.top_add_36s_36s_36_2_1_Adder_6_U.ain_s0  = \add_36s_36s_36_2_1_U11.top_add_36s_36s_36_2_1_Adder_6_U.a ;
assign \add_36s_36s_36_2_1_U11.top_add_36s_36s_36_2_1_Adder_6_U.bin_s0  = \add_36s_36s_36_2_1_U11.top_add_36s_36s_36_2_1_Adder_6_U.b ;
assign \add_36s_36s_36_2_1_U11.top_add_36s_36s_36_2_1_Adder_6_U.s  = { \add_36s_36s_36_2_1_U11.top_add_36s_36s_36_2_1_Adder_6_U.fas_s2 , \add_36s_36s_36_2_1_U11.top_add_36s_36s_36_2_1_Adder_6_U.sum_s1  };
assign \add_36s_36s_36_2_1_U11.top_add_36s_36s_36_2_1_Adder_6_U.u2.a  = \add_36s_36s_36_2_1_U11.top_add_36s_36s_36_2_1_Adder_6_U.ain_s1 ;
assign \add_36s_36s_36_2_1_U11.top_add_36s_36s_36_2_1_Adder_6_U.u2.b  = \add_36s_36s_36_2_1_U11.top_add_36s_36s_36_2_1_Adder_6_U.bin_s1 ;
assign \add_36s_36s_36_2_1_U11.top_add_36s_36s_36_2_1_Adder_6_U.u2.cin  = \add_36s_36s_36_2_1_U11.top_add_36s_36s_36_2_1_Adder_6_U.carry_s1 ;
assign \add_36s_36s_36_2_1_U11.top_add_36s_36s_36_2_1_Adder_6_U.facout_s2  = \add_36s_36s_36_2_1_U11.top_add_36s_36s_36_2_1_Adder_6_U.u2.cout ;
assign \add_36s_36s_36_2_1_U11.top_add_36s_36s_36_2_1_Adder_6_U.fas_s2  = \add_36s_36s_36_2_1_U11.top_add_36s_36s_36_2_1_Adder_6_U.u2.s ;
assign \add_36s_36s_36_2_1_U11.top_add_36s_36s_36_2_1_Adder_6_U.u1.a  = \add_36s_36s_36_2_1_U11.top_add_36s_36s_36_2_1_Adder_6_U.a [17:0];
assign \add_36s_36s_36_2_1_U11.top_add_36s_36s_36_2_1_Adder_6_U.u1.b  = \add_36s_36s_36_2_1_U11.top_add_36s_36s_36_2_1_Adder_6_U.b [17:0];
assign \add_36s_36s_36_2_1_U11.top_add_36s_36s_36_2_1_Adder_6_U.u1.cin  = 1'h0;
assign \add_36s_36s_36_2_1_U11.top_add_36s_36s_36_2_1_Adder_6_U.facout_s1  = \add_36s_36s_36_2_1_U11.top_add_36s_36s_36_2_1_Adder_6_U.u1.cout ;
assign \add_36s_36s_36_2_1_U11.top_add_36s_36s_36_2_1_Adder_6_U.fas_s1  = \add_36s_36s_36_2_1_U11.top_add_36s_36s_36_2_1_Adder_6_U.u1.s ;
assign \add_36s_36s_36_2_1_U11.top_add_36s_36s_36_2_1_Adder_6_U.a  = \add_36s_36s_36_2_1_U11.din0 ;
assign \add_36s_36s_36_2_1_U11.top_add_36s_36s_36_2_1_Adder_6_U.b  = \add_36s_36s_36_2_1_U11.din1 ;
assign \add_36s_36s_36_2_1_U11.top_add_36s_36s_36_2_1_Adder_6_U.ce  = \add_36s_36s_36_2_1_U11.ce ;
assign \add_36s_36s_36_2_1_U11.top_add_36s_36s_36_2_1_Adder_6_U.clk  = \add_36s_36s_36_2_1_U11.clk ;
assign \add_36s_36s_36_2_1_U11.top_add_36s_36s_36_2_1_Adder_6_U.reset  = \add_36s_36s_36_2_1_U11.reset ;
assign \add_36s_36s_36_2_1_U11.dout  = \add_36s_36s_36_2_1_U11.top_add_36s_36s_36_2_1_Adder_6_U.s ;
assign \add_36s_36s_36_2_1_U11.ce  = 1'h1;
assign \add_36s_36s_36_2_1_U11.clk  = ap_clk;
assign \add_36s_36s_36_2_1_U11.din0  = { op_25_V_reg_1122[31], op_25_V_reg_1122, 3'h0 };
assign \add_36s_36s_36_2_1_U11.din1  = { op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12 };
assign grp_fu_522_p2 = \add_36s_36s_36_2_1_U11.dout ;
assign \add_36s_36s_36_2_1_U11.reset  = ap_rst;
assign \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_13_U.ain_s0  = \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_13_U.a ;
assign \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_13_U.bin_s0  = \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_13_U.b ;
assign \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_13_U.s  = { \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_13_U.fas_s2 , \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_13_U.sum_s1  };
assign \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_13_U.u2.a  = \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_13_U.ain_s1 ;
assign \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_13_U.u2.b  = \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_13_U.bin_s1 ;
assign \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_13_U.u2.cin  = \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_13_U.carry_s1 ;
assign \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_13_U.facout_s2  = \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_13_U.u2.cout ;
assign \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_13_U.fas_s2  = \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_13_U.u2.s ;
assign \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_13_U.u1.a  = \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_13_U.a [16:0];
assign \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_13_U.u1.b  = \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_13_U.b [16:0];
assign \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_13_U.u1.cin  = 1'h0;
assign \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_13_U.facout_s1  = \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_13_U.u1.cout ;
assign \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_13_U.fas_s1  = \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_13_U.u1.s ;
assign \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_13_U.a  = \add_34s_34s_34_2_1_U23.din0 ;
assign \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_13_U.b  = \add_34s_34s_34_2_1_U23.din1 ;
assign \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_13_U.ce  = \add_34s_34s_34_2_1_U23.ce ;
assign \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_13_U.clk  = \add_34s_34s_34_2_1_U23.clk ;
assign \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_13_U.reset  = \add_34s_34s_34_2_1_U23.reset ;
assign \add_34s_34s_34_2_1_U23.dout  = \add_34s_34s_34_2_1_U23.top_add_34s_34s_34_2_1_Adder_13_U.s ;
assign \add_34s_34s_34_2_1_U23.ce  = 1'h1;
assign \add_34s_34s_34_2_1_U23.clk  = ap_clk;
assign \add_34s_34s_34_2_1_U23.din0  = { ret_V_27_reg_1404[31], ret_V_27_reg_1404, 1'h0 };
assign \add_34s_34s_34_2_1_U23.din1  = { op_19_V_reg_1398[3], op_19_V_reg_1398[3], op_19_V_reg_1398[3], op_19_V_reg_1398[3], op_19_V_reg_1398[3], op_19_V_reg_1398[3], op_19_V_reg_1398[3], op_19_V_reg_1398[3], op_19_V_reg_1398[3], op_19_V_reg_1398[3], op_19_V_reg_1398[3], op_19_V_reg_1398[3], op_19_V_reg_1398[3], op_19_V_reg_1398[3], op_19_V_reg_1398[3], op_19_V_reg_1398[3], op_19_V_reg_1398[3], op_19_V_reg_1398[3], op_19_V_reg_1398[3], op_19_V_reg_1398[3], op_19_V_reg_1398[3], op_19_V_reg_1398[3], op_19_V_reg_1398[3], op_19_V_reg_1398[3], op_19_V_reg_1398[3], op_19_V_reg_1398[3], op_19_V_reg_1398[3], op_19_V_reg_1398[3], op_19_V_reg_1398[3], op_19_V_reg_1398[3], op_19_V_reg_1398 };
assign grp_fu_931_p2 = \add_34s_34s_34_2_1_U23.dout ;
assign \add_34s_34s_34_2_1_U23.reset  = ap_rst;
assign \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_13_U.ain_s0  = \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_13_U.a ;
assign \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_13_U.bin_s0  = \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_13_U.b ;
assign \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_13_U.s  = { \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_13_U.fas_s2 , \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_13_U.sum_s1  };
assign \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_13_U.u2.a  = \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_13_U.ain_s1 ;
assign \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_13_U.u2.b  = \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_13_U.bin_s1 ;
assign \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_13_U.u2.cin  = \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_13_U.carry_s1 ;
assign \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_13_U.facout_s2  = \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_13_U.u2.cout ;
assign \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_13_U.fas_s2  = \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_13_U.u2.s ;
assign \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_13_U.u1.a  = \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_13_U.a [16:0];
assign \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_13_U.u1.b  = \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_13_U.b [16:0];
assign \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_13_U.u1.cin  = 1'h0;
assign \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_13_U.facout_s1  = \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_13_U.u1.cout ;
assign \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_13_U.fas_s1  = \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_13_U.u1.s ;
assign \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_13_U.a  = \add_34s_34s_34_2_1_U20.din0 ;
assign \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_13_U.b  = \add_34s_34s_34_2_1_U20.din1 ;
assign \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_13_U.ce  = \add_34s_34s_34_2_1_U20.ce ;
assign \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_13_U.clk  = \add_34s_34s_34_2_1_U20.clk ;
assign \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_13_U.reset  = \add_34s_34s_34_2_1_U20.reset ;
assign \add_34s_34s_34_2_1_U20.dout  = \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_13_U.s ;
assign \add_34s_34s_34_2_1_U20.ce  = 1'h1;
assign \add_34s_34s_34_2_1_U20.clk  = ap_clk;
assign \add_34s_34s_34_2_1_U20.din0  = { op_29_V_reg_1296[31], op_29_V_reg_1296, 1'h0 };
assign \add_34s_34s_34_2_1_U20.din1  = { op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17 };
assign grp_fu_768_p2 = \add_34s_34s_34_2_1_U20.dout ;
assign \add_34s_34s_34_2_1_U20.reset  = ap_rst;
assign \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_11_U.ain_s0  = \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_11_U.a ;
assign \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_11_U.bin_s0  = \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_11_U.b ;
assign \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_11_U.s  = { \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_11_U.fas_s2 , \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_11_U.sum_s1  };
assign \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_11_U.u2.a  = \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_11_U.ain_s1 ;
assign \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_11_U.u2.b  = \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_11_U.bin_s1 ;
assign \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_11_U.u2.cin  = \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_11_U.carry_s1 ;
assign \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_11_U.facout_s2  = \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_11_U.u2.cout ;
assign \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_11_U.fas_s2  = \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_11_U.u2.s ;
assign \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_11_U.u1.a  = \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_11_U.a [15:0];
assign \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_11_U.u1.b  = \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_11_U.b [15:0];
assign \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_11_U.u1.cin  = 1'h0;
assign \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_11_U.facout_s1  = \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_11_U.u1.cout ;
assign \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_11_U.fas_s1  = \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_11_U.u1.s ;
assign \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_11_U.a  = \add_32s_32ns_32_2_1_U18.din0 ;
assign \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_11_U.b  = \add_32s_32ns_32_2_1_U18.din1 ;
assign \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_11_U.ce  = \add_32s_32ns_32_2_1_U18.ce ;
assign \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_11_U.clk  = \add_32s_32ns_32_2_1_U18.clk ;
assign \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_11_U.reset  = \add_32s_32ns_32_2_1_U18.reset ;
assign \add_32s_32ns_32_2_1_U18.dout  = \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_11_U.s ;
assign \add_32s_32ns_32_2_1_U18.ce  = 1'h1;
assign \add_32s_32ns_32_2_1_U18.clk  = ap_clk;
assign \add_32s_32ns_32_2_1_U18.din0  = { add_ln69_reg_1276[9], add_ln69_reg_1276[9], add_ln69_reg_1276[9], add_ln69_reg_1276[9], add_ln69_reg_1276[9], add_ln69_reg_1276[9], add_ln69_reg_1276[9], add_ln69_reg_1276[9], add_ln69_reg_1276[9], add_ln69_reg_1276[9], add_ln69_reg_1276[9], add_ln69_reg_1276[9], add_ln69_reg_1276[9], add_ln69_reg_1276[9], add_ln69_reg_1276[9], add_ln69_reg_1276[9], add_ln69_reg_1276[9], add_ln69_reg_1276[9], add_ln69_reg_1276[9], add_ln69_reg_1276[9], add_ln69_reg_1276[9], add_ln69_reg_1276[9], add_ln69_reg_1276 };
assign \add_32s_32ns_32_2_1_U18.din1  = ret_V_24_reg_1271;
assign grp_fu_732_p2 = \add_32s_32ns_32_2_1_U18.dout ;
assign \add_32s_32ns_32_2_1_U18.reset  = ap_rst;
assign \add_32ns_32s_32_2_1_U6.top_add_32ns_32s_32_2_1_Adder_5_U.ain_s0  = \add_32ns_32s_32_2_1_U6.top_add_32ns_32s_32_2_1_Adder_5_U.a ;
assign \add_32ns_32s_32_2_1_U6.top_add_32ns_32s_32_2_1_Adder_5_U.bin_s0  = \add_32ns_32s_32_2_1_U6.top_add_32ns_32s_32_2_1_Adder_5_U.b ;
assign \add_32ns_32s_32_2_1_U6.top_add_32ns_32s_32_2_1_Adder_5_U.s  = { \add_32ns_32s_32_2_1_U6.top_add_32ns_32s_32_2_1_Adder_5_U.fas_s2 , \add_32ns_32s_32_2_1_U6.top_add_32ns_32s_32_2_1_Adder_5_U.sum_s1  };
assign \add_32ns_32s_32_2_1_U6.top_add_32ns_32s_32_2_1_Adder_5_U.u2.a  = \add_32ns_32s_32_2_1_U6.top_add_32ns_32s_32_2_1_Adder_5_U.ain_s1 ;
assign \add_32ns_32s_32_2_1_U6.top_add_32ns_32s_32_2_1_Adder_5_U.u2.b  = \add_32ns_32s_32_2_1_U6.top_add_32ns_32s_32_2_1_Adder_5_U.bin_s1 ;
assign \add_32ns_32s_32_2_1_U6.top_add_32ns_32s_32_2_1_Adder_5_U.u2.cin  = \add_32ns_32s_32_2_1_U6.top_add_32ns_32s_32_2_1_Adder_5_U.carry_s1 ;
assign \add_32ns_32s_32_2_1_U6.top_add_32ns_32s_32_2_1_Adder_5_U.facout_s2  = \add_32ns_32s_32_2_1_U6.top_add_32ns_32s_32_2_1_Adder_5_U.u2.cout ;
assign \add_32ns_32s_32_2_1_U6.top_add_32ns_32s_32_2_1_Adder_5_U.fas_s2  = \add_32ns_32s_32_2_1_U6.top_add_32ns_32s_32_2_1_Adder_5_U.u2.s ;
assign \add_32ns_32s_32_2_1_U6.top_add_32ns_32s_32_2_1_Adder_5_U.u1.a  = \add_32ns_32s_32_2_1_U6.top_add_32ns_32s_32_2_1_Adder_5_U.a [15:0];
assign \add_32ns_32s_32_2_1_U6.top_add_32ns_32s_32_2_1_Adder_5_U.u1.b  = \add_32ns_32s_32_2_1_U6.top_add_32ns_32s_32_2_1_Adder_5_U.b [15:0];
assign \add_32ns_32s_32_2_1_U6.top_add_32ns_32s_32_2_1_Adder_5_U.u1.cin  = 1'h0;
assign \add_32ns_32s_32_2_1_U6.top_add_32ns_32s_32_2_1_Adder_5_U.facout_s1  = \add_32ns_32s_32_2_1_U6.top_add_32ns_32s_32_2_1_Adder_5_U.u1.cout ;
assign \add_32ns_32s_32_2_1_U6.top_add_32ns_32s_32_2_1_Adder_5_U.fas_s1  = \add_32ns_32s_32_2_1_U6.top_add_32ns_32s_32_2_1_Adder_5_U.u1.s ;
assign \add_32ns_32s_32_2_1_U6.top_add_32ns_32s_32_2_1_Adder_5_U.a  = \add_32ns_32s_32_2_1_U6.din0 ;
assign \add_32ns_32s_32_2_1_U6.top_add_32ns_32s_32_2_1_Adder_5_U.b  = \add_32ns_32s_32_2_1_U6.din1 ;
assign \add_32ns_32s_32_2_1_U6.top_add_32ns_32s_32_2_1_Adder_5_U.ce  = \add_32ns_32s_32_2_1_U6.ce ;
assign \add_32ns_32s_32_2_1_U6.top_add_32ns_32s_32_2_1_Adder_5_U.clk  = \add_32ns_32s_32_2_1_U6.clk ;
assign \add_32ns_32s_32_2_1_U6.top_add_32ns_32s_32_2_1_Adder_5_U.reset  = \add_32ns_32s_32_2_1_U6.reset ;
assign \add_32ns_32s_32_2_1_U6.dout  = \add_32ns_32s_32_2_1_U6.top_add_32ns_32s_32_2_1_Adder_5_U.s ;
assign \add_32ns_32s_32_2_1_U6.ce  = 1'h1;
assign \add_32ns_32s_32_2_1_U6.clk  = ap_clk;
assign \add_32ns_32s_32_2_1_U6.din0  = ret_V_18_reg_1065;
assign \add_32ns_32s_32_2_1_U6.din1  = { op_8[3], op_8[3], op_8[3], op_8[3], op_8[3], op_8[3], op_8[3], op_8[3], op_8[3], op_8[3], op_8[3], op_8[3], op_8[3], op_8[3], op_8[3], op_8[3], op_8[3], op_8[3], op_8[3], op_8[3], op_8[3], op_8[3], op_8[3], op_8[3], op_8[3], op_8[3], op_8[3], op_8[3], op_8 };
assign grp_fu_406_p2 = \add_32ns_32s_32_2_1_U6.dout ;
assign \add_32ns_32s_32_2_1_U6.reset  = ap_rst;
assign \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_5_U.ain_s0  = \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_5_U.a ;
assign \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_5_U.bin_s0  = \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_5_U.b ;
assign \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_5_U.s  = { \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_5_U.fas_s2 , \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_5_U.sum_s1  };
assign \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_5_U.u2.a  = \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_5_U.ain_s1 ;
assign \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_5_U.u2.b  = \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_5_U.bin_s1 ;
assign \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_5_U.u2.cin  = \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_5_U.carry_s1 ;
assign \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_5_U.facout_s2  = \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_5_U.u2.cout ;
assign \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_5_U.fas_s2  = \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_5_U.u2.s ;
assign \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_5_U.u1.a  = \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_5_U.a [15:0];
assign \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_5_U.u1.b  = \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_5_U.b [15:0];
assign \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_5_U.u1.cin  = 1'h0;
assign \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_5_U.facout_s1  = \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_5_U.u1.cout ;
assign \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_5_U.fas_s1  = \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_5_U.u1.s ;
assign \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_5_U.a  = \add_32ns_32s_32_2_1_U22.din0 ;
assign \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_5_U.b  = \add_32ns_32s_32_2_1_U22.din1 ;
assign \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_5_U.ce  = \add_32ns_32s_32_2_1_U22.ce ;
assign \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_5_U.clk  = \add_32ns_32s_32_2_1_U22.clk ;
assign \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_5_U.reset  = \add_32ns_32s_32_2_1_U22.reset ;
assign \add_32ns_32s_32_2_1_U22.dout  = \add_32ns_32s_32_2_1_U22.top_add_32ns_32s_32_2_1_Adder_5_U.s ;
assign \add_32ns_32s_32_2_1_U22.ce  = 1'h1;
assign \add_32ns_32s_32_2_1_U22.clk  = ap_clk;
assign \add_32ns_32s_32_2_1_U22.din0  = ret_V_26_reg_1383;
assign \add_32ns_32s_32_2_1_U22.din1  = { op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18 };
assign grp_fu_892_p2 = \add_32ns_32s_32_2_1_U22.dout ;
assign \add_32ns_32s_32_2_1_U22.reset  = ap_rst;
assign \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_5_U.ain_s0  = \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_5_U.a ;
assign \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_5_U.bin_s0  = \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_5_U.b ;
assign \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_5_U.s  = { \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_5_U.fas_s2 , \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_5_U.sum_s1  };
assign \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_5_U.u2.a  = \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_5_U.ain_s1 ;
assign \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_5_U.u2.b  = \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_5_U.bin_s1 ;
assign \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_5_U.u2.cin  = \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_5_U.carry_s1 ;
assign \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_5_U.facout_s2  = \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_5_U.u2.cout ;
assign \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_5_U.fas_s2  = \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_5_U.u2.s ;
assign \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_5_U.u1.a  = \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_5_U.a [15:0];
assign \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_5_U.u1.b  = \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_5_U.b [15:0];
assign \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_5_U.u1.cin  = 1'h0;
assign \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_5_U.facout_s1  = \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_5_U.u1.cout ;
assign \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_5_U.fas_s1  = \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_5_U.u1.s ;
assign \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_5_U.a  = \add_32ns_32s_32_2_1_U16.din0 ;
assign \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_5_U.b  = \add_32ns_32s_32_2_1_U16.din1 ;
assign \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_5_U.ce  = \add_32ns_32s_32_2_1_U16.ce ;
assign \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_5_U.clk  = \add_32ns_32s_32_2_1_U16.clk ;
assign \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_5_U.reset  = \add_32ns_32s_32_2_1_U16.reset ;
assign \add_32ns_32s_32_2_1_U16.dout  = \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_5_U.s ;
assign \add_32ns_32s_32_2_1_U16.ce  = 1'h1;
assign \add_32ns_32s_32_2_1_U16.clk  = ap_clk;
assign \add_32ns_32s_32_2_1_U16.din0  = ret_V_23_reg_1206;
assign \add_32ns_32s_32_2_1_U16.din1  = { op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13 };
assign grp_fu_659_p2 = \add_32ns_32s_32_2_1_U16.dout ;
assign \add_32ns_32s_32_2_1_U16.reset  = ap_rst;
assign \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_4_U.ain_s0  = \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_4_U.a ;
assign \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_4_U.bin_s0  = \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_4_U.b ;
assign \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_4_U.s  = { \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_4_U.fas_s2 , \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_4_U.sum_s1  };
assign \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.a  = \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_4_U.ain_s1 ;
assign \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.b  = \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_4_U.bin_s1 ;
assign \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.cin  = \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_4_U.carry_s1 ;
assign \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_4_U.facout_s2  = \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.cout ;
assign \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_4_U.fas_s2  = \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.s ;
assign \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.a  = \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_4_U.a [15:0];
assign \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.b  = \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_4_U.b [15:0];
assign \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.cin  = 1'h0;
assign \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_4_U.facout_s1  = \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.cout ;
assign \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_4_U.fas_s1  = \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.s ;
assign \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_4_U.a  = \add_32ns_32ns_32_2_1_U9.din0 ;
assign \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_4_U.b  = \add_32ns_32ns_32_2_1_U9.din1 ;
assign \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_4_U.ce  = \add_32ns_32ns_32_2_1_U9.ce ;
assign \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_4_U.clk  = \add_32ns_32ns_32_2_1_U9.clk ;
assign \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_4_U.reset  = \add_32ns_32ns_32_2_1_U9.reset ;
assign \add_32ns_32ns_32_2_1_U9.dout  = \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_4_U.s ;
assign \add_32ns_32ns_32_2_1_U9.ce  = 1'h1;
assign \add_32ns_32ns_32_2_1_U9.clk  = ap_clk;
assign \add_32ns_32ns_32_2_1_U9.din0  = ret_V_21_reg_1112;
assign \add_32ns_32ns_32_2_1_U9.din1  = { 24'h000000, op_10 };
assign grp_fu_480_p2 = \add_32ns_32ns_32_2_1_U9.dout ;
assign \add_32ns_32ns_32_2_1_U9.reset  = ap_rst;
assign \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.ain_s0  = \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.a ;
assign \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.bin_s0  = \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.b ;
assign \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.s  = { \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.fas_s2 , \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.sum_s1  };
assign \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.a  = \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.ain_s1 ;
assign \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.b  = \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.bin_s1 ;
assign \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.cin  = \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.carry_s1 ;
assign \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.facout_s2  = \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.cout ;
assign \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.fas_s2  = \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.s ;
assign \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.a  = \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.a [15:0];
assign \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.b  = \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.b [15:0];
assign \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.cin  = 1'h0;
assign \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.facout_s1  = \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.cout ;
assign \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.fas_s1  = \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.s ;
assign \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.a  = \add_32ns_32ns_32_2_1_U8.din0 ;
assign \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.b  = \add_32ns_32ns_32_2_1_U8.din1 ;
assign \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.ce  = \add_32ns_32ns_32_2_1_U8.ce ;
assign \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.clk  = \add_32ns_32ns_32_2_1_U8.clk ;
assign \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.reset  = \add_32ns_32ns_32_2_1_U8.reset ;
assign \add_32ns_32ns_32_2_1_U8.dout  = \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.s ;
assign \add_32ns_32ns_32_2_1_U8.ce  = 1'h1;
assign \add_32ns_32ns_32_2_1_U8.clk  = ap_clk;
assign \add_32ns_32ns_32_2_1_U8.din0  = ret_V_8_cast_reg_1100;
assign \add_32ns_32ns_32_2_1_U8.din1  = 32'd1;
assign grp_fu_452_p2 = \add_32ns_32ns_32_2_1_U8.dout ;
assign \add_32ns_32ns_32_2_1_U8.reset  = ap_rst;
assign \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.ain_s0  = \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.a ;
assign \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.bin_s0  = \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.b ;
assign \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.s  = { \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.fas_s2 , \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.sum_s1  };
assign \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.a  = \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.ain_s1 ;
assign \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.b  = \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.bin_s1 ;
assign \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.cin  = \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.carry_s1 ;
assign \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.facout_s2  = \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.cout ;
assign \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.fas_s2  = \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.s ;
assign \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.a  = \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.a [15:0];
assign \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.b  = \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.b [15:0];
assign \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.cin  = 1'h0;
assign \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.facout_s1  = \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.cout ;
assign \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.fas_s1  = \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.s ;
assign \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.a  = \add_32ns_32ns_32_2_1_U5.din0 ;
assign \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.b  = \add_32ns_32ns_32_2_1_U5.din1 ;
assign \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.ce  = \add_32ns_32ns_32_2_1_U5.ce ;
assign \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.clk  = \add_32ns_32ns_32_2_1_U5.clk ;
assign \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.reset  = \add_32ns_32ns_32_2_1_U5.reset ;
assign \add_32ns_32ns_32_2_1_U5.dout  = \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.s ;
assign \add_32ns_32ns_32_2_1_U5.ce  = 1'h1;
assign \add_32ns_32ns_32_2_1_U5.clk  = ap_clk;
assign \add_32ns_32ns_32_2_1_U5.din0  = ret_V_4_cast_reg_1053;
assign \add_32ns_32ns_32_2_1_U5.din1  = 32'd1;
assign grp_fu_378_p2 = \add_32ns_32ns_32_2_1_U5.dout ;
assign \add_32ns_32ns_32_2_1_U5.reset  = ap_rst;
assign \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_4_U.ain_s0  = \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_4_U.a ;
assign \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_4_U.bin_s0  = \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_4_U.b ;
assign \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_4_U.s  = { \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_4_U.fas_s2 , \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_4_U.sum_s1  };
assign \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.a  = \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_4_U.ain_s1 ;
assign \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.b  = \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_4_U.bin_s1 ;
assign \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.cin  = \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_4_U.carry_s1 ;
assign \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_4_U.facout_s2  = \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.cout ;
assign \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_4_U.fas_s2  = \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.s ;
assign \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.a  = \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_4_U.a [15:0];
assign \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.b  = \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_4_U.b [15:0];
assign \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.cin  = 1'h0;
assign \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_4_U.facout_s1  = \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.cout ;
assign \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_4_U.fas_s1  = \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.s ;
assign \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_4_U.a  = \add_32ns_32ns_32_2_1_U24.din0 ;
assign \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_4_U.b  = \add_32ns_32ns_32_2_1_U24.din1 ;
assign \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_4_U.ce  = \add_32ns_32ns_32_2_1_U24.ce ;
assign \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_4_U.clk  = \add_32ns_32ns_32_2_1_U24.clk ;
assign \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_4_U.reset  = \add_32ns_32ns_32_2_1_U24.reset ;
assign \add_32ns_32ns_32_2_1_U24.dout  = \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_4_U.s ;
assign \add_32ns_32ns_32_2_1_U24.ce  = 1'h1;
assign \add_32ns_32ns_32_2_1_U24.clk  = ap_clk;
assign \add_32ns_32ns_32_2_1_U24.din0  = ret_V_24_cast_reg_1424;
assign \add_32ns_32ns_32_2_1_U24.din1  = 32'd1;
assign grp_fu_947_p2 = \add_32ns_32ns_32_2_1_U24.dout ;
assign \add_32ns_32ns_32_2_1_U24.reset  = ap_rst;
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_4_U.ain_s0  = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_4_U.a ;
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_4_U.bin_s0  = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_4_U.b ;
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_4_U.s  = { \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_4_U.fas_s2 , \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_4_U.sum_s1  };
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.a  = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_4_U.ain_s1 ;
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.b  = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_4_U.bin_s1 ;
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.cin  = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_4_U.carry_s1 ;
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_4_U.facout_s2  = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.cout ;
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_4_U.fas_s2  = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.s ;
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.a  = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_4_U.a [15:0];
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.b  = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_4_U.b [15:0];
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.cin  = 1'h0;
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_4_U.facout_s1  = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.cout ;
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_4_U.fas_s1  = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.s ;
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_4_U.a  = \add_32ns_32ns_32_2_1_U21.din0 ;
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_4_U.b  = \add_32ns_32ns_32_2_1_U21.din1 ;
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_4_U.ce  = \add_32ns_32ns_32_2_1_U21.ce ;
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_4_U.clk  = \add_32ns_32ns_32_2_1_U21.clk ;
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_4_U.reset  = \add_32ns_32ns_32_2_1_U21.reset ;
assign \add_32ns_32ns_32_2_1_U21.dout  = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_4_U.s ;
assign \add_32ns_32ns_32_2_1_U21.ce  = 1'h1;
assign \add_32ns_32ns_32_2_1_U21.clk  = ap_clk;
assign \add_32ns_32ns_32_2_1_U21.din0  = ret_V_21_cast_reg_1341;
assign \add_32ns_32ns_32_2_1_U21.din1  = 32'd1;
assign grp_fu_798_p2 = \add_32ns_32ns_32_2_1_U21.dout ;
assign \add_32ns_32ns_32_2_1_U21.reset  = ap_rst;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_4_U.ain_s0  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_4_U.a ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_4_U.bin_s0  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_4_U.b ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_4_U.s  = { \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_4_U.fas_s2 , \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_4_U.sum_s1  };
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.a  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_4_U.ain_s1 ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.b  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_4_U.bin_s1 ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.cin  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_4_U.carry_s1 ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_4_U.facout_s2  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.cout ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_4_U.fas_s2  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.s ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.a  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_4_U.a [15:0];
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.b  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_4_U.b [15:0];
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.cin  = 1'h0;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_4_U.facout_s1  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.cout ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_4_U.fas_s1  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.s ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_4_U.a  = \add_32ns_32ns_32_2_1_U12.din0 ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_4_U.b  = \add_32ns_32ns_32_2_1_U12.din1 ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_4_U.ce  = \add_32ns_32ns_32_2_1_U12.ce ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_4_U.clk  = \add_32ns_32ns_32_2_1_U12.clk ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_4_U.reset  = \add_32ns_32ns_32_2_1_U12.reset ;
assign \add_32ns_32ns_32_2_1_U12.dout  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_4_U.s ;
assign \add_32ns_32ns_32_2_1_U12.ce  = 1'h1;
assign \add_32ns_32ns_32_2_1_U12.clk  = ap_clk;
assign \add_32ns_32ns_32_2_1_U12.din0  = ret_V_14_cast_reg_1172;
assign \add_32ns_32ns_32_2_1_U12.din1  = 32'd1;
assign grp_fu_584_p2 = \add_32ns_32ns_32_2_1_U12.dout ;
assign \add_32ns_32ns_32_2_1_U12.reset  = ap_rst;
assign \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_10_U.ain_s0  = \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_10_U.a ;
assign \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_10_U.bin_s0  = \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_10_U.b ;
assign \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_10_U.s  = { \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_10_U.fas_s2 , \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_10_U.sum_s1  };
assign \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_10_U.u2.a  = \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_10_U.ain_s1 ;
assign \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_10_U.u2.b  = \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_10_U.bin_s1 ;
assign \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_10_U.u2.cin  = \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_10_U.carry_s1 ;
assign \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_10_U.facout_s2  = \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_10_U.u2.cout ;
assign \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_10_U.fas_s2  = \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_10_U.u2.s ;
assign \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_10_U.u1.a  = \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_10_U.a [4:0];
assign \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_10_U.u1.b  = \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_10_U.b [4:0];
assign \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_10_U.u1.cin  = 1'h0;
assign \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_10_U.facout_s1  = \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_10_U.u1.cout ;
assign \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_10_U.fas_s1  = \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_10_U.u1.s ;
assign \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_10_U.a  = \add_10s_10ns_10_2_1_U17.din0 ;
assign \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_10_U.b  = \add_10s_10ns_10_2_1_U17.din1 ;
assign \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_10_U.ce  = \add_10s_10ns_10_2_1_U17.ce ;
assign \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_10_U.clk  = \add_10s_10ns_10_2_1_U17.clk ;
assign \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_10_U.reset  = \add_10s_10ns_10_2_1_U17.reset ;
assign \add_10s_10ns_10_2_1_U17.dout  = \add_10s_10ns_10_2_1_U17.top_add_10s_10ns_10_2_1_Adder_10_U.s ;
assign \add_10s_10ns_10_2_1_U17.ce  = 1'h1;
assign \add_10s_10ns_10_2_1_U17.clk  = ap_clk;
assign \add_10s_10ns_10_2_1_U17.din0  = { op_16[7], op_16[7], op_16 };
assign \add_10s_10ns_10_2_1_U17.din1  = { 2'h0, op_15 };
assign grp_fu_672_p2 = \add_10s_10ns_10_2_1_U17.dout ;
assign \add_10s_10ns_10_2_1_U17.reset  = ap_rst;
endmodule


// Machine B:
// Processed by function `add_clk_enable_signal` in `verilog_tricks.py`.
// Processed by function `remove_reset_signal` in `verilog_tricks.py`.
module top_B (
  ap_clk,
  ap_start,
  ap_done,
  ap_idle,
  ap_ready,
  op_0,
  op_1,
  op_2,
  op_4,
  op_5,
  op_6,
  op_8,
  op_9,
  op_10,
  op_12,
  op_13,
  op_14,
  op_15,
  op_16,
  op_17,
  op_18,
  op_32,
  op_32_ap_vld,
clk_enable
);
input clk_enable;


input ap_clk;
wire ap_rst;
assign ap_rst = op_32_ap_vld;
input ap_start;
input op_0;
input [3:0] op_1;
input [7:0] op_10;
input [3:0] op_12;
input [7:0] op_13;
input [1:0] op_14;
input [7:0] op_15;
input [7:0] op_16;
input [3:0] op_17;
input [1:0] op_18;
input [3:0] op_2;
input [15:0] op_4;
input [7:0] op_5;
input [15:0] op_6;
input [3:0] op_8;
input [3:0] op_9;
output ap_done;
output ap_idle;
output ap_ready;
output [31:0] op_32;
output op_32_ap_vld;


reg [9:0] add_ln69_reg_1088;
reg and_ln786_reg_1149;
reg [8:0] ap_CS_fsm = 9'h001;
reg deleted_zeros_reg_1144;
reg icmp_ln410_reg_1078;
reg icmp_ln851_1_reg_1041;
reg icmp_ln851_2_reg_1063;
reg [31:0] op_23_V_reg_1046;
reg [31:0] op_25_V_reg_1068;
reg p_Result_11_reg_1098;
reg p_Result_13_reg_1107;
reg p_Result_14_reg_1119;
reg [3:0] p_Val2_5_reg_1113;
reg [43:0] ret_V_17_reg_1029;
reg [35:0] ret_V_20_reg_1051;
reg [31:0] ret_V_21_cast_reg_1132;
reg [31:0] ret_V_23_reg_1083;
reg [33:0] ret_V_25_reg_1127;
reg [31:0] ret_V_27_reg_1159;
reg [31:0] ret_V_4_cast_reg_1034;
reg [31:0] ret_V_8_cast_reg_1056;
reg [4:0] ret_reg_1024;
reg [3:0] select_ln340_reg_1154;
reg [7:0] trunc_ln_reg_1073;
reg xor_ln416_reg_1139;
wire [9:0] _000_;
wire _001_;
wire [8:0] _002_;
wire _003_;
wire _004_;
wire _005_;
wire _006_;
wire [31:0] _007_;
wire [31:0] _008_;
wire _009_;
wire _010_;
wire _011_;
wire [3:0] _012_;
wire [43:0] _013_;
wire [35:0] _014_;
wire [31:0] _015_;
wire [31:0] _016_;
wire [33:0] _017_;
wire [31:0] _018_;
wire [31:0] _019_;
wire [31:0] _020_;
wire [4:0] _021_;
wire [3:0] _022_;
wire [7:0] _023_;
wire _024_;
wire [1:0] _025_;
wire _026_;
wire _027_;
wire _028_;
wire _029_;
wire _030_;
wire _031_;
wire _032_;
wire _033_;
wire _034_;
wire _035_;
wire _036_;
wire _037_;
wire _038_;
wire _039_;
wire _040_;
wire _041_;
wire _042_;
wire _043_;
wire Range1_all_zeros_fu_824_p2;
wire [7:0] add_ln1192_1_fu_676_p2;
wire [31:0] add_ln691_1_fu_393_p2;
wire [31:0] add_ln691_2_fu_469_p2;
wire [31:0] add_ln691_3_fu_606_p2;
wire [31:0] add_ln691_4_fu_909_p2;
wire [31:0] add_ln691_5_fu_1001_p2;
wire [6:0] add_ln691_fu_322_p2;
wire [9:0] add_ln69_fu_636_p2;
wire and_ln412_fu_740_p2;
wire and_ln785_1_fu_947_p2;
wire and_ln785_fu_938_p2;
wire and_ln786_fu_875_p2;
wire [16:0] and_ln_fu_541_p4;
wire ap_CS_fsm_state1;
wire ap_CS_fsm_state2;
wire ap_CS_fsm_state3;
wire ap_CS_fsm_state4;
wire ap_CS_fsm_state5;
wire ap_CS_fsm_state6;
wire ap_CS_fsm_state7;
wire ap_CS_fsm_state8;
wire ap_CS_fsm_state9;
wire [8:0] ap_NS_fsm;
wire ap_clk;
wire ap_done;
wire ap_idle;
wire ap_ready;
wire ap_rst;
wire ap_start;
wire carry_1_fu_819_p2;
wire deleted_ones_fu_836_p3;
wire deleted_zeros_fu_829_p3;
wire icmp_ln410_fu_551_p2;
wire icmp_ln851_1_fu_380_p2;
wire icmp_ln851_2_fu_456_p2;
wire icmp_ln851_3_fu_600_p2;
wire icmp_ln851_fu_316_p2;
wire neg_src_fu_853_p2;
wire op_0;
wire [3:0] op_1;
wire [7:0] op_10;
wire [7:0] op_11_V_fu_645_p2;
wire [3:0] op_12;
wire [7:0] op_13;
wire [1:0] op_14;
wire [7:0] op_15;
wire [7:0] op_16;
wire [3:0] op_17;
wire [1:0] op_18;
wire [3:0] op_19_V_fu_952_p3;
wire [3:0] op_2;
wire [31:0] op_23_V_fu_415_p2;
wire [31:0] op_25_V_fu_491_p2;
wire [31:0] op_29_V_fu_776_p2;
wire [31:0] op_32;
wire op_32_ap_vld;
wire [15:0] op_4;
wire [7:0] op_5;
wire [15:0] op_6;
wire [3:0] op_8;
wire [3:0] op_9;
wire or_ln340_1_fu_886_p2;
wire or_ln340_fu_880_p2;
wire or_ln412_fu_734_p2;
wire or_ln781_fu_848_p2;
wire or_ln785_1_fu_942_p2;
wire or_ln785_fu_864_p2;
wire overflow_fu_869_p2;
wire p_Result_10_fu_989_p3;
wire p_Result_12_fu_708_p3;
wire p_Result_1_fu_386_p3;
wire p_Result_5_fu_700_p3;
wire p_Result_7_fu_462_p3;
wire p_Result_8_fu_588_p3;
wire p_Result_9_fu_899_p3;
wire p_Result_s_fu_304_p3;
wire [3:0] p_Val2_4_fu_690_p4;
wire [3:0] p_Val2_5_fu_750_p2;
wire r_fu_720_p2;
wire [31:0] ret_V_14_cast_fu_578_p4;
wire [8:0] ret_V_15_fu_284_p2;
wire [16:0] ret_V_16_fu_513_p2;
wire [43:0] ret_V_17_fu_360_p2;
wire [31:0] ret_V_18_fu_404_p3;
wire [8:0] ret_V_19_fu_670_p2;
wire [35:0] ret_V_20_fu_436_p2;
wire [31:0] ret_V_21_fu_480_p3;
wire [35:0] ret_V_22_fu_572_p2;
wire [31:0] ret_V_23_fu_620_p3;
wire [31:0] ret_V_24_cast_fu_979_p4;
wire [31:0] ret_V_24_fu_768_p2;
wire [33:0] ret_V_25_fu_798_p2;
wire [31:0] ret_V_26_fu_921_p3;
wire [31:0] ret_V_27_fu_932_p2;
wire [33:0] ret_V_28_fu_973_p2;
wire [4:0] ret_fu_263_p2;
wire [32:0] rhs_10_fu_786_p3;
wire [32:0] rhs_13_fu_962_p3;
wire [7:0] rhs_1_fu_273_p3;
wire [9:0] rhs_2_fu_501_p3;
wire [6:0] rhs_3_fu_654_p3;
wire [34:0] rhs_5_fu_425_p3;
wire [34:0] rhs_7_fu_561_p3;
wire [4:0] select_ln215_fu_251_p3;
wire [3:0] select_ln340_fu_892_p3;
wire [6:0] select_ln353_fu_340_p3;
wire [31:0] select_ln850_1_fu_398_p3;
wire [31:0] select_ln850_2_fu_474_p3;
wire [31:0] select_ln850_3_fu_612_p3;
wire [31:0] select_ln850_4_fu_914_p3;
wire [31:0] select_ln850_5_fu_1007_p3;
wire [6:0] select_ln850_fu_332_p3;
wire [33:0] sext_ln1192_10_fu_969_p1;
wire [8:0] sext_ln1192_1_fu_280_p1;
wire [43:0] sext_ln1192_2_fu_356_p1;
wire [8:0] sext_ln1192_3_fu_662_p1;
wire [7:0] sext_ln1192_4_fu_666_p1;
wire [35:0] sext_ln1192_5_fu_432_p1;
wire [35:0] sext_ln1192_6_fu_568_p1;
wire [31:0] sext_ln1192_7_fu_764_p1;
wire [33:0] sext_ln1192_8_fu_794_p1;
wire [31:0] sext_ln1192_9_fu_928_p1;
wire [7:0] sext_ln1192_fu_269_p0;
wire [8:0] sext_ln1192_fu_269_p1;
wire [4:0] sext_ln215_fu_259_p1;
wire [9:0] sext_ln69_1_fu_632_p1;
wire [31:0] sext_ln69_2_fu_773_p1;
wire [31:0] sext_ln69_fu_411_p1;
wire [15:0] sext_ln703_1_fu_328_p0;
wire [43:0] sext_ln703_1_fu_328_p1;
wire [8:0] sext_ln703_2_fu_650_p1;
wire [3:0] sext_ln703_3_fu_421_p0;
wire [35:0] sext_ln703_3_fu_421_p1;
wire [3:0] sext_ln703_4_fu_557_p0;
wire [35:0] sext_ln703_4_fu_557_p1;
wire [3:0] sext_ln703_5_fu_782_p0;
wire [33:0] sext_ln703_5_fu_782_p1;
wire [33:0] sext_ln703_6_fu_958_p1;
wire [16:0] sext_ln703_fu_497_p1;
wire [6:0] sext_ln850_fu_300_p1;
wire [5:0] tmp_1_fu_290_p4;
wire [17:0] tmp_2_fu_348_p3;
wire tmp_fu_529_p3;
wire trunc_ln410_fu_537_p1;
wire [2:0] trunc_ln718_fu_716_p1;
wire [15:0] trunc_ln851_1_fu_376_p0;
wire [10:0] trunc_ln851_1_fu_376_p1;
wire [3:0] trunc_ln851_2_fu_452_p0;
wire [2:0] trunc_ln851_2_fu_452_p1;
wire [3:0] trunc_ln851_3_fu_596_p0;
wire [2:0] trunc_ln851_3_fu_596_p1;
wire [3:0] trunc_ln851_4_fu_906_p0;
wire trunc_ln851_4_fu_906_p1;
wire trunc_ln851_5_fu_997_p1;
wire [7:0] trunc_ln851_fu_312_p0;
wire [2:0] trunc_ln851_fu_312_p1;
wire xor_ln416_fu_814_p2;
wire xor_ln781_fu_843_p2;
wire xor_ln785_fu_858_p2;
wire [16:0] zext_ln1193_fu_509_p1;
wire [3:0] zext_ln415_1_fu_746_p1;
wire [7:0] zext_ln415_fu_642_p1;
wire [9:0] zext_ln69_1_fu_628_p1;
wire [31:0] zext_ln69_fu_487_p1;


assign add_ln1192_1_fu_676_p2 = $signed({ op_14, 5'h00 }) + $signed(op_11_V_fu_645_p2);
assign add_ln691_1_fu_393_p2 = ret_V_4_cast_reg_1034 + 1'h1;
assign add_ln691_2_fu_469_p2 = ret_V_8_cast_reg_1056 + 1'h1;
assign add_ln691_3_fu_606_p2 = ret_V_22_fu_572_p2[34:3] + 1'h1;
assign add_ln691_4_fu_909_p2 = ret_V_21_cast_reg_1132 + 1'h1;
assign add_ln691_5_fu_1001_p2 = ret_V_28_fu_973_p2[32:1] + 1'h1;
assign add_ln691_fu_322_p2 = $signed(ret_V_15_fu_284_p2[8:3]) + $signed(2'h1);
assign add_ln69_fu_636_p2 = $signed(op_16) + $signed({ 1'h0, op_15 });
assign op_11_V_fu_645_p2 = trunc_ln_reg_1073 + icmp_ln410_reg_1078;
assign op_23_V_fu_415_p2 = $signed(ret_V_18_fu_404_p3) + $signed(op_8);
assign op_25_V_fu_491_p2 = ret_V_21_fu_480_p3 + op_10;
assign op_29_V_fu_776_p2 = $signed(add_ln69_reg_1088) + $signed(ret_V_24_fu_768_p2);
assign p_Val2_5_fu_750_p2 = add_ln1192_1_fu_676_p2[7:4] + and_ln412_fu_740_p2;
assign ret_V_15_fu_284_p2 = $signed({ ret_reg_1024, 3'h0 }) + $signed(op_5);
assign { ret_V_17_fu_360_p2[43], ret_V_17_fu_360_p2[17:0] } = $signed({ select_ln353_fu_340_p3, 11'h000 }) + $signed(op_6);
assign ret_V_19_fu_670_p2 = $signed({ op_14, 5'h00 }) + $signed(op_11_V_fu_645_p2);
assign ret_V_20_fu_436_p2 = $signed({ op_23_V_reg_1046, 3'h0 }) + $signed(op_9);
assign ret_V_22_fu_572_p2 = $signed({ op_25_V_reg_1068, 3'h0 }) + $signed(op_12);
assign ret_V_24_fu_768_p2 = $signed(ret_V_23_reg_1083) + $signed(op_13);
assign ret_V_25_fu_798_p2 = $signed({ op_29_V_fu_776_p2, 1'h0 }) + $signed(op_17);
assign ret_V_27_fu_932_p2 = $signed(ret_V_26_fu_921_p3) + $signed(op_18);
assign ret_V_28_fu_973_p2 = $signed({ ret_V_27_reg_1159, 1'h0 }) + $signed(op_19_V_fu_952_p3);
assign ret_fu_263_p2 = $signed(op_2) + $signed(select_ln215_fu_251_p3);
assign _026_ = ap_CS_fsm[0] & _028_;
assign _027_ = ap_CS_fsm[0] & ap_start;
assign and_ln412_fu_740_p2 = op_11_V_fu_645_p2[3] & or_ln412_fu_734_p2;
assign and_ln785_1_fu_947_p2 = or_ln785_1_fu_942_p2 & and_ln786_reg_1149;
assign and_ln785_fu_938_p2 = xor_ln416_reg_1139 & deleted_zeros_reg_1144;
assign and_ln786_fu_875_p2 = p_Result_14_reg_1119 & deleted_ones_fu_836_p3;
assign carry_1_fu_819_p2 = xor_ln416_fu_814_p2 & p_Result_13_reg_1107;
assign neg_src_fu_853_p2 = p_Result_11_reg_1098 & or_ln781_fu_848_p2;
assign overflow_fu_869_p2 = or_ln785_fu_864_p2 & Range1_all_zeros_fu_824_p2;
assign Range1_all_zeros_fu_824_p2 = ~ p_Result_11_reg_1098;
assign xor_ln416_fu_814_p2 = ~ p_Result_14_reg_1119;
assign xor_ln781_fu_843_p2 = ~ p_Result_13_reg_1107;
assign xor_ln785_fu_858_p2 = ~ deleted_zeros_fu_829_p3;
assign _028_ = ~ ap_start;
assign _029_ = { ret_V_16_fu_513_p2[16], ret_V_16_fu_513_p2[0] } == 1'h1;
assign _030_ = | op_6[10:0];
assign _031_ = | op_9[2:0];
assign _032_ = | op_12[2:0];
assign _033_ = | op_5[2:0];
assign _034_ = | op_11_V_fu_645_p2[2:0];
assign or_ln340_1_fu_886_p2 = or_ln340_fu_880_p2 | neg_src_fu_853_p2;
assign or_ln340_fu_880_p2 = overflow_fu_869_p2 | and_ln786_fu_875_p2;
assign or_ln412_fu_734_p2 = r_fu_720_p2 | add_ln1192_1_fu_676_p2[4];
assign or_ln781_fu_848_p2 = xor_ln781_fu_843_p2 | p_Result_14_reg_1119;
assign or_ln785_1_fu_942_p2 = p_Result_11_reg_1098 | and_ln785_fu_938_p2;
assign or_ln785_fu_864_p2 = xor_ln785_fu_858_p2 | p_Result_14_reg_1119;
always @(posedge ap_clk)
ret_reg_1024 <= _021_;
always @(posedge ap_clk)
p_Result_11_reg_1098 <= _009_;
always @(posedge ap_clk)
p_Result_13_reg_1107 <= _010_;
always @(posedge ap_clk)
p_Val2_5_reg_1113 <= _012_;
always @(posedge ap_clk)
p_Result_14_reg_1119 <= _011_;
always @(posedge ap_clk)
ret_V_25_reg_1127 <= _017_;
always @(posedge ap_clk)
ret_V_21_cast_reg_1132 <= _015_;
always @(posedge ap_clk)
op_25_V_reg_1068 <= _008_;
always @(posedge ap_clk)
op_23_V_reg_1046 <= _007_;
always @(posedge ap_clk)
ret_V_20_reg_1051 <= _014_;
always @(posedge ap_clk)
ret_V_8_cast_reg_1056 <= _020_;
always @(posedge ap_clk)
icmp_ln851_2_reg_1063 <= _006_;
always @(posedge ap_clk)
ret_V_17_reg_1029 <= _013_;
always @(posedge ap_clk)
ret_V_4_cast_reg_1034 <= _019_;
always @(posedge ap_clk)
icmp_ln851_1_reg_1041 <= _005_;
always @(posedge ap_clk)
xor_ln416_reg_1139 <= _024_;
always @(posedge ap_clk)
deleted_zeros_reg_1144 <= _003_;
always @(posedge ap_clk)
and_ln786_reg_1149 <= _001_;
always @(posedge ap_clk)
select_ln340_reg_1154 <= _022_;
always @(posedge ap_clk)
ret_V_27_reg_1159 <= _018_;
always @(posedge ap_clk)
trunc_ln_reg_1073 <= _023_;
always @(posedge ap_clk)
icmp_ln410_reg_1078 <= _004_;
always @(posedge ap_clk)
ret_V_23_reg_1083 <= _016_;
always @(posedge ap_clk)
add_ln69_reg_1088 <= _000_;
always @(posedge ap_clk)
ap_CS_fsm <= _002_;
assign _025_ = _027_ ? 2'h2 : 2'h1;
assign _035_ = ap_CS_fsm == 1'h1;
function [8:0] _120_;
input [8:0] a;
input [80:0] b;
input [8:0] s;
case (s)
9'b000000001:
_120_ = b[8:0];
9'b000000010:
_120_ = b[17:9];
9'b000000100:
_120_ = b[26:18];
9'b000001000:
_120_ = b[35:27];
9'b000010000:
_120_ = b[44:36];
9'b000100000:
_120_ = b[53:45];
9'b001000000:
_120_ = b[62:54];
9'b010000000:
_120_ = b[71:63];
9'b100000000:
_120_ = b[80:72];
9'b000000000:
_120_ = a;
default:
_120_ = 9'bx;
endcase
endfunction
assign ap_NS_fsm = _120_(9'hxxx, { 7'h00, _025_, 72'h020202020202020001 }, { _035_, _043_, _042_, _041_, _040_, _039_, _038_, _037_, _036_ });
assign _036_ = ap_CS_fsm == 9'h100;
assign _037_ = ap_CS_fsm == 8'h80;
assign _038_ = ap_CS_fsm == 7'h40;
assign _039_ = ap_CS_fsm == 6'h20;
assign _040_ = ap_CS_fsm == 5'h10;
assign _041_ = ap_CS_fsm == 4'h8;
assign _042_ = ap_CS_fsm == 3'h4;
assign _043_ = ap_CS_fsm == 2'h2;
assign op_32_ap_vld = ap_CS_fsm[8] ? 1'h1 : 1'h0;
assign ap_idle = _026_ ? 1'h1 : 1'h0;
assign _021_ = ap_CS_fsm[0] ? ret_fu_263_p2 : ret_reg_1024;
assign _015_ = ap_CS_fsm[6] ? ret_V_25_fu_798_p2[32:1] : ret_V_21_cast_reg_1132;
assign _017_ = ap_CS_fsm[6] ? ret_V_25_fu_798_p2 : ret_V_25_reg_1127;
assign _011_ = ap_CS_fsm[6] ? p_Val2_5_fu_750_p2[3] : p_Result_14_reg_1119;
assign _012_ = ap_CS_fsm[6] ? p_Val2_5_fu_750_p2 : p_Val2_5_reg_1113;
assign _010_ = ap_CS_fsm[6] ? add_ln1192_1_fu_676_p2[7] : p_Result_13_reg_1107;
assign _009_ = ap_CS_fsm[6] ? ret_V_19_fu_670_p2[8] : p_Result_11_reg_1098;
assign _008_ = ap_CS_fsm[4] ? op_25_V_fu_491_p2 : op_25_V_reg_1068;
assign _007_ = ap_CS_fsm[2] ? op_23_V_fu_415_p2 : op_23_V_reg_1046;
assign _006_ = ap_CS_fsm[3] ? icmp_ln851_2_fu_456_p2 : icmp_ln851_2_reg_1063;
assign _020_ = ap_CS_fsm[3] ? ret_V_20_fu_436_p2[34:3] : ret_V_8_cast_reg_1056;
assign _014_ = ap_CS_fsm[3] ? ret_V_20_fu_436_p2 : ret_V_20_reg_1051;
assign _005_ = ap_CS_fsm[1] ? icmp_ln851_1_fu_380_p2 : icmp_ln851_1_reg_1041;
assign _019_ = ap_CS_fsm[1] ? { ret_V_17_fu_360_p2[43], ret_V_17_fu_360_p2[43], ret_V_17_fu_360_p2[43], ret_V_17_fu_360_p2[43], ret_V_17_fu_360_p2[43], ret_V_17_fu_360_p2[43], ret_V_17_fu_360_p2[43], ret_V_17_fu_360_p2[43], ret_V_17_fu_360_p2[43], ret_V_17_fu_360_p2[43], ret_V_17_fu_360_p2[43], ret_V_17_fu_360_p2[43], ret_V_17_fu_360_p2[43], ret_V_17_fu_360_p2[43], ret_V_17_fu_360_p2[43], ret_V_17_fu_360_p2[43], ret_V_17_fu_360_p2[43], ret_V_17_fu_360_p2[43], ret_V_17_fu_360_p2[43], ret_V_17_fu_360_p2[43], ret_V_17_fu_360_p2[43], ret_V_17_fu_360_p2[43], ret_V_17_fu_360_p2[43], ret_V_17_fu_360_p2[43], ret_V_17_fu_360_p2[43], ret_V_17_fu_360_p2[17:11] } : ret_V_4_cast_reg_1034;
assign _013_ = ap_CS_fsm[1] ? { ret_V_17_fu_360_p2[43], ret_V_17_fu_360_p2[43], ret_V_17_fu_360_p2[43], ret_V_17_fu_360_p2[43], ret_V_17_fu_360_p2[43], ret_V_17_fu_360_p2[43], ret_V_17_fu_360_p2[43], ret_V_17_fu_360_p2[43], ret_V_17_fu_360_p2[43], ret_V_17_fu_360_p2[43], ret_V_17_fu_360_p2[43], ret_V_17_fu_360_p2[43], ret_V_17_fu_360_p2[43], ret_V_17_fu_360_p2[43], ret_V_17_fu_360_p2[43], ret_V_17_fu_360_p2[43], ret_V_17_fu_360_p2[43], ret_V_17_fu_360_p2[43], ret_V_17_fu_360_p2[43], ret_V_17_fu_360_p2[43], ret_V_17_fu_360_p2[43], ret_V_17_fu_360_p2[43], ret_V_17_fu_360_p2[43], ret_V_17_fu_360_p2[43], ret_V_17_fu_360_p2[43], ret_V_17_fu_360_p2[43], ret_V_17_fu_360_p2[17:0] } : ret_V_17_reg_1029;
assign _018_ = ap_CS_fsm[7] ? ret_V_27_fu_932_p2 : ret_V_27_reg_1159;
assign _022_ = ap_CS_fsm[7] ? select_ln340_fu_892_p3 : select_ln340_reg_1154;
assign _001_ = ap_CS_fsm[7] ? and_ln786_fu_875_p2 : and_ln786_reg_1149;
assign _003_ = ap_CS_fsm[7] ? deleted_zeros_fu_829_p3 : deleted_zeros_reg_1144;
assign _024_ = ap_CS_fsm[7] ? xor_ln416_fu_814_p2 : xor_ln416_reg_1139;
assign _000_ = ap_CS_fsm[5] ? add_ln69_fu_636_p2 : add_ln69_reg_1088;
assign _016_ = ap_CS_fsm[5] ? ret_V_23_fu_620_p3 : ret_V_23_reg_1083;
assign _004_ = ap_CS_fsm[5] ? icmp_ln410_fu_551_p2 : icmp_ln410_reg_1078;
assign _023_ = ap_CS_fsm[5] ? ret_V_16_fu_513_p2[8:1] : trunc_ln_reg_1073;
assign _002_ = ap_rst ? 9'h001 : ap_NS_fsm;
assign ret_V_16_fu_513_p2 = $signed(op_4) - $signed({ 1'h0, op_1, 6'h00 });
assign deleted_ones_fu_836_p3 = carry_1_fu_819_p2 ? Range1_all_zeros_fu_824_p2 : p_Result_11_reg_1098;
assign deleted_zeros_fu_829_p3 = carry_1_fu_819_p2 ? p_Result_11_reg_1098 : Range1_all_zeros_fu_824_p2;
assign icmp_ln410_fu_551_p2 = _029_ ? 1'h1 : 1'h0;
assign icmp_ln851_1_fu_380_p2 = _030_ ? 1'h1 : 1'h0;
assign icmp_ln851_2_fu_456_p2 = _031_ ? 1'h1 : 1'h0;
assign icmp_ln851_3_fu_600_p2 = _032_ ? 1'h1 : 1'h0;
assign icmp_ln851_fu_316_p2 = _033_ ? 1'h1 : 1'h0;
assign op_19_V_fu_952_p3 = and_ln785_1_fu_947_p2 ? p_Val2_5_reg_1113 : select_ln340_reg_1154;
assign op_32 = ret_V_28_fu_973_p2[33] ? select_ln850_5_fu_1007_p3 : ret_V_28_fu_973_p2[32:1];
assign r_fu_720_p2 = _034_ ? 1'h1 : 1'h0;
assign ret_V_18_fu_404_p3 = ret_V_17_reg_1029[43] ? select_ln850_1_fu_398_p3 : ret_V_4_cast_reg_1034;
assign ret_V_21_fu_480_p3 = ret_V_20_reg_1051[35] ? select_ln850_2_fu_474_p3 : ret_V_8_cast_reg_1056;
assign ret_V_23_fu_620_p3 = ret_V_22_fu_572_p2[35] ? select_ln850_3_fu_612_p3 : ret_V_22_fu_572_p2[34:3];
assign ret_V_26_fu_921_p3 = ret_V_25_reg_1127[33] ? select_ln850_4_fu_914_p3 : ret_V_21_cast_reg_1132;
assign select_ln215_fu_251_p3 = op_0 ? 5'h1f : 5'h00;
assign select_ln340_fu_892_p3 = or_ln340_1_fu_886_p2 ? 4'h0 : p_Val2_5_reg_1113;
assign select_ln353_fu_340_p3 = ret_V_15_fu_284_p2[8] ? select_ln850_fu_332_p3 : { 2'h0, ret_V_15_fu_284_p2[7:3] };
assign select_ln850_1_fu_398_p3 = icmp_ln851_1_reg_1041 ? add_ln691_1_fu_393_p2 : ret_V_4_cast_reg_1034;
assign select_ln850_2_fu_474_p3 = icmp_ln851_2_reg_1063 ? add_ln691_2_fu_469_p2 : ret_V_8_cast_reg_1056;
assign select_ln850_3_fu_612_p3 = icmp_ln851_3_fu_600_p2 ? add_ln691_3_fu_606_p2 : ret_V_22_fu_572_p2[34:3];
assign select_ln850_4_fu_914_p3 = op_17[0] ? add_ln691_4_fu_909_p2 : ret_V_21_cast_reg_1132;
assign select_ln850_5_fu_1007_p3 = op_19_V_fu_952_p3[0] ? add_ln691_5_fu_1001_p2 : ret_V_28_fu_973_p2[32:1];
assign select_ln850_fu_332_p3 = icmp_ln851_fu_316_p2 ? add_ln691_fu_322_p2 : { 2'h3, ret_V_15_fu_284_p2[7:3] };
assign and_ln_fu_541_p4 = { ret_V_16_fu_513_p2[16], 15'h0000, ret_V_16_fu_513_p2[0] };
assign ap_CS_fsm_state1 = ap_CS_fsm[0];
assign ap_CS_fsm_state2 = ap_CS_fsm[1];
assign ap_CS_fsm_state3 = ap_CS_fsm[2];
assign ap_CS_fsm_state4 = ap_CS_fsm[3];
assign ap_CS_fsm_state5 = ap_CS_fsm[4];
assign ap_CS_fsm_state6 = ap_CS_fsm[5];
assign ap_CS_fsm_state7 = ap_CS_fsm[6];
assign ap_CS_fsm_state8 = ap_CS_fsm[7];
assign ap_CS_fsm_state9 = ap_CS_fsm[8];
assign ap_done = op_32_ap_vld;
assign ap_ready = op_32_ap_vld;
assign p_Result_10_fu_989_p3 = ret_V_28_fu_973_p2[33];
assign p_Result_12_fu_708_p3 = op_11_V_fu_645_p2[3];
assign p_Result_1_fu_386_p3 = ret_V_17_reg_1029[43];
assign p_Result_5_fu_700_p3 = add_ln1192_1_fu_676_p2[4];
assign p_Result_7_fu_462_p3 = ret_V_20_reg_1051[35];
assign p_Result_8_fu_588_p3 = ret_V_22_fu_572_p2[35];
assign p_Result_9_fu_899_p3 = ret_V_25_reg_1127[33];
assign p_Result_s_fu_304_p3 = ret_V_15_fu_284_p2[8];
assign p_Val2_4_fu_690_p4 = add_ln1192_1_fu_676_p2[7:4];
assign ret_V_14_cast_fu_578_p4 = ret_V_22_fu_572_p2[34:3];
assign ret_V_17_fu_360_p2[42:18] = { ret_V_17_fu_360_p2[43], ret_V_17_fu_360_p2[43], ret_V_17_fu_360_p2[43], ret_V_17_fu_360_p2[43], ret_V_17_fu_360_p2[43], ret_V_17_fu_360_p2[43], ret_V_17_fu_360_p2[43], ret_V_17_fu_360_p2[43], ret_V_17_fu_360_p2[43], ret_V_17_fu_360_p2[43], ret_V_17_fu_360_p2[43], ret_V_17_fu_360_p2[43], ret_V_17_fu_360_p2[43], ret_V_17_fu_360_p2[43], ret_V_17_fu_360_p2[43], ret_V_17_fu_360_p2[43], ret_V_17_fu_360_p2[43], ret_V_17_fu_360_p2[43], ret_V_17_fu_360_p2[43], ret_V_17_fu_360_p2[43], ret_V_17_fu_360_p2[43], ret_V_17_fu_360_p2[43], ret_V_17_fu_360_p2[43], ret_V_17_fu_360_p2[43], ret_V_17_fu_360_p2[43] };
assign ret_V_24_cast_fu_979_p4 = ret_V_28_fu_973_p2[32:1];
assign rhs_10_fu_786_p3 = { op_29_V_fu_776_p2, 1'h0 };
assign rhs_13_fu_962_p3 = { ret_V_27_reg_1159, 1'h0 };
assign rhs_1_fu_273_p3 = { ret_reg_1024, 3'h0 };
assign rhs_2_fu_501_p3 = { op_1, 6'h00 };
assign rhs_3_fu_654_p3 = { op_14, 5'h00 };
assign rhs_5_fu_425_p3 = { op_23_V_reg_1046, 3'h0 };
assign rhs_7_fu_561_p3 = { op_25_V_reg_1068, 3'h0 };
assign sext_ln1192_10_fu_969_p1 = { ret_V_27_reg_1159[31], ret_V_27_reg_1159, 1'h0 };
assign sext_ln1192_1_fu_280_p1 = { ret_reg_1024[4], ret_reg_1024, 3'h0 };
assign sext_ln1192_2_fu_356_p1 = { select_ln353_fu_340_p3[6], select_ln353_fu_340_p3[6], select_ln353_fu_340_p3[6], select_ln353_fu_340_p3[6], select_ln353_fu_340_p3[6], select_ln353_fu_340_p3[6], select_ln353_fu_340_p3[6], select_ln353_fu_340_p3[6], select_ln353_fu_340_p3[6], select_ln353_fu_340_p3[6], select_ln353_fu_340_p3[6], select_ln353_fu_340_p3[6], select_ln353_fu_340_p3[6], select_ln353_fu_340_p3[6], select_ln353_fu_340_p3[6], select_ln353_fu_340_p3[6], select_ln353_fu_340_p3[6], select_ln353_fu_340_p3[6], select_ln353_fu_340_p3[6], select_ln353_fu_340_p3[6], select_ln353_fu_340_p3[6], select_ln353_fu_340_p3[6], select_ln353_fu_340_p3[6], select_ln353_fu_340_p3[6], select_ln353_fu_340_p3[6], select_ln353_fu_340_p3[6], select_ln353_fu_340_p3, 11'h000 };
assign sext_ln1192_3_fu_662_p1 = { op_14[1], op_14[1], op_14, 5'h00 };
assign sext_ln1192_4_fu_666_p1 = { op_14[1], op_14, 5'h00 };
assign sext_ln1192_5_fu_432_p1 = { op_23_V_reg_1046[31], op_23_V_reg_1046, 3'h0 };
assign sext_ln1192_6_fu_568_p1 = { op_25_V_reg_1068[31], op_25_V_reg_1068, 3'h0 };
assign sext_ln1192_7_fu_764_p1 = { op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13 };
assign sext_ln1192_8_fu_794_p1 = { op_29_V_fu_776_p2[31], op_29_V_fu_776_p2, 1'h0 };
assign sext_ln1192_9_fu_928_p1 = { op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18 };
assign sext_ln1192_fu_269_p0 = op_5;
assign sext_ln1192_fu_269_p1 = { op_5[7], op_5 };
assign sext_ln215_fu_259_p1 = { op_2[3], op_2 };
assign sext_ln69_1_fu_632_p1 = { op_16[7], op_16[7], op_16 };
assign sext_ln69_2_fu_773_p1 = { add_ln69_reg_1088[9], add_ln69_reg_1088[9], add_ln69_reg_1088[9], add_ln69_reg_1088[9], add_ln69_reg_1088[9], add_ln69_reg_1088[9], add_ln69_reg_1088[9], add_ln69_reg_1088[9], add_ln69_reg_1088[9], add_ln69_reg_1088[9], add_ln69_reg_1088[9], add_ln69_reg_1088[9], add_ln69_reg_1088[9], add_ln69_reg_1088[9], add_ln69_reg_1088[9], add_ln69_reg_1088[9], add_ln69_reg_1088[9], add_ln69_reg_1088[9], add_ln69_reg_1088[9], add_ln69_reg_1088[9], add_ln69_reg_1088[9], add_ln69_reg_1088[9], add_ln69_reg_1088 };
assign sext_ln69_fu_411_p1 = { op_8[3], op_8[3], op_8[3], op_8[3], op_8[3], op_8[3], op_8[3], op_8[3], op_8[3], op_8[3], op_8[3], op_8[3], op_8[3], op_8[3], op_8[3], op_8[3], op_8[3], op_8[3], op_8[3], op_8[3], op_8[3], op_8[3], op_8[3], op_8[3], op_8[3], op_8[3], op_8[3], op_8[3], op_8 };
assign sext_ln703_1_fu_328_p0 = op_6;
assign sext_ln703_1_fu_328_p1 = { op_6[15], op_6[15], op_6[15], op_6[15], op_6[15], op_6[15], op_6[15], op_6[15], op_6[15], op_6[15], op_6[15], op_6[15], op_6[15], op_6[15], op_6[15], op_6[15], op_6[15], op_6[15], op_6[15], op_6[15], op_6[15], op_6[15], op_6[15], op_6[15], op_6[15], op_6[15], op_6[15], op_6[15], op_6 };
assign sext_ln703_2_fu_650_p1 = { op_11_V_fu_645_p2[7], op_11_V_fu_645_p2 };
assign sext_ln703_3_fu_421_p0 = op_9;
assign sext_ln703_3_fu_421_p1 = { op_9[3], op_9[3], op_9[3], op_9[3], op_9[3], op_9[3], op_9[3], op_9[3], op_9[3], op_9[3], op_9[3], op_9[3], op_9[3], op_9[3], op_9[3], op_9[3], op_9[3], op_9[3], op_9[3], op_9[3], op_9[3], op_9[3], op_9[3], op_9[3], op_9[3], op_9[3], op_9[3], op_9[3], op_9[3], op_9[3], op_9[3], op_9[3], op_9 };
assign sext_ln703_4_fu_557_p0 = op_12;
assign sext_ln703_4_fu_557_p1 = { op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12 };
assign sext_ln703_5_fu_782_p0 = op_17;
assign sext_ln703_5_fu_782_p1 = { op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17 };
assign sext_ln703_6_fu_958_p1 = { op_19_V_fu_952_p3[3], op_19_V_fu_952_p3[3], op_19_V_fu_952_p3[3], op_19_V_fu_952_p3[3], op_19_V_fu_952_p3[3], op_19_V_fu_952_p3[3], op_19_V_fu_952_p3[3], op_19_V_fu_952_p3[3], op_19_V_fu_952_p3[3], op_19_V_fu_952_p3[3], op_19_V_fu_952_p3[3], op_19_V_fu_952_p3[3], op_19_V_fu_952_p3[3], op_19_V_fu_952_p3[3], op_19_V_fu_952_p3[3], op_19_V_fu_952_p3[3], op_19_V_fu_952_p3[3], op_19_V_fu_952_p3[3], op_19_V_fu_952_p3[3], op_19_V_fu_952_p3[3], op_19_V_fu_952_p3[3], op_19_V_fu_952_p3[3], op_19_V_fu_952_p3[3], op_19_V_fu_952_p3[3], op_19_V_fu_952_p3[3], op_19_V_fu_952_p3[3], op_19_V_fu_952_p3[3], op_19_V_fu_952_p3[3], op_19_V_fu_952_p3[3], op_19_V_fu_952_p3[3], op_19_V_fu_952_p3 };
assign sext_ln703_fu_497_p1 = { op_4[15], op_4 };
assign sext_ln850_fu_300_p1 = { ret_V_15_fu_284_p2[8], ret_V_15_fu_284_p2[8:3] };
assign tmp_1_fu_290_p4 = ret_V_15_fu_284_p2[8:3];
assign tmp_2_fu_348_p3 = { select_ln353_fu_340_p3, 11'h000 };
assign tmp_fu_529_p3 = ret_V_16_fu_513_p2[16];
assign trunc_ln410_fu_537_p1 = ret_V_16_fu_513_p2[0];
assign trunc_ln718_fu_716_p1 = op_11_V_fu_645_p2[2:0];
assign trunc_ln851_1_fu_376_p0 = op_6;
assign trunc_ln851_1_fu_376_p1 = op_6[10:0];
assign trunc_ln851_2_fu_452_p0 = op_9;
assign trunc_ln851_2_fu_452_p1 = op_9[2:0];
assign trunc_ln851_3_fu_596_p0 = op_12;
assign trunc_ln851_3_fu_596_p1 = op_12[2:0];
assign trunc_ln851_4_fu_906_p0 = op_17;
assign trunc_ln851_4_fu_906_p1 = op_17[0];
assign trunc_ln851_5_fu_997_p1 = op_19_V_fu_952_p3[0];
assign trunc_ln851_fu_312_p0 = op_5;
assign trunc_ln851_fu_312_p1 = op_5[2:0];
assign zext_ln1193_fu_509_p1 = { 7'h00, op_1, 6'h00 };
assign zext_ln415_1_fu_746_p1 = { 3'h0, and_ln412_fu_740_p2 };
assign zext_ln415_fu_642_p1 = { 7'h00, icmp_ln410_reg_1078 };
assign zext_ln69_1_fu_628_p1 = { 2'h0, op_15 };
assign zext_ln69_fu_487_p1 = { 24'h000000, op_10 };
endmodule


// Product machine:
module top_A_times_top_B (ap_start, op_0, op_1, op_10, op_12, op_13, op_14, op_15, op_16, op_17, op_18, op_2, op_4, op_5, op_6, op_8, op_9, ap_clk, unsafe_signal);
input ap_start;
input op_0;
input [3:0] op_1;
input [7:0] op_10;
input [3:0] op_12;
input [7:0] op_13;
input [1:0] op_14;
input [7:0] op_15;
input [7:0] op_16;
input [3:0] op_17;
input [1:0] op_18;
input [3:0] op_2;
input [15:0] op_4;
input [7:0] op_5;
input [15:0] op_6;
input [3:0] op_8;
input [3:0] op_9;
input ap_clk;
output unsafe_signal;
reg _setup;
initial _setup = 1'b0;
always @ (posedge ap_clk) _setup <= 1'b1;
reg ap_start_internal;
always @ (posedge ap_clk) if (!_setup) ap_start_internal <= ap_start;
reg op_0_internal;
always @ (posedge ap_clk) if (!_setup) op_0_internal <= op_0;
reg [3:0] op_1_internal;
always @ (posedge ap_clk) if (!_setup) op_1_internal <= op_1;
reg [7:0] op_10_internal;
always @ (posedge ap_clk) if (!_setup) op_10_internal <= op_10;
reg [3:0] op_12_internal;
always @ (posedge ap_clk) if (!_setup) op_12_internal <= op_12;
reg [7:0] op_13_internal;
always @ (posedge ap_clk) if (!_setup) op_13_internal <= op_13;
reg [1:0] op_14_internal;
always @ (posedge ap_clk) if (!_setup) op_14_internal <= op_14;
reg [7:0] op_15_internal;
always @ (posedge ap_clk) if (!_setup) op_15_internal <= op_15;
reg [7:0] op_16_internal;
always @ (posedge ap_clk) if (!_setup) op_16_internal <= op_16;
reg [3:0] op_17_internal;
always @ (posedge ap_clk) if (!_setup) op_17_internal <= op_17;
reg [1:0] op_18_internal;
always @ (posedge ap_clk) if (!_setup) op_18_internal <= op_18;
reg [3:0] op_2_internal;
always @ (posedge ap_clk) if (!_setup) op_2_internal <= op_2;
reg [15:0] op_4_internal;
always @ (posedge ap_clk) if (!_setup) op_4_internal <= op_4;
reg [7:0] op_5_internal;
always @ (posedge ap_clk) if (!_setup) op_5_internal <= op_5;
reg [15:0] op_6_internal;
always @ (posedge ap_clk) if (!_setup) op_6_internal <= op_6;
reg [3:0] op_8_internal;
always @ (posedge ap_clk) if (!_setup) op_8_internal <= op_8;
reg [3:0] op_9_internal;
always @ (posedge ap_clk) if (!_setup) op_9_internal <= op_9;
wire ap_done_A;
wire ap_done_B;
wire ap_done_eq;
assign ap_done_eq = ap_done_A == ap_done_B;
wire ap_idle_A;
wire ap_idle_B;
wire ap_idle_eq;
assign ap_idle_eq = ap_idle_A == ap_idle_B;
wire ap_ready_A;
wire ap_ready_B;
wire ap_ready_eq;
assign ap_ready_eq = ap_ready_A == ap_ready_B;
wire [31:0] op_32_A;
wire [31:0] op_32_B;
wire op_32_eq;
assign op_32_eq = op_32_A == op_32_B;
wire op_32_ap_vld_A;
wire op_32_ap_vld_B;
wire clk_enable_A;
wire clk_enable_B;
assign clk_enable_A = _setup & (~op_32_ap_vld_A | op_32_ap_vld_B);
assign clk_enable_B = _setup;
wire divergent;
assign divergent = ~(ap_done_eq & ap_idle_eq & ap_ready_eq & op_32_eq);
assign unsafe_signal = op_32_ap_vld_A & op_32_ap_vld_B & divergent;
top_A instance_A (
    .ap_clk(ap_clk),
    .clk_enable(clk_enable_A),
    .ap_start(ap_start_internal),
    .op_0(op_0_internal),
    .op_1(op_1_internal),
    .op_10(op_10_internal),
    .op_12(op_12_internal),
    .op_13(op_13_internal),
    .op_14(op_14_internal),
    .op_15(op_15_internal),
    .op_16(op_16_internal),
    .op_17(op_17_internal),
    .op_18(op_18_internal),
    .op_2(op_2_internal),
    .op_4(op_4_internal),
    .op_5(op_5_internal),
    .op_6(op_6_internal),
    .op_8(op_8_internal),
    .op_9(op_9_internal),
    .ap_done(ap_done_A),
    .ap_idle(ap_idle_A),
    .ap_ready(ap_ready_A),
    .op_32(op_32_A),
    .op_32_ap_vld(op_32_ap_vld_A)
);
top_B instance_B (
    .ap_clk(ap_clk),
    .clk_enable(clk_enable_B),
    .ap_start(ap_start_internal),
    .op_0(op_0_internal),
    .op_1(op_1_internal),
    .op_10(op_10_internal),
    .op_12(op_12_internal),
    .op_13(op_13_internal),
    .op_14(op_14_internal),
    .op_15(op_15_internal),
    .op_16(op_16_internal),
    .op_17(op_17_internal),
    .op_18(op_18_internal),
    .op_2(op_2_internal),
    .op_4(op_4_internal),
    .op_5(op_5_internal),
    .op_6(op_6_internal),
    .op_8(op_8_internal),
    .op_9(op_9_internal),
    .ap_done(ap_done_B),
    .ap_idle(ap_idle_B),
    .ap_ready(ap_ready_B),
    .op_32(op_32_B),
    .op_32_ap_vld(op_32_ap_vld_B)
);
endmodule
