// Processed by function `construct_kairos` in `verilog_tricks.py`.
// Machine A:
// Processed by function `add_clk_enable_signal` in `verilog_tricks.py`.
// Processed by function `remove_reset_signal` in `verilog_tricks.py`.
module top_A (
  ap_clk,
  ap_start,
  ap_done,
  ap_idle,
  ap_ready,
  op_0,
  op_1,
  op_2,
  op_3,
  op_4,
  op_6,
  op_10,
  op_11,
  op_12,
  op_30,
  op_30_ap_vld,
clk_enable
);
input clk_enable;


input ap_clk;
wire ap_rst;
assign ap_rst = op_30_ap_vld;
input ap_start;
input [3:0] op_0;
input [7:0] op_1;
input [7:0] op_10;
input [7:0] op_11;
input [7:0] op_12;
input [7:0] op_2;
input [31:0] op_3;
input [3:0] op_4;
input [1:0] op_6;
output ap_done;
output ap_idle;
output ap_ready;
output [31:0] op_30;
output op_30_ap_vld;


reg [5:0] \add_11s_11s_11_2_1_U2.top_add_11s_11s_11_2_1_Adder_1_U.ain_s1 ;
reg [5:0] \add_11s_11s_11_2_1_U2.top_add_11s_11s_11_2_1_Adder_1_U.bin_s1 ;
reg \add_11s_11s_11_2_1_U2.top_add_11s_11s_11_2_1_Adder_1_U.carry_s1 ;
reg [4:0] \add_11s_11s_11_2_1_U2.top_add_11s_11s_11_2_1_Adder_1_U.sum_s1 ;
reg \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.ain_s1 ;
reg \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.bin_s1 ;
reg \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.carry_s1 ;
reg \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.sum_s1 ;
reg \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_0_U.ain_s1 ;
reg \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_0_U.bin_s1 ;
reg \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_0_U.carry_s1 ;
reg \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_0_U.sum_s1 ;
reg [16:0] \add_33ns_33s_33_2_1_U5.top_add_33ns_33s_33_2_1_Adder_3_U.ain_s1 ;
reg [16:0] \add_33ns_33s_33_2_1_U5.top_add_33ns_33s_33_2_1_Adder_3_U.bin_s1 ;
reg \add_33ns_33s_33_2_1_U5.top_add_33ns_33s_33_2_1_Adder_3_U.carry_s1 ;
reg [15:0] \add_33ns_33s_33_2_1_U5.top_add_33ns_33s_33_2_1_Adder_3_U.sum_s1 ;
reg [1:0] \add_3ns_3ns_3_2_1_U13.top_add_3ns_3ns_3_2_1_Adder_9_U.ain_s1 ;
reg [1:0] \add_3ns_3ns_3_2_1_U13.top_add_3ns_3ns_3_2_1_Adder_9_U.bin_s1 ;
reg \add_3ns_3ns_3_2_1_U13.top_add_3ns_3ns_3_2_1_Adder_9_U.carry_s1 ;
reg \add_3ns_3ns_3_2_1_U13.top_add_3ns_3ns_3_2_1_Adder_9_U.sum_s1 ;
reg [1:0] \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.ain_s1 ;
reg [1:0] \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.bin_s1 ;
reg \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.carry_s1 ;
reg [1:0] \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.sum_s1 ;
reg [1:0] \add_4s_4s_4_2_1_U16.top_add_4s_4s_4_2_1_Adder_12_U.ain_s1 ;
reg [1:0] \add_4s_4s_4_2_1_U16.top_add_4s_4s_4_2_1_Adder_12_U.bin_s1 ;
reg \add_4s_4s_4_2_1_U16.top_add_4s_4s_4_2_1_Adder_12_U.carry_s1 ;
reg [1:0] \add_4s_4s_4_2_1_U16.top_add_4s_4s_4_2_1_Adder_12_U.sum_s1 ;
reg [2:0] \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_5_U.ain_s1 ;
reg [2:0] \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_5_U.bin_s1 ;
reg \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_5_U.carry_s1 ;
reg [1:0] \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_5_U.sum_s1 ;
reg [2:0] \add_6ns_6s_6_2_1_U15.top_add_6ns_6s_6_2_1_Adder_11_U.ain_s1 ;
reg [2:0] \add_6ns_6s_6_2_1_U15.top_add_6ns_6s_6_2_1_Adder_11_U.bin_s1 ;
reg \add_6ns_6s_6_2_1_U15.top_add_6ns_6s_6_2_1_Adder_11_U.carry_s1 ;
reg [2:0] \add_6ns_6s_6_2_1_U15.top_add_6ns_6s_6_2_1_Adder_11_U.sum_s1 ;
reg [2:0] \add_6s_6ns_6_2_1_U18.top_add_6s_6ns_6_2_1_Adder_14_U.ain_s1 ;
reg [2:0] \add_6s_6ns_6_2_1_U18.top_add_6s_6ns_6_2_1_Adder_14_U.bin_s1 ;
reg \add_6s_6ns_6_2_1_U18.top_add_6s_6ns_6_2_1_Adder_14_U.carry_s1 ;
reg [2:0] \add_6s_6ns_6_2_1_U18.top_add_6s_6ns_6_2_1_Adder_14_U.sum_s1 ;
reg [3:0] \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_8_U.ain_s1 ;
reg [3:0] \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_8_U.bin_s1 ;
reg \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_8_U.carry_s1 ;
reg [2:0] \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_8_U.sum_s1 ;
reg [3:0] \add_7s_7s_7_2_1_U10.top_add_7s_7s_7_2_1_Adder_6_U.ain_s1 ;
reg [3:0] \add_7s_7s_7_2_1_U10.top_add_7s_7s_7_2_1_Adder_6_U.bin_s1 ;
reg \add_7s_7s_7_2_1_U10.top_add_7s_7s_7_2_1_Adder_6_U.carry_s1 ;
reg [2:0] \add_7s_7s_7_2_1_U10.top_add_7s_7s_7_2_1_Adder_6_U.sum_s1 ;
reg [4:0] \add_9ns_9ns_9_2_1_U17.top_add_9ns_9ns_9_2_1_Adder_13_U.ain_s1 ;
reg [4:0] \add_9ns_9ns_9_2_1_U17.top_add_9ns_9ns_9_2_1_Adder_13_U.bin_s1 ;
reg \add_9ns_9ns_9_2_1_U17.top_add_9ns_9ns_9_2_1_Adder_13_U.carry_s1 ;
reg [3:0] \add_9ns_9ns_9_2_1_U17.top_add_9ns_9ns_9_2_1_Adder_13_U.sum_s1 ;
reg [4:0] \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_15_U.ain_s1 ;
reg [4:0] \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_15_U.bin_s1 ;
reg \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_15_U.carry_s1 ;
reg [3:0] \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_15_U.sum_s1 ;
reg [4:0] \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_10_U.ain_s1 ;
reg [4:0] \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_10_U.bin_s1 ;
reg \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_10_U.carry_s1 ;
reg [3:0] \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_10_U.sum_s1 ;
reg [6:0] add_ln691_reg_897;
reg [8:0] add_ln69_1_reg_977;
reg [5:0] add_ln69_2_reg_962;
reg [3:0] add_ln69_3_reg_967;
reg [5:0] add_ln69_4_reg_982;
reg [8:0] add_ln69_reg_957;
reg [18:0] ap_CS_fsm = 19'h00001;
reg icmp_ln851_1_reg_736;
reg icmp_ln851_2_reg_670;
reg icmp_ln851_3_reg_882;
reg icmp_ln851_reg_701;
reg [31:0] \lshr_32ns_32s_32_7_1_U9.din1_cast_array[0] ;
reg [31:0] \lshr_32ns_32s_32_7_1_U9.din1_cast_array[1] ;
reg [31:0] \lshr_32ns_32s_32_7_1_U9.din1_cast_array[2] ;
reg [31:0] \lshr_32ns_32s_32_7_1_U9.din1_cast_array[3] ;
reg [31:0] \lshr_32ns_32s_32_7_1_U9.din1_cast_array[4] ;
reg [31:0] \lshr_32ns_32s_32_7_1_U9.din1_cast_array[5] ;
reg [31:0] \lshr_32ns_32s_32_7_1_U9.dout_array[0] ;
reg [31:0] \lshr_32ns_32s_32_7_1_U9.dout_array[1] ;
reg [31:0] \lshr_32ns_32s_32_7_1_U9.dout_array[2] ;
reg [31:0] \lshr_32ns_32s_32_7_1_U9.dout_array[3] ;
reg [31:0] \lshr_32ns_32s_32_7_1_U9.dout_array[4] ;
reg [31:0] \lshr_32ns_32s_32_7_1_U9.dout_array[5] ;
reg [3:0] op_15_V_reg_907;
reg p_Result_1_reg_730;
reg [2:0] ret_V_13_reg_863;
reg [2:0] ret_V_14_reg_902;
reg [2:0] ret_V_15_reg_917;
reg [3:0] ret_V_16_reg_792;
reg [10:0] ret_V_18_reg_711;
reg [1:0] ret_V_19_reg_802;
reg [32:0] ret_V_20_reg_770;
reg ret_V_21_reg_807;
reg [6:0] ret_V_22_reg_848;
reg [6:0] ret_V_23_reg_912;
reg [8:0] ret_V_24_reg_858;
reg [3:0] ret_V_25_reg_813;
reg [4:0] ret_V_2_reg_797;
reg [3:0] ret_V_3_cast5_reg_758;
reg [1:0] ret_V_3_cast_reg_723;
reg [1:0] ret_V_3_reg_765;
reg [1:0] ret_V_7_reg_663;
reg [1:0] ret_V_8_reg_675;
reg [1:0] ret_V_9_reg_680;
reg [4:0] ret_V_reg_716;
reg [8:0] select_ln69_reg_952;
reg [8:0] select_ln703_reg_823;
reg [4:0] select_ln850_7_reg_818;
reg [6:0] sext_ln850_reg_875;
reg [31:0] \shl_32ns_32s_32_7_1_U8.din1_cast_array[0] ;
reg [31:0] \shl_32ns_32s_32_7_1_U8.din1_cast_array[1] ;
reg [31:0] \shl_32ns_32s_32_7_1_U8.din1_cast_array[2] ;
reg [31:0] \shl_32ns_32s_32_7_1_U8.din1_cast_array[3] ;
reg [31:0] \shl_32ns_32s_32_7_1_U8.din1_cast_array[4] ;
reg [31:0] \shl_32ns_32s_32_7_1_U8.din1_cast_array[5] ;
reg [31:0] \shl_32ns_32s_32_7_1_U8.dout_array[0] ;
reg [31:0] \shl_32ns_32s_32_7_1_U8.dout_array[1] ;
reg [31:0] \shl_32ns_32s_32_7_1_U8.dout_array[2] ;
reg [31:0] \shl_32ns_32s_32_7_1_U8.dout_array[3] ;
reg [31:0] \shl_32ns_32s_32_7_1_U8.dout_array[4] ;
reg [31:0] \shl_32ns_32s_32_7_1_U8.dout_array[5] ;
reg [1:0] \sub_3ns_3s_3_2_1_U3.top_sub_3ns_3s_3_2_1_Adder_2_U.ain_s1 ;
reg [1:0] \sub_3ns_3s_3_2_1_U3.top_sub_3ns_3s_3_2_1_Adder_2_U.bin_s1 ;
reg \sub_3ns_3s_3_2_1_U3.top_sub_3ns_3s_3_2_1_Adder_2_U.carry_s1 ;
reg \sub_3ns_3s_3_2_1_U3.top_sub_3ns_3s_3_2_1_Adder_2_U.sum_s1 ;
reg [4:0] \sub_9ns_9s_9_2_1_U11.top_sub_9ns_9s_9_2_1_Adder_7_U.ain_s1 ;
reg [4:0] \sub_9ns_9s_9_2_1_U11.top_sub_9ns_9s_9_2_1_Adder_7_U.bin_s1 ;
reg \sub_9ns_9s_9_2_1_U11.top_sub_9ns_9s_9_2_1_Adder_7_U.carry_s1 ;
reg [3:0] \sub_9ns_9s_9_2_1_U11.top_sub_9ns_9s_9_2_1_Adder_7_U.sum_s1 ;
reg [2:0] sub_ln1497_reg_753;
reg [5:0] tmp_1_reg_853;
reg tmp_4_reg_686;
reg [3:0] trunc_ln1497_1_reg_892;
reg [3:0] trunc_ln1497_reg_887;
reg [5:0] trunc_ln851_4_reg_870;
wire [6:0] _000_;
wire [8:0] _001_;
wire [5:0] _002_;
wire [3:0] _003_;
wire [5:0] _004_;
wire [8:0] _005_;
wire [18:0] _006_;
wire _007_;
wire _008_;
wire _009_;
wire _010_;
wire [3:0] _011_;
wire _012_;
wire [2:0] _013_;
wire [2:0] _014_;
wire [2:0] _015_;
wire [3:0] _016_;
wire [10:0] _017_;
wire [1:0] _018_;
wire [32:0] _019_;
wire _020_;
wire [6:0] _021_;
wire [6:0] _022_;
wire [8:0] _023_;
wire [3:0] _024_;
wire [4:0] _025_;
wire [3:0] _026_;
wire [1:0] _027_;
wire [1:0] _028_;
wire [1:0] _029_;
wire [1:0] _030_;
wire [1:0] _031_;
wire [4:0] _032_;
wire [1:0] _033_;
wire [2:0] _034_;
wire [4:0] _035_;
wire [6:0] _036_;
wire [2:0] _037_;
wire [5:0] _038_;
wire _039_;
wire [3:0] _040_;
wire [3:0] _041_;
wire [5:0] _042_;
wire [1:0] _043_;
wire _044_;
wire _045_;
wire _046_;
wire _047_;
wire _048_;
wire _049_;
wire _050_;
wire _051_;
wire _052_;
wire _053_;
wire _054_;
wire _055_;
wire _056_;
wire [5:0] _057_;
wire [5:0] _058_;
wire _059_;
wire [4:0] _060_;
wire [5:0] _061_;
wire [6:0] _062_;
wire _063_;
wire _064_;
wire _065_;
wire _066_;
wire [1:0] _067_;
wire [1:0] _068_;
wire _069_;
wire _070_;
wire _071_;
wire _072_;
wire [1:0] _073_;
wire [1:0] _074_;
wire [16:0] _075_;
wire [16:0] _076_;
wire _077_;
wire [15:0] _078_;
wire [16:0] _079_;
wire [17:0] _080_;
wire [1:0] _081_;
wire [1:0] _082_;
wire _083_;
wire _084_;
wire [1:0] _085_;
wire [2:0] _086_;
wire [1:0] _087_;
wire [1:0] _088_;
wire _089_;
wire [1:0] _090_;
wire [2:0] _091_;
wire [2:0] _092_;
wire [1:0] _093_;
wire [1:0] _094_;
wire _095_;
wire [1:0] _096_;
wire [2:0] _097_;
wire [2:0] _098_;
wire [2:0] _099_;
wire [2:0] _100_;
wire _101_;
wire [1:0] _102_;
wire [2:0] _103_;
wire [3:0] _104_;
wire [2:0] _105_;
wire [2:0] _106_;
wire _107_;
wire [2:0] _108_;
wire [3:0] _109_;
wire [3:0] _110_;
wire [2:0] _111_;
wire [2:0] _112_;
wire _113_;
wire [2:0] _114_;
wire [3:0] _115_;
wire [3:0] _116_;
wire [3:0] _117_;
wire [3:0] _118_;
wire _119_;
wire [2:0] _120_;
wire [3:0] _121_;
wire [4:0] _122_;
wire [3:0] _123_;
wire [3:0] _124_;
wire _125_;
wire [2:0] _126_;
wire [3:0] _127_;
wire [4:0] _128_;
wire [4:0] _129_;
wire [4:0] _130_;
wire _131_;
wire [3:0] _132_;
wire [4:0] _133_;
wire [5:0] _134_;
wire [4:0] _135_;
wire [4:0] _136_;
wire _137_;
wire [3:0] _138_;
wire [4:0] _139_;
wire [5:0] _140_;
wire [4:0] _141_;
wire [4:0] _142_;
wire _143_;
wire [3:0] _144_;
wire [4:0] _145_;
wire [5:0] _146_;
wire [31:0] _147_;
wire [31:0] _148_;
wire [31:0] _149_;
wire [31:0] _150_;
wire [31:0] _151_;
wire [31:0] _152_;
wire [31:0] _153_;
wire [31:0] _154_;
wire [31:0] _155_;
wire [31:0] _156_;
wire [31:0] _157_;
wire [31:0] _158_;
wire [31:0] _159_;
wire [31:0] _160_;
wire [31:0] _161_;
wire [31:0] _162_;
wire [31:0] _163_;
wire [31:0] _164_;
wire [31:0] _165_;
wire [31:0] _166_;
wire [31:0] _167_;
wire [31:0] _168_;
wire [31:0] _169_;
wire [31:0] _170_;
wire [31:0] _171_;
wire [31:0] _172_;
wire [31:0] _173_;
wire [31:0] _174_;
wire [31:0] _175_;
wire [31:0] _176_;
wire [31:0] _177_;
wire [31:0] _178_;
wire [31:0] _179_;
wire [31:0] _180_;
wire [31:0] _181_;
wire [31:0] _182_;
wire [31:0] _183_;
wire [31:0] _184_;
wire [31:0] _185_;
wire [31:0] _186_;
wire [31:0] _187_;
wire [31:0] _188_;
wire [31:0] _189_;
wire [31:0] _190_;
wire [31:0] _191_;
wire [31:0] _192_;
wire [31:0] _193_;
wire [31:0] _194_;
wire [31:0] _195_;
wire [31:0] _196_;
wire [31:0] _197_;
wire [31:0] _198_;
wire [31:0] _199_;
wire [31:0] _200_;
wire [31:0] _201_;
wire [31:0] _202_;
wire [31:0] _203_;
wire [31:0] _204_;
wire [31:0] _205_;
wire [31:0] _206_;
wire [1:0] _207_;
wire [1:0] _208_;
wire _209_;
wire _210_;
wire [1:0] _211_;
wire [2:0] _212_;
wire [4:0] _213_;
wire [4:0] _214_;
wire _215_;
wire [3:0] _216_;
wire [4:0] _217_;
wire [5:0] _218_;
wire _219_;
wire _220_;
wire _221_;
wire _222_;
wire _223_;
wire _224_;
wire _225_;
wire _226_;
wire _227_;
wire _228_;
wire _229_;
wire _230_;
wire _231_;
wire _232_;
wire _233_;
wire _234_;
wire _235_;
wire _236_;
wire _237_;
wire \add_11s_11s_11_2_1_U2.ce ;
wire \add_11s_11s_11_2_1_U2.clk ;
wire [10:0] \add_11s_11s_11_2_1_U2.din0 ;
wire [10:0] \add_11s_11s_11_2_1_U2.din1 ;
wire [10:0] \add_11s_11s_11_2_1_U2.dout ;
wire \add_11s_11s_11_2_1_U2.reset ;
wire [10:0] \add_11s_11s_11_2_1_U2.top_add_11s_11s_11_2_1_Adder_1_U.a ;
wire [10:0] \add_11s_11s_11_2_1_U2.top_add_11s_11s_11_2_1_Adder_1_U.ain_s0 ;
wire [10:0] \add_11s_11s_11_2_1_U2.top_add_11s_11s_11_2_1_Adder_1_U.b ;
wire [10:0] \add_11s_11s_11_2_1_U2.top_add_11s_11s_11_2_1_Adder_1_U.bin_s0 ;
wire \add_11s_11s_11_2_1_U2.top_add_11s_11s_11_2_1_Adder_1_U.ce ;
wire \add_11s_11s_11_2_1_U2.top_add_11s_11s_11_2_1_Adder_1_U.clk ;
wire \add_11s_11s_11_2_1_U2.top_add_11s_11s_11_2_1_Adder_1_U.facout_s1 ;
wire \add_11s_11s_11_2_1_U2.top_add_11s_11s_11_2_1_Adder_1_U.facout_s2 ;
wire [4:0] \add_11s_11s_11_2_1_U2.top_add_11s_11s_11_2_1_Adder_1_U.fas_s1 ;
wire [5:0] \add_11s_11s_11_2_1_U2.top_add_11s_11s_11_2_1_Adder_1_U.fas_s2 ;
wire \add_11s_11s_11_2_1_U2.top_add_11s_11s_11_2_1_Adder_1_U.reset ;
wire [10:0] \add_11s_11s_11_2_1_U2.top_add_11s_11s_11_2_1_Adder_1_U.s ;
wire [4:0] \add_11s_11s_11_2_1_U2.top_add_11s_11s_11_2_1_Adder_1_U.u1.a ;
wire [4:0] \add_11s_11s_11_2_1_U2.top_add_11s_11s_11_2_1_Adder_1_U.u1.b ;
wire \add_11s_11s_11_2_1_U2.top_add_11s_11s_11_2_1_Adder_1_U.u1.cin ;
wire \add_11s_11s_11_2_1_U2.top_add_11s_11s_11_2_1_Adder_1_U.u1.cout ;
wire [4:0] \add_11s_11s_11_2_1_U2.top_add_11s_11s_11_2_1_Adder_1_U.u1.s ;
wire [5:0] \add_11s_11s_11_2_1_U2.top_add_11s_11s_11_2_1_Adder_1_U.u2.a ;
wire [5:0] \add_11s_11s_11_2_1_U2.top_add_11s_11s_11_2_1_Adder_1_U.u2.b ;
wire \add_11s_11s_11_2_1_U2.top_add_11s_11s_11_2_1_Adder_1_U.u2.cin ;
wire \add_11s_11s_11_2_1_U2.top_add_11s_11s_11_2_1_Adder_1_U.u2.cout ;
wire [5:0] \add_11s_11s_11_2_1_U2.top_add_11s_11s_11_2_1_Adder_1_U.u2.s ;
wire \add_2ns_2ns_2_2_1_U1.ce ;
wire \add_2ns_2ns_2_2_1_U1.clk ;
wire [1:0] \add_2ns_2ns_2_2_1_U1.din0 ;
wire [1:0] \add_2ns_2ns_2_2_1_U1.din1 ;
wire [1:0] \add_2ns_2ns_2_2_1_U1.dout ;
wire \add_2ns_2ns_2_2_1_U1.reset ;
wire [1:0] \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.a ;
wire [1:0] \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.ain_s0 ;
wire [1:0] \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.b ;
wire [1:0] \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.bin_s0 ;
wire \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.ce ;
wire \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.clk ;
wire \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.facout_s1 ;
wire \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.facout_s2 ;
wire \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.fas_s1 ;
wire \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.fas_s2 ;
wire \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.reset ;
wire [1:0] \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.s ;
wire \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.u1.a ;
wire \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.u1.b ;
wire \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.u1.cin ;
wire \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.u1.cout ;
wire \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.u1.s ;
wire \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.u2.a ;
wire \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.u2.b ;
wire \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.u2.cin ;
wire \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.u2.cout ;
wire \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.u2.s ;
wire \add_2ns_2ns_2_2_1_U4.ce ;
wire \add_2ns_2ns_2_2_1_U4.clk ;
wire [1:0] \add_2ns_2ns_2_2_1_U4.din0 ;
wire [1:0] \add_2ns_2ns_2_2_1_U4.din1 ;
wire [1:0] \add_2ns_2ns_2_2_1_U4.dout ;
wire \add_2ns_2ns_2_2_1_U4.reset ;
wire [1:0] \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_0_U.a ;
wire [1:0] \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_0_U.ain_s0 ;
wire [1:0] \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_0_U.b ;
wire [1:0] \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_0_U.bin_s0 ;
wire \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_0_U.ce ;
wire \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_0_U.clk ;
wire \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_0_U.facout_s1 ;
wire \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_0_U.facout_s2 ;
wire \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_0_U.fas_s1 ;
wire \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_0_U.fas_s2 ;
wire \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_0_U.reset ;
wire [1:0] \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_0_U.s ;
wire \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_0_U.u1.a ;
wire \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_0_U.u1.b ;
wire \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_0_U.u1.cin ;
wire \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_0_U.u1.cout ;
wire \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_0_U.u1.s ;
wire \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_0_U.u2.a ;
wire \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_0_U.u2.b ;
wire \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_0_U.u2.cin ;
wire \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_0_U.u2.cout ;
wire \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_0_U.u2.s ;
wire \add_33ns_33s_33_2_1_U5.ce ;
wire \add_33ns_33s_33_2_1_U5.clk ;
wire [32:0] \add_33ns_33s_33_2_1_U5.din0 ;
wire [32:0] \add_33ns_33s_33_2_1_U5.din1 ;
wire [32:0] \add_33ns_33s_33_2_1_U5.dout ;
wire \add_33ns_33s_33_2_1_U5.reset ;
wire [32:0] \add_33ns_33s_33_2_1_U5.top_add_33ns_33s_33_2_1_Adder_3_U.a ;
wire [32:0] \add_33ns_33s_33_2_1_U5.top_add_33ns_33s_33_2_1_Adder_3_U.ain_s0 ;
wire [32:0] \add_33ns_33s_33_2_1_U5.top_add_33ns_33s_33_2_1_Adder_3_U.b ;
wire [32:0] \add_33ns_33s_33_2_1_U5.top_add_33ns_33s_33_2_1_Adder_3_U.bin_s0 ;
wire \add_33ns_33s_33_2_1_U5.top_add_33ns_33s_33_2_1_Adder_3_U.ce ;
wire \add_33ns_33s_33_2_1_U5.top_add_33ns_33s_33_2_1_Adder_3_U.clk ;
wire \add_33ns_33s_33_2_1_U5.top_add_33ns_33s_33_2_1_Adder_3_U.facout_s1 ;
wire \add_33ns_33s_33_2_1_U5.top_add_33ns_33s_33_2_1_Adder_3_U.facout_s2 ;
wire [15:0] \add_33ns_33s_33_2_1_U5.top_add_33ns_33s_33_2_1_Adder_3_U.fas_s1 ;
wire [16:0] \add_33ns_33s_33_2_1_U5.top_add_33ns_33s_33_2_1_Adder_3_U.fas_s2 ;
wire \add_33ns_33s_33_2_1_U5.top_add_33ns_33s_33_2_1_Adder_3_U.reset ;
wire [32:0] \add_33ns_33s_33_2_1_U5.top_add_33ns_33s_33_2_1_Adder_3_U.s ;
wire [15:0] \add_33ns_33s_33_2_1_U5.top_add_33ns_33s_33_2_1_Adder_3_U.u1.a ;
wire [15:0] \add_33ns_33s_33_2_1_U5.top_add_33ns_33s_33_2_1_Adder_3_U.u1.b ;
wire \add_33ns_33s_33_2_1_U5.top_add_33ns_33s_33_2_1_Adder_3_U.u1.cin ;
wire \add_33ns_33s_33_2_1_U5.top_add_33ns_33s_33_2_1_Adder_3_U.u1.cout ;
wire [15:0] \add_33ns_33s_33_2_1_U5.top_add_33ns_33s_33_2_1_Adder_3_U.u1.s ;
wire [16:0] \add_33ns_33s_33_2_1_U5.top_add_33ns_33s_33_2_1_Adder_3_U.u2.a ;
wire [16:0] \add_33ns_33s_33_2_1_U5.top_add_33ns_33s_33_2_1_Adder_3_U.u2.b ;
wire \add_33ns_33s_33_2_1_U5.top_add_33ns_33s_33_2_1_Adder_3_U.u2.cin ;
wire \add_33ns_33s_33_2_1_U5.top_add_33ns_33s_33_2_1_Adder_3_U.u2.cout ;
wire [16:0] \add_33ns_33s_33_2_1_U5.top_add_33ns_33s_33_2_1_Adder_3_U.u2.s ;
wire \add_3ns_3ns_3_2_1_U13.ce ;
wire \add_3ns_3ns_3_2_1_U13.clk ;
wire [2:0] \add_3ns_3ns_3_2_1_U13.din0 ;
wire [2:0] \add_3ns_3ns_3_2_1_U13.din1 ;
wire [2:0] \add_3ns_3ns_3_2_1_U13.dout ;
wire \add_3ns_3ns_3_2_1_U13.reset ;
wire [2:0] \add_3ns_3ns_3_2_1_U13.top_add_3ns_3ns_3_2_1_Adder_9_U.a ;
wire [2:0] \add_3ns_3ns_3_2_1_U13.top_add_3ns_3ns_3_2_1_Adder_9_U.ain_s0 ;
wire [2:0] \add_3ns_3ns_3_2_1_U13.top_add_3ns_3ns_3_2_1_Adder_9_U.b ;
wire [2:0] \add_3ns_3ns_3_2_1_U13.top_add_3ns_3ns_3_2_1_Adder_9_U.bin_s0 ;
wire \add_3ns_3ns_3_2_1_U13.top_add_3ns_3ns_3_2_1_Adder_9_U.ce ;
wire \add_3ns_3ns_3_2_1_U13.top_add_3ns_3ns_3_2_1_Adder_9_U.clk ;
wire \add_3ns_3ns_3_2_1_U13.top_add_3ns_3ns_3_2_1_Adder_9_U.facout_s1 ;
wire \add_3ns_3ns_3_2_1_U13.top_add_3ns_3ns_3_2_1_Adder_9_U.facout_s2 ;
wire \add_3ns_3ns_3_2_1_U13.top_add_3ns_3ns_3_2_1_Adder_9_U.fas_s1 ;
wire [1:0] \add_3ns_3ns_3_2_1_U13.top_add_3ns_3ns_3_2_1_Adder_9_U.fas_s2 ;
wire \add_3ns_3ns_3_2_1_U13.top_add_3ns_3ns_3_2_1_Adder_9_U.reset ;
wire [2:0] \add_3ns_3ns_3_2_1_U13.top_add_3ns_3ns_3_2_1_Adder_9_U.s ;
wire \add_3ns_3ns_3_2_1_U13.top_add_3ns_3ns_3_2_1_Adder_9_U.u1.a ;
wire \add_3ns_3ns_3_2_1_U13.top_add_3ns_3ns_3_2_1_Adder_9_U.u1.b ;
wire \add_3ns_3ns_3_2_1_U13.top_add_3ns_3ns_3_2_1_Adder_9_U.u1.cin ;
wire \add_3ns_3ns_3_2_1_U13.top_add_3ns_3ns_3_2_1_Adder_9_U.u1.cout ;
wire \add_3ns_3ns_3_2_1_U13.top_add_3ns_3ns_3_2_1_Adder_9_U.u1.s ;
wire [1:0] \add_3ns_3ns_3_2_1_U13.top_add_3ns_3ns_3_2_1_Adder_9_U.u2.a ;
wire [1:0] \add_3ns_3ns_3_2_1_U13.top_add_3ns_3ns_3_2_1_Adder_9_U.u2.b ;
wire \add_3ns_3ns_3_2_1_U13.top_add_3ns_3ns_3_2_1_Adder_9_U.u2.cin ;
wire \add_3ns_3ns_3_2_1_U13.top_add_3ns_3ns_3_2_1_Adder_9_U.u2.cout ;
wire [1:0] \add_3ns_3ns_3_2_1_U13.top_add_3ns_3ns_3_2_1_Adder_9_U.u2.s ;
wire \add_4ns_4ns_4_2_1_U6.ce ;
wire \add_4ns_4ns_4_2_1_U6.clk ;
wire [3:0] \add_4ns_4ns_4_2_1_U6.din0 ;
wire [3:0] \add_4ns_4ns_4_2_1_U6.din1 ;
wire [3:0] \add_4ns_4ns_4_2_1_U6.dout ;
wire \add_4ns_4ns_4_2_1_U6.reset ;
wire [3:0] \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.a ;
wire [3:0] \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.ain_s0 ;
wire [3:0] \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.b ;
wire [3:0] \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.bin_s0 ;
wire \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.ce ;
wire \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.clk ;
wire \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.facout_s1 ;
wire \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.facout_s2 ;
wire [1:0] \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.fas_s1 ;
wire [1:0] \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.fas_s2 ;
wire \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.reset ;
wire [3:0] \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.s ;
wire [1:0] \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.u1.a ;
wire [1:0] \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.u1.b ;
wire \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.u1.cin ;
wire \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.u1.cout ;
wire [1:0] \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.u1.s ;
wire [1:0] \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.u2.a ;
wire [1:0] \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.u2.b ;
wire \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.u2.cin ;
wire \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.u2.cout ;
wire [1:0] \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.u2.s ;
wire \add_4s_4s_4_2_1_U16.ce ;
wire \add_4s_4s_4_2_1_U16.clk ;
wire [3:0] \add_4s_4s_4_2_1_U16.din0 ;
wire [3:0] \add_4s_4s_4_2_1_U16.din1 ;
wire [3:0] \add_4s_4s_4_2_1_U16.dout ;
wire \add_4s_4s_4_2_1_U16.reset ;
wire [3:0] \add_4s_4s_4_2_1_U16.top_add_4s_4s_4_2_1_Adder_12_U.a ;
wire [3:0] \add_4s_4s_4_2_1_U16.top_add_4s_4s_4_2_1_Adder_12_U.ain_s0 ;
wire [3:0] \add_4s_4s_4_2_1_U16.top_add_4s_4s_4_2_1_Adder_12_U.b ;
wire [3:0] \add_4s_4s_4_2_1_U16.top_add_4s_4s_4_2_1_Adder_12_U.bin_s0 ;
wire \add_4s_4s_4_2_1_U16.top_add_4s_4s_4_2_1_Adder_12_U.ce ;
wire \add_4s_4s_4_2_1_U16.top_add_4s_4s_4_2_1_Adder_12_U.clk ;
wire \add_4s_4s_4_2_1_U16.top_add_4s_4s_4_2_1_Adder_12_U.facout_s1 ;
wire \add_4s_4s_4_2_1_U16.top_add_4s_4s_4_2_1_Adder_12_U.facout_s2 ;
wire [1:0] \add_4s_4s_4_2_1_U16.top_add_4s_4s_4_2_1_Adder_12_U.fas_s1 ;
wire [1:0] \add_4s_4s_4_2_1_U16.top_add_4s_4s_4_2_1_Adder_12_U.fas_s2 ;
wire \add_4s_4s_4_2_1_U16.top_add_4s_4s_4_2_1_Adder_12_U.reset ;
wire [3:0] \add_4s_4s_4_2_1_U16.top_add_4s_4s_4_2_1_Adder_12_U.s ;
wire [1:0] \add_4s_4s_4_2_1_U16.top_add_4s_4s_4_2_1_Adder_12_U.u1.a ;
wire [1:0] \add_4s_4s_4_2_1_U16.top_add_4s_4s_4_2_1_Adder_12_U.u1.b ;
wire \add_4s_4s_4_2_1_U16.top_add_4s_4s_4_2_1_Adder_12_U.u1.cin ;
wire \add_4s_4s_4_2_1_U16.top_add_4s_4s_4_2_1_Adder_12_U.u1.cout ;
wire [1:0] \add_4s_4s_4_2_1_U16.top_add_4s_4s_4_2_1_Adder_12_U.u1.s ;
wire [1:0] \add_4s_4s_4_2_1_U16.top_add_4s_4s_4_2_1_Adder_12_U.u2.a ;
wire [1:0] \add_4s_4s_4_2_1_U16.top_add_4s_4s_4_2_1_Adder_12_U.u2.b ;
wire \add_4s_4s_4_2_1_U16.top_add_4s_4s_4_2_1_Adder_12_U.u2.cin ;
wire \add_4s_4s_4_2_1_U16.top_add_4s_4s_4_2_1_Adder_12_U.u2.cout ;
wire [1:0] \add_4s_4s_4_2_1_U16.top_add_4s_4s_4_2_1_Adder_12_U.u2.s ;
wire \add_5ns_5ns_5_2_1_U7.ce ;
wire \add_5ns_5ns_5_2_1_U7.clk ;
wire [4:0] \add_5ns_5ns_5_2_1_U7.din0 ;
wire [4:0] \add_5ns_5ns_5_2_1_U7.din1 ;
wire [4:0] \add_5ns_5ns_5_2_1_U7.dout ;
wire \add_5ns_5ns_5_2_1_U7.reset ;
wire [4:0] \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_5_U.a ;
wire [4:0] \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_5_U.ain_s0 ;
wire [4:0] \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_5_U.b ;
wire [4:0] \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_5_U.bin_s0 ;
wire \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_5_U.ce ;
wire \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_5_U.clk ;
wire \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_5_U.facout_s1 ;
wire \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_5_U.facout_s2 ;
wire [1:0] \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_5_U.fas_s1 ;
wire [2:0] \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_5_U.fas_s2 ;
wire \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_5_U.reset ;
wire [4:0] \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_5_U.s ;
wire [1:0] \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_5_U.u1.a ;
wire [1:0] \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_5_U.u1.b ;
wire \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_5_U.u1.cin ;
wire \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_5_U.u1.cout ;
wire [1:0] \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_5_U.u1.s ;
wire [2:0] \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_5_U.u2.a ;
wire [2:0] \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_5_U.u2.b ;
wire \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_5_U.u2.cin ;
wire \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_5_U.u2.cout ;
wire [2:0] \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_5_U.u2.s ;
wire \add_6ns_6s_6_2_1_U15.ce ;
wire \add_6ns_6s_6_2_1_U15.clk ;
wire [5:0] \add_6ns_6s_6_2_1_U15.din0 ;
wire [5:0] \add_6ns_6s_6_2_1_U15.din1 ;
wire [5:0] \add_6ns_6s_6_2_1_U15.dout ;
wire \add_6ns_6s_6_2_1_U15.reset ;
wire [5:0] \add_6ns_6s_6_2_1_U15.top_add_6ns_6s_6_2_1_Adder_11_U.a ;
wire [5:0] \add_6ns_6s_6_2_1_U15.top_add_6ns_6s_6_2_1_Adder_11_U.ain_s0 ;
wire [5:0] \add_6ns_6s_6_2_1_U15.top_add_6ns_6s_6_2_1_Adder_11_U.b ;
wire [5:0] \add_6ns_6s_6_2_1_U15.top_add_6ns_6s_6_2_1_Adder_11_U.bin_s0 ;
wire \add_6ns_6s_6_2_1_U15.top_add_6ns_6s_6_2_1_Adder_11_U.ce ;
wire \add_6ns_6s_6_2_1_U15.top_add_6ns_6s_6_2_1_Adder_11_U.clk ;
wire \add_6ns_6s_6_2_1_U15.top_add_6ns_6s_6_2_1_Adder_11_U.facout_s1 ;
wire \add_6ns_6s_6_2_1_U15.top_add_6ns_6s_6_2_1_Adder_11_U.facout_s2 ;
wire [2:0] \add_6ns_6s_6_2_1_U15.top_add_6ns_6s_6_2_1_Adder_11_U.fas_s1 ;
wire [2:0] \add_6ns_6s_6_2_1_U15.top_add_6ns_6s_6_2_1_Adder_11_U.fas_s2 ;
wire \add_6ns_6s_6_2_1_U15.top_add_6ns_6s_6_2_1_Adder_11_U.reset ;
wire [5:0] \add_6ns_6s_6_2_1_U15.top_add_6ns_6s_6_2_1_Adder_11_U.s ;
wire [2:0] \add_6ns_6s_6_2_1_U15.top_add_6ns_6s_6_2_1_Adder_11_U.u1.a ;
wire [2:0] \add_6ns_6s_6_2_1_U15.top_add_6ns_6s_6_2_1_Adder_11_U.u1.b ;
wire \add_6ns_6s_6_2_1_U15.top_add_6ns_6s_6_2_1_Adder_11_U.u1.cin ;
wire \add_6ns_6s_6_2_1_U15.top_add_6ns_6s_6_2_1_Adder_11_U.u1.cout ;
wire [2:0] \add_6ns_6s_6_2_1_U15.top_add_6ns_6s_6_2_1_Adder_11_U.u1.s ;
wire [2:0] \add_6ns_6s_6_2_1_U15.top_add_6ns_6s_6_2_1_Adder_11_U.u2.a ;
wire [2:0] \add_6ns_6s_6_2_1_U15.top_add_6ns_6s_6_2_1_Adder_11_U.u2.b ;
wire \add_6ns_6s_6_2_1_U15.top_add_6ns_6s_6_2_1_Adder_11_U.u2.cin ;
wire \add_6ns_6s_6_2_1_U15.top_add_6ns_6s_6_2_1_Adder_11_U.u2.cout ;
wire [2:0] \add_6ns_6s_6_2_1_U15.top_add_6ns_6s_6_2_1_Adder_11_U.u2.s ;
wire \add_6s_6ns_6_2_1_U18.ce ;
wire \add_6s_6ns_6_2_1_U18.clk ;
wire [5:0] \add_6s_6ns_6_2_1_U18.din0 ;
wire [5:0] \add_6s_6ns_6_2_1_U18.din1 ;
wire [5:0] \add_6s_6ns_6_2_1_U18.dout ;
wire \add_6s_6ns_6_2_1_U18.reset ;
wire [5:0] \add_6s_6ns_6_2_1_U18.top_add_6s_6ns_6_2_1_Adder_14_U.a ;
wire [5:0] \add_6s_6ns_6_2_1_U18.top_add_6s_6ns_6_2_1_Adder_14_U.ain_s0 ;
wire [5:0] \add_6s_6ns_6_2_1_U18.top_add_6s_6ns_6_2_1_Adder_14_U.b ;
wire [5:0] \add_6s_6ns_6_2_1_U18.top_add_6s_6ns_6_2_1_Adder_14_U.bin_s0 ;
wire \add_6s_6ns_6_2_1_U18.top_add_6s_6ns_6_2_1_Adder_14_U.ce ;
wire \add_6s_6ns_6_2_1_U18.top_add_6s_6ns_6_2_1_Adder_14_U.clk ;
wire \add_6s_6ns_6_2_1_U18.top_add_6s_6ns_6_2_1_Adder_14_U.facout_s1 ;
wire \add_6s_6ns_6_2_1_U18.top_add_6s_6ns_6_2_1_Adder_14_U.facout_s2 ;
wire [2:0] \add_6s_6ns_6_2_1_U18.top_add_6s_6ns_6_2_1_Adder_14_U.fas_s1 ;
wire [2:0] \add_6s_6ns_6_2_1_U18.top_add_6s_6ns_6_2_1_Adder_14_U.fas_s2 ;
wire \add_6s_6ns_6_2_1_U18.top_add_6s_6ns_6_2_1_Adder_14_U.reset ;
wire [5:0] \add_6s_6ns_6_2_1_U18.top_add_6s_6ns_6_2_1_Adder_14_U.s ;
wire [2:0] \add_6s_6ns_6_2_1_U18.top_add_6s_6ns_6_2_1_Adder_14_U.u1.a ;
wire [2:0] \add_6s_6ns_6_2_1_U18.top_add_6s_6ns_6_2_1_Adder_14_U.u1.b ;
wire \add_6s_6ns_6_2_1_U18.top_add_6s_6ns_6_2_1_Adder_14_U.u1.cin ;
wire \add_6s_6ns_6_2_1_U18.top_add_6s_6ns_6_2_1_Adder_14_U.u1.cout ;
wire [2:0] \add_6s_6ns_6_2_1_U18.top_add_6s_6ns_6_2_1_Adder_14_U.u1.s ;
wire [2:0] \add_6s_6ns_6_2_1_U18.top_add_6s_6ns_6_2_1_Adder_14_U.u2.a ;
wire [2:0] \add_6s_6ns_6_2_1_U18.top_add_6s_6ns_6_2_1_Adder_14_U.u2.b ;
wire \add_6s_6ns_6_2_1_U18.top_add_6s_6ns_6_2_1_Adder_14_U.u2.cin ;
wire \add_6s_6ns_6_2_1_U18.top_add_6s_6ns_6_2_1_Adder_14_U.u2.cout ;
wire [2:0] \add_6s_6ns_6_2_1_U18.top_add_6s_6ns_6_2_1_Adder_14_U.u2.s ;
wire \add_7s_7ns_7_2_1_U12.ce ;
wire \add_7s_7ns_7_2_1_U12.clk ;
wire [6:0] \add_7s_7ns_7_2_1_U12.din0 ;
wire [6:0] \add_7s_7ns_7_2_1_U12.din1 ;
wire [6:0] \add_7s_7ns_7_2_1_U12.dout ;
wire \add_7s_7ns_7_2_1_U12.reset ;
wire [6:0] \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_8_U.a ;
wire [6:0] \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_8_U.ain_s0 ;
wire [6:0] \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_8_U.b ;
wire [6:0] \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_8_U.bin_s0 ;
wire \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_8_U.ce ;
wire \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_8_U.clk ;
wire \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_8_U.facout_s1 ;
wire \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_8_U.facout_s2 ;
wire [2:0] \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_8_U.fas_s1 ;
wire [3:0] \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_8_U.fas_s2 ;
wire \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_8_U.reset ;
wire [6:0] \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_8_U.s ;
wire [2:0] \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_8_U.u1.a ;
wire [2:0] \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_8_U.u1.b ;
wire \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_8_U.u1.cin ;
wire \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_8_U.u1.cout ;
wire [2:0] \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_8_U.u1.s ;
wire [3:0] \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_8_U.u2.a ;
wire [3:0] \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_8_U.u2.b ;
wire \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_8_U.u2.cin ;
wire \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_8_U.u2.cout ;
wire [3:0] \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_8_U.u2.s ;
wire \add_7s_7s_7_2_1_U10.ce ;
wire \add_7s_7s_7_2_1_U10.clk ;
wire [6:0] \add_7s_7s_7_2_1_U10.din0 ;
wire [6:0] \add_7s_7s_7_2_1_U10.din1 ;
wire [6:0] \add_7s_7s_7_2_1_U10.dout ;
wire \add_7s_7s_7_2_1_U10.reset ;
wire [6:0] \add_7s_7s_7_2_1_U10.top_add_7s_7s_7_2_1_Adder_6_U.a ;
wire [6:0] \add_7s_7s_7_2_1_U10.top_add_7s_7s_7_2_1_Adder_6_U.ain_s0 ;
wire [6:0] \add_7s_7s_7_2_1_U10.top_add_7s_7s_7_2_1_Adder_6_U.b ;
wire [6:0] \add_7s_7s_7_2_1_U10.top_add_7s_7s_7_2_1_Adder_6_U.bin_s0 ;
wire \add_7s_7s_7_2_1_U10.top_add_7s_7s_7_2_1_Adder_6_U.ce ;
wire \add_7s_7s_7_2_1_U10.top_add_7s_7s_7_2_1_Adder_6_U.clk ;
wire \add_7s_7s_7_2_1_U10.top_add_7s_7s_7_2_1_Adder_6_U.facout_s1 ;
wire \add_7s_7s_7_2_1_U10.top_add_7s_7s_7_2_1_Adder_6_U.facout_s2 ;
wire [2:0] \add_7s_7s_7_2_1_U10.top_add_7s_7s_7_2_1_Adder_6_U.fas_s1 ;
wire [3:0] \add_7s_7s_7_2_1_U10.top_add_7s_7s_7_2_1_Adder_6_U.fas_s2 ;
wire \add_7s_7s_7_2_1_U10.top_add_7s_7s_7_2_1_Adder_6_U.reset ;
wire [6:0] \add_7s_7s_7_2_1_U10.top_add_7s_7s_7_2_1_Adder_6_U.s ;
wire [2:0] \add_7s_7s_7_2_1_U10.top_add_7s_7s_7_2_1_Adder_6_U.u1.a ;
wire [2:0] \add_7s_7s_7_2_1_U10.top_add_7s_7s_7_2_1_Adder_6_U.u1.b ;
wire \add_7s_7s_7_2_1_U10.top_add_7s_7s_7_2_1_Adder_6_U.u1.cin ;
wire \add_7s_7s_7_2_1_U10.top_add_7s_7s_7_2_1_Adder_6_U.u1.cout ;
wire [2:0] \add_7s_7s_7_2_1_U10.top_add_7s_7s_7_2_1_Adder_6_U.u1.s ;
wire [3:0] \add_7s_7s_7_2_1_U10.top_add_7s_7s_7_2_1_Adder_6_U.u2.a ;
wire [3:0] \add_7s_7s_7_2_1_U10.top_add_7s_7s_7_2_1_Adder_6_U.u2.b ;
wire \add_7s_7s_7_2_1_U10.top_add_7s_7s_7_2_1_Adder_6_U.u2.cin ;
wire \add_7s_7s_7_2_1_U10.top_add_7s_7s_7_2_1_Adder_6_U.u2.cout ;
wire [3:0] \add_7s_7s_7_2_1_U10.top_add_7s_7s_7_2_1_Adder_6_U.u2.s ;
wire \add_9ns_9ns_9_2_1_U17.ce ;
wire \add_9ns_9ns_9_2_1_U17.clk ;
wire [8:0] \add_9ns_9ns_9_2_1_U17.din0 ;
wire [8:0] \add_9ns_9ns_9_2_1_U17.din1 ;
wire [8:0] \add_9ns_9ns_9_2_1_U17.dout ;
wire \add_9ns_9ns_9_2_1_U17.reset ;
wire [8:0] \add_9ns_9ns_9_2_1_U17.top_add_9ns_9ns_9_2_1_Adder_13_U.a ;
wire [8:0] \add_9ns_9ns_9_2_1_U17.top_add_9ns_9ns_9_2_1_Adder_13_U.ain_s0 ;
wire [8:0] \add_9ns_9ns_9_2_1_U17.top_add_9ns_9ns_9_2_1_Adder_13_U.b ;
wire [8:0] \add_9ns_9ns_9_2_1_U17.top_add_9ns_9ns_9_2_1_Adder_13_U.bin_s0 ;
wire \add_9ns_9ns_9_2_1_U17.top_add_9ns_9ns_9_2_1_Adder_13_U.ce ;
wire \add_9ns_9ns_9_2_1_U17.top_add_9ns_9ns_9_2_1_Adder_13_U.clk ;
wire \add_9ns_9ns_9_2_1_U17.top_add_9ns_9ns_9_2_1_Adder_13_U.facout_s1 ;
wire \add_9ns_9ns_9_2_1_U17.top_add_9ns_9ns_9_2_1_Adder_13_U.facout_s2 ;
wire [3:0] \add_9ns_9ns_9_2_1_U17.top_add_9ns_9ns_9_2_1_Adder_13_U.fas_s1 ;
wire [4:0] \add_9ns_9ns_9_2_1_U17.top_add_9ns_9ns_9_2_1_Adder_13_U.fas_s2 ;
wire \add_9ns_9ns_9_2_1_U17.top_add_9ns_9ns_9_2_1_Adder_13_U.reset ;
wire [8:0] \add_9ns_9ns_9_2_1_U17.top_add_9ns_9ns_9_2_1_Adder_13_U.s ;
wire [3:0] \add_9ns_9ns_9_2_1_U17.top_add_9ns_9ns_9_2_1_Adder_13_U.u1.a ;
wire [3:0] \add_9ns_9ns_9_2_1_U17.top_add_9ns_9ns_9_2_1_Adder_13_U.u1.b ;
wire \add_9ns_9ns_9_2_1_U17.top_add_9ns_9ns_9_2_1_Adder_13_U.u1.cin ;
wire \add_9ns_9ns_9_2_1_U17.top_add_9ns_9ns_9_2_1_Adder_13_U.u1.cout ;
wire [3:0] \add_9ns_9ns_9_2_1_U17.top_add_9ns_9ns_9_2_1_Adder_13_U.u1.s ;
wire [4:0] \add_9ns_9ns_9_2_1_U17.top_add_9ns_9ns_9_2_1_Adder_13_U.u2.a ;
wire [4:0] \add_9ns_9ns_9_2_1_U17.top_add_9ns_9ns_9_2_1_Adder_13_U.u2.b ;
wire \add_9ns_9ns_9_2_1_U17.top_add_9ns_9ns_9_2_1_Adder_13_U.u2.cin ;
wire \add_9ns_9ns_9_2_1_U17.top_add_9ns_9ns_9_2_1_Adder_13_U.u2.cout ;
wire [4:0] \add_9ns_9ns_9_2_1_U17.top_add_9ns_9ns_9_2_1_Adder_13_U.u2.s ;
wire \add_9s_9ns_9_2_1_U19.ce ;
wire \add_9s_9ns_9_2_1_U19.clk ;
wire [8:0] \add_9s_9ns_9_2_1_U19.din0 ;
wire [8:0] \add_9s_9ns_9_2_1_U19.din1 ;
wire [8:0] \add_9s_9ns_9_2_1_U19.dout ;
wire \add_9s_9ns_9_2_1_U19.reset ;
wire [8:0] \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_15_U.a ;
wire [8:0] \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_15_U.ain_s0 ;
wire [8:0] \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_15_U.b ;
wire [8:0] \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_15_U.bin_s0 ;
wire \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_15_U.ce ;
wire \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_15_U.clk ;
wire \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_15_U.facout_s1 ;
wire \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_15_U.facout_s2 ;
wire [3:0] \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_15_U.fas_s1 ;
wire [4:0] \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_15_U.fas_s2 ;
wire \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_15_U.reset ;
wire [8:0] \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_15_U.s ;
wire [3:0] \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_15_U.u1.a ;
wire [3:0] \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_15_U.u1.b ;
wire \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_15_U.u1.cin ;
wire \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_15_U.u1.cout ;
wire [3:0] \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_15_U.u1.s ;
wire [4:0] \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_15_U.u2.a ;
wire [4:0] \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_15_U.u2.b ;
wire \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_15_U.u2.cin ;
wire \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_15_U.u2.cout ;
wire [4:0] \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_15_U.u2.s ;
wire \add_9s_9s_9_2_1_U14.ce ;
wire \add_9s_9s_9_2_1_U14.clk ;
wire [8:0] \add_9s_9s_9_2_1_U14.din0 ;
wire [8:0] \add_9s_9s_9_2_1_U14.din1 ;
wire [8:0] \add_9s_9s_9_2_1_U14.dout ;
wire \add_9s_9s_9_2_1_U14.reset ;
wire [8:0] \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_10_U.a ;
wire [8:0] \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_10_U.ain_s0 ;
wire [8:0] \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_10_U.b ;
wire [8:0] \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_10_U.bin_s0 ;
wire \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_10_U.ce ;
wire \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_10_U.clk ;
wire \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_10_U.facout_s1 ;
wire \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_10_U.facout_s2 ;
wire [3:0] \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_10_U.fas_s1 ;
wire [4:0] \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_10_U.fas_s2 ;
wire \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_10_U.reset ;
wire [8:0] \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_10_U.s ;
wire [3:0] \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_10_U.u1.a ;
wire [3:0] \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_10_U.u1.b ;
wire \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_10_U.u1.cin ;
wire \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_10_U.u1.cout ;
wire [3:0] \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_10_U.u1.s ;
wire [4:0] \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_10_U.u2.a ;
wire [4:0] \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_10_U.u2.b ;
wire \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_10_U.u2.cin ;
wire \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_10_U.u2.cout ;
wire [4:0] \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_10_U.u2.s ;
wire and_ln353_fu_412_p2;
wire ap_CS_fsm_state1;
wire ap_CS_fsm_state10;
wire ap_CS_fsm_state11;
wire ap_CS_fsm_state12;
wire ap_CS_fsm_state13;
wire ap_CS_fsm_state14;
wire ap_CS_fsm_state15;
wire ap_CS_fsm_state16;
wire ap_CS_fsm_state17;
wire ap_CS_fsm_state18;
wire ap_CS_fsm_state19;
wire ap_CS_fsm_state2;
wire ap_CS_fsm_state3;
wire ap_CS_fsm_state4;
wire ap_CS_fsm_state5;
wire ap_CS_fsm_state6;
wire ap_CS_fsm_state7;
wire ap_CS_fsm_state8;
wire ap_CS_fsm_state9;
wire [18:0] ap_NS_fsm;
wire ap_clk;
wire ap_done;
wire ap_idle;
wire ap_ready;
wire ap_rst;
wire ap_start;
wire [31:0] conv_i482_fu_363_p1;
wire [1:0] grp_fu_199_p0;
wire [1:0] grp_fu_199_p2;
wire [10:0] grp_fu_248_p0;
wire [10:0] grp_fu_248_p1;
wire [10:0] grp_fu_248_p2;
wire [2:0] grp_fu_267_p1;
wire [2:0] grp_fu_267_p2;
wire [1:0] grp_fu_311_p0;
wire [1:0] grp_fu_311_p2;
wire [32:0] grp_fu_333_p0;
wire [32:0] grp_fu_333_p1;
wire [32:0] grp_fu_333_p2;
wire [3:0] grp_fu_349_p0;
wire [3:0] grp_fu_349_p2;
wire [4:0] grp_fu_355_p2;
wire [31:0] grp_fu_367_p1;
wire [31:0] grp_fu_367_p2;
wire [31:0] grp_fu_376_p1;
wire [31:0] grp_fu_376_p2;
wire [6:0] grp_fu_476_p0;
wire [6:0] grp_fu_476_p1;
wire [6:0] grp_fu_476_p2;
wire [8:0] grp_fu_485_p1;
wire [8:0] grp_fu_485_p2;
wire [6:0] grp_fu_517_p0;
wire [6:0] grp_fu_517_p2;
wire [2:0] grp_fu_528_p2;
wire [8:0] grp_fu_607_p0;
wire [8:0] grp_fu_607_p1;
wire [8:0] grp_fu_607_p2;
wire [5:0] grp_fu_613_p0;
wire [5:0] grp_fu_613_p1;
wire [5:0] grp_fu_613_p2;
wire [3:0] grp_fu_619_p0;
wire [3:0] grp_fu_619_p1;
wire [3:0] grp_fu_619_p2;
wire [8:0] grp_fu_632_p2;
wire [5:0] grp_fu_639_p0;
wire [5:0] grp_fu_639_p2;
wire [8:0] grp_fu_647_p0;
wire [8:0] grp_fu_647_p2;
wire icmp_ln851_1_fu_305_p2;
wire icmp_ln851_2_fu_193_p2;
wire icmp_ln851_3_fu_523_p2;
wire icmp_ln851_fu_258_p2;
wire [9:0] lhs_fu_232_p3;
wire \lshr_32ns_32s_32_7_1_U9.ce ;
wire \lshr_32ns_32s_32_7_1_U9.clk ;
wire [31:0] \lshr_32ns_32s_32_7_1_U9.din0 ;
wire [31:0] \lshr_32ns_32s_32_7_1_U9.din1 ;
wire [31:0] \lshr_32ns_32s_32_7_1_U9.din1_cast ;
wire [31:0] \lshr_32ns_32s_32_7_1_U9.din1_mask ;
wire [31:0] \lshr_32ns_32s_32_7_1_U9.dout ;
wire \lshr_32ns_32s_32_7_1_U9.reset ;
wire [3:0] op_0;
wire [7:0] op_1;
wire [7:0] op_10;
wire [7:0] op_11;
wire [7:0] op_12;
wire [3:0] op_15_V_fu_541_p3;
wire [7:0] op_2;
wire [31:0] op_3;
wire [31:0] op_30;
wire op_30_ap_vld;
wire [3:0] op_4;
wire [1:0] op_6;
wire [31:0] p_Result_1_fu_293_p1;
wire p_Result_2_fu_400_p3;
wire [7:0] p_Result_3_fu_205_p1;
wire p_Result_3_fu_205_p3;
wire p_Result_4_fu_546_p3;
wire p_Result_5_fu_569_p3;
wire p_Result_s_fu_435_p3;
wire [2:0] ret_V_15_fu_581_p3;
wire [1:0] ret_V_19_fu_387_p3;
wire ret_V_21_fu_418_p2;
wire [6:0] ret_V_23_fu_562_p3;
wire [3:0] ret_V_25_fu_429_p3;
wire [31:0] ret_V_3_cast5_fu_339_p1;
wire [31:0] ret_V_3_cast_fu_283_p1;
wire [7:0] ret_V_7_fu_179_p1;
wire [1:0] ret_V_9_fu_217_p3;
wire [5:0] rhs_1_fu_465_p3;
wire [20:0] rhs_fu_321_p3;
wire [1:0] select_ln69_fu_625_p3;
wire [8:0] select_ln703_fu_454_p3;
wire [1:0] select_ln850_1_fu_212_p3;
wire [4:0] select_ln850_3_fu_442_p3;
wire [6:0] select_ln850_4_fu_556_p3;
wire [2:0] select_ln850_5_fu_576_p3;
wire [3:0] select_ln850_6_fu_424_p3;
wire [4:0] select_ln850_7_fu_447_p3;
wire [1:0] select_ln850_fu_382_p3;
wire [1:0] sext_ln1192_1_fu_461_p0;
wire [31:0] sext_ln703_1_fu_317_p0;
wire [7:0] sext_ln703_2_fu_482_p0;
wire [7:0] sext_ln703_fu_244_p0;
wire [6:0] sext_ln850_fu_514_p1;
wire \shl_32ns_32s_32_7_1_U8.ce ;
wire \shl_32ns_32s_32_7_1_U8.clk ;
wire [31:0] \shl_32ns_32s_32_7_1_U8.din0 ;
wire [31:0] \shl_32ns_32s_32_7_1_U8.din1 ;
wire [31:0] \shl_32ns_32s_32_7_1_U8.din1_cast ;
wire [31:0] \shl_32ns_32s_32_7_1_U8.din1_mask ;
wire [31:0] \shl_32ns_32s_32_7_1_U8.dout ;
wire \shl_32ns_32s_32_7_1_U8.reset ;
wire \sub_3ns_3s_3_2_1_U3.ce ;
wire \sub_3ns_3s_3_2_1_U3.clk ;
wire [2:0] \sub_3ns_3s_3_2_1_U3.din0 ;
wire [2:0] \sub_3ns_3s_3_2_1_U3.din1 ;
wire [2:0] \sub_3ns_3s_3_2_1_U3.dout ;
wire \sub_3ns_3s_3_2_1_U3.reset ;
wire [2:0] \sub_3ns_3s_3_2_1_U3.top_sub_3ns_3s_3_2_1_Adder_2_U.a ;
wire [2:0] \sub_3ns_3s_3_2_1_U3.top_sub_3ns_3s_3_2_1_Adder_2_U.ain_s0 ;
wire [2:0] \sub_3ns_3s_3_2_1_U3.top_sub_3ns_3s_3_2_1_Adder_2_U.b ;
wire [2:0] \sub_3ns_3s_3_2_1_U3.top_sub_3ns_3s_3_2_1_Adder_2_U.bin_s0 ;
wire \sub_3ns_3s_3_2_1_U3.top_sub_3ns_3s_3_2_1_Adder_2_U.ce ;
wire \sub_3ns_3s_3_2_1_U3.top_sub_3ns_3s_3_2_1_Adder_2_U.clk ;
wire \sub_3ns_3s_3_2_1_U3.top_sub_3ns_3s_3_2_1_Adder_2_U.facout_s1 ;
wire \sub_3ns_3s_3_2_1_U3.top_sub_3ns_3s_3_2_1_Adder_2_U.facout_s2 ;
wire \sub_3ns_3s_3_2_1_U3.top_sub_3ns_3s_3_2_1_Adder_2_U.fas_s1 ;
wire [1:0] \sub_3ns_3s_3_2_1_U3.top_sub_3ns_3s_3_2_1_Adder_2_U.fas_s2 ;
wire \sub_3ns_3s_3_2_1_U3.top_sub_3ns_3s_3_2_1_Adder_2_U.reset ;
wire [2:0] \sub_3ns_3s_3_2_1_U3.top_sub_3ns_3s_3_2_1_Adder_2_U.s ;
wire \sub_3ns_3s_3_2_1_U3.top_sub_3ns_3s_3_2_1_Adder_2_U.u1.a ;
wire \sub_3ns_3s_3_2_1_U3.top_sub_3ns_3s_3_2_1_Adder_2_U.u1.b ;
wire \sub_3ns_3s_3_2_1_U3.top_sub_3ns_3s_3_2_1_Adder_2_U.u1.cin ;
wire \sub_3ns_3s_3_2_1_U3.top_sub_3ns_3s_3_2_1_Adder_2_U.u1.cout ;
wire \sub_3ns_3s_3_2_1_U3.top_sub_3ns_3s_3_2_1_Adder_2_U.u1.s ;
wire [1:0] \sub_3ns_3s_3_2_1_U3.top_sub_3ns_3s_3_2_1_Adder_2_U.u2.a ;
wire [1:0] \sub_3ns_3s_3_2_1_U3.top_sub_3ns_3s_3_2_1_Adder_2_U.u2.b ;
wire \sub_3ns_3s_3_2_1_U3.top_sub_3ns_3s_3_2_1_Adder_2_U.u2.cin ;
wire \sub_3ns_3s_3_2_1_U3.top_sub_3ns_3s_3_2_1_Adder_2_U.u2.cout ;
wire [1:0] \sub_3ns_3s_3_2_1_U3.top_sub_3ns_3s_3_2_1_Adder_2_U.u2.s ;
wire \sub_9ns_9s_9_2_1_U11.ce ;
wire \sub_9ns_9s_9_2_1_U11.clk ;
wire [8:0] \sub_9ns_9s_9_2_1_U11.din0 ;
wire [8:0] \sub_9ns_9s_9_2_1_U11.din1 ;
wire [8:0] \sub_9ns_9s_9_2_1_U11.dout ;
wire \sub_9ns_9s_9_2_1_U11.reset ;
wire [8:0] \sub_9ns_9s_9_2_1_U11.top_sub_9ns_9s_9_2_1_Adder_7_U.a ;
wire [8:0] \sub_9ns_9s_9_2_1_U11.top_sub_9ns_9s_9_2_1_Adder_7_U.ain_s0 ;
wire [8:0] \sub_9ns_9s_9_2_1_U11.top_sub_9ns_9s_9_2_1_Adder_7_U.b ;
wire [8:0] \sub_9ns_9s_9_2_1_U11.top_sub_9ns_9s_9_2_1_Adder_7_U.bin_s0 ;
wire \sub_9ns_9s_9_2_1_U11.top_sub_9ns_9s_9_2_1_Adder_7_U.ce ;
wire \sub_9ns_9s_9_2_1_U11.top_sub_9ns_9s_9_2_1_Adder_7_U.clk ;
wire \sub_9ns_9s_9_2_1_U11.top_sub_9ns_9s_9_2_1_Adder_7_U.facout_s1 ;
wire \sub_9ns_9s_9_2_1_U11.top_sub_9ns_9s_9_2_1_Adder_7_U.facout_s2 ;
wire [3:0] \sub_9ns_9s_9_2_1_U11.top_sub_9ns_9s_9_2_1_Adder_7_U.fas_s1 ;
wire [4:0] \sub_9ns_9s_9_2_1_U11.top_sub_9ns_9s_9_2_1_Adder_7_U.fas_s2 ;
wire \sub_9ns_9s_9_2_1_U11.top_sub_9ns_9s_9_2_1_Adder_7_U.reset ;
wire [8:0] \sub_9ns_9s_9_2_1_U11.top_sub_9ns_9s_9_2_1_Adder_7_U.s ;
wire [3:0] \sub_9ns_9s_9_2_1_U11.top_sub_9ns_9s_9_2_1_Adder_7_U.u1.a ;
wire [3:0] \sub_9ns_9s_9_2_1_U11.top_sub_9ns_9s_9_2_1_Adder_7_U.u1.b ;
wire \sub_9ns_9s_9_2_1_U11.top_sub_9ns_9s_9_2_1_Adder_7_U.u1.cin ;
wire \sub_9ns_9s_9_2_1_U11.top_sub_9ns_9s_9_2_1_Adder_7_U.u1.cout ;
wire [3:0] \sub_9ns_9s_9_2_1_U11.top_sub_9ns_9s_9_2_1_Adder_7_U.u1.s ;
wire [4:0] \sub_9ns_9s_9_2_1_U11.top_sub_9ns_9s_9_2_1_Adder_7_U.u2.a ;
wire [4:0] \sub_9ns_9s_9_2_1_U11.top_sub_9ns_9s_9_2_1_Adder_7_U.u2.b ;
wire \sub_9ns_9s_9_2_1_U11.top_sub_9ns_9s_9_2_1_Adder_7_U.u2.cin ;
wire \sub_9ns_9s_9_2_1_U11.top_sub_9ns_9s_9_2_1_Adder_7_U.u2.cout ;
wire [4:0] \sub_9ns_9s_9_2_1_U11.top_sub_9ns_9s_9_2_1_Adder_7_U.u2.s ;
wire tmp_fu_393_p3;
wire [3:0] trunc_ln1497_1_fu_537_p1;
wire [3:0] trunc_ln1497_fu_533_p1;
wire [31:0] trunc_ln851_1_fu_301_p0;
wire [16:0] trunc_ln851_1_fu_301_p1;
wire [7:0] trunc_ln851_2_fu_189_p0;
wire [5:0] trunc_ln851_2_fu_189_p1;
wire [1:0] trunc_ln851_3_fu_553_p0;
wire trunc_ln851_3_fu_553_p1;
wire [5:0] trunc_ln851_4_fu_510_p1;
wire [7:0] trunc_ln851_fu_254_p0;
wire [5:0] trunc_ln851_fu_254_p1;
wire xor_ln850_fu_407_p2;


assign _044_ = _050_ & ap_CS_fsm[6];
assign _045_ = tmp_4_reg_686 & ap_CS_fsm[4];
assign _046_ = _051_ & ap_CS_fsm[11];
assign _047_ = tmp_4_reg_686 & ap_CS_fsm[11];
assign _048_ = _052_ & ap_CS_fsm[0];
assign _049_ = ap_start & ap_CS_fsm[0];
assign and_ln353_fu_412_p2 = xor_ln850_fu_407_p2 & ret_V_20_reg_770[32];
assign xor_ln850_fu_407_p2 = ~ icmp_ln851_1_reg_736;
assign _050_ = ~ icmp_ln851_reg_701;
assign _051_ = ~ tmp_4_reg_686;
assign _052_ = ~ ap_start;
assign _053_ = ! op_3[16:0];
assign _054_ = ! op_11[5:0];
assign _055_ = ! trunc_ln851_4_reg_870;
assign _056_ = ! op_1[5:0];
always @(posedge \add_11s_11s_11_2_1_U2.top_add_11s_11s_11_2_1_Adder_1_U.clk )
\add_11s_11s_11_2_1_U2.top_add_11s_11s_11_2_1_Adder_1_U.bin_s1  <= _058_;
always @(posedge \add_11s_11s_11_2_1_U2.top_add_11s_11s_11_2_1_Adder_1_U.clk )
\add_11s_11s_11_2_1_U2.top_add_11s_11s_11_2_1_Adder_1_U.ain_s1  <= _057_;
always @(posedge \add_11s_11s_11_2_1_U2.top_add_11s_11s_11_2_1_Adder_1_U.clk )
\add_11s_11s_11_2_1_U2.top_add_11s_11s_11_2_1_Adder_1_U.sum_s1  <= _060_;
always @(posedge \add_11s_11s_11_2_1_U2.top_add_11s_11s_11_2_1_Adder_1_U.clk )
\add_11s_11s_11_2_1_U2.top_add_11s_11s_11_2_1_Adder_1_U.carry_s1  <= _059_;
assign _058_ = \add_11s_11s_11_2_1_U2.top_add_11s_11s_11_2_1_Adder_1_U.ce  ? \add_11s_11s_11_2_1_U2.top_add_11s_11s_11_2_1_Adder_1_U.b [10:5] : \add_11s_11s_11_2_1_U2.top_add_11s_11s_11_2_1_Adder_1_U.bin_s1 ;
assign _057_ = \add_11s_11s_11_2_1_U2.top_add_11s_11s_11_2_1_Adder_1_U.ce  ? \add_11s_11s_11_2_1_U2.top_add_11s_11s_11_2_1_Adder_1_U.a [10:5] : \add_11s_11s_11_2_1_U2.top_add_11s_11s_11_2_1_Adder_1_U.ain_s1 ;
assign _059_ = \add_11s_11s_11_2_1_U2.top_add_11s_11s_11_2_1_Adder_1_U.ce  ? \add_11s_11s_11_2_1_U2.top_add_11s_11s_11_2_1_Adder_1_U.facout_s1  : \add_11s_11s_11_2_1_U2.top_add_11s_11s_11_2_1_Adder_1_U.carry_s1 ;
assign _060_ = \add_11s_11s_11_2_1_U2.top_add_11s_11s_11_2_1_Adder_1_U.ce  ? \add_11s_11s_11_2_1_U2.top_add_11s_11s_11_2_1_Adder_1_U.fas_s1  : \add_11s_11s_11_2_1_U2.top_add_11s_11s_11_2_1_Adder_1_U.sum_s1 ;
assign _061_ = \add_11s_11s_11_2_1_U2.top_add_11s_11s_11_2_1_Adder_1_U.u1.a  + \add_11s_11s_11_2_1_U2.top_add_11s_11s_11_2_1_Adder_1_U.u1.b ;
assign { \add_11s_11s_11_2_1_U2.top_add_11s_11s_11_2_1_Adder_1_U.u1.cout , \add_11s_11s_11_2_1_U2.top_add_11s_11s_11_2_1_Adder_1_U.u1.s  } = _061_ + \add_11s_11s_11_2_1_U2.top_add_11s_11s_11_2_1_Adder_1_U.u1.cin ;
assign _062_ = \add_11s_11s_11_2_1_U2.top_add_11s_11s_11_2_1_Adder_1_U.u2.a  + \add_11s_11s_11_2_1_U2.top_add_11s_11s_11_2_1_Adder_1_U.u2.b ;
assign { \add_11s_11s_11_2_1_U2.top_add_11s_11s_11_2_1_Adder_1_U.u2.cout , \add_11s_11s_11_2_1_U2.top_add_11s_11s_11_2_1_Adder_1_U.u2.s  } = _062_ + \add_11s_11s_11_2_1_U2.top_add_11s_11s_11_2_1_Adder_1_U.u2.cin ;
always @(posedge \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.clk )
\add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.bin_s1  <= _064_;
always @(posedge \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.clk )
\add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.ain_s1  <= _063_;
always @(posedge \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.clk )
\add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.sum_s1  <= _066_;
always @(posedge \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.clk )
\add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.carry_s1  <= _065_;
assign _064_ = \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.ce  ? \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.b [1] : \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.bin_s1 ;
assign _063_ = \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.ce  ? \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.a [1] : \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.ain_s1 ;
assign _065_ = \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.ce  ? \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.facout_s1  : \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.carry_s1 ;
assign _066_ = \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.ce  ? \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.fas_s1  : \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.sum_s1 ;
assign _067_ = \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.u1.a  + \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.u1.b ;
assign { \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.u1.cout , \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.u1.s  } = _067_ + \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.u1.cin ;
assign _068_ = \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.u2.a  + \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.u2.b ;
assign { \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.u2.cout , \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.u2.s  } = _068_ + \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.u2.cin ;
always @(posedge \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_0_U.clk )
\add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_0_U.bin_s1  <= _070_;
always @(posedge \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_0_U.clk )
\add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_0_U.ain_s1  <= _069_;
always @(posedge \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_0_U.clk )
\add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_0_U.sum_s1  <= _072_;
always @(posedge \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_0_U.clk )
\add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_0_U.carry_s1  <= _071_;
assign _070_ = \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_0_U.ce  ? \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_0_U.b [1] : \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_0_U.bin_s1 ;
assign _069_ = \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_0_U.ce  ? \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_0_U.a [1] : \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_0_U.ain_s1 ;
assign _071_ = \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_0_U.ce  ? \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_0_U.facout_s1  : \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_0_U.carry_s1 ;
assign _072_ = \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_0_U.ce  ? \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_0_U.fas_s1  : \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_0_U.sum_s1 ;
assign _073_ = \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_0_U.u1.a  + \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_0_U.u1.b ;
assign { \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_0_U.u1.cout , \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_0_U.u1.s  } = _073_ + \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_0_U.u1.cin ;
assign _074_ = \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_0_U.u2.a  + \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_0_U.u2.b ;
assign { \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_0_U.u2.cout , \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_0_U.u2.s  } = _074_ + \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_0_U.u2.cin ;
always @(posedge \add_33ns_33s_33_2_1_U5.top_add_33ns_33s_33_2_1_Adder_3_U.clk )
\add_33ns_33s_33_2_1_U5.top_add_33ns_33s_33_2_1_Adder_3_U.bin_s1  <= _076_;
always @(posedge \add_33ns_33s_33_2_1_U5.top_add_33ns_33s_33_2_1_Adder_3_U.clk )
\add_33ns_33s_33_2_1_U5.top_add_33ns_33s_33_2_1_Adder_3_U.ain_s1  <= _075_;
always @(posedge \add_33ns_33s_33_2_1_U5.top_add_33ns_33s_33_2_1_Adder_3_U.clk )
\add_33ns_33s_33_2_1_U5.top_add_33ns_33s_33_2_1_Adder_3_U.sum_s1  <= _078_;
always @(posedge \add_33ns_33s_33_2_1_U5.top_add_33ns_33s_33_2_1_Adder_3_U.clk )
\add_33ns_33s_33_2_1_U5.top_add_33ns_33s_33_2_1_Adder_3_U.carry_s1  <= _077_;
assign _076_ = \add_33ns_33s_33_2_1_U5.top_add_33ns_33s_33_2_1_Adder_3_U.ce  ? \add_33ns_33s_33_2_1_U5.top_add_33ns_33s_33_2_1_Adder_3_U.b [32:16] : \add_33ns_33s_33_2_1_U5.top_add_33ns_33s_33_2_1_Adder_3_U.bin_s1 ;
assign _075_ = \add_33ns_33s_33_2_1_U5.top_add_33ns_33s_33_2_1_Adder_3_U.ce  ? \add_33ns_33s_33_2_1_U5.top_add_33ns_33s_33_2_1_Adder_3_U.a [32:16] : \add_33ns_33s_33_2_1_U5.top_add_33ns_33s_33_2_1_Adder_3_U.ain_s1 ;
assign _077_ = \add_33ns_33s_33_2_1_U5.top_add_33ns_33s_33_2_1_Adder_3_U.ce  ? \add_33ns_33s_33_2_1_U5.top_add_33ns_33s_33_2_1_Adder_3_U.facout_s1  : \add_33ns_33s_33_2_1_U5.top_add_33ns_33s_33_2_1_Adder_3_U.carry_s1 ;
assign _078_ = \add_33ns_33s_33_2_1_U5.top_add_33ns_33s_33_2_1_Adder_3_U.ce  ? \add_33ns_33s_33_2_1_U5.top_add_33ns_33s_33_2_1_Adder_3_U.fas_s1  : \add_33ns_33s_33_2_1_U5.top_add_33ns_33s_33_2_1_Adder_3_U.sum_s1 ;
assign _079_ = \add_33ns_33s_33_2_1_U5.top_add_33ns_33s_33_2_1_Adder_3_U.u1.a  + \add_33ns_33s_33_2_1_U5.top_add_33ns_33s_33_2_1_Adder_3_U.u1.b ;
assign { \add_33ns_33s_33_2_1_U5.top_add_33ns_33s_33_2_1_Adder_3_U.u1.cout , \add_33ns_33s_33_2_1_U5.top_add_33ns_33s_33_2_1_Adder_3_U.u1.s  } = _079_ + \add_33ns_33s_33_2_1_U5.top_add_33ns_33s_33_2_1_Adder_3_U.u1.cin ;
assign _080_ = \add_33ns_33s_33_2_1_U5.top_add_33ns_33s_33_2_1_Adder_3_U.u2.a  + \add_33ns_33s_33_2_1_U5.top_add_33ns_33s_33_2_1_Adder_3_U.u2.b ;
assign { \add_33ns_33s_33_2_1_U5.top_add_33ns_33s_33_2_1_Adder_3_U.u2.cout , \add_33ns_33s_33_2_1_U5.top_add_33ns_33s_33_2_1_Adder_3_U.u2.s  } = _080_ + \add_33ns_33s_33_2_1_U5.top_add_33ns_33s_33_2_1_Adder_3_U.u2.cin ;
always @(posedge \add_3ns_3ns_3_2_1_U13.top_add_3ns_3ns_3_2_1_Adder_9_U.clk )
\add_3ns_3ns_3_2_1_U13.top_add_3ns_3ns_3_2_1_Adder_9_U.bin_s1  <= _082_;
always @(posedge \add_3ns_3ns_3_2_1_U13.top_add_3ns_3ns_3_2_1_Adder_9_U.clk )
\add_3ns_3ns_3_2_1_U13.top_add_3ns_3ns_3_2_1_Adder_9_U.ain_s1  <= _081_;
always @(posedge \add_3ns_3ns_3_2_1_U13.top_add_3ns_3ns_3_2_1_Adder_9_U.clk )
\add_3ns_3ns_3_2_1_U13.top_add_3ns_3ns_3_2_1_Adder_9_U.sum_s1  <= _084_;
always @(posedge \add_3ns_3ns_3_2_1_U13.top_add_3ns_3ns_3_2_1_Adder_9_U.clk )
\add_3ns_3ns_3_2_1_U13.top_add_3ns_3ns_3_2_1_Adder_9_U.carry_s1  <= _083_;
assign _082_ = \add_3ns_3ns_3_2_1_U13.top_add_3ns_3ns_3_2_1_Adder_9_U.ce  ? \add_3ns_3ns_3_2_1_U13.top_add_3ns_3ns_3_2_1_Adder_9_U.b [2:1] : \add_3ns_3ns_3_2_1_U13.top_add_3ns_3ns_3_2_1_Adder_9_U.bin_s1 ;
assign _081_ = \add_3ns_3ns_3_2_1_U13.top_add_3ns_3ns_3_2_1_Adder_9_U.ce  ? \add_3ns_3ns_3_2_1_U13.top_add_3ns_3ns_3_2_1_Adder_9_U.a [2:1] : \add_3ns_3ns_3_2_1_U13.top_add_3ns_3ns_3_2_1_Adder_9_U.ain_s1 ;
assign _083_ = \add_3ns_3ns_3_2_1_U13.top_add_3ns_3ns_3_2_1_Adder_9_U.ce  ? \add_3ns_3ns_3_2_1_U13.top_add_3ns_3ns_3_2_1_Adder_9_U.facout_s1  : \add_3ns_3ns_3_2_1_U13.top_add_3ns_3ns_3_2_1_Adder_9_U.carry_s1 ;
assign _084_ = \add_3ns_3ns_3_2_1_U13.top_add_3ns_3ns_3_2_1_Adder_9_U.ce  ? \add_3ns_3ns_3_2_1_U13.top_add_3ns_3ns_3_2_1_Adder_9_U.fas_s1  : \add_3ns_3ns_3_2_1_U13.top_add_3ns_3ns_3_2_1_Adder_9_U.sum_s1 ;
assign _085_ = \add_3ns_3ns_3_2_1_U13.top_add_3ns_3ns_3_2_1_Adder_9_U.u1.a  + \add_3ns_3ns_3_2_1_U13.top_add_3ns_3ns_3_2_1_Adder_9_U.u1.b ;
assign { \add_3ns_3ns_3_2_1_U13.top_add_3ns_3ns_3_2_1_Adder_9_U.u1.cout , \add_3ns_3ns_3_2_1_U13.top_add_3ns_3ns_3_2_1_Adder_9_U.u1.s  } = _085_ + \add_3ns_3ns_3_2_1_U13.top_add_3ns_3ns_3_2_1_Adder_9_U.u1.cin ;
assign _086_ = \add_3ns_3ns_3_2_1_U13.top_add_3ns_3ns_3_2_1_Adder_9_U.u2.a  + \add_3ns_3ns_3_2_1_U13.top_add_3ns_3ns_3_2_1_Adder_9_U.u2.b ;
assign { \add_3ns_3ns_3_2_1_U13.top_add_3ns_3ns_3_2_1_Adder_9_U.u2.cout , \add_3ns_3ns_3_2_1_U13.top_add_3ns_3ns_3_2_1_Adder_9_U.u2.s  } = _086_ + \add_3ns_3ns_3_2_1_U13.top_add_3ns_3ns_3_2_1_Adder_9_U.u2.cin ;
always @(posedge \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.clk )
\add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.bin_s1  <= _088_;
always @(posedge \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.clk )
\add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.ain_s1  <= _087_;
always @(posedge \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.clk )
\add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.sum_s1  <= _090_;
always @(posedge \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.clk )
\add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.carry_s1  <= _089_;
assign _088_ = \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.ce  ? \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.b [3:2] : \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.bin_s1 ;
assign _087_ = \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.ce  ? \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.a [3:2] : \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.ain_s1 ;
assign _089_ = \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.ce  ? \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.facout_s1  : \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.carry_s1 ;
assign _090_ = \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.ce  ? \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.fas_s1  : \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.sum_s1 ;
assign _091_ = \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.u1.a  + \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.u1.b ;
assign { \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.u1.cout , \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.u1.s  } = _091_ + \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.u1.cin ;
assign _092_ = \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.u2.a  + \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.u2.b ;
assign { \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.u2.cout , \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.u2.s  } = _092_ + \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.u2.cin ;
always @(posedge \add_4s_4s_4_2_1_U16.top_add_4s_4s_4_2_1_Adder_12_U.clk )
\add_4s_4s_4_2_1_U16.top_add_4s_4s_4_2_1_Adder_12_U.bin_s1  <= _094_;
always @(posedge \add_4s_4s_4_2_1_U16.top_add_4s_4s_4_2_1_Adder_12_U.clk )
\add_4s_4s_4_2_1_U16.top_add_4s_4s_4_2_1_Adder_12_U.ain_s1  <= _093_;
always @(posedge \add_4s_4s_4_2_1_U16.top_add_4s_4s_4_2_1_Adder_12_U.clk )
\add_4s_4s_4_2_1_U16.top_add_4s_4s_4_2_1_Adder_12_U.sum_s1  <= _096_;
always @(posedge \add_4s_4s_4_2_1_U16.top_add_4s_4s_4_2_1_Adder_12_U.clk )
\add_4s_4s_4_2_1_U16.top_add_4s_4s_4_2_1_Adder_12_U.carry_s1  <= _095_;
assign _094_ = \add_4s_4s_4_2_1_U16.top_add_4s_4s_4_2_1_Adder_12_U.ce  ? \add_4s_4s_4_2_1_U16.top_add_4s_4s_4_2_1_Adder_12_U.b [3:2] : \add_4s_4s_4_2_1_U16.top_add_4s_4s_4_2_1_Adder_12_U.bin_s1 ;
assign _093_ = \add_4s_4s_4_2_1_U16.top_add_4s_4s_4_2_1_Adder_12_U.ce  ? \add_4s_4s_4_2_1_U16.top_add_4s_4s_4_2_1_Adder_12_U.a [3:2] : \add_4s_4s_4_2_1_U16.top_add_4s_4s_4_2_1_Adder_12_U.ain_s1 ;
assign _095_ = \add_4s_4s_4_2_1_U16.top_add_4s_4s_4_2_1_Adder_12_U.ce  ? \add_4s_4s_4_2_1_U16.top_add_4s_4s_4_2_1_Adder_12_U.facout_s1  : \add_4s_4s_4_2_1_U16.top_add_4s_4s_4_2_1_Adder_12_U.carry_s1 ;
assign _096_ = \add_4s_4s_4_2_1_U16.top_add_4s_4s_4_2_1_Adder_12_U.ce  ? \add_4s_4s_4_2_1_U16.top_add_4s_4s_4_2_1_Adder_12_U.fas_s1  : \add_4s_4s_4_2_1_U16.top_add_4s_4s_4_2_1_Adder_12_U.sum_s1 ;
assign _097_ = \add_4s_4s_4_2_1_U16.top_add_4s_4s_4_2_1_Adder_12_U.u1.a  + \add_4s_4s_4_2_1_U16.top_add_4s_4s_4_2_1_Adder_12_U.u1.b ;
assign { \add_4s_4s_4_2_1_U16.top_add_4s_4s_4_2_1_Adder_12_U.u1.cout , \add_4s_4s_4_2_1_U16.top_add_4s_4s_4_2_1_Adder_12_U.u1.s  } = _097_ + \add_4s_4s_4_2_1_U16.top_add_4s_4s_4_2_1_Adder_12_U.u1.cin ;
assign _098_ = \add_4s_4s_4_2_1_U16.top_add_4s_4s_4_2_1_Adder_12_U.u2.a  + \add_4s_4s_4_2_1_U16.top_add_4s_4s_4_2_1_Adder_12_U.u2.b ;
assign { \add_4s_4s_4_2_1_U16.top_add_4s_4s_4_2_1_Adder_12_U.u2.cout , \add_4s_4s_4_2_1_U16.top_add_4s_4s_4_2_1_Adder_12_U.u2.s  } = _098_ + \add_4s_4s_4_2_1_U16.top_add_4s_4s_4_2_1_Adder_12_U.u2.cin ;
always @(posedge \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_5_U.clk )
\add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_5_U.bin_s1  <= _100_;
always @(posedge \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_5_U.clk )
\add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_5_U.ain_s1  <= _099_;
always @(posedge \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_5_U.clk )
\add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_5_U.sum_s1  <= _102_;
always @(posedge \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_5_U.clk )
\add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_5_U.carry_s1  <= _101_;
assign _100_ = \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_5_U.ce  ? \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_5_U.b [4:2] : \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_5_U.bin_s1 ;
assign _099_ = \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_5_U.ce  ? \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_5_U.a [4:2] : \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_5_U.ain_s1 ;
assign _101_ = \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_5_U.ce  ? \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_5_U.facout_s1  : \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_5_U.carry_s1 ;
assign _102_ = \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_5_U.ce  ? \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_5_U.fas_s1  : \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_5_U.sum_s1 ;
assign _103_ = \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_5_U.u1.a  + \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_5_U.u1.b ;
assign { \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_5_U.u1.cout , \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_5_U.u1.s  } = _103_ + \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_5_U.u1.cin ;
assign _104_ = \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_5_U.u2.a  + \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_5_U.u2.b ;
assign { \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_5_U.u2.cout , \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_5_U.u2.s  } = _104_ + \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_5_U.u2.cin ;
always @(posedge \add_6ns_6s_6_2_1_U15.top_add_6ns_6s_6_2_1_Adder_11_U.clk )
\add_6ns_6s_6_2_1_U15.top_add_6ns_6s_6_2_1_Adder_11_U.bin_s1  <= _106_;
always @(posedge \add_6ns_6s_6_2_1_U15.top_add_6ns_6s_6_2_1_Adder_11_U.clk )
\add_6ns_6s_6_2_1_U15.top_add_6ns_6s_6_2_1_Adder_11_U.ain_s1  <= _105_;
always @(posedge \add_6ns_6s_6_2_1_U15.top_add_6ns_6s_6_2_1_Adder_11_U.clk )
\add_6ns_6s_6_2_1_U15.top_add_6ns_6s_6_2_1_Adder_11_U.sum_s1  <= _108_;
always @(posedge \add_6ns_6s_6_2_1_U15.top_add_6ns_6s_6_2_1_Adder_11_U.clk )
\add_6ns_6s_6_2_1_U15.top_add_6ns_6s_6_2_1_Adder_11_U.carry_s1  <= _107_;
assign _106_ = \add_6ns_6s_6_2_1_U15.top_add_6ns_6s_6_2_1_Adder_11_U.ce  ? \add_6ns_6s_6_2_1_U15.top_add_6ns_6s_6_2_1_Adder_11_U.b [5:3] : \add_6ns_6s_6_2_1_U15.top_add_6ns_6s_6_2_1_Adder_11_U.bin_s1 ;
assign _105_ = \add_6ns_6s_6_2_1_U15.top_add_6ns_6s_6_2_1_Adder_11_U.ce  ? \add_6ns_6s_6_2_1_U15.top_add_6ns_6s_6_2_1_Adder_11_U.a [5:3] : \add_6ns_6s_6_2_1_U15.top_add_6ns_6s_6_2_1_Adder_11_U.ain_s1 ;
assign _107_ = \add_6ns_6s_6_2_1_U15.top_add_6ns_6s_6_2_1_Adder_11_U.ce  ? \add_6ns_6s_6_2_1_U15.top_add_6ns_6s_6_2_1_Adder_11_U.facout_s1  : \add_6ns_6s_6_2_1_U15.top_add_6ns_6s_6_2_1_Adder_11_U.carry_s1 ;
assign _108_ = \add_6ns_6s_6_2_1_U15.top_add_6ns_6s_6_2_1_Adder_11_U.ce  ? \add_6ns_6s_6_2_1_U15.top_add_6ns_6s_6_2_1_Adder_11_U.fas_s1  : \add_6ns_6s_6_2_1_U15.top_add_6ns_6s_6_2_1_Adder_11_U.sum_s1 ;
assign _109_ = \add_6ns_6s_6_2_1_U15.top_add_6ns_6s_6_2_1_Adder_11_U.u1.a  + \add_6ns_6s_6_2_1_U15.top_add_6ns_6s_6_2_1_Adder_11_U.u1.b ;
assign { \add_6ns_6s_6_2_1_U15.top_add_6ns_6s_6_2_1_Adder_11_U.u1.cout , \add_6ns_6s_6_2_1_U15.top_add_6ns_6s_6_2_1_Adder_11_U.u1.s  } = _109_ + \add_6ns_6s_6_2_1_U15.top_add_6ns_6s_6_2_1_Adder_11_U.u1.cin ;
assign _110_ = \add_6ns_6s_6_2_1_U15.top_add_6ns_6s_6_2_1_Adder_11_U.u2.a  + \add_6ns_6s_6_2_1_U15.top_add_6ns_6s_6_2_1_Adder_11_U.u2.b ;
assign { \add_6ns_6s_6_2_1_U15.top_add_6ns_6s_6_2_1_Adder_11_U.u2.cout , \add_6ns_6s_6_2_1_U15.top_add_6ns_6s_6_2_1_Adder_11_U.u2.s  } = _110_ + \add_6ns_6s_6_2_1_U15.top_add_6ns_6s_6_2_1_Adder_11_U.u2.cin ;
always @(posedge \add_6s_6ns_6_2_1_U18.top_add_6s_6ns_6_2_1_Adder_14_U.clk )
\add_6s_6ns_6_2_1_U18.top_add_6s_6ns_6_2_1_Adder_14_U.bin_s1  <= _112_;
always @(posedge \add_6s_6ns_6_2_1_U18.top_add_6s_6ns_6_2_1_Adder_14_U.clk )
\add_6s_6ns_6_2_1_U18.top_add_6s_6ns_6_2_1_Adder_14_U.ain_s1  <= _111_;
always @(posedge \add_6s_6ns_6_2_1_U18.top_add_6s_6ns_6_2_1_Adder_14_U.clk )
\add_6s_6ns_6_2_1_U18.top_add_6s_6ns_6_2_1_Adder_14_U.sum_s1  <= _114_;
always @(posedge \add_6s_6ns_6_2_1_U18.top_add_6s_6ns_6_2_1_Adder_14_U.clk )
\add_6s_6ns_6_2_1_U18.top_add_6s_6ns_6_2_1_Adder_14_U.carry_s1  <= _113_;
assign _112_ = \add_6s_6ns_6_2_1_U18.top_add_6s_6ns_6_2_1_Adder_14_U.ce  ? \add_6s_6ns_6_2_1_U18.top_add_6s_6ns_6_2_1_Adder_14_U.b [5:3] : \add_6s_6ns_6_2_1_U18.top_add_6s_6ns_6_2_1_Adder_14_U.bin_s1 ;
assign _111_ = \add_6s_6ns_6_2_1_U18.top_add_6s_6ns_6_2_1_Adder_14_U.ce  ? \add_6s_6ns_6_2_1_U18.top_add_6s_6ns_6_2_1_Adder_14_U.a [5:3] : \add_6s_6ns_6_2_1_U18.top_add_6s_6ns_6_2_1_Adder_14_U.ain_s1 ;
assign _113_ = \add_6s_6ns_6_2_1_U18.top_add_6s_6ns_6_2_1_Adder_14_U.ce  ? \add_6s_6ns_6_2_1_U18.top_add_6s_6ns_6_2_1_Adder_14_U.facout_s1  : \add_6s_6ns_6_2_1_U18.top_add_6s_6ns_6_2_1_Adder_14_U.carry_s1 ;
assign _114_ = \add_6s_6ns_6_2_1_U18.top_add_6s_6ns_6_2_1_Adder_14_U.ce  ? \add_6s_6ns_6_2_1_U18.top_add_6s_6ns_6_2_1_Adder_14_U.fas_s1  : \add_6s_6ns_6_2_1_U18.top_add_6s_6ns_6_2_1_Adder_14_U.sum_s1 ;
assign _115_ = \add_6s_6ns_6_2_1_U18.top_add_6s_6ns_6_2_1_Adder_14_U.u1.a  + \add_6s_6ns_6_2_1_U18.top_add_6s_6ns_6_2_1_Adder_14_U.u1.b ;
assign { \add_6s_6ns_6_2_1_U18.top_add_6s_6ns_6_2_1_Adder_14_U.u1.cout , \add_6s_6ns_6_2_1_U18.top_add_6s_6ns_6_2_1_Adder_14_U.u1.s  } = _115_ + \add_6s_6ns_6_2_1_U18.top_add_6s_6ns_6_2_1_Adder_14_U.u1.cin ;
assign _116_ = \add_6s_6ns_6_2_1_U18.top_add_6s_6ns_6_2_1_Adder_14_U.u2.a  + \add_6s_6ns_6_2_1_U18.top_add_6s_6ns_6_2_1_Adder_14_U.u2.b ;
assign { \add_6s_6ns_6_2_1_U18.top_add_6s_6ns_6_2_1_Adder_14_U.u2.cout , \add_6s_6ns_6_2_1_U18.top_add_6s_6ns_6_2_1_Adder_14_U.u2.s  } = _116_ + \add_6s_6ns_6_2_1_U18.top_add_6s_6ns_6_2_1_Adder_14_U.u2.cin ;
always @(posedge \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_8_U.clk )
\add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_8_U.bin_s1  <= _118_;
always @(posedge \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_8_U.clk )
\add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_8_U.ain_s1  <= _117_;
always @(posedge \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_8_U.clk )
\add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_8_U.sum_s1  <= _120_;
always @(posedge \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_8_U.clk )
\add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_8_U.carry_s1  <= _119_;
assign _118_ = \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_8_U.ce  ? \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_8_U.b [6:3] : \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_8_U.bin_s1 ;
assign _117_ = \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_8_U.ce  ? \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_8_U.a [6:3] : \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_8_U.ain_s1 ;
assign _119_ = \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_8_U.ce  ? \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_8_U.facout_s1  : \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_8_U.carry_s1 ;
assign _120_ = \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_8_U.ce  ? \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_8_U.fas_s1  : \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_8_U.sum_s1 ;
assign _121_ = \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_8_U.u1.a  + \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_8_U.u1.b ;
assign { \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_8_U.u1.cout , \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_8_U.u1.s  } = _121_ + \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_8_U.u1.cin ;
assign _122_ = \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_8_U.u2.a  + \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_8_U.u2.b ;
assign { \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_8_U.u2.cout , \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_8_U.u2.s  } = _122_ + \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_8_U.u2.cin ;
always @(posedge \add_7s_7s_7_2_1_U10.top_add_7s_7s_7_2_1_Adder_6_U.clk )
\add_7s_7s_7_2_1_U10.top_add_7s_7s_7_2_1_Adder_6_U.bin_s1  <= _124_;
always @(posedge \add_7s_7s_7_2_1_U10.top_add_7s_7s_7_2_1_Adder_6_U.clk )
\add_7s_7s_7_2_1_U10.top_add_7s_7s_7_2_1_Adder_6_U.ain_s1  <= _123_;
always @(posedge \add_7s_7s_7_2_1_U10.top_add_7s_7s_7_2_1_Adder_6_U.clk )
\add_7s_7s_7_2_1_U10.top_add_7s_7s_7_2_1_Adder_6_U.sum_s1  <= _126_;
always @(posedge \add_7s_7s_7_2_1_U10.top_add_7s_7s_7_2_1_Adder_6_U.clk )
\add_7s_7s_7_2_1_U10.top_add_7s_7s_7_2_1_Adder_6_U.carry_s1  <= _125_;
assign _124_ = \add_7s_7s_7_2_1_U10.top_add_7s_7s_7_2_1_Adder_6_U.ce  ? \add_7s_7s_7_2_1_U10.top_add_7s_7s_7_2_1_Adder_6_U.b [6:3] : \add_7s_7s_7_2_1_U10.top_add_7s_7s_7_2_1_Adder_6_U.bin_s1 ;
assign _123_ = \add_7s_7s_7_2_1_U10.top_add_7s_7s_7_2_1_Adder_6_U.ce  ? \add_7s_7s_7_2_1_U10.top_add_7s_7s_7_2_1_Adder_6_U.a [6:3] : \add_7s_7s_7_2_1_U10.top_add_7s_7s_7_2_1_Adder_6_U.ain_s1 ;
assign _125_ = \add_7s_7s_7_2_1_U10.top_add_7s_7s_7_2_1_Adder_6_U.ce  ? \add_7s_7s_7_2_1_U10.top_add_7s_7s_7_2_1_Adder_6_U.facout_s1  : \add_7s_7s_7_2_1_U10.top_add_7s_7s_7_2_1_Adder_6_U.carry_s1 ;
assign _126_ = \add_7s_7s_7_2_1_U10.top_add_7s_7s_7_2_1_Adder_6_U.ce  ? \add_7s_7s_7_2_1_U10.top_add_7s_7s_7_2_1_Adder_6_U.fas_s1  : \add_7s_7s_7_2_1_U10.top_add_7s_7s_7_2_1_Adder_6_U.sum_s1 ;
assign _127_ = \add_7s_7s_7_2_1_U10.top_add_7s_7s_7_2_1_Adder_6_U.u1.a  + \add_7s_7s_7_2_1_U10.top_add_7s_7s_7_2_1_Adder_6_U.u1.b ;
assign { \add_7s_7s_7_2_1_U10.top_add_7s_7s_7_2_1_Adder_6_U.u1.cout , \add_7s_7s_7_2_1_U10.top_add_7s_7s_7_2_1_Adder_6_U.u1.s  } = _127_ + \add_7s_7s_7_2_1_U10.top_add_7s_7s_7_2_1_Adder_6_U.u1.cin ;
assign _128_ = \add_7s_7s_7_2_1_U10.top_add_7s_7s_7_2_1_Adder_6_U.u2.a  + \add_7s_7s_7_2_1_U10.top_add_7s_7s_7_2_1_Adder_6_U.u2.b ;
assign { \add_7s_7s_7_2_1_U10.top_add_7s_7s_7_2_1_Adder_6_U.u2.cout , \add_7s_7s_7_2_1_U10.top_add_7s_7s_7_2_1_Adder_6_U.u2.s  } = _128_ + \add_7s_7s_7_2_1_U10.top_add_7s_7s_7_2_1_Adder_6_U.u2.cin ;
always @(posedge \add_9ns_9ns_9_2_1_U17.top_add_9ns_9ns_9_2_1_Adder_13_U.clk )
\add_9ns_9ns_9_2_1_U17.top_add_9ns_9ns_9_2_1_Adder_13_U.bin_s1  <= _130_;
always @(posedge \add_9ns_9ns_9_2_1_U17.top_add_9ns_9ns_9_2_1_Adder_13_U.clk )
\add_9ns_9ns_9_2_1_U17.top_add_9ns_9ns_9_2_1_Adder_13_U.ain_s1  <= _129_;
always @(posedge \add_9ns_9ns_9_2_1_U17.top_add_9ns_9ns_9_2_1_Adder_13_U.clk )
\add_9ns_9ns_9_2_1_U17.top_add_9ns_9ns_9_2_1_Adder_13_U.sum_s1  <= _132_;
always @(posedge \add_9ns_9ns_9_2_1_U17.top_add_9ns_9ns_9_2_1_Adder_13_U.clk )
\add_9ns_9ns_9_2_1_U17.top_add_9ns_9ns_9_2_1_Adder_13_U.carry_s1  <= _131_;
assign _130_ = \add_9ns_9ns_9_2_1_U17.top_add_9ns_9ns_9_2_1_Adder_13_U.ce  ? \add_9ns_9ns_9_2_1_U17.top_add_9ns_9ns_9_2_1_Adder_13_U.b [8:4] : \add_9ns_9ns_9_2_1_U17.top_add_9ns_9ns_9_2_1_Adder_13_U.bin_s1 ;
assign _129_ = \add_9ns_9ns_9_2_1_U17.top_add_9ns_9ns_9_2_1_Adder_13_U.ce  ? \add_9ns_9ns_9_2_1_U17.top_add_9ns_9ns_9_2_1_Adder_13_U.a [8:4] : \add_9ns_9ns_9_2_1_U17.top_add_9ns_9ns_9_2_1_Adder_13_U.ain_s1 ;
assign _131_ = \add_9ns_9ns_9_2_1_U17.top_add_9ns_9ns_9_2_1_Adder_13_U.ce  ? \add_9ns_9ns_9_2_1_U17.top_add_9ns_9ns_9_2_1_Adder_13_U.facout_s1  : \add_9ns_9ns_9_2_1_U17.top_add_9ns_9ns_9_2_1_Adder_13_U.carry_s1 ;
assign _132_ = \add_9ns_9ns_9_2_1_U17.top_add_9ns_9ns_9_2_1_Adder_13_U.ce  ? \add_9ns_9ns_9_2_1_U17.top_add_9ns_9ns_9_2_1_Adder_13_U.fas_s1  : \add_9ns_9ns_9_2_1_U17.top_add_9ns_9ns_9_2_1_Adder_13_U.sum_s1 ;
assign _133_ = \add_9ns_9ns_9_2_1_U17.top_add_9ns_9ns_9_2_1_Adder_13_U.u1.a  + \add_9ns_9ns_9_2_1_U17.top_add_9ns_9ns_9_2_1_Adder_13_U.u1.b ;
assign { \add_9ns_9ns_9_2_1_U17.top_add_9ns_9ns_9_2_1_Adder_13_U.u1.cout , \add_9ns_9ns_9_2_1_U17.top_add_9ns_9ns_9_2_1_Adder_13_U.u1.s  } = _133_ + \add_9ns_9ns_9_2_1_U17.top_add_9ns_9ns_9_2_1_Adder_13_U.u1.cin ;
assign _134_ = \add_9ns_9ns_9_2_1_U17.top_add_9ns_9ns_9_2_1_Adder_13_U.u2.a  + \add_9ns_9ns_9_2_1_U17.top_add_9ns_9ns_9_2_1_Adder_13_U.u2.b ;
assign { \add_9ns_9ns_9_2_1_U17.top_add_9ns_9ns_9_2_1_Adder_13_U.u2.cout , \add_9ns_9ns_9_2_1_U17.top_add_9ns_9ns_9_2_1_Adder_13_U.u2.s  } = _134_ + \add_9ns_9ns_9_2_1_U17.top_add_9ns_9ns_9_2_1_Adder_13_U.u2.cin ;
always @(posedge \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_15_U.clk )
\add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_15_U.bin_s1  <= _136_;
always @(posedge \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_15_U.clk )
\add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_15_U.ain_s1  <= _135_;
always @(posedge \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_15_U.clk )
\add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_15_U.sum_s1  <= _138_;
always @(posedge \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_15_U.clk )
\add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_15_U.carry_s1  <= _137_;
assign _136_ = \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_15_U.ce  ? \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_15_U.b [8:4] : \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_15_U.bin_s1 ;
assign _135_ = \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_15_U.ce  ? \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_15_U.a [8:4] : \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_15_U.ain_s1 ;
assign _137_ = \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_15_U.ce  ? \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_15_U.facout_s1  : \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_15_U.carry_s1 ;
assign _138_ = \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_15_U.ce  ? \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_15_U.fas_s1  : \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_15_U.sum_s1 ;
assign _139_ = \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_15_U.u1.a  + \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_15_U.u1.b ;
assign { \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_15_U.u1.cout , \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_15_U.u1.s  } = _139_ + \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_15_U.u1.cin ;
assign _140_ = \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_15_U.u2.a  + \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_15_U.u2.b ;
assign { \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_15_U.u2.cout , \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_15_U.u2.s  } = _140_ + \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_15_U.u2.cin ;
always @(posedge \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_10_U.clk )
\add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_10_U.bin_s1  <= _142_;
always @(posedge \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_10_U.clk )
\add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_10_U.ain_s1  <= _141_;
always @(posedge \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_10_U.clk )
\add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_10_U.sum_s1  <= _144_;
always @(posedge \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_10_U.clk )
\add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_10_U.carry_s1  <= _143_;
assign _142_ = \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_10_U.ce  ? \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_10_U.b [8:4] : \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_10_U.bin_s1 ;
assign _141_ = \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_10_U.ce  ? \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_10_U.a [8:4] : \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_10_U.ain_s1 ;
assign _143_ = \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_10_U.ce  ? \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_10_U.facout_s1  : \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_10_U.carry_s1 ;
assign _144_ = \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_10_U.ce  ? \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_10_U.fas_s1  : \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_10_U.sum_s1 ;
assign _145_ = \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_10_U.u1.a  + \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_10_U.u1.b ;
assign { \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_10_U.u1.cout , \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_10_U.u1.s  } = _145_ + \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_10_U.u1.cin ;
assign _146_ = \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_10_U.u2.a  + \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_10_U.u2.b ;
assign { \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_10_U.u2.cout , \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_10_U.u2.s  } = _146_ + \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_10_U.u2.cin ;
always @(posedge \lshr_32ns_32s_32_7_1_U9.clk )
\lshr_32ns_32s_32_7_1_U9.dout_array[5]  <= _158_;
always @(posedge \lshr_32ns_32s_32_7_1_U9.clk )
\lshr_32ns_32s_32_7_1_U9.din1_cast_array[5]  <= _152_;
always @(posedge \lshr_32ns_32s_32_7_1_U9.clk )
\lshr_32ns_32s_32_7_1_U9.dout_array[4]  <= _157_;
always @(posedge \lshr_32ns_32s_32_7_1_U9.clk )
\lshr_32ns_32s_32_7_1_U9.din1_cast_array[4]  <= _151_;
always @(posedge \lshr_32ns_32s_32_7_1_U9.clk )
\lshr_32ns_32s_32_7_1_U9.dout_array[3]  <= _156_;
always @(posedge \lshr_32ns_32s_32_7_1_U9.clk )
\lshr_32ns_32s_32_7_1_U9.din1_cast_array[3]  <= _150_;
always @(posedge \lshr_32ns_32s_32_7_1_U9.clk )
\lshr_32ns_32s_32_7_1_U9.dout_array[2]  <= _155_;
always @(posedge \lshr_32ns_32s_32_7_1_U9.clk )
\lshr_32ns_32s_32_7_1_U9.din1_cast_array[2]  <= _149_;
always @(posedge \lshr_32ns_32s_32_7_1_U9.clk )
\lshr_32ns_32s_32_7_1_U9.dout_array[1]  <= _154_;
always @(posedge \lshr_32ns_32s_32_7_1_U9.clk )
\lshr_32ns_32s_32_7_1_U9.din1_cast_array[1]  <= _148_;
always @(posedge \lshr_32ns_32s_32_7_1_U9.clk )
\lshr_32ns_32s_32_7_1_U9.dout_array[0]  <= _153_;
always @(posedge \lshr_32ns_32s_32_7_1_U9.clk )
\lshr_32ns_32s_32_7_1_U9.din1_cast_array[0]  <= _147_;
assign _159_ = \lshr_32ns_32s_32_7_1_U9.ce  ? \lshr_32ns_32s_32_7_1_U9.din1_cast_array[4]  : \lshr_32ns_32s_32_7_1_U9.din1_cast_array[5] ;
assign _152_ = \lshr_32ns_32s_32_7_1_U9.reset  ? 32'd0 : _159_;
assign _160_ = \lshr_32ns_32s_32_7_1_U9.ce  ? _176_ : \lshr_32ns_32s_32_7_1_U9.dout_array[5] ;
assign _158_ = \lshr_32ns_32s_32_7_1_U9.reset  ? 32'd0 : _160_;
assign _161_ = \lshr_32ns_32s_32_7_1_U9.ce  ? \lshr_32ns_32s_32_7_1_U9.din1_cast_array[3]  : \lshr_32ns_32s_32_7_1_U9.din1_cast_array[4] ;
assign _151_ = \lshr_32ns_32s_32_7_1_U9.reset  ? 32'd0 : _161_;
assign _162_ = \lshr_32ns_32s_32_7_1_U9.ce  ? _175_ : \lshr_32ns_32s_32_7_1_U9.dout_array[4] ;
assign _157_ = \lshr_32ns_32s_32_7_1_U9.reset  ? 32'd0 : _162_;
assign _163_ = \lshr_32ns_32s_32_7_1_U9.ce  ? \lshr_32ns_32s_32_7_1_U9.din1_cast_array[2]  : \lshr_32ns_32s_32_7_1_U9.din1_cast_array[3] ;
assign _150_ = \lshr_32ns_32s_32_7_1_U9.reset  ? 32'd0 : _163_;
assign _164_ = \lshr_32ns_32s_32_7_1_U9.ce  ? _174_ : \lshr_32ns_32s_32_7_1_U9.dout_array[3] ;
assign _156_ = \lshr_32ns_32s_32_7_1_U9.reset  ? 32'd0 : _164_;
assign _165_ = \lshr_32ns_32s_32_7_1_U9.ce  ? \lshr_32ns_32s_32_7_1_U9.din1_cast_array[1]  : \lshr_32ns_32s_32_7_1_U9.din1_cast_array[2] ;
assign _149_ = \lshr_32ns_32s_32_7_1_U9.reset  ? 32'd0 : _165_;
assign _166_ = \lshr_32ns_32s_32_7_1_U9.ce  ? _173_ : \lshr_32ns_32s_32_7_1_U9.dout_array[2] ;
assign _155_ = \lshr_32ns_32s_32_7_1_U9.reset  ? 32'd0 : _166_;
assign _167_ = \lshr_32ns_32s_32_7_1_U9.ce  ? \lshr_32ns_32s_32_7_1_U9.din1_cast_array[0]  : \lshr_32ns_32s_32_7_1_U9.din1_cast_array[1] ;
assign _148_ = \lshr_32ns_32s_32_7_1_U9.reset  ? 32'd0 : _167_;
assign _168_ = \lshr_32ns_32s_32_7_1_U9.ce  ? _172_ : \lshr_32ns_32s_32_7_1_U9.dout_array[1] ;
assign _154_ = \lshr_32ns_32s_32_7_1_U9.reset  ? 32'd0 : _168_;
assign _169_ = \lshr_32ns_32s_32_7_1_U9.ce  ? \lshr_32ns_32s_32_7_1_U9.din1  : \lshr_32ns_32s_32_7_1_U9.din1_cast_array[0] ;
assign _147_ = \lshr_32ns_32s_32_7_1_U9.reset  ? 32'd0 : _169_;
assign _170_ = \lshr_32ns_32s_32_7_1_U9.ce  ? _171_ : \lshr_32ns_32s_32_7_1_U9.dout_array[0] ;
assign _153_ = \lshr_32ns_32s_32_7_1_U9.reset  ? 32'd0 : _170_;
assign _171_ = \lshr_32ns_32s_32_7_1_U9.din0  >> { \lshr_32ns_32s_32_7_1_U9.din1 [31:30], 30'h00000000 };
assign _172_ = \lshr_32ns_32s_32_7_1_U9.dout_array[0]  >> { \lshr_32ns_32s_32_7_1_U9.din1_cast_array[0] [29:25], 25'h0000000 };
assign _173_ = \lshr_32ns_32s_32_7_1_U9.dout_array[1]  >> { \lshr_32ns_32s_32_7_1_U9.din1_cast_array[1] [24:20], 20'h00000 };
assign _174_ = \lshr_32ns_32s_32_7_1_U9.dout_array[2]  >> { \lshr_32ns_32s_32_7_1_U9.din1_cast_array[2] [19:15], 15'h0000 };
assign _175_ = \lshr_32ns_32s_32_7_1_U9.dout_array[3]  >> { \lshr_32ns_32s_32_7_1_U9.din1_cast_array[3] [14:10], 10'h000 };
assign _176_ = \lshr_32ns_32s_32_7_1_U9.dout_array[4]  >> { \lshr_32ns_32s_32_7_1_U9.din1_cast_array[4] [9:5], 5'h00 };
assign \lshr_32ns_32s_32_7_1_U9.dout  = \lshr_32ns_32s_32_7_1_U9.dout_array[5]  >> \lshr_32ns_32s_32_7_1_U9.din1_cast_array[5] [4:0];
always @(posedge \shl_32ns_32s_32_7_1_U8.clk )
\shl_32ns_32s_32_7_1_U8.dout_array[5]  <= _188_;
always @(posedge \shl_32ns_32s_32_7_1_U8.clk )
\shl_32ns_32s_32_7_1_U8.din1_cast_array[5]  <= _182_;
always @(posedge \shl_32ns_32s_32_7_1_U8.clk )
\shl_32ns_32s_32_7_1_U8.dout_array[4]  <= _187_;
always @(posedge \shl_32ns_32s_32_7_1_U8.clk )
\shl_32ns_32s_32_7_1_U8.din1_cast_array[4]  <= _181_;
always @(posedge \shl_32ns_32s_32_7_1_U8.clk )
\shl_32ns_32s_32_7_1_U8.dout_array[3]  <= _186_;
always @(posedge \shl_32ns_32s_32_7_1_U8.clk )
\shl_32ns_32s_32_7_1_U8.din1_cast_array[3]  <= _180_;
always @(posedge \shl_32ns_32s_32_7_1_U8.clk )
\shl_32ns_32s_32_7_1_U8.dout_array[2]  <= _185_;
always @(posedge \shl_32ns_32s_32_7_1_U8.clk )
\shl_32ns_32s_32_7_1_U8.din1_cast_array[2]  <= _179_;
always @(posedge \shl_32ns_32s_32_7_1_U8.clk )
\shl_32ns_32s_32_7_1_U8.dout_array[1]  <= _184_;
always @(posedge \shl_32ns_32s_32_7_1_U8.clk )
\shl_32ns_32s_32_7_1_U8.din1_cast_array[1]  <= _178_;
always @(posedge \shl_32ns_32s_32_7_1_U8.clk )
\shl_32ns_32s_32_7_1_U8.dout_array[0]  <= _183_;
always @(posedge \shl_32ns_32s_32_7_1_U8.clk )
\shl_32ns_32s_32_7_1_U8.din1_cast_array[0]  <= _177_;
assign _189_ = \shl_32ns_32s_32_7_1_U8.ce  ? \shl_32ns_32s_32_7_1_U8.din1_cast_array[4]  : \shl_32ns_32s_32_7_1_U8.din1_cast_array[5] ;
assign _182_ = \shl_32ns_32s_32_7_1_U8.reset  ? 32'd0 : _189_;
assign _190_ = \shl_32ns_32s_32_7_1_U8.ce  ? _206_ : \shl_32ns_32s_32_7_1_U8.dout_array[5] ;
assign _188_ = \shl_32ns_32s_32_7_1_U8.reset  ? 32'd0 : _190_;
assign _191_ = \shl_32ns_32s_32_7_1_U8.ce  ? \shl_32ns_32s_32_7_1_U8.din1_cast_array[3]  : \shl_32ns_32s_32_7_1_U8.din1_cast_array[4] ;
assign _181_ = \shl_32ns_32s_32_7_1_U8.reset  ? 32'd0 : _191_;
assign _192_ = \shl_32ns_32s_32_7_1_U8.ce  ? _205_ : \shl_32ns_32s_32_7_1_U8.dout_array[4] ;
assign _187_ = \shl_32ns_32s_32_7_1_U8.reset  ? 32'd0 : _192_;
assign _193_ = \shl_32ns_32s_32_7_1_U8.ce  ? \shl_32ns_32s_32_7_1_U8.din1_cast_array[2]  : \shl_32ns_32s_32_7_1_U8.din1_cast_array[3] ;
assign _180_ = \shl_32ns_32s_32_7_1_U8.reset  ? 32'd0 : _193_;
assign _194_ = \shl_32ns_32s_32_7_1_U8.ce  ? _204_ : \shl_32ns_32s_32_7_1_U8.dout_array[3] ;
assign _186_ = \shl_32ns_32s_32_7_1_U8.reset  ? 32'd0 : _194_;
assign _195_ = \shl_32ns_32s_32_7_1_U8.ce  ? \shl_32ns_32s_32_7_1_U8.din1_cast_array[1]  : \shl_32ns_32s_32_7_1_U8.din1_cast_array[2] ;
assign _179_ = \shl_32ns_32s_32_7_1_U8.reset  ? 32'd0 : _195_;
assign _196_ = \shl_32ns_32s_32_7_1_U8.ce  ? _203_ : \shl_32ns_32s_32_7_1_U8.dout_array[2] ;
assign _185_ = \shl_32ns_32s_32_7_1_U8.reset  ? 32'd0 : _196_;
assign _197_ = \shl_32ns_32s_32_7_1_U8.ce  ? \shl_32ns_32s_32_7_1_U8.din1_cast_array[0]  : \shl_32ns_32s_32_7_1_U8.din1_cast_array[1] ;
assign _178_ = \shl_32ns_32s_32_7_1_U8.reset  ? 32'd0 : _197_;
assign _198_ = \shl_32ns_32s_32_7_1_U8.ce  ? _202_ : \shl_32ns_32s_32_7_1_U8.dout_array[1] ;
assign _184_ = \shl_32ns_32s_32_7_1_U8.reset  ? 32'd0 : _198_;
assign _199_ = \shl_32ns_32s_32_7_1_U8.ce  ? \shl_32ns_32s_32_7_1_U8.din1  : \shl_32ns_32s_32_7_1_U8.din1_cast_array[0] ;
assign _177_ = \shl_32ns_32s_32_7_1_U8.reset  ? 32'd0 : _199_;
assign _200_ = \shl_32ns_32s_32_7_1_U8.ce  ? _201_ : \shl_32ns_32s_32_7_1_U8.dout_array[0] ;
assign _183_ = \shl_32ns_32s_32_7_1_U8.reset  ? 32'd0 : _200_;
assign _201_ = \shl_32ns_32s_32_7_1_U8.din0  << { \shl_32ns_32s_32_7_1_U8.din1 [31:30], 30'h00000000 };
assign _202_ = \shl_32ns_32s_32_7_1_U8.dout_array[0]  << { \shl_32ns_32s_32_7_1_U8.din1_cast_array[0] [29:25], 25'h0000000 };
assign _203_ = \shl_32ns_32s_32_7_1_U8.dout_array[1]  << { \shl_32ns_32s_32_7_1_U8.din1_cast_array[1] [24:20], 20'h00000 };
assign _204_ = \shl_32ns_32s_32_7_1_U8.dout_array[2]  << { \shl_32ns_32s_32_7_1_U8.din1_cast_array[2] [19:15], 15'h0000 };
assign _205_ = \shl_32ns_32s_32_7_1_U8.dout_array[3]  << { \shl_32ns_32s_32_7_1_U8.din1_cast_array[3] [14:10], 10'h000 };
assign _206_ = \shl_32ns_32s_32_7_1_U8.dout_array[4]  << { \shl_32ns_32s_32_7_1_U8.din1_cast_array[4] [9:5], 5'h00 };
assign \shl_32ns_32s_32_7_1_U8.dout  = \shl_32ns_32s_32_7_1_U8.dout_array[5]  << \shl_32ns_32s_32_7_1_U8.din1_cast_array[5] [4:0];
assign \sub_3ns_3s_3_2_1_U3.top_sub_3ns_3s_3_2_1_Adder_2_U.bin_s0  = ~ \sub_3ns_3s_3_2_1_U3.top_sub_3ns_3s_3_2_1_Adder_2_U.b ;
always @(posedge \sub_3ns_3s_3_2_1_U3.top_sub_3ns_3s_3_2_1_Adder_2_U.clk )
\sub_3ns_3s_3_2_1_U3.top_sub_3ns_3s_3_2_1_Adder_2_U.bin_s1  <= _208_;
always @(posedge \sub_3ns_3s_3_2_1_U3.top_sub_3ns_3s_3_2_1_Adder_2_U.clk )
\sub_3ns_3s_3_2_1_U3.top_sub_3ns_3s_3_2_1_Adder_2_U.ain_s1  <= _207_;
always @(posedge \sub_3ns_3s_3_2_1_U3.top_sub_3ns_3s_3_2_1_Adder_2_U.clk )
\sub_3ns_3s_3_2_1_U3.top_sub_3ns_3s_3_2_1_Adder_2_U.sum_s1  <= _210_;
always @(posedge \sub_3ns_3s_3_2_1_U3.top_sub_3ns_3s_3_2_1_Adder_2_U.clk )
\sub_3ns_3s_3_2_1_U3.top_sub_3ns_3s_3_2_1_Adder_2_U.carry_s1  <= _209_;
assign _208_ = \sub_3ns_3s_3_2_1_U3.top_sub_3ns_3s_3_2_1_Adder_2_U.ce  ? \sub_3ns_3s_3_2_1_U3.top_sub_3ns_3s_3_2_1_Adder_2_U.bin_s0 [2:1] : \sub_3ns_3s_3_2_1_U3.top_sub_3ns_3s_3_2_1_Adder_2_U.bin_s1 ;
assign _207_ = \sub_3ns_3s_3_2_1_U3.top_sub_3ns_3s_3_2_1_Adder_2_U.ce  ? \sub_3ns_3s_3_2_1_U3.top_sub_3ns_3s_3_2_1_Adder_2_U.a [2:1] : \sub_3ns_3s_3_2_1_U3.top_sub_3ns_3s_3_2_1_Adder_2_U.ain_s1 ;
assign _209_ = \sub_3ns_3s_3_2_1_U3.top_sub_3ns_3s_3_2_1_Adder_2_U.ce  ? \sub_3ns_3s_3_2_1_U3.top_sub_3ns_3s_3_2_1_Adder_2_U.facout_s1  : \sub_3ns_3s_3_2_1_U3.top_sub_3ns_3s_3_2_1_Adder_2_U.carry_s1 ;
assign _210_ = \sub_3ns_3s_3_2_1_U3.top_sub_3ns_3s_3_2_1_Adder_2_U.ce  ? \sub_3ns_3s_3_2_1_U3.top_sub_3ns_3s_3_2_1_Adder_2_U.fas_s1  : \sub_3ns_3s_3_2_1_U3.top_sub_3ns_3s_3_2_1_Adder_2_U.sum_s1 ;
assign _211_ = \sub_3ns_3s_3_2_1_U3.top_sub_3ns_3s_3_2_1_Adder_2_U.u1.a  + \sub_3ns_3s_3_2_1_U3.top_sub_3ns_3s_3_2_1_Adder_2_U.u1.b ;
assign { \sub_3ns_3s_3_2_1_U3.top_sub_3ns_3s_3_2_1_Adder_2_U.u1.cout , \sub_3ns_3s_3_2_1_U3.top_sub_3ns_3s_3_2_1_Adder_2_U.u1.s  } = _211_ + \sub_3ns_3s_3_2_1_U3.top_sub_3ns_3s_3_2_1_Adder_2_U.u1.cin ;
assign _212_ = \sub_3ns_3s_3_2_1_U3.top_sub_3ns_3s_3_2_1_Adder_2_U.u2.a  + \sub_3ns_3s_3_2_1_U3.top_sub_3ns_3s_3_2_1_Adder_2_U.u2.b ;
assign { \sub_3ns_3s_3_2_1_U3.top_sub_3ns_3s_3_2_1_Adder_2_U.u2.cout , \sub_3ns_3s_3_2_1_U3.top_sub_3ns_3s_3_2_1_Adder_2_U.u2.s  } = _212_ + \sub_3ns_3s_3_2_1_U3.top_sub_3ns_3s_3_2_1_Adder_2_U.u2.cin ;
assign \sub_9ns_9s_9_2_1_U11.top_sub_9ns_9s_9_2_1_Adder_7_U.bin_s0  = ~ \sub_9ns_9s_9_2_1_U11.top_sub_9ns_9s_9_2_1_Adder_7_U.b ;
always @(posedge \sub_9ns_9s_9_2_1_U11.top_sub_9ns_9s_9_2_1_Adder_7_U.clk )
\sub_9ns_9s_9_2_1_U11.top_sub_9ns_9s_9_2_1_Adder_7_U.bin_s1  <= _214_;
always @(posedge \sub_9ns_9s_9_2_1_U11.top_sub_9ns_9s_9_2_1_Adder_7_U.clk )
\sub_9ns_9s_9_2_1_U11.top_sub_9ns_9s_9_2_1_Adder_7_U.ain_s1  <= _213_;
always @(posedge \sub_9ns_9s_9_2_1_U11.top_sub_9ns_9s_9_2_1_Adder_7_U.clk )
\sub_9ns_9s_9_2_1_U11.top_sub_9ns_9s_9_2_1_Adder_7_U.sum_s1  <= _216_;
always @(posedge \sub_9ns_9s_9_2_1_U11.top_sub_9ns_9s_9_2_1_Adder_7_U.clk )
\sub_9ns_9s_9_2_1_U11.top_sub_9ns_9s_9_2_1_Adder_7_U.carry_s1  <= _215_;
assign _214_ = \sub_9ns_9s_9_2_1_U11.top_sub_9ns_9s_9_2_1_Adder_7_U.ce  ? \sub_9ns_9s_9_2_1_U11.top_sub_9ns_9s_9_2_1_Adder_7_U.bin_s0 [8:4] : \sub_9ns_9s_9_2_1_U11.top_sub_9ns_9s_9_2_1_Adder_7_U.bin_s1 ;
assign _213_ = \sub_9ns_9s_9_2_1_U11.top_sub_9ns_9s_9_2_1_Adder_7_U.ce  ? \sub_9ns_9s_9_2_1_U11.top_sub_9ns_9s_9_2_1_Adder_7_U.a [8:4] : \sub_9ns_9s_9_2_1_U11.top_sub_9ns_9s_9_2_1_Adder_7_U.ain_s1 ;
assign _215_ = \sub_9ns_9s_9_2_1_U11.top_sub_9ns_9s_9_2_1_Adder_7_U.ce  ? \sub_9ns_9s_9_2_1_U11.top_sub_9ns_9s_9_2_1_Adder_7_U.facout_s1  : \sub_9ns_9s_9_2_1_U11.top_sub_9ns_9s_9_2_1_Adder_7_U.carry_s1 ;
assign _216_ = \sub_9ns_9s_9_2_1_U11.top_sub_9ns_9s_9_2_1_Adder_7_U.ce  ? \sub_9ns_9s_9_2_1_U11.top_sub_9ns_9s_9_2_1_Adder_7_U.fas_s1  : \sub_9ns_9s_9_2_1_U11.top_sub_9ns_9s_9_2_1_Adder_7_U.sum_s1 ;
assign _217_ = \sub_9ns_9s_9_2_1_U11.top_sub_9ns_9s_9_2_1_Adder_7_U.u1.a  + \sub_9ns_9s_9_2_1_U11.top_sub_9ns_9s_9_2_1_Adder_7_U.u1.b ;
assign { \sub_9ns_9s_9_2_1_U11.top_sub_9ns_9s_9_2_1_Adder_7_U.u1.cout , \sub_9ns_9s_9_2_1_U11.top_sub_9ns_9s_9_2_1_Adder_7_U.u1.s  } = _217_ + \sub_9ns_9s_9_2_1_U11.top_sub_9ns_9s_9_2_1_Adder_7_U.u1.cin ;
assign _218_ = \sub_9ns_9s_9_2_1_U11.top_sub_9ns_9s_9_2_1_Adder_7_U.u2.a  + \sub_9ns_9s_9_2_1_U11.top_sub_9ns_9s_9_2_1_Adder_7_U.u2.b ;
assign { \sub_9ns_9s_9_2_1_U11.top_sub_9ns_9s_9_2_1_Adder_7_U.u2.cout , \sub_9ns_9s_9_2_1_U11.top_sub_9ns_9s_9_2_1_Adder_7_U.u2.s  } = _218_ + \sub_9ns_9s_9_2_1_U11.top_sub_9ns_9s_9_2_1_Adder_7_U.u2.cin ;
always @(posedge ap_clk)
select_ln703_reg_823[5:0] <= 6'h00;
always @(posedge ap_clk)
select_ln69_reg_952[8:2] <= 7'h00;
always @(posedge ap_clk)
trunc_ln1497_reg_887 <= _041_;
always @(posedge ap_clk)
trunc_ln1497_1_reg_892 <= _040_;
always @(posedge ap_clk)
sub_ln1497_reg_753 <= _037_;
always @(posedge ap_clk)
select_ln850_7_reg_818 <= _035_;
always @(posedge ap_clk)
select_ln703_reg_823[8:6] <= _034_;
always @(posedge ap_clk)
ret_V_9_reg_680 <= _031_;
always @(posedge ap_clk)
tmp_4_reg_686 <= _039_;
always @(posedge ap_clk)
ret_V_8_reg_675 <= _030_;
always @(posedge ap_clk)
ret_V_2_reg_797 <= _025_;
always @(posedge ap_clk)
ret_V_19_reg_802 <= _018_;
always @(posedge ap_clk)
ret_V_21_reg_807 <= _020_;
always @(posedge ap_clk)
ret_V_25_reg_813 <= _024_;
always @(posedge ap_clk)
ret_V_3_reg_765 <= _028_;
always @(posedge ap_clk)
ret_V_20_reg_770 <= _019_;
always @(posedge ap_clk)
ret_V_16_reg_792 <= _016_;
always @(posedge ap_clk)
ret_V_22_reg_848 <= _021_;
always @(posedge ap_clk)
tmp_1_reg_853 <= _038_;
always @(posedge ap_clk)
ret_V_24_reg_858 <= _023_;
always @(posedge ap_clk)
ret_V_13_reg_863 <= _013_;
always @(posedge ap_clk)
trunc_ln851_4_reg_870 <= _042_;
always @(posedge ap_clk)
op_15_V_reg_907 <= _011_;
always @(posedge ap_clk)
ret_V_23_reg_912 <= _022_;
always @(posedge ap_clk)
ret_V_15_reg_917 <= _015_;
always @(posedge ap_clk)
icmp_ln851_reg_701 <= _010_;
always @(posedge ap_clk)
sext_ln850_reg_875 <= _036_;
always @(posedge ap_clk)
icmp_ln851_3_reg_882 <= _009_;
always @(posedge ap_clk)
ret_V_7_reg_663 <= _029_;
always @(posedge ap_clk)
icmp_ln851_2_reg_670 <= _008_;
always @(posedge ap_clk)
ret_V_18_reg_711 <= _017_;
always @(posedge ap_clk)
ret_V_reg_716 <= _032_;
always @(posedge ap_clk)
ret_V_3_cast_reg_723 <= _027_;
always @(posedge ap_clk)
p_Result_1_reg_730 <= _012_;
always @(posedge ap_clk)
icmp_ln851_1_reg_736 <= _007_;
always @(posedge ap_clk)
ret_V_3_cast5_reg_758 <= _026_;
always @(posedge ap_clk)
select_ln69_reg_952[1:0] <= _033_;
always @(posedge ap_clk)
add_ln69_reg_957 <= _005_;
always @(posedge ap_clk)
add_ln69_2_reg_962 <= _002_;
always @(posedge ap_clk)
add_ln69_3_reg_967 <= _003_;
always @(posedge ap_clk)
add_ln69_1_reg_977 <= _001_;
always @(posedge ap_clk)
add_ln69_4_reg_982 <= _004_;
always @(posedge ap_clk)
add_ln691_reg_897 <= _000_;
always @(posedge ap_clk)
ret_V_14_reg_902 <= _014_;
always @(posedge ap_clk)
ap_CS_fsm <= _006_;
assign _043_ = _049_ ? 2'h2 : 2'h1;
assign _219_ = ap_CS_fsm == 1'h1;
function [18:0] _592_;
input [18:0] a;
input [360:0] b;
input [18:0] s;
case (s)
19'b0000000000000000001:
_592_ = b[18:0];
19'b0000000000000000010:
_592_ = b[37:19];
19'b0000000000000000100:
_592_ = b[56:38];
19'b0000000000000001000:
_592_ = b[75:57];
19'b0000000000000010000:
_592_ = b[94:76];
19'b0000000000000100000:
_592_ = b[113:95];
19'b0000000000001000000:
_592_ = b[132:114];
19'b0000000000010000000:
_592_ = b[151:133];
19'b0000000000100000000:
_592_ = b[170:152];
19'b0000000001000000000:
_592_ = b[189:171];
19'b0000000010000000000:
_592_ = b[208:190];
19'b0000000100000000000:
_592_ = b[227:209];
19'b0000001000000000000:
_592_ = b[246:228];
19'b0000010000000000000:
_592_ = b[265:247];
19'b0000100000000000000:
_592_ = b[284:266];
19'b0001000000000000000:
_592_ = b[303:285];
19'b0010000000000000000:
_592_ = b[322:304];
19'b0100000000000000000:
_592_ = b[341:323];
19'b1000000000000000000:
_592_ = b[360:342];
19'b0000000000000000000:
_592_ = a;
default:
_592_ = 19'bx;
endcase
endfunction
assign ap_NS_fsm = _592_(19'hxxxxx, { 17'h00000, _043_, 342'h00002000080002000080002000080002000080002000080002000080002000080002000080002000000001 }, { _219_, _237_, _236_, _235_, _234_, _233_, _232_, _231_, _230_, _229_, _228_, _227_, _226_, _225_, _224_, _223_, _222_, _221_, _220_ });
assign _220_ = ap_CS_fsm == 19'h40000;
assign _221_ = ap_CS_fsm == 18'h20000;
assign _222_ = ap_CS_fsm == 17'h10000;
assign _223_ = ap_CS_fsm == 16'h8000;
assign _224_ = ap_CS_fsm == 15'h4000;
assign _225_ = ap_CS_fsm == 14'h2000;
assign _226_ = ap_CS_fsm == 13'h1000;
assign _227_ = ap_CS_fsm == 12'h800;
assign _228_ = ap_CS_fsm == 11'h400;
assign _229_ = ap_CS_fsm == 10'h200;
assign _230_ = ap_CS_fsm == 9'h100;
assign _231_ = ap_CS_fsm == 8'h80;
assign _232_ = ap_CS_fsm == 7'h40;
assign _233_ = ap_CS_fsm == 6'h20;
assign _234_ = ap_CS_fsm == 5'h10;
assign _235_ = ap_CS_fsm == 4'h8;
assign _236_ = ap_CS_fsm == 3'h4;
assign _237_ = ap_CS_fsm == 2'h2;
assign op_30_ap_vld = ap_CS_fsm[18] ? 1'h1 : 1'h0;
assign ap_idle = _048_ ? 1'h1 : 1'h0;
assign _041_ = _047_ ? grp_fu_376_p2[3:0] : trunc_ln1497_reg_887;
assign _040_ = _046_ ? grp_fu_367_p2[3:0] : trunc_ln1497_1_reg_892;
assign _037_ = _045_ ? grp_fu_267_p2 : sub_ln1497_reg_753;
assign _034_ = ap_CS_fsm[7] ? select_ln703_fu_454_p3[8:6] : select_ln703_reg_823[8:6];
assign _035_ = ap_CS_fsm[7] ? select_ln850_7_fu_447_p3 : select_ln850_7_reg_818;
assign _039_ = ap_CS_fsm[2] ? ret_V_9_fu_217_p3[1] : tmp_4_reg_686;
assign _031_ = ap_CS_fsm[2] ? ret_V_9_fu_217_p3 : ret_V_9_reg_680;
assign _030_ = ap_CS_fsm[1] ? grp_fu_199_p2 : ret_V_8_reg_675;
assign _025_ = _044_ ? grp_fu_355_p2 : ret_V_2_reg_797;
assign _024_ = ap_CS_fsm[6] ? ret_V_25_fu_429_p3 : ret_V_25_reg_813;
assign _020_ = ap_CS_fsm[6] ? ret_V_21_fu_418_p2 : ret_V_21_reg_807;
assign _018_ = ap_CS_fsm[6] ? ret_V_19_fu_387_p3 : ret_V_19_reg_802;
assign _016_ = ap_CS_fsm[5] ? grp_fu_349_p2 : ret_V_16_reg_792;
assign _019_ = ap_CS_fsm[5] ? grp_fu_333_p2 : ret_V_20_reg_770;
assign _028_ = ap_CS_fsm[5] ? grp_fu_311_p2 : ret_V_3_reg_765;
assign _042_ = ap_CS_fsm[9] ? grp_fu_485_p2[5:0] : trunc_ln851_4_reg_870;
assign _013_ = ap_CS_fsm[9] ? grp_fu_485_p2[8:6] : ret_V_13_reg_863;
assign _023_ = ap_CS_fsm[9] ? grp_fu_485_p2 : ret_V_24_reg_858;
assign _038_ = ap_CS_fsm[9] ? grp_fu_476_p2[6:1] : tmp_1_reg_853;
assign _021_ = ap_CS_fsm[9] ? grp_fu_476_p2 : ret_V_22_reg_848;
assign _015_ = ap_CS_fsm[12] ? ret_V_15_fu_581_p3 : ret_V_15_reg_917;
assign _022_ = ap_CS_fsm[12] ? ret_V_23_fu_562_p3 : ret_V_23_reg_912;
assign _011_ = ap_CS_fsm[12] ? op_15_V_fu_541_p3 : op_15_V_reg_907;
assign _010_ = ap_CS_fsm[3] ? icmp_ln851_fu_258_p2 : icmp_ln851_reg_701;
assign _009_ = ap_CS_fsm[10] ? icmp_ln851_3_fu_523_p2 : icmp_ln851_3_reg_882;
assign _036_ = ap_CS_fsm[10] ? { tmp_1_reg_853[5], tmp_1_reg_853 } : sext_ln850_reg_875;
assign _008_ = ap_CS_fsm[0] ? icmp_ln851_2_fu_193_p2 : icmp_ln851_2_reg_670;
assign _029_ = ap_CS_fsm[0] ? op_11[7:6] : ret_V_7_reg_663;
assign _026_ = ap_CS_fsm[4] ? op_3[20:17] : ret_V_3_cast5_reg_758;
assign _007_ = ap_CS_fsm[4] ? icmp_ln851_1_fu_305_p2 : icmp_ln851_1_reg_736;
assign _012_ = ap_CS_fsm[4] ? op_3[31] : p_Result_1_reg_730;
assign _027_ = ap_CS_fsm[4] ? op_3[18:17] : ret_V_3_cast_reg_723;
assign _032_ = ap_CS_fsm[4] ? grp_fu_248_p2[10:6] : ret_V_reg_716;
assign _017_ = ap_CS_fsm[4] ? grp_fu_248_p2 : ret_V_18_reg_711;
assign _003_ = ap_CS_fsm[14] ? grp_fu_619_p2 : add_ln69_3_reg_967;
assign _002_ = ap_CS_fsm[14] ? grp_fu_613_p2 : add_ln69_2_reg_962;
assign _005_ = ap_CS_fsm[14] ? grp_fu_607_p2 : add_ln69_reg_957;
assign _033_ = ap_CS_fsm[14] ? select_ln69_fu_625_p3 : select_ln69_reg_952[1:0];
assign _004_ = ap_CS_fsm[16] ? grp_fu_639_p2 : add_ln69_4_reg_982;
assign _001_ = ap_CS_fsm[16] ? grp_fu_632_p2 : add_ln69_1_reg_977;
assign _014_ = ap_CS_fsm[11] ? grp_fu_528_p2 : ret_V_14_reg_902;
assign _000_ = ap_CS_fsm[11] ? grp_fu_517_p2 : add_ln691_reg_897;
assign _006_ = ap_rst ? 19'h00001 : ap_NS_fsm;
assign icmp_ln851_1_fu_305_p2 = _053_ ? 1'h1 : 1'h0;
assign icmp_ln851_2_fu_193_p2 = _054_ ? 1'h1 : 1'h0;
assign icmp_ln851_3_fu_523_p2 = _055_ ? 1'h1 : 1'h0;
assign icmp_ln851_fu_258_p2 = _056_ ? 1'h1 : 1'h0;
assign op_15_V_fu_541_p3 = tmp_4_reg_686 ? trunc_ln1497_reg_887 : trunc_ln1497_1_reg_892;
assign ret_V_15_fu_581_p3 = ret_V_24_reg_858[8] ? select_ln850_5_fu_576_p3 : ret_V_13_reg_863;
assign ret_V_19_fu_387_p3 = p_Result_1_reg_730 ? select_ln850_fu_382_p3 : ret_V_3_cast_reg_723;
assign ret_V_23_fu_562_p3 = ret_V_22_reg_848[6] ? select_ln850_4_fu_556_p3 : sext_ln850_reg_875;
assign ret_V_25_fu_429_p3 = p_Result_1_reg_730 ? select_ln850_6_fu_424_p3 : ret_V_3_cast5_reg_758;
assign ret_V_9_fu_217_p3 = op_11[7] ? select_ln850_1_fu_212_p3 : ret_V_7_reg_663;
assign select_ln69_fu_625_p3 = ret_V_21_reg_807 ? 2'h1 : 2'h2;
assign select_ln703_fu_454_p3 = ret_V_21_reg_807 ? 9'h1c0 : 9'h000;
assign select_ln850_1_fu_212_p3 = icmp_ln851_2_reg_670 ? ret_V_7_reg_663 : ret_V_8_reg_675;
assign select_ln850_3_fu_442_p3 = icmp_ln851_reg_701 ? ret_V_reg_716 : ret_V_2_reg_797;
assign select_ln850_4_fu_556_p3 = op_6[0] ? add_ln691_reg_897 : sext_ln850_reg_875;
assign select_ln850_5_fu_576_p3 = icmp_ln851_3_reg_882 ? ret_V_13_reg_863 : ret_V_14_reg_902;
assign select_ln850_6_fu_424_p3 = icmp_ln851_1_reg_736 ? ret_V_3_cast5_reg_758 : ret_V_16_reg_792;
assign select_ln850_7_fu_447_p3 = ret_V_18_reg_711[10] ? select_ln850_3_fu_442_p3 : ret_V_reg_716;
assign select_ln850_fu_382_p3 = icmp_ln851_1_reg_736 ? ret_V_3_cast_reg_723 : ret_V_3_reg_765;
assign ret_V_21_fu_418_p2 = ret_V_20_reg_770[17] ^ and_ln353_fu_412_p2;
assign ap_CS_fsm_state1 = ap_CS_fsm[0];
assign ap_CS_fsm_state10 = ap_CS_fsm[9];
assign ap_CS_fsm_state11 = ap_CS_fsm[10];
assign ap_CS_fsm_state12 = ap_CS_fsm[11];
assign ap_CS_fsm_state13 = ap_CS_fsm[12];
assign ap_CS_fsm_state14 = ap_CS_fsm[13];
assign ap_CS_fsm_state15 = ap_CS_fsm[14];
assign ap_CS_fsm_state16 = ap_CS_fsm[15];
assign ap_CS_fsm_state17 = ap_CS_fsm[16];
assign ap_CS_fsm_state18 = ap_CS_fsm[17];
assign ap_CS_fsm_state19 = ap_CS_fsm[18];
assign ap_CS_fsm_state2 = ap_CS_fsm[1];
assign ap_CS_fsm_state3 = ap_CS_fsm[2];
assign ap_CS_fsm_state4 = ap_CS_fsm[3];
assign ap_CS_fsm_state5 = ap_CS_fsm[4];
assign ap_CS_fsm_state6 = ap_CS_fsm[5];
assign ap_CS_fsm_state7 = ap_CS_fsm[6];
assign ap_CS_fsm_state8 = ap_CS_fsm[7];
assign ap_CS_fsm_state9 = ap_CS_fsm[8];
assign ap_done = op_30_ap_vld;
assign ap_ready = op_30_ap_vld;
assign conv_i482_fu_363_p1 = { 24'h000000, op_2 };
assign grp_fu_199_p0 = op_11[7:6];
assign grp_fu_248_p0 = { op_0[3], op_0, 6'h00 };
assign grp_fu_248_p1 = { op_1[7], op_1[7], op_1[7], op_1 };
assign grp_fu_267_p1 = { ret_V_9_reg_680[1], ret_V_9_reg_680 };
assign grp_fu_311_p0 = op_3[18:17];
assign grp_fu_333_p0 = { 12'h000, op_4, 17'h00000 };
assign grp_fu_333_p1 = { op_3[31], op_3 };
assign grp_fu_349_p0 = op_3[20:17];
assign grp_fu_367_p1 = { ret_V_9_reg_680[1], ret_V_9_reg_680[1], ret_V_9_reg_680[1], ret_V_9_reg_680[1], ret_V_9_reg_680[1], ret_V_9_reg_680[1], ret_V_9_reg_680[1], ret_V_9_reg_680[1], ret_V_9_reg_680[1], ret_V_9_reg_680[1], ret_V_9_reg_680[1], ret_V_9_reg_680[1], ret_V_9_reg_680[1], ret_V_9_reg_680[1], ret_V_9_reg_680[1], ret_V_9_reg_680[1], ret_V_9_reg_680[1], ret_V_9_reg_680[1], ret_V_9_reg_680[1], ret_V_9_reg_680[1], ret_V_9_reg_680[1], ret_V_9_reg_680[1], ret_V_9_reg_680[1], ret_V_9_reg_680[1], ret_V_9_reg_680[1], ret_V_9_reg_680[1], ret_V_9_reg_680[1], ret_V_9_reg_680[1], ret_V_9_reg_680[1], ret_V_9_reg_680[1], ret_V_9_reg_680 };
assign grp_fu_376_p1 = { sub_ln1497_reg_753[2], sub_ln1497_reg_753[2], sub_ln1497_reg_753[2], sub_ln1497_reg_753[2], sub_ln1497_reg_753[2], sub_ln1497_reg_753[2], sub_ln1497_reg_753[2], sub_ln1497_reg_753[2], sub_ln1497_reg_753[2], sub_ln1497_reg_753[2], sub_ln1497_reg_753[2], sub_ln1497_reg_753[2], sub_ln1497_reg_753[2], sub_ln1497_reg_753[2], sub_ln1497_reg_753[2], sub_ln1497_reg_753[2], sub_ln1497_reg_753[2], sub_ln1497_reg_753[2], sub_ln1497_reg_753[2], sub_ln1497_reg_753[2], sub_ln1497_reg_753[2], sub_ln1497_reg_753[2], sub_ln1497_reg_753[2], sub_ln1497_reg_753[2], sub_ln1497_reg_753[2], sub_ln1497_reg_753[2], sub_ln1497_reg_753[2], sub_ln1497_reg_753[2], sub_ln1497_reg_753[2], sub_ln1497_reg_753 };
assign grp_fu_476_p0 = { select_ln850_7_reg_818[4], select_ln850_7_reg_818, 1'h0 };
assign grp_fu_476_p1 = { op_6[1], op_6[1], op_6[1], op_6[1], op_6[1], op_6 };
assign grp_fu_485_p1 = { op_11[7], op_11 };
assign grp_fu_517_p0 = { tmp_1_reg_853[5], tmp_1_reg_853 };
assign grp_fu_607_p0 = { ret_V_23_reg_912[6], ret_V_23_reg_912[6], ret_V_23_reg_912 };
assign grp_fu_607_p1 = { op_12[7], op_12 };
assign grp_fu_613_p0 = { 2'h0, op_15_V_reg_907 };
assign grp_fu_613_p1 = { ret_V_25_reg_813[3], ret_V_25_reg_813[3], ret_V_25_reg_813 };
assign grp_fu_619_p0 = { ret_V_15_reg_917[2], ret_V_15_reg_917 };
assign grp_fu_619_p1 = { ret_V_19_reg_802[1], ret_V_19_reg_802[1], ret_V_19_reg_802 };
assign grp_fu_639_p0 = { add_ln69_3_reg_967[3], add_ln69_3_reg_967[3], add_ln69_3_reg_967 };
assign grp_fu_647_p0 = { add_ln69_4_reg_982[5], add_ln69_4_reg_982[5], add_ln69_4_reg_982[5], add_ln69_4_reg_982 };
assign lhs_fu_232_p3 = { op_0, 6'h00 };
assign op_30 = { grp_fu_647_p2[8], grp_fu_647_p2[8], grp_fu_647_p2[8], grp_fu_647_p2[8], grp_fu_647_p2[8], grp_fu_647_p2[8], grp_fu_647_p2[8], grp_fu_647_p2[8], grp_fu_647_p2[8], grp_fu_647_p2[8], grp_fu_647_p2[8], grp_fu_647_p2[8], grp_fu_647_p2[8], grp_fu_647_p2[8], grp_fu_647_p2[8], grp_fu_647_p2[8], grp_fu_647_p2[8], grp_fu_647_p2[8], grp_fu_647_p2[8], grp_fu_647_p2[8], grp_fu_647_p2[8], grp_fu_647_p2[8], grp_fu_647_p2[8], grp_fu_647_p2 };
assign p_Result_1_fu_293_p1 = op_3;
assign p_Result_2_fu_400_p3 = ret_V_20_reg_770[32];
assign p_Result_3_fu_205_p1 = op_11;
assign p_Result_3_fu_205_p3 = op_11[7];
assign p_Result_4_fu_546_p3 = ret_V_22_reg_848[6];
assign p_Result_5_fu_569_p3 = ret_V_24_reg_858[8];
assign p_Result_s_fu_435_p3 = ret_V_18_reg_711[10];
assign ret_V_3_cast5_fu_339_p1 = op_3;
assign ret_V_3_cast_fu_283_p1 = op_3;
assign ret_V_7_fu_179_p1 = op_11;
assign rhs_1_fu_465_p3 = { select_ln850_7_reg_818, 1'h0 };
assign rhs_fu_321_p3 = { op_4, 17'h00000 };
assign sext_ln1192_1_fu_461_p0 = op_6;
assign sext_ln703_1_fu_317_p0 = op_3;
assign sext_ln703_2_fu_482_p0 = op_11;
assign sext_ln703_fu_244_p0 = op_1;
assign sext_ln850_fu_514_p1 = { tmp_1_reg_853[5], tmp_1_reg_853 };
assign tmp_fu_393_p3 = ret_V_20_reg_770[17];
assign trunc_ln1497_1_fu_537_p1 = grp_fu_367_p2[3:0];
assign trunc_ln1497_fu_533_p1 = grp_fu_376_p2[3:0];
assign trunc_ln851_1_fu_301_p0 = op_3;
assign trunc_ln851_1_fu_301_p1 = op_3[16:0];
assign trunc_ln851_2_fu_189_p0 = op_11;
assign trunc_ln851_2_fu_189_p1 = op_11[5:0];
assign trunc_ln851_3_fu_553_p0 = op_6;
assign trunc_ln851_3_fu_553_p1 = op_6[0];
assign trunc_ln851_4_fu_510_p1 = grp_fu_485_p2[5:0];
assign trunc_ln851_fu_254_p0 = op_1;
assign trunc_ln851_fu_254_p1 = op_1[5:0];
assign \sub_9ns_9s_9_2_1_U11.top_sub_9ns_9s_9_2_1_Adder_7_U.ain_s0  = \sub_9ns_9s_9_2_1_U11.top_sub_9ns_9s_9_2_1_Adder_7_U.a ;
assign \sub_9ns_9s_9_2_1_U11.top_sub_9ns_9s_9_2_1_Adder_7_U.s  = { \sub_9ns_9s_9_2_1_U11.top_sub_9ns_9s_9_2_1_Adder_7_U.fas_s2 , \sub_9ns_9s_9_2_1_U11.top_sub_9ns_9s_9_2_1_Adder_7_U.sum_s1  };
assign \sub_9ns_9s_9_2_1_U11.top_sub_9ns_9s_9_2_1_Adder_7_U.u2.a  = \sub_9ns_9s_9_2_1_U11.top_sub_9ns_9s_9_2_1_Adder_7_U.ain_s1 ;
assign \sub_9ns_9s_9_2_1_U11.top_sub_9ns_9s_9_2_1_Adder_7_U.u2.b  = \sub_9ns_9s_9_2_1_U11.top_sub_9ns_9s_9_2_1_Adder_7_U.bin_s1 ;
assign \sub_9ns_9s_9_2_1_U11.top_sub_9ns_9s_9_2_1_Adder_7_U.u2.cin  = \sub_9ns_9s_9_2_1_U11.top_sub_9ns_9s_9_2_1_Adder_7_U.carry_s1 ;
assign \sub_9ns_9s_9_2_1_U11.top_sub_9ns_9s_9_2_1_Adder_7_U.facout_s2  = \sub_9ns_9s_9_2_1_U11.top_sub_9ns_9s_9_2_1_Adder_7_U.u2.cout ;
assign \sub_9ns_9s_9_2_1_U11.top_sub_9ns_9s_9_2_1_Adder_7_U.fas_s2  = \sub_9ns_9s_9_2_1_U11.top_sub_9ns_9s_9_2_1_Adder_7_U.u2.s ;
assign \sub_9ns_9s_9_2_1_U11.top_sub_9ns_9s_9_2_1_Adder_7_U.u1.a  = \sub_9ns_9s_9_2_1_U11.top_sub_9ns_9s_9_2_1_Adder_7_U.a [3:0];
assign \sub_9ns_9s_9_2_1_U11.top_sub_9ns_9s_9_2_1_Adder_7_U.u1.b  = \sub_9ns_9s_9_2_1_U11.top_sub_9ns_9s_9_2_1_Adder_7_U.bin_s0 [3:0];
assign \sub_9ns_9s_9_2_1_U11.top_sub_9ns_9s_9_2_1_Adder_7_U.u1.cin  = 1'h1;
assign \sub_9ns_9s_9_2_1_U11.top_sub_9ns_9s_9_2_1_Adder_7_U.facout_s1  = \sub_9ns_9s_9_2_1_U11.top_sub_9ns_9s_9_2_1_Adder_7_U.u1.cout ;
assign \sub_9ns_9s_9_2_1_U11.top_sub_9ns_9s_9_2_1_Adder_7_U.fas_s1  = \sub_9ns_9s_9_2_1_U11.top_sub_9ns_9s_9_2_1_Adder_7_U.u1.s ;
assign \sub_9ns_9s_9_2_1_U11.top_sub_9ns_9s_9_2_1_Adder_7_U.a  = \sub_9ns_9s_9_2_1_U11.din0 ;
assign \sub_9ns_9s_9_2_1_U11.top_sub_9ns_9s_9_2_1_Adder_7_U.b  = \sub_9ns_9s_9_2_1_U11.din1 ;
assign \sub_9ns_9s_9_2_1_U11.top_sub_9ns_9s_9_2_1_Adder_7_U.ce  = \sub_9ns_9s_9_2_1_U11.ce ;
assign \sub_9ns_9s_9_2_1_U11.top_sub_9ns_9s_9_2_1_Adder_7_U.clk  = \sub_9ns_9s_9_2_1_U11.clk ;
assign \sub_9ns_9s_9_2_1_U11.top_sub_9ns_9s_9_2_1_Adder_7_U.reset  = \sub_9ns_9s_9_2_1_U11.reset ;
assign \sub_9ns_9s_9_2_1_U11.dout  = \sub_9ns_9s_9_2_1_U11.top_sub_9ns_9s_9_2_1_Adder_7_U.s ;
assign \sub_9ns_9s_9_2_1_U11.ce  = 1'h1;
assign \sub_9ns_9s_9_2_1_U11.clk  = ap_clk;
assign \sub_9ns_9s_9_2_1_U11.din0  = select_ln703_reg_823;
assign \sub_9ns_9s_9_2_1_U11.din1  = { op_11[7], op_11 };
assign grp_fu_485_p2 = \sub_9ns_9s_9_2_1_U11.dout ;
assign \sub_9ns_9s_9_2_1_U11.reset  = ap_rst;
assign \sub_3ns_3s_3_2_1_U3.top_sub_3ns_3s_3_2_1_Adder_2_U.ain_s0  = \sub_3ns_3s_3_2_1_U3.top_sub_3ns_3s_3_2_1_Adder_2_U.a ;
assign \sub_3ns_3s_3_2_1_U3.top_sub_3ns_3s_3_2_1_Adder_2_U.s  = { \sub_3ns_3s_3_2_1_U3.top_sub_3ns_3s_3_2_1_Adder_2_U.fas_s2 , \sub_3ns_3s_3_2_1_U3.top_sub_3ns_3s_3_2_1_Adder_2_U.sum_s1  };
assign \sub_3ns_3s_3_2_1_U3.top_sub_3ns_3s_3_2_1_Adder_2_U.u2.a  = \sub_3ns_3s_3_2_1_U3.top_sub_3ns_3s_3_2_1_Adder_2_U.ain_s1 ;
assign \sub_3ns_3s_3_2_1_U3.top_sub_3ns_3s_3_2_1_Adder_2_U.u2.b  = \sub_3ns_3s_3_2_1_U3.top_sub_3ns_3s_3_2_1_Adder_2_U.bin_s1 ;
assign \sub_3ns_3s_3_2_1_U3.top_sub_3ns_3s_3_2_1_Adder_2_U.u2.cin  = \sub_3ns_3s_3_2_1_U3.top_sub_3ns_3s_3_2_1_Adder_2_U.carry_s1 ;
assign \sub_3ns_3s_3_2_1_U3.top_sub_3ns_3s_3_2_1_Adder_2_U.facout_s2  = \sub_3ns_3s_3_2_1_U3.top_sub_3ns_3s_3_2_1_Adder_2_U.u2.cout ;
assign \sub_3ns_3s_3_2_1_U3.top_sub_3ns_3s_3_2_1_Adder_2_U.fas_s2  = \sub_3ns_3s_3_2_1_U3.top_sub_3ns_3s_3_2_1_Adder_2_U.u2.s ;
assign \sub_3ns_3s_3_2_1_U3.top_sub_3ns_3s_3_2_1_Adder_2_U.u1.a  = \sub_3ns_3s_3_2_1_U3.top_sub_3ns_3s_3_2_1_Adder_2_U.a [0];
assign \sub_3ns_3s_3_2_1_U3.top_sub_3ns_3s_3_2_1_Adder_2_U.u1.b  = \sub_3ns_3s_3_2_1_U3.top_sub_3ns_3s_3_2_1_Adder_2_U.bin_s0 [0];
assign \sub_3ns_3s_3_2_1_U3.top_sub_3ns_3s_3_2_1_Adder_2_U.u1.cin  = 1'h1;
assign \sub_3ns_3s_3_2_1_U3.top_sub_3ns_3s_3_2_1_Adder_2_U.facout_s1  = \sub_3ns_3s_3_2_1_U3.top_sub_3ns_3s_3_2_1_Adder_2_U.u1.cout ;
assign \sub_3ns_3s_3_2_1_U3.top_sub_3ns_3s_3_2_1_Adder_2_U.fas_s1  = \sub_3ns_3s_3_2_1_U3.top_sub_3ns_3s_3_2_1_Adder_2_U.u1.s ;
assign \sub_3ns_3s_3_2_1_U3.top_sub_3ns_3s_3_2_1_Adder_2_U.a  = \sub_3ns_3s_3_2_1_U3.din0 ;
assign \sub_3ns_3s_3_2_1_U3.top_sub_3ns_3s_3_2_1_Adder_2_U.b  = \sub_3ns_3s_3_2_1_U3.din1 ;
assign \sub_3ns_3s_3_2_1_U3.top_sub_3ns_3s_3_2_1_Adder_2_U.ce  = \sub_3ns_3s_3_2_1_U3.ce ;
assign \sub_3ns_3s_3_2_1_U3.top_sub_3ns_3s_3_2_1_Adder_2_U.clk  = \sub_3ns_3s_3_2_1_U3.clk ;
assign \sub_3ns_3s_3_2_1_U3.top_sub_3ns_3s_3_2_1_Adder_2_U.reset  = \sub_3ns_3s_3_2_1_U3.reset ;
assign \sub_3ns_3s_3_2_1_U3.dout  = \sub_3ns_3s_3_2_1_U3.top_sub_3ns_3s_3_2_1_Adder_2_U.s ;
assign \sub_3ns_3s_3_2_1_U3.ce  = 1'h1;
assign \sub_3ns_3s_3_2_1_U3.clk  = ap_clk;
assign \sub_3ns_3s_3_2_1_U3.din0  = 3'h0;
assign \sub_3ns_3s_3_2_1_U3.din1  = { ret_V_9_reg_680[1], ret_V_9_reg_680 };
assign grp_fu_267_p2 = \sub_3ns_3s_3_2_1_U3.dout ;
assign \sub_3ns_3s_3_2_1_U3.reset  = ap_rst;
assign \shl_32ns_32s_32_7_1_U8.din1_cast  = \shl_32ns_32s_32_7_1_U8.din1 ;
assign \shl_32ns_32s_32_7_1_U8.din1_mask  = 32'd31;
assign \shl_32ns_32s_32_7_1_U8.ce  = 1'h1;
assign \shl_32ns_32s_32_7_1_U8.clk  = ap_clk;
assign \shl_32ns_32s_32_7_1_U8.din0  = { 24'h000000, op_2 };
assign \shl_32ns_32s_32_7_1_U8.din1  = { ret_V_9_reg_680[1], ret_V_9_reg_680[1], ret_V_9_reg_680[1], ret_V_9_reg_680[1], ret_V_9_reg_680[1], ret_V_9_reg_680[1], ret_V_9_reg_680[1], ret_V_9_reg_680[1], ret_V_9_reg_680[1], ret_V_9_reg_680[1], ret_V_9_reg_680[1], ret_V_9_reg_680[1], ret_V_9_reg_680[1], ret_V_9_reg_680[1], ret_V_9_reg_680[1], ret_V_9_reg_680[1], ret_V_9_reg_680[1], ret_V_9_reg_680[1], ret_V_9_reg_680[1], ret_V_9_reg_680[1], ret_V_9_reg_680[1], ret_V_9_reg_680[1], ret_V_9_reg_680[1], ret_V_9_reg_680[1], ret_V_9_reg_680[1], ret_V_9_reg_680[1], ret_V_9_reg_680[1], ret_V_9_reg_680[1], ret_V_9_reg_680[1], ret_V_9_reg_680[1], ret_V_9_reg_680 };
assign grp_fu_367_p2 = \shl_32ns_32s_32_7_1_U8.dout ;
assign \shl_32ns_32s_32_7_1_U8.reset  = ap_rst;
assign \lshr_32ns_32s_32_7_1_U9.din1_cast  = \lshr_32ns_32s_32_7_1_U9.din1 ;
assign \lshr_32ns_32s_32_7_1_U9.din1_mask  = 32'd31;
assign \lshr_32ns_32s_32_7_1_U9.ce  = 1'h1;
assign \lshr_32ns_32s_32_7_1_U9.clk  = ap_clk;
assign \lshr_32ns_32s_32_7_1_U9.din0  = { 24'h000000, op_2 };
assign \lshr_32ns_32s_32_7_1_U9.din1  = { sub_ln1497_reg_753[2], sub_ln1497_reg_753[2], sub_ln1497_reg_753[2], sub_ln1497_reg_753[2], sub_ln1497_reg_753[2], sub_ln1497_reg_753[2], sub_ln1497_reg_753[2], sub_ln1497_reg_753[2], sub_ln1497_reg_753[2], sub_ln1497_reg_753[2], sub_ln1497_reg_753[2], sub_ln1497_reg_753[2], sub_ln1497_reg_753[2], sub_ln1497_reg_753[2], sub_ln1497_reg_753[2], sub_ln1497_reg_753[2], sub_ln1497_reg_753[2], sub_ln1497_reg_753[2], sub_ln1497_reg_753[2], sub_ln1497_reg_753[2], sub_ln1497_reg_753[2], sub_ln1497_reg_753[2], sub_ln1497_reg_753[2], sub_ln1497_reg_753[2], sub_ln1497_reg_753[2], sub_ln1497_reg_753[2], sub_ln1497_reg_753[2], sub_ln1497_reg_753[2], sub_ln1497_reg_753[2], sub_ln1497_reg_753 };
assign grp_fu_376_p2 = \lshr_32ns_32s_32_7_1_U9.dout ;
assign \lshr_32ns_32s_32_7_1_U9.reset  = ap_rst;
assign \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_10_U.ain_s0  = \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_10_U.a ;
assign \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_10_U.bin_s0  = \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_10_U.b ;
assign \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_10_U.s  = { \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_10_U.fas_s2 , \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_10_U.sum_s1  };
assign \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_10_U.u2.a  = \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_10_U.ain_s1 ;
assign \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_10_U.u2.b  = \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_10_U.bin_s1 ;
assign \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_10_U.u2.cin  = \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_10_U.carry_s1 ;
assign \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_10_U.facout_s2  = \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_10_U.u2.cout ;
assign \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_10_U.fas_s2  = \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_10_U.u2.s ;
assign \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_10_U.u1.a  = \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_10_U.a [3:0];
assign \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_10_U.u1.b  = \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_10_U.b [3:0];
assign \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_10_U.u1.cin  = 1'h0;
assign \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_10_U.facout_s1  = \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_10_U.u1.cout ;
assign \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_10_U.fas_s1  = \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_10_U.u1.s ;
assign \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_10_U.a  = \add_9s_9s_9_2_1_U14.din0 ;
assign \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_10_U.b  = \add_9s_9s_9_2_1_U14.din1 ;
assign \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_10_U.ce  = \add_9s_9s_9_2_1_U14.ce ;
assign \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_10_U.clk  = \add_9s_9s_9_2_1_U14.clk ;
assign \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_10_U.reset  = \add_9s_9s_9_2_1_U14.reset ;
assign \add_9s_9s_9_2_1_U14.dout  = \add_9s_9s_9_2_1_U14.top_add_9s_9s_9_2_1_Adder_10_U.s ;
assign \add_9s_9s_9_2_1_U14.ce  = 1'h1;
assign \add_9s_9s_9_2_1_U14.clk  = ap_clk;
assign \add_9s_9s_9_2_1_U14.din0  = { ret_V_23_reg_912[6], ret_V_23_reg_912[6], ret_V_23_reg_912 };
assign \add_9s_9s_9_2_1_U14.din1  = { op_12[7], op_12 };
assign grp_fu_607_p2 = \add_9s_9s_9_2_1_U14.dout ;
assign \add_9s_9s_9_2_1_U14.reset  = ap_rst;
assign \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_15_U.ain_s0  = \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_15_U.a ;
assign \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_15_U.bin_s0  = \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_15_U.b ;
assign \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_15_U.s  = { \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_15_U.fas_s2 , \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_15_U.sum_s1  };
assign \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_15_U.u2.a  = \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_15_U.ain_s1 ;
assign \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_15_U.u2.b  = \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_15_U.bin_s1 ;
assign \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_15_U.u2.cin  = \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_15_U.carry_s1 ;
assign \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_15_U.facout_s2  = \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_15_U.u2.cout ;
assign \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_15_U.fas_s2  = \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_15_U.u2.s ;
assign \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_15_U.u1.a  = \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_15_U.a [3:0];
assign \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_15_U.u1.b  = \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_15_U.b [3:0];
assign \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_15_U.u1.cin  = 1'h0;
assign \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_15_U.facout_s1  = \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_15_U.u1.cout ;
assign \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_15_U.fas_s1  = \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_15_U.u1.s ;
assign \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_15_U.a  = \add_9s_9ns_9_2_1_U19.din0 ;
assign \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_15_U.b  = \add_9s_9ns_9_2_1_U19.din1 ;
assign \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_15_U.ce  = \add_9s_9ns_9_2_1_U19.ce ;
assign \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_15_U.clk  = \add_9s_9ns_9_2_1_U19.clk ;
assign \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_15_U.reset  = \add_9s_9ns_9_2_1_U19.reset ;
assign \add_9s_9ns_9_2_1_U19.dout  = \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_15_U.s ;
assign \add_9s_9ns_9_2_1_U19.ce  = 1'h1;
assign \add_9s_9ns_9_2_1_U19.clk  = ap_clk;
assign \add_9s_9ns_9_2_1_U19.din0  = { add_ln69_4_reg_982[5], add_ln69_4_reg_982[5], add_ln69_4_reg_982[5], add_ln69_4_reg_982 };
assign \add_9s_9ns_9_2_1_U19.din1  = add_ln69_1_reg_977;
assign grp_fu_647_p2 = \add_9s_9ns_9_2_1_U19.dout ;
assign \add_9s_9ns_9_2_1_U19.reset  = ap_rst;
assign \add_9ns_9ns_9_2_1_U17.top_add_9ns_9ns_9_2_1_Adder_13_U.ain_s0  = \add_9ns_9ns_9_2_1_U17.top_add_9ns_9ns_9_2_1_Adder_13_U.a ;
assign \add_9ns_9ns_9_2_1_U17.top_add_9ns_9ns_9_2_1_Adder_13_U.bin_s0  = \add_9ns_9ns_9_2_1_U17.top_add_9ns_9ns_9_2_1_Adder_13_U.b ;
assign \add_9ns_9ns_9_2_1_U17.top_add_9ns_9ns_9_2_1_Adder_13_U.s  = { \add_9ns_9ns_9_2_1_U17.top_add_9ns_9ns_9_2_1_Adder_13_U.fas_s2 , \add_9ns_9ns_9_2_1_U17.top_add_9ns_9ns_9_2_1_Adder_13_U.sum_s1  };
assign \add_9ns_9ns_9_2_1_U17.top_add_9ns_9ns_9_2_1_Adder_13_U.u2.a  = \add_9ns_9ns_9_2_1_U17.top_add_9ns_9ns_9_2_1_Adder_13_U.ain_s1 ;
assign \add_9ns_9ns_9_2_1_U17.top_add_9ns_9ns_9_2_1_Adder_13_U.u2.b  = \add_9ns_9ns_9_2_1_U17.top_add_9ns_9ns_9_2_1_Adder_13_U.bin_s1 ;
assign \add_9ns_9ns_9_2_1_U17.top_add_9ns_9ns_9_2_1_Adder_13_U.u2.cin  = \add_9ns_9ns_9_2_1_U17.top_add_9ns_9ns_9_2_1_Adder_13_U.carry_s1 ;
assign \add_9ns_9ns_9_2_1_U17.top_add_9ns_9ns_9_2_1_Adder_13_U.facout_s2  = \add_9ns_9ns_9_2_1_U17.top_add_9ns_9ns_9_2_1_Adder_13_U.u2.cout ;
assign \add_9ns_9ns_9_2_1_U17.top_add_9ns_9ns_9_2_1_Adder_13_U.fas_s2  = \add_9ns_9ns_9_2_1_U17.top_add_9ns_9ns_9_2_1_Adder_13_U.u2.s ;
assign \add_9ns_9ns_9_2_1_U17.top_add_9ns_9ns_9_2_1_Adder_13_U.u1.a  = \add_9ns_9ns_9_2_1_U17.top_add_9ns_9ns_9_2_1_Adder_13_U.a [3:0];
assign \add_9ns_9ns_9_2_1_U17.top_add_9ns_9ns_9_2_1_Adder_13_U.u1.b  = \add_9ns_9ns_9_2_1_U17.top_add_9ns_9ns_9_2_1_Adder_13_U.b [3:0];
assign \add_9ns_9ns_9_2_1_U17.top_add_9ns_9ns_9_2_1_Adder_13_U.u1.cin  = 1'h0;
assign \add_9ns_9ns_9_2_1_U17.top_add_9ns_9ns_9_2_1_Adder_13_U.facout_s1  = \add_9ns_9ns_9_2_1_U17.top_add_9ns_9ns_9_2_1_Adder_13_U.u1.cout ;
assign \add_9ns_9ns_9_2_1_U17.top_add_9ns_9ns_9_2_1_Adder_13_U.fas_s1  = \add_9ns_9ns_9_2_1_U17.top_add_9ns_9ns_9_2_1_Adder_13_U.u1.s ;
assign \add_9ns_9ns_9_2_1_U17.top_add_9ns_9ns_9_2_1_Adder_13_U.a  = \add_9ns_9ns_9_2_1_U17.din0 ;
assign \add_9ns_9ns_9_2_1_U17.top_add_9ns_9ns_9_2_1_Adder_13_U.b  = \add_9ns_9ns_9_2_1_U17.din1 ;
assign \add_9ns_9ns_9_2_1_U17.top_add_9ns_9ns_9_2_1_Adder_13_U.ce  = \add_9ns_9ns_9_2_1_U17.ce ;
assign \add_9ns_9ns_9_2_1_U17.top_add_9ns_9ns_9_2_1_Adder_13_U.clk  = \add_9ns_9ns_9_2_1_U17.clk ;
assign \add_9ns_9ns_9_2_1_U17.top_add_9ns_9ns_9_2_1_Adder_13_U.reset  = \add_9ns_9ns_9_2_1_U17.reset ;
assign \add_9ns_9ns_9_2_1_U17.dout  = \add_9ns_9ns_9_2_1_U17.top_add_9ns_9ns_9_2_1_Adder_13_U.s ;
assign \add_9ns_9ns_9_2_1_U17.ce  = 1'h1;
assign \add_9ns_9ns_9_2_1_U17.clk  = ap_clk;
assign \add_9ns_9ns_9_2_1_U17.din0  = add_ln69_reg_957;
assign \add_9ns_9ns_9_2_1_U17.din1  = select_ln69_reg_952;
assign grp_fu_632_p2 = \add_9ns_9ns_9_2_1_U17.dout ;
assign \add_9ns_9ns_9_2_1_U17.reset  = ap_rst;
assign \add_7s_7s_7_2_1_U10.top_add_7s_7s_7_2_1_Adder_6_U.ain_s0  = \add_7s_7s_7_2_1_U10.top_add_7s_7s_7_2_1_Adder_6_U.a ;
assign \add_7s_7s_7_2_1_U10.top_add_7s_7s_7_2_1_Adder_6_U.bin_s0  = \add_7s_7s_7_2_1_U10.top_add_7s_7s_7_2_1_Adder_6_U.b ;
assign \add_7s_7s_7_2_1_U10.top_add_7s_7s_7_2_1_Adder_6_U.s  = { \add_7s_7s_7_2_1_U10.top_add_7s_7s_7_2_1_Adder_6_U.fas_s2 , \add_7s_7s_7_2_1_U10.top_add_7s_7s_7_2_1_Adder_6_U.sum_s1  };
assign \add_7s_7s_7_2_1_U10.top_add_7s_7s_7_2_1_Adder_6_U.u2.a  = \add_7s_7s_7_2_1_U10.top_add_7s_7s_7_2_1_Adder_6_U.ain_s1 ;
assign \add_7s_7s_7_2_1_U10.top_add_7s_7s_7_2_1_Adder_6_U.u2.b  = \add_7s_7s_7_2_1_U10.top_add_7s_7s_7_2_1_Adder_6_U.bin_s1 ;
assign \add_7s_7s_7_2_1_U10.top_add_7s_7s_7_2_1_Adder_6_U.u2.cin  = \add_7s_7s_7_2_1_U10.top_add_7s_7s_7_2_1_Adder_6_U.carry_s1 ;
assign \add_7s_7s_7_2_1_U10.top_add_7s_7s_7_2_1_Adder_6_U.facout_s2  = \add_7s_7s_7_2_1_U10.top_add_7s_7s_7_2_1_Adder_6_U.u2.cout ;
assign \add_7s_7s_7_2_1_U10.top_add_7s_7s_7_2_1_Adder_6_U.fas_s2  = \add_7s_7s_7_2_1_U10.top_add_7s_7s_7_2_1_Adder_6_U.u2.s ;
assign \add_7s_7s_7_2_1_U10.top_add_7s_7s_7_2_1_Adder_6_U.u1.a  = \add_7s_7s_7_2_1_U10.top_add_7s_7s_7_2_1_Adder_6_U.a [2:0];
assign \add_7s_7s_7_2_1_U10.top_add_7s_7s_7_2_1_Adder_6_U.u1.b  = \add_7s_7s_7_2_1_U10.top_add_7s_7s_7_2_1_Adder_6_U.b [2:0];
assign \add_7s_7s_7_2_1_U10.top_add_7s_7s_7_2_1_Adder_6_U.u1.cin  = 1'h0;
assign \add_7s_7s_7_2_1_U10.top_add_7s_7s_7_2_1_Adder_6_U.facout_s1  = \add_7s_7s_7_2_1_U10.top_add_7s_7s_7_2_1_Adder_6_U.u1.cout ;
assign \add_7s_7s_7_2_1_U10.top_add_7s_7s_7_2_1_Adder_6_U.fas_s1  = \add_7s_7s_7_2_1_U10.top_add_7s_7s_7_2_1_Adder_6_U.u1.s ;
assign \add_7s_7s_7_2_1_U10.top_add_7s_7s_7_2_1_Adder_6_U.a  = \add_7s_7s_7_2_1_U10.din0 ;
assign \add_7s_7s_7_2_1_U10.top_add_7s_7s_7_2_1_Adder_6_U.b  = \add_7s_7s_7_2_1_U10.din1 ;
assign \add_7s_7s_7_2_1_U10.top_add_7s_7s_7_2_1_Adder_6_U.ce  = \add_7s_7s_7_2_1_U10.ce ;
assign \add_7s_7s_7_2_1_U10.top_add_7s_7s_7_2_1_Adder_6_U.clk  = \add_7s_7s_7_2_1_U10.clk ;
assign \add_7s_7s_7_2_1_U10.top_add_7s_7s_7_2_1_Adder_6_U.reset  = \add_7s_7s_7_2_1_U10.reset ;
assign \add_7s_7s_7_2_1_U10.dout  = \add_7s_7s_7_2_1_U10.top_add_7s_7s_7_2_1_Adder_6_U.s ;
assign \add_7s_7s_7_2_1_U10.ce  = 1'h1;
assign \add_7s_7s_7_2_1_U10.clk  = ap_clk;
assign \add_7s_7s_7_2_1_U10.din0  = { select_ln850_7_reg_818[4], select_ln850_7_reg_818, 1'h0 };
assign \add_7s_7s_7_2_1_U10.din1  = { op_6[1], op_6[1], op_6[1], op_6[1], op_6[1], op_6 };
assign grp_fu_476_p2 = \add_7s_7s_7_2_1_U10.dout ;
assign \add_7s_7s_7_2_1_U10.reset  = ap_rst;
assign \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_8_U.ain_s0  = \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_8_U.a ;
assign \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_8_U.bin_s0  = \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_8_U.b ;
assign \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_8_U.s  = { \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_8_U.fas_s2 , \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_8_U.sum_s1  };
assign \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_8_U.u2.a  = \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_8_U.ain_s1 ;
assign \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_8_U.u2.b  = \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_8_U.bin_s1 ;
assign \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_8_U.u2.cin  = \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_8_U.carry_s1 ;
assign \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_8_U.facout_s2  = \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_8_U.u2.cout ;
assign \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_8_U.fas_s2  = \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_8_U.u2.s ;
assign \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_8_U.u1.a  = \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_8_U.a [2:0];
assign \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_8_U.u1.b  = \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_8_U.b [2:0];
assign \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_8_U.u1.cin  = 1'h0;
assign \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_8_U.facout_s1  = \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_8_U.u1.cout ;
assign \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_8_U.fas_s1  = \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_8_U.u1.s ;
assign \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_8_U.a  = \add_7s_7ns_7_2_1_U12.din0 ;
assign \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_8_U.b  = \add_7s_7ns_7_2_1_U12.din1 ;
assign \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_8_U.ce  = \add_7s_7ns_7_2_1_U12.ce ;
assign \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_8_U.clk  = \add_7s_7ns_7_2_1_U12.clk ;
assign \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_8_U.reset  = \add_7s_7ns_7_2_1_U12.reset ;
assign \add_7s_7ns_7_2_1_U12.dout  = \add_7s_7ns_7_2_1_U12.top_add_7s_7ns_7_2_1_Adder_8_U.s ;
assign \add_7s_7ns_7_2_1_U12.ce  = 1'h1;
assign \add_7s_7ns_7_2_1_U12.clk  = ap_clk;
assign \add_7s_7ns_7_2_1_U12.din0  = { tmp_1_reg_853[5], tmp_1_reg_853 };
assign \add_7s_7ns_7_2_1_U12.din1  = 7'h01;
assign grp_fu_517_p2 = \add_7s_7ns_7_2_1_U12.dout ;
assign \add_7s_7ns_7_2_1_U12.reset  = ap_rst;
assign \add_6s_6ns_6_2_1_U18.top_add_6s_6ns_6_2_1_Adder_14_U.ain_s0  = \add_6s_6ns_6_2_1_U18.top_add_6s_6ns_6_2_1_Adder_14_U.a ;
assign \add_6s_6ns_6_2_1_U18.top_add_6s_6ns_6_2_1_Adder_14_U.bin_s0  = \add_6s_6ns_6_2_1_U18.top_add_6s_6ns_6_2_1_Adder_14_U.b ;
assign \add_6s_6ns_6_2_1_U18.top_add_6s_6ns_6_2_1_Adder_14_U.s  = { \add_6s_6ns_6_2_1_U18.top_add_6s_6ns_6_2_1_Adder_14_U.fas_s2 , \add_6s_6ns_6_2_1_U18.top_add_6s_6ns_6_2_1_Adder_14_U.sum_s1  };
assign \add_6s_6ns_6_2_1_U18.top_add_6s_6ns_6_2_1_Adder_14_U.u2.a  = \add_6s_6ns_6_2_1_U18.top_add_6s_6ns_6_2_1_Adder_14_U.ain_s1 ;
assign \add_6s_6ns_6_2_1_U18.top_add_6s_6ns_6_2_1_Adder_14_U.u2.b  = \add_6s_6ns_6_2_1_U18.top_add_6s_6ns_6_2_1_Adder_14_U.bin_s1 ;
assign \add_6s_6ns_6_2_1_U18.top_add_6s_6ns_6_2_1_Adder_14_U.u2.cin  = \add_6s_6ns_6_2_1_U18.top_add_6s_6ns_6_2_1_Adder_14_U.carry_s1 ;
assign \add_6s_6ns_6_2_1_U18.top_add_6s_6ns_6_2_1_Adder_14_U.facout_s2  = \add_6s_6ns_6_2_1_U18.top_add_6s_6ns_6_2_1_Adder_14_U.u2.cout ;
assign \add_6s_6ns_6_2_1_U18.top_add_6s_6ns_6_2_1_Adder_14_U.fas_s2  = \add_6s_6ns_6_2_1_U18.top_add_6s_6ns_6_2_1_Adder_14_U.u2.s ;
assign \add_6s_6ns_6_2_1_U18.top_add_6s_6ns_6_2_1_Adder_14_U.u1.a  = \add_6s_6ns_6_2_1_U18.top_add_6s_6ns_6_2_1_Adder_14_U.a [2:0];
assign \add_6s_6ns_6_2_1_U18.top_add_6s_6ns_6_2_1_Adder_14_U.u1.b  = \add_6s_6ns_6_2_1_U18.top_add_6s_6ns_6_2_1_Adder_14_U.b [2:0];
assign \add_6s_6ns_6_2_1_U18.top_add_6s_6ns_6_2_1_Adder_14_U.u1.cin  = 1'h0;
assign \add_6s_6ns_6_2_1_U18.top_add_6s_6ns_6_2_1_Adder_14_U.facout_s1  = \add_6s_6ns_6_2_1_U18.top_add_6s_6ns_6_2_1_Adder_14_U.u1.cout ;
assign \add_6s_6ns_6_2_1_U18.top_add_6s_6ns_6_2_1_Adder_14_U.fas_s1  = \add_6s_6ns_6_2_1_U18.top_add_6s_6ns_6_2_1_Adder_14_U.u1.s ;
assign \add_6s_6ns_6_2_1_U18.top_add_6s_6ns_6_2_1_Adder_14_U.a  = \add_6s_6ns_6_2_1_U18.din0 ;
assign \add_6s_6ns_6_2_1_U18.top_add_6s_6ns_6_2_1_Adder_14_U.b  = \add_6s_6ns_6_2_1_U18.din1 ;
assign \add_6s_6ns_6_2_1_U18.top_add_6s_6ns_6_2_1_Adder_14_U.ce  = \add_6s_6ns_6_2_1_U18.ce ;
assign \add_6s_6ns_6_2_1_U18.top_add_6s_6ns_6_2_1_Adder_14_U.clk  = \add_6s_6ns_6_2_1_U18.clk ;
assign \add_6s_6ns_6_2_1_U18.top_add_6s_6ns_6_2_1_Adder_14_U.reset  = \add_6s_6ns_6_2_1_U18.reset ;
assign \add_6s_6ns_6_2_1_U18.dout  = \add_6s_6ns_6_2_1_U18.top_add_6s_6ns_6_2_1_Adder_14_U.s ;
assign \add_6s_6ns_6_2_1_U18.ce  = 1'h1;
assign \add_6s_6ns_6_2_1_U18.clk  = ap_clk;
assign \add_6s_6ns_6_2_1_U18.din0  = { add_ln69_3_reg_967[3], add_ln69_3_reg_967[3], add_ln69_3_reg_967 };
assign \add_6s_6ns_6_2_1_U18.din1  = add_ln69_2_reg_962;
assign grp_fu_639_p2 = \add_6s_6ns_6_2_1_U18.dout ;
assign \add_6s_6ns_6_2_1_U18.reset  = ap_rst;
assign \add_6ns_6s_6_2_1_U15.top_add_6ns_6s_6_2_1_Adder_11_U.ain_s0  = \add_6ns_6s_6_2_1_U15.top_add_6ns_6s_6_2_1_Adder_11_U.a ;
assign \add_6ns_6s_6_2_1_U15.top_add_6ns_6s_6_2_1_Adder_11_U.bin_s0  = \add_6ns_6s_6_2_1_U15.top_add_6ns_6s_6_2_1_Adder_11_U.b ;
assign \add_6ns_6s_6_2_1_U15.top_add_6ns_6s_6_2_1_Adder_11_U.s  = { \add_6ns_6s_6_2_1_U15.top_add_6ns_6s_6_2_1_Adder_11_U.fas_s2 , \add_6ns_6s_6_2_1_U15.top_add_6ns_6s_6_2_1_Adder_11_U.sum_s1  };
assign \add_6ns_6s_6_2_1_U15.top_add_6ns_6s_6_2_1_Adder_11_U.u2.a  = \add_6ns_6s_6_2_1_U15.top_add_6ns_6s_6_2_1_Adder_11_U.ain_s1 ;
assign \add_6ns_6s_6_2_1_U15.top_add_6ns_6s_6_2_1_Adder_11_U.u2.b  = \add_6ns_6s_6_2_1_U15.top_add_6ns_6s_6_2_1_Adder_11_U.bin_s1 ;
assign \add_6ns_6s_6_2_1_U15.top_add_6ns_6s_6_2_1_Adder_11_U.u2.cin  = \add_6ns_6s_6_2_1_U15.top_add_6ns_6s_6_2_1_Adder_11_U.carry_s1 ;
assign \add_6ns_6s_6_2_1_U15.top_add_6ns_6s_6_2_1_Adder_11_U.facout_s2  = \add_6ns_6s_6_2_1_U15.top_add_6ns_6s_6_2_1_Adder_11_U.u2.cout ;
assign \add_6ns_6s_6_2_1_U15.top_add_6ns_6s_6_2_1_Adder_11_U.fas_s2  = \add_6ns_6s_6_2_1_U15.top_add_6ns_6s_6_2_1_Adder_11_U.u2.s ;
assign \add_6ns_6s_6_2_1_U15.top_add_6ns_6s_6_2_1_Adder_11_U.u1.a  = \add_6ns_6s_6_2_1_U15.top_add_6ns_6s_6_2_1_Adder_11_U.a [2:0];
assign \add_6ns_6s_6_2_1_U15.top_add_6ns_6s_6_2_1_Adder_11_U.u1.b  = \add_6ns_6s_6_2_1_U15.top_add_6ns_6s_6_2_1_Adder_11_U.b [2:0];
assign \add_6ns_6s_6_2_1_U15.top_add_6ns_6s_6_2_1_Adder_11_U.u1.cin  = 1'h0;
assign \add_6ns_6s_6_2_1_U15.top_add_6ns_6s_6_2_1_Adder_11_U.facout_s1  = \add_6ns_6s_6_2_1_U15.top_add_6ns_6s_6_2_1_Adder_11_U.u1.cout ;
assign \add_6ns_6s_6_2_1_U15.top_add_6ns_6s_6_2_1_Adder_11_U.fas_s1  = \add_6ns_6s_6_2_1_U15.top_add_6ns_6s_6_2_1_Adder_11_U.u1.s ;
assign \add_6ns_6s_6_2_1_U15.top_add_6ns_6s_6_2_1_Adder_11_U.a  = \add_6ns_6s_6_2_1_U15.din0 ;
assign \add_6ns_6s_6_2_1_U15.top_add_6ns_6s_6_2_1_Adder_11_U.b  = \add_6ns_6s_6_2_1_U15.din1 ;
assign \add_6ns_6s_6_2_1_U15.top_add_6ns_6s_6_2_1_Adder_11_U.ce  = \add_6ns_6s_6_2_1_U15.ce ;
assign \add_6ns_6s_6_2_1_U15.top_add_6ns_6s_6_2_1_Adder_11_U.clk  = \add_6ns_6s_6_2_1_U15.clk ;
assign \add_6ns_6s_6_2_1_U15.top_add_6ns_6s_6_2_1_Adder_11_U.reset  = \add_6ns_6s_6_2_1_U15.reset ;
assign \add_6ns_6s_6_2_1_U15.dout  = \add_6ns_6s_6_2_1_U15.top_add_6ns_6s_6_2_1_Adder_11_U.s ;
assign \add_6ns_6s_6_2_1_U15.ce  = 1'h1;
assign \add_6ns_6s_6_2_1_U15.clk  = ap_clk;
assign \add_6ns_6s_6_2_1_U15.din0  = { 2'h0, op_15_V_reg_907 };
assign \add_6ns_6s_6_2_1_U15.din1  = { ret_V_25_reg_813[3], ret_V_25_reg_813[3], ret_V_25_reg_813 };
assign grp_fu_613_p2 = \add_6ns_6s_6_2_1_U15.dout ;
assign \add_6ns_6s_6_2_1_U15.reset  = ap_rst;
assign \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_5_U.ain_s0  = \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_5_U.a ;
assign \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_5_U.bin_s0  = \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_5_U.b ;
assign \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_5_U.s  = { \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_5_U.fas_s2 , \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_5_U.sum_s1  };
assign \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_5_U.u2.a  = \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_5_U.ain_s1 ;
assign \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_5_U.u2.b  = \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_5_U.bin_s1 ;
assign \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_5_U.u2.cin  = \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_5_U.carry_s1 ;
assign \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_5_U.facout_s2  = \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_5_U.u2.cout ;
assign \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_5_U.fas_s2  = \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_5_U.u2.s ;
assign \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_5_U.u1.a  = \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_5_U.a [1:0];
assign \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_5_U.u1.b  = \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_5_U.b [1:0];
assign \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_5_U.u1.cin  = 1'h0;
assign \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_5_U.facout_s1  = \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_5_U.u1.cout ;
assign \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_5_U.fas_s1  = \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_5_U.u1.s ;
assign \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_5_U.a  = \add_5ns_5ns_5_2_1_U7.din0 ;
assign \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_5_U.b  = \add_5ns_5ns_5_2_1_U7.din1 ;
assign \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_5_U.ce  = \add_5ns_5ns_5_2_1_U7.ce ;
assign \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_5_U.clk  = \add_5ns_5ns_5_2_1_U7.clk ;
assign \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_5_U.reset  = \add_5ns_5ns_5_2_1_U7.reset ;
assign \add_5ns_5ns_5_2_1_U7.dout  = \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_5_U.s ;
assign \add_5ns_5ns_5_2_1_U7.ce  = 1'h1;
assign \add_5ns_5ns_5_2_1_U7.clk  = ap_clk;
assign \add_5ns_5ns_5_2_1_U7.din0  = ret_V_reg_716;
assign \add_5ns_5ns_5_2_1_U7.din1  = 5'h01;
assign grp_fu_355_p2 = \add_5ns_5ns_5_2_1_U7.dout ;
assign \add_5ns_5ns_5_2_1_U7.reset  = ap_rst;
assign \add_4s_4s_4_2_1_U16.top_add_4s_4s_4_2_1_Adder_12_U.ain_s0  = \add_4s_4s_4_2_1_U16.top_add_4s_4s_4_2_1_Adder_12_U.a ;
assign \add_4s_4s_4_2_1_U16.top_add_4s_4s_4_2_1_Adder_12_U.bin_s0  = \add_4s_4s_4_2_1_U16.top_add_4s_4s_4_2_1_Adder_12_U.b ;
assign \add_4s_4s_4_2_1_U16.top_add_4s_4s_4_2_1_Adder_12_U.s  = { \add_4s_4s_4_2_1_U16.top_add_4s_4s_4_2_1_Adder_12_U.fas_s2 , \add_4s_4s_4_2_1_U16.top_add_4s_4s_4_2_1_Adder_12_U.sum_s1  };
assign \add_4s_4s_4_2_1_U16.top_add_4s_4s_4_2_1_Adder_12_U.u2.a  = \add_4s_4s_4_2_1_U16.top_add_4s_4s_4_2_1_Adder_12_U.ain_s1 ;
assign \add_4s_4s_4_2_1_U16.top_add_4s_4s_4_2_1_Adder_12_U.u2.b  = \add_4s_4s_4_2_1_U16.top_add_4s_4s_4_2_1_Adder_12_U.bin_s1 ;
assign \add_4s_4s_4_2_1_U16.top_add_4s_4s_4_2_1_Adder_12_U.u2.cin  = \add_4s_4s_4_2_1_U16.top_add_4s_4s_4_2_1_Adder_12_U.carry_s1 ;
assign \add_4s_4s_4_2_1_U16.top_add_4s_4s_4_2_1_Adder_12_U.facout_s2  = \add_4s_4s_4_2_1_U16.top_add_4s_4s_4_2_1_Adder_12_U.u2.cout ;
assign \add_4s_4s_4_2_1_U16.top_add_4s_4s_4_2_1_Adder_12_U.fas_s2  = \add_4s_4s_4_2_1_U16.top_add_4s_4s_4_2_1_Adder_12_U.u2.s ;
assign \add_4s_4s_4_2_1_U16.top_add_4s_4s_4_2_1_Adder_12_U.u1.a  = \add_4s_4s_4_2_1_U16.top_add_4s_4s_4_2_1_Adder_12_U.a [1:0];
assign \add_4s_4s_4_2_1_U16.top_add_4s_4s_4_2_1_Adder_12_U.u1.b  = \add_4s_4s_4_2_1_U16.top_add_4s_4s_4_2_1_Adder_12_U.b [1:0];
assign \add_4s_4s_4_2_1_U16.top_add_4s_4s_4_2_1_Adder_12_U.u1.cin  = 1'h0;
assign \add_4s_4s_4_2_1_U16.top_add_4s_4s_4_2_1_Adder_12_U.facout_s1  = \add_4s_4s_4_2_1_U16.top_add_4s_4s_4_2_1_Adder_12_U.u1.cout ;
assign \add_4s_4s_4_2_1_U16.top_add_4s_4s_4_2_1_Adder_12_U.fas_s1  = \add_4s_4s_4_2_1_U16.top_add_4s_4s_4_2_1_Adder_12_U.u1.s ;
assign \add_4s_4s_4_2_1_U16.top_add_4s_4s_4_2_1_Adder_12_U.a  = \add_4s_4s_4_2_1_U16.din0 ;
assign \add_4s_4s_4_2_1_U16.top_add_4s_4s_4_2_1_Adder_12_U.b  = \add_4s_4s_4_2_1_U16.din1 ;
assign \add_4s_4s_4_2_1_U16.top_add_4s_4s_4_2_1_Adder_12_U.ce  = \add_4s_4s_4_2_1_U16.ce ;
assign \add_4s_4s_4_2_1_U16.top_add_4s_4s_4_2_1_Adder_12_U.clk  = \add_4s_4s_4_2_1_U16.clk ;
assign \add_4s_4s_4_2_1_U16.top_add_4s_4s_4_2_1_Adder_12_U.reset  = \add_4s_4s_4_2_1_U16.reset ;
assign \add_4s_4s_4_2_1_U16.dout  = \add_4s_4s_4_2_1_U16.top_add_4s_4s_4_2_1_Adder_12_U.s ;
assign \add_4s_4s_4_2_1_U16.ce  = 1'h1;
assign \add_4s_4s_4_2_1_U16.clk  = ap_clk;
assign \add_4s_4s_4_2_1_U16.din0  = { ret_V_15_reg_917[2], ret_V_15_reg_917 };
assign \add_4s_4s_4_2_1_U16.din1  = { ret_V_19_reg_802[1], ret_V_19_reg_802[1], ret_V_19_reg_802 };
assign grp_fu_619_p2 = \add_4s_4s_4_2_1_U16.dout ;
assign \add_4s_4s_4_2_1_U16.reset  = ap_rst;
assign \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.ain_s0  = \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.a ;
assign \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.bin_s0  = \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.b ;
assign \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.s  = { \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.fas_s2 , \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.sum_s1  };
assign \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.u2.a  = \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.ain_s1 ;
assign \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.u2.b  = \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.bin_s1 ;
assign \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.u2.cin  = \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.carry_s1 ;
assign \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.facout_s2  = \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.u2.cout ;
assign \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.fas_s2  = \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.u2.s ;
assign \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.u1.a  = \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.a [1:0];
assign \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.u1.b  = \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.b [1:0];
assign \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.u1.cin  = 1'h0;
assign \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.facout_s1  = \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.u1.cout ;
assign \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.fas_s1  = \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.u1.s ;
assign \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.a  = \add_4ns_4ns_4_2_1_U6.din0 ;
assign \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.b  = \add_4ns_4ns_4_2_1_U6.din1 ;
assign \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.ce  = \add_4ns_4ns_4_2_1_U6.ce ;
assign \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.clk  = \add_4ns_4ns_4_2_1_U6.clk ;
assign \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.reset  = \add_4ns_4ns_4_2_1_U6.reset ;
assign \add_4ns_4ns_4_2_1_U6.dout  = \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.s ;
assign \add_4ns_4ns_4_2_1_U6.ce  = 1'h1;
assign \add_4ns_4ns_4_2_1_U6.clk  = ap_clk;
assign \add_4ns_4ns_4_2_1_U6.din0  = op_3[20:17];
assign \add_4ns_4ns_4_2_1_U6.din1  = 4'h1;
assign grp_fu_349_p2 = \add_4ns_4ns_4_2_1_U6.dout ;
assign \add_4ns_4ns_4_2_1_U6.reset  = ap_rst;
assign \add_3ns_3ns_3_2_1_U13.top_add_3ns_3ns_3_2_1_Adder_9_U.ain_s0  = \add_3ns_3ns_3_2_1_U13.top_add_3ns_3ns_3_2_1_Adder_9_U.a ;
assign \add_3ns_3ns_3_2_1_U13.top_add_3ns_3ns_3_2_1_Adder_9_U.bin_s0  = \add_3ns_3ns_3_2_1_U13.top_add_3ns_3ns_3_2_1_Adder_9_U.b ;
assign \add_3ns_3ns_3_2_1_U13.top_add_3ns_3ns_3_2_1_Adder_9_U.s  = { \add_3ns_3ns_3_2_1_U13.top_add_3ns_3ns_3_2_1_Adder_9_U.fas_s2 , \add_3ns_3ns_3_2_1_U13.top_add_3ns_3ns_3_2_1_Adder_9_U.sum_s1  };
assign \add_3ns_3ns_3_2_1_U13.top_add_3ns_3ns_3_2_1_Adder_9_U.u2.a  = \add_3ns_3ns_3_2_1_U13.top_add_3ns_3ns_3_2_1_Adder_9_U.ain_s1 ;
assign \add_3ns_3ns_3_2_1_U13.top_add_3ns_3ns_3_2_1_Adder_9_U.u2.b  = \add_3ns_3ns_3_2_1_U13.top_add_3ns_3ns_3_2_1_Adder_9_U.bin_s1 ;
assign \add_3ns_3ns_3_2_1_U13.top_add_3ns_3ns_3_2_1_Adder_9_U.u2.cin  = \add_3ns_3ns_3_2_1_U13.top_add_3ns_3ns_3_2_1_Adder_9_U.carry_s1 ;
assign \add_3ns_3ns_3_2_1_U13.top_add_3ns_3ns_3_2_1_Adder_9_U.facout_s2  = \add_3ns_3ns_3_2_1_U13.top_add_3ns_3ns_3_2_1_Adder_9_U.u2.cout ;
assign \add_3ns_3ns_3_2_1_U13.top_add_3ns_3ns_3_2_1_Adder_9_U.fas_s2  = \add_3ns_3ns_3_2_1_U13.top_add_3ns_3ns_3_2_1_Adder_9_U.u2.s ;
assign \add_3ns_3ns_3_2_1_U13.top_add_3ns_3ns_3_2_1_Adder_9_U.u1.a  = \add_3ns_3ns_3_2_1_U13.top_add_3ns_3ns_3_2_1_Adder_9_U.a [0];
assign \add_3ns_3ns_3_2_1_U13.top_add_3ns_3ns_3_2_1_Adder_9_U.u1.b  = \add_3ns_3ns_3_2_1_U13.top_add_3ns_3ns_3_2_1_Adder_9_U.b [0];
assign \add_3ns_3ns_3_2_1_U13.top_add_3ns_3ns_3_2_1_Adder_9_U.u1.cin  = 1'h0;
assign \add_3ns_3ns_3_2_1_U13.top_add_3ns_3ns_3_2_1_Adder_9_U.facout_s1  = \add_3ns_3ns_3_2_1_U13.top_add_3ns_3ns_3_2_1_Adder_9_U.u1.cout ;
assign \add_3ns_3ns_3_2_1_U13.top_add_3ns_3ns_3_2_1_Adder_9_U.fas_s1  = \add_3ns_3ns_3_2_1_U13.top_add_3ns_3ns_3_2_1_Adder_9_U.u1.s ;
assign \add_3ns_3ns_3_2_1_U13.top_add_3ns_3ns_3_2_1_Adder_9_U.a  = \add_3ns_3ns_3_2_1_U13.din0 ;
assign \add_3ns_3ns_3_2_1_U13.top_add_3ns_3ns_3_2_1_Adder_9_U.b  = \add_3ns_3ns_3_2_1_U13.din1 ;
assign \add_3ns_3ns_3_2_1_U13.top_add_3ns_3ns_3_2_1_Adder_9_U.ce  = \add_3ns_3ns_3_2_1_U13.ce ;
assign \add_3ns_3ns_3_2_1_U13.top_add_3ns_3ns_3_2_1_Adder_9_U.clk  = \add_3ns_3ns_3_2_1_U13.clk ;
assign \add_3ns_3ns_3_2_1_U13.top_add_3ns_3ns_3_2_1_Adder_9_U.reset  = \add_3ns_3ns_3_2_1_U13.reset ;
assign \add_3ns_3ns_3_2_1_U13.dout  = \add_3ns_3ns_3_2_1_U13.top_add_3ns_3ns_3_2_1_Adder_9_U.s ;
assign \add_3ns_3ns_3_2_1_U13.ce  = 1'h1;
assign \add_3ns_3ns_3_2_1_U13.clk  = ap_clk;
assign \add_3ns_3ns_3_2_1_U13.din0  = ret_V_13_reg_863;
assign \add_3ns_3ns_3_2_1_U13.din1  = 3'h1;
assign grp_fu_528_p2 = \add_3ns_3ns_3_2_1_U13.dout ;
assign \add_3ns_3ns_3_2_1_U13.reset  = ap_rst;
assign \add_33ns_33s_33_2_1_U5.top_add_33ns_33s_33_2_1_Adder_3_U.ain_s0  = \add_33ns_33s_33_2_1_U5.top_add_33ns_33s_33_2_1_Adder_3_U.a ;
assign \add_33ns_33s_33_2_1_U5.top_add_33ns_33s_33_2_1_Adder_3_U.bin_s0  = \add_33ns_33s_33_2_1_U5.top_add_33ns_33s_33_2_1_Adder_3_U.b ;
assign \add_33ns_33s_33_2_1_U5.top_add_33ns_33s_33_2_1_Adder_3_U.s  = { \add_33ns_33s_33_2_1_U5.top_add_33ns_33s_33_2_1_Adder_3_U.fas_s2 , \add_33ns_33s_33_2_1_U5.top_add_33ns_33s_33_2_1_Adder_3_U.sum_s1  };
assign \add_33ns_33s_33_2_1_U5.top_add_33ns_33s_33_2_1_Adder_3_U.u2.a  = \add_33ns_33s_33_2_1_U5.top_add_33ns_33s_33_2_1_Adder_3_U.ain_s1 ;
assign \add_33ns_33s_33_2_1_U5.top_add_33ns_33s_33_2_1_Adder_3_U.u2.b  = \add_33ns_33s_33_2_1_U5.top_add_33ns_33s_33_2_1_Adder_3_U.bin_s1 ;
assign \add_33ns_33s_33_2_1_U5.top_add_33ns_33s_33_2_1_Adder_3_U.u2.cin  = \add_33ns_33s_33_2_1_U5.top_add_33ns_33s_33_2_1_Adder_3_U.carry_s1 ;
assign \add_33ns_33s_33_2_1_U5.top_add_33ns_33s_33_2_1_Adder_3_U.facout_s2  = \add_33ns_33s_33_2_1_U5.top_add_33ns_33s_33_2_1_Adder_3_U.u2.cout ;
assign \add_33ns_33s_33_2_1_U5.top_add_33ns_33s_33_2_1_Adder_3_U.fas_s2  = \add_33ns_33s_33_2_1_U5.top_add_33ns_33s_33_2_1_Adder_3_U.u2.s ;
assign \add_33ns_33s_33_2_1_U5.top_add_33ns_33s_33_2_1_Adder_3_U.u1.a  = \add_33ns_33s_33_2_1_U5.top_add_33ns_33s_33_2_1_Adder_3_U.a [15:0];
assign \add_33ns_33s_33_2_1_U5.top_add_33ns_33s_33_2_1_Adder_3_U.u1.b  = \add_33ns_33s_33_2_1_U5.top_add_33ns_33s_33_2_1_Adder_3_U.b [15:0];
assign \add_33ns_33s_33_2_1_U5.top_add_33ns_33s_33_2_1_Adder_3_U.u1.cin  = 1'h0;
assign \add_33ns_33s_33_2_1_U5.top_add_33ns_33s_33_2_1_Adder_3_U.facout_s1  = \add_33ns_33s_33_2_1_U5.top_add_33ns_33s_33_2_1_Adder_3_U.u1.cout ;
assign \add_33ns_33s_33_2_1_U5.top_add_33ns_33s_33_2_1_Adder_3_U.fas_s1  = \add_33ns_33s_33_2_1_U5.top_add_33ns_33s_33_2_1_Adder_3_U.u1.s ;
assign \add_33ns_33s_33_2_1_U5.top_add_33ns_33s_33_2_1_Adder_3_U.a  = \add_33ns_33s_33_2_1_U5.din0 ;
assign \add_33ns_33s_33_2_1_U5.top_add_33ns_33s_33_2_1_Adder_3_U.b  = \add_33ns_33s_33_2_1_U5.din1 ;
assign \add_33ns_33s_33_2_1_U5.top_add_33ns_33s_33_2_1_Adder_3_U.ce  = \add_33ns_33s_33_2_1_U5.ce ;
assign \add_33ns_33s_33_2_1_U5.top_add_33ns_33s_33_2_1_Adder_3_U.clk  = \add_33ns_33s_33_2_1_U5.clk ;
assign \add_33ns_33s_33_2_1_U5.top_add_33ns_33s_33_2_1_Adder_3_U.reset  = \add_33ns_33s_33_2_1_U5.reset ;
assign \add_33ns_33s_33_2_1_U5.dout  = \add_33ns_33s_33_2_1_U5.top_add_33ns_33s_33_2_1_Adder_3_U.s ;
assign \add_33ns_33s_33_2_1_U5.ce  = 1'h1;
assign \add_33ns_33s_33_2_1_U5.clk  = ap_clk;
assign \add_33ns_33s_33_2_1_U5.din0  = { 12'h000, op_4, 17'h00000 };
assign \add_33ns_33s_33_2_1_U5.din1  = { op_3[31], op_3 };
assign grp_fu_333_p2 = \add_33ns_33s_33_2_1_U5.dout ;
assign \add_33ns_33s_33_2_1_U5.reset  = ap_rst;
assign \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_0_U.ain_s0  = \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_0_U.a ;
assign \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_0_U.bin_s0  = \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_0_U.b ;
assign \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_0_U.s  = { \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_0_U.fas_s2 , \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_0_U.sum_s1  };
assign \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_0_U.u2.a  = \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_0_U.ain_s1 ;
assign \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_0_U.u2.b  = \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_0_U.bin_s1 ;
assign \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_0_U.u2.cin  = \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_0_U.carry_s1 ;
assign \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_0_U.facout_s2  = \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_0_U.u2.cout ;
assign \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_0_U.fas_s2  = \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_0_U.u2.s ;
assign \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_0_U.u1.a  = \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_0_U.a [0];
assign \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_0_U.u1.b  = \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_0_U.b [0];
assign \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_0_U.u1.cin  = 1'h0;
assign \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_0_U.facout_s1  = \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_0_U.u1.cout ;
assign \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_0_U.fas_s1  = \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_0_U.u1.s ;
assign \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_0_U.a  = \add_2ns_2ns_2_2_1_U4.din0 ;
assign \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_0_U.b  = \add_2ns_2ns_2_2_1_U4.din1 ;
assign \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_0_U.ce  = \add_2ns_2ns_2_2_1_U4.ce ;
assign \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_0_U.clk  = \add_2ns_2ns_2_2_1_U4.clk ;
assign \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_0_U.reset  = \add_2ns_2ns_2_2_1_U4.reset ;
assign \add_2ns_2ns_2_2_1_U4.dout  = \add_2ns_2ns_2_2_1_U4.top_add_2ns_2ns_2_2_1_Adder_0_U.s ;
assign \add_2ns_2ns_2_2_1_U4.ce  = 1'h1;
assign \add_2ns_2ns_2_2_1_U4.clk  = ap_clk;
assign \add_2ns_2ns_2_2_1_U4.din0  = op_3[18:17];
assign \add_2ns_2ns_2_2_1_U4.din1  = 2'h1;
assign grp_fu_311_p2 = \add_2ns_2ns_2_2_1_U4.dout ;
assign \add_2ns_2ns_2_2_1_U4.reset  = ap_rst;
assign \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.ain_s0  = \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.a ;
assign \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.bin_s0  = \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.b ;
assign \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.s  = { \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.fas_s2 , \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.sum_s1  };
assign \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.u2.a  = \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.ain_s1 ;
assign \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.u2.b  = \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.bin_s1 ;
assign \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.u2.cin  = \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.carry_s1 ;
assign \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.facout_s2  = \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.u2.cout ;
assign \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.fas_s2  = \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.u2.s ;
assign \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.u1.a  = \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.a [0];
assign \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.u1.b  = \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.b [0];
assign \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.u1.cin  = 1'h0;
assign \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.facout_s1  = \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.u1.cout ;
assign \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.fas_s1  = \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.u1.s ;
assign \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.a  = \add_2ns_2ns_2_2_1_U1.din0 ;
assign \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.b  = \add_2ns_2ns_2_2_1_U1.din1 ;
assign \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.ce  = \add_2ns_2ns_2_2_1_U1.ce ;
assign \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.clk  = \add_2ns_2ns_2_2_1_U1.clk ;
assign \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.reset  = \add_2ns_2ns_2_2_1_U1.reset ;
assign \add_2ns_2ns_2_2_1_U1.dout  = \add_2ns_2ns_2_2_1_U1.top_add_2ns_2ns_2_2_1_Adder_0_U.s ;
assign \add_2ns_2ns_2_2_1_U1.ce  = 1'h1;
assign \add_2ns_2ns_2_2_1_U1.clk  = ap_clk;
assign \add_2ns_2ns_2_2_1_U1.din0  = op_11[7:6];
assign \add_2ns_2ns_2_2_1_U1.din1  = 2'h1;
assign grp_fu_199_p2 = \add_2ns_2ns_2_2_1_U1.dout ;
assign \add_2ns_2ns_2_2_1_U1.reset  = ap_rst;
assign \add_11s_11s_11_2_1_U2.top_add_11s_11s_11_2_1_Adder_1_U.ain_s0  = \add_11s_11s_11_2_1_U2.top_add_11s_11s_11_2_1_Adder_1_U.a ;
assign \add_11s_11s_11_2_1_U2.top_add_11s_11s_11_2_1_Adder_1_U.bin_s0  = \add_11s_11s_11_2_1_U2.top_add_11s_11s_11_2_1_Adder_1_U.b ;
assign \add_11s_11s_11_2_1_U2.top_add_11s_11s_11_2_1_Adder_1_U.s  = { \add_11s_11s_11_2_1_U2.top_add_11s_11s_11_2_1_Adder_1_U.fas_s2 , \add_11s_11s_11_2_1_U2.top_add_11s_11s_11_2_1_Adder_1_U.sum_s1  };
assign \add_11s_11s_11_2_1_U2.top_add_11s_11s_11_2_1_Adder_1_U.u2.a  = \add_11s_11s_11_2_1_U2.top_add_11s_11s_11_2_1_Adder_1_U.ain_s1 ;
assign \add_11s_11s_11_2_1_U2.top_add_11s_11s_11_2_1_Adder_1_U.u2.b  = \add_11s_11s_11_2_1_U2.top_add_11s_11s_11_2_1_Adder_1_U.bin_s1 ;
assign \add_11s_11s_11_2_1_U2.top_add_11s_11s_11_2_1_Adder_1_U.u2.cin  = \add_11s_11s_11_2_1_U2.top_add_11s_11s_11_2_1_Adder_1_U.carry_s1 ;
assign \add_11s_11s_11_2_1_U2.top_add_11s_11s_11_2_1_Adder_1_U.facout_s2  = \add_11s_11s_11_2_1_U2.top_add_11s_11s_11_2_1_Adder_1_U.u2.cout ;
assign \add_11s_11s_11_2_1_U2.top_add_11s_11s_11_2_1_Adder_1_U.fas_s2  = \add_11s_11s_11_2_1_U2.top_add_11s_11s_11_2_1_Adder_1_U.u2.s ;
assign \add_11s_11s_11_2_1_U2.top_add_11s_11s_11_2_1_Adder_1_U.u1.a  = \add_11s_11s_11_2_1_U2.top_add_11s_11s_11_2_1_Adder_1_U.a [4:0];
assign \add_11s_11s_11_2_1_U2.top_add_11s_11s_11_2_1_Adder_1_U.u1.b  = \add_11s_11s_11_2_1_U2.top_add_11s_11s_11_2_1_Adder_1_U.b [4:0];
assign \add_11s_11s_11_2_1_U2.top_add_11s_11s_11_2_1_Adder_1_U.u1.cin  = 1'h0;
assign \add_11s_11s_11_2_1_U2.top_add_11s_11s_11_2_1_Adder_1_U.facout_s1  = \add_11s_11s_11_2_1_U2.top_add_11s_11s_11_2_1_Adder_1_U.u1.cout ;
assign \add_11s_11s_11_2_1_U2.top_add_11s_11s_11_2_1_Adder_1_U.fas_s1  = \add_11s_11s_11_2_1_U2.top_add_11s_11s_11_2_1_Adder_1_U.u1.s ;
assign \add_11s_11s_11_2_1_U2.top_add_11s_11s_11_2_1_Adder_1_U.a  = \add_11s_11s_11_2_1_U2.din0 ;
assign \add_11s_11s_11_2_1_U2.top_add_11s_11s_11_2_1_Adder_1_U.b  = \add_11s_11s_11_2_1_U2.din1 ;
assign \add_11s_11s_11_2_1_U2.top_add_11s_11s_11_2_1_Adder_1_U.ce  = \add_11s_11s_11_2_1_U2.ce ;
assign \add_11s_11s_11_2_1_U2.top_add_11s_11s_11_2_1_Adder_1_U.clk  = \add_11s_11s_11_2_1_U2.clk ;
assign \add_11s_11s_11_2_1_U2.top_add_11s_11s_11_2_1_Adder_1_U.reset  = \add_11s_11s_11_2_1_U2.reset ;
assign \add_11s_11s_11_2_1_U2.dout  = \add_11s_11s_11_2_1_U2.top_add_11s_11s_11_2_1_Adder_1_U.s ;
assign \add_11s_11s_11_2_1_U2.ce  = 1'h1;
assign \add_11s_11s_11_2_1_U2.clk  = ap_clk;
assign \add_11s_11s_11_2_1_U2.din0  = { op_0[3], op_0, 6'h00 };
assign \add_11s_11s_11_2_1_U2.din1  = { op_1[7], op_1[7], op_1[7], op_1 };
assign grp_fu_248_p2 = \add_11s_11s_11_2_1_U2.dout ;
assign \add_11s_11s_11_2_1_U2.reset  = ap_rst;
endmodule


// Machine B:
// Processed by function `add_clk_enable_signal` in `verilog_tricks.py`.
// Processed by function `remove_reset_signal` in `verilog_tricks.py`.
module top_B (
  ap_clk,
  ap_start,
  ap_done,
  ap_idle,
  ap_ready,
  op_0,
  op_1,
  op_2,
  op_3,
  op_4,
  op_6,
  op_10,
  op_11,
  op_12,
  op_30,
  op_30_ap_vld,
clk_enable
);
input clk_enable;


input ap_clk;
wire ap_rst;
assign ap_rst = op_30_ap_vld;
input ap_start;
input [3:0] op_0;
input [7:0] op_1;
input [7:0] op_10;
input [7:0] op_11;
input [7:0] op_12;
input [7:0] op_2;
input [31:0] op_3;
input [3:0] op_4;
input [1:0] op_6;
output ap_done;
output ap_idle;
output ap_ready;
output [31:0] op_30;
output op_30_ap_vld;


reg [3:0] add_ln69_3_reg_749;
reg [5:0] add_ln69_4_reg_759;
reg [8:0] add_ln69_reg_754;
reg [3:0] ap_CS_fsm = 4'h1;
reg [3:0] op_15_V_reg_734;
reg [1:0] ret_V_19_reg_706;
reg ret_V_21_reg_711;
reg [6:0] ret_V_22_reg_739;
reg [3:0] ret_V_25_reg_724;
reg [1:0] ret_V_9_reg_717;
reg [5:0] tmp_1_reg_744;
wire [3:0] _000_;
wire [5:0] _001_;
wire [8:0] _002_;
wire [3:0] _003_;
wire [3:0] _004_;
wire [1:0] _005_;
wire _006_;
wire [6:0] _007_;
wire [3:0] _008_;
wire [1:0] _009_;
wire [5:0] _010_;
wire [1:0] _011_;
wire _012_;
wire _013_;
wire _014_;
wire _015_;
wire _016_;
wire _017_;
wire _018_;
wire _019_;
wire _020_;
wire _021_;
wire _022_;
wire [6:0] add_ln691_fu_618_p2;
wire [8:0] add_ln69_1_fu_682_p2;
wire [5:0] add_ln69_2_fu_660_p2;
wire [3:0] add_ln69_3_fu_599_p2;
wire [5:0] add_ln69_4_fu_669_p2;
wire [8:0] add_ln69_5_fu_690_p2;
wire [8:0] add_ln69_fu_654_p2;
wire and_ln353_fu_273_p2;
wire ap_CS_fsm_state1;
wire ap_CS_fsm_state2;
wire ap_CS_fsm_state3;
wire ap_CS_fsm_state4;
wire [3:0] ap_NS_fsm;
wire ap_clk;
wire ap_done;
wire ap_idle;
wire ap_ready;
wire ap_rst;
wire ap_start;
wire [31:0] conv_i482_fu_436_p1;
wire icmp_ln851_1_fu_201_p2;
wire icmp_ln851_2_fu_307_p2;
wire icmp_ln851_3_fu_564_p2;
wire icmp_ln851_fu_411_p2;
wire [9:0] lhs_fu_367_p3;
wire [31:0] lshr_ln1497_fu_456_p2;
wire [3:0] op_0;
wire [7:0] op_1;
wire [7:0] op_10;
wire [7:0] op_11;
wire [7:0] op_12;
wire [3:0] op_15_V_fu_470_p3;
wire [7:0] op_2;
wire [31:0] op_3;
wire [31:0] op_30;
wire op_30_ap_vld;
wire [3:0] op_4;
wire [1:0] op_6;
wire [31:0] p_Result_1_fu_189_p1;
wire p_Result_1_fu_189_p3;
wire p_Result_2_fu_259_p3;
wire [7:0] p_Result_3_fu_295_p1;
wire p_Result_3_fu_295_p3;
wire p_Result_4_fu_608_p3;
wire p_Result_5_fu_552_p3;
wire p_Result_s_fu_399_p3;
wire [2:0] ret_V_13_fu_542_p4;
wire [2:0] ret_V_14_fu_570_p2;
wire [2:0] ret_V_15_fu_584_p3;
wire [3:0] ret_V_16_fu_345_p2;
wire [10:0] ret_V_18_fu_383_p2;
wire [1:0] ret_V_19_fu_221_p3;
wire [32:0] ret_V_20_fu_245_p2;
wire ret_V_21_fu_279_p2;
wire [6:0] ret_V_22_fu_510_p2;
wire [6:0] ret_V_23_fu_632_p3;
wire [8:0] ret_V_24_fu_536_p2;
wire [3:0] ret_V_25_fu_359_p3;
wire [4:0] ret_V_2_fu_417_p2;
wire [31:0] ret_V_3_cast5_fu_335_p1;
wire [3:0] ret_V_3_cast5_fu_335_p4;
wire [31:0] ret_V_3_cast_fu_179_p1;
wire [1:0] ret_V_3_cast_fu_179_p4;
wire [1:0] ret_V_3_fu_207_p2;
wire [7:0] ret_V_7_fu_285_p1;
wire [1:0] ret_V_7_fu_285_p4;
wire [1:0] ret_V_8_fu_313_p2;
wire [1:0] ret_V_9_fu_327_p3;
wire [4:0] ret_V_fu_389_p4;
wire [5:0] rhs_1_fu_498_p3;
wire [20:0] rhs_fu_233_p3;
wire [1:0] select_ln69_fu_675_p3;
wire [8:0] select_ln703_fu_526_p3;
wire [1:0] select_ln850_1_fu_319_p3;
wire [4:0] select_ln850_3_fu_482_p3;
wire [6:0] select_ln850_4_fu_624_p3;
wire [2:0] select_ln850_5_fu_576_p3;
wire [3:0] select_ln850_6_fu_351_p3;
wire [4:0] select_ln850_7_fu_490_p3;
wire [1:0] select_ln850_fu_213_p3;
wire [1:0] sext_ln1192_1_fu_478_p0;
wire [6:0] sext_ln1192_1_fu_478_p1;
wire [6:0] sext_ln1192_2_fu_506_p1;
wire [10:0] sext_ln1192_fu_375_p1;
wire [3:0] sext_ln1193_fu_592_p1;
wire [31:0] sext_ln1497_1_fu_452_p1;
wire [2:0] sext_ln1497_fu_426_p1;
wire [8:0] sext_ln27_fu_644_p1;
wire [31:0] sext_ln545_fu_423_p1;
wire [3:0] sext_ln69_1_fu_595_p1;
wire [5:0] sext_ln69_2_fu_666_p1;
wire [8:0] sext_ln69_3_fu_687_p1;
wire [5:0] sext_ln69_fu_651_p1;
wire [31:0] sext_ln703_1_fu_229_p0;
wire [32:0] sext_ln703_1_fu_229_p1;
wire [7:0] sext_ln703_2_fu_533_p0;
wire [8:0] sext_ln703_2_fu_533_p1;
wire [7:0] sext_ln703_fu_379_p0;
wire [10:0] sext_ln703_fu_379_p1;
wire [8:0] sext_ln831_fu_640_p1;
wire [6:0] sext_ln850_fu_605_p1;
wire [31:0] shl_ln1497_fu_440_p2;
wire [2:0] sub_ln1497_fu_446_p2;
wire tmp_4_fu_429_p3;
wire tmp_fu_251_p3;
wire [3:0] trunc_ln1497_1_fu_466_p1;
wire [3:0] trunc_ln1497_fu_462_p1;
wire [31:0] trunc_ln851_1_fu_197_p0;
wire [16:0] trunc_ln851_1_fu_197_p1;
wire [7:0] trunc_ln851_2_fu_303_p0;
wire [5:0] trunc_ln851_2_fu_303_p1;
wire [1:0] trunc_ln851_3_fu_615_p0;
wire trunc_ln851_3_fu_615_p1;
wire [5:0] trunc_ln851_4_fu_560_p1;
wire [7:0] trunc_ln851_fu_407_p0;
wire [5:0] trunc_ln851_fu_407_p1;
wire xor_ln850_fu_267_p2;
wire [32:0] zext_ln1192_fu_241_p1;
wire [5:0] zext_ln27_fu_648_p1;


assign add_ln691_fu_618_p2 = $signed(tmp_1_reg_744) + $signed(2'h1);
assign add_ln69_1_fu_682_p2 = add_ln69_reg_754 + { 7'h00, select_ln69_fu_675_p3 };
assign add_ln69_2_fu_660_p2 = $signed({ 1'h0, op_15_V_reg_734 }) + $signed(ret_V_25_reg_724);
assign add_ln69_3_fu_599_p2 = $signed(ret_V_15_fu_584_p3) + $signed(ret_V_19_reg_706);
assign add_ln69_4_fu_669_p2 = $signed(add_ln69_3_reg_749) + $signed(add_ln69_2_fu_660_p2);
assign add_ln69_5_fu_690_p2 = $signed(add_ln69_4_reg_759) + $signed(add_ln69_1_fu_682_p2);
assign add_ln69_fu_654_p2 = $signed(ret_V_23_fu_632_p3) + $signed(op_12);
assign ret_V_14_fu_570_p2 = ret_V_24_fu_536_p2[8:6] + 1'h1;
assign ret_V_16_fu_345_p2 = op_3[20:17] + 1'h1;
assign ret_V_18_fu_383_p2 = $signed({ op_0, 6'h00 }) + $signed(op_1);
assign ret_V_20_fu_245_p2 = $signed({ 1'h0, op_4, 17'h00000 }) + $signed(op_3);
assign ret_V_22_fu_510_p2 = $signed({ select_ln850_7_fu_490_p3, 1'h0 }) + $signed(op_6);
assign ret_V_2_fu_417_p2 = ret_V_18_fu_383_p2[10:6] + 1'h1;
assign ret_V_3_fu_207_p2 = op_3[18:17] + 1'h1;
assign ret_V_8_fu_313_p2 = op_11[7:6] + 1'h1;
assign _012_ = _014_ & ap_CS_fsm[0];
assign _013_ = ap_start & ap_CS_fsm[0];
assign and_ln353_fu_273_p2 = xor_ln850_fu_267_p2 & ret_V_20_fu_245_p2[32];
assign xor_ln850_fu_267_p2 = ~ icmp_ln851_1_fu_201_p2;
assign _014_ = ~ ap_start;
assign _015_ = ! op_3[16:0];
assign _016_ = ! op_11[5:0];
assign _017_ = ! ret_V_24_fu_536_p2[5:0];
assign _018_ = ! op_1[5:0];
always @(posedge ap_clk)
ret_V_19_reg_706 <= _005_;
always @(posedge ap_clk)
ret_V_21_reg_711 <= _006_;
always @(posedge ap_clk)
ret_V_9_reg_717 <= _009_;
always @(posedge ap_clk)
ret_V_25_reg_724 <= _008_;
always @(posedge ap_clk)
add_ln69_reg_754 <= _002_;
always @(posedge ap_clk)
add_ln69_4_reg_759 <= _001_;
always @(posedge ap_clk)
op_15_V_reg_734 <= _004_;
always @(posedge ap_clk)
ret_V_22_reg_739 <= _007_;
always @(posedge ap_clk)
tmp_1_reg_744 <= _010_;
always @(posedge ap_clk)
add_ln69_3_reg_749 <= _000_;
always @(posedge ap_clk)
ap_CS_fsm <= _003_;
assign op_30_ap_vld = ap_CS_fsm[3] ? 1'h1 : 1'h0;
assign ap_idle = _012_ ? 1'h1 : 1'h0;
assign _008_ = ap_CS_fsm[0] ? ret_V_25_fu_359_p3 : ret_V_25_reg_724;
assign _009_ = ap_CS_fsm[0] ? ret_V_9_fu_327_p3 : ret_V_9_reg_717;
assign _006_ = ap_CS_fsm[0] ? ret_V_21_fu_279_p2 : ret_V_21_reg_711;
assign _005_ = ap_CS_fsm[0] ? ret_V_19_fu_221_p3 : ret_V_19_reg_706;
assign _001_ = ap_CS_fsm[2] ? add_ln69_4_fu_669_p2 : add_ln69_4_reg_759;
assign _002_ = ap_CS_fsm[2] ? add_ln69_fu_654_p2 : add_ln69_reg_754;
assign _000_ = ap_CS_fsm[1] ? add_ln69_3_fu_599_p2 : add_ln69_3_reg_749;
assign _010_ = ap_CS_fsm[1] ? ret_V_22_fu_510_p2[6:1] : tmp_1_reg_744;
assign _007_ = ap_CS_fsm[1] ? ret_V_22_fu_510_p2 : ret_V_22_reg_739;
assign _004_ = ap_CS_fsm[1] ? op_15_V_fu_470_p3 : op_15_V_reg_734;
assign _003_ = ap_rst ? 4'h1 : ap_NS_fsm;
assign _011_ = _013_ ? 2'h2 : 2'h1;
assign _019_ = ap_CS_fsm == 1'h1;
function [3:0] _073_;
input [3:0] a;
input [15:0] b;
input [3:0] s;
case (s)
4'b0001:
_073_ = b[3:0];
4'b0010:
_073_ = b[7:4];
4'b0100:
_073_ = b[11:8];
4'b1000:
_073_ = b[15:12];
4'b0000:
_073_ = a;
default:
_073_ = 4'bx;
endcase
endfunction
assign ap_NS_fsm = _073_(4'hx, { 2'h0, _011_, 12'h481 }, { _019_, _022_, _021_, _020_ });
assign _020_ = ap_CS_fsm == 4'h8;
assign _021_ = ap_CS_fsm == 3'h4;
assign _022_ = ap_CS_fsm == 2'h2;
assign trunc_ln1497_1_fu_466_p1 = op_2 << { ret_V_9_reg_717[1], ret_V_9_reg_717[1], ret_V_9_reg_717[1], ret_V_9_reg_717[1], ret_V_9_reg_717[1], ret_V_9_reg_717[1], ret_V_9_reg_717[1], ret_V_9_reg_717[1], ret_V_9_reg_717[1], ret_V_9_reg_717[1], ret_V_9_reg_717[1], ret_V_9_reg_717[1], ret_V_9_reg_717[1], ret_V_9_reg_717[1], ret_V_9_reg_717[1], ret_V_9_reg_717[1], ret_V_9_reg_717[1], ret_V_9_reg_717[1], ret_V_9_reg_717[1], ret_V_9_reg_717[1], ret_V_9_reg_717[1], ret_V_9_reg_717[1], ret_V_9_reg_717[1], ret_V_9_reg_717[1], ret_V_9_reg_717[1], ret_V_9_reg_717[1], ret_V_9_reg_717[1], ret_V_9_reg_717[1], ret_V_9_reg_717[1], ret_V_9_reg_717[1], ret_V_9_reg_717 };
assign trunc_ln1497_fu_462_p1 = op_2 >> { sub_ln1497_fu_446_p2[2], sub_ln1497_fu_446_p2[2], sub_ln1497_fu_446_p2[2], sub_ln1497_fu_446_p2[2], sub_ln1497_fu_446_p2[2], sub_ln1497_fu_446_p2[2], sub_ln1497_fu_446_p2[2], sub_ln1497_fu_446_p2[2], sub_ln1497_fu_446_p2[2], sub_ln1497_fu_446_p2[2], sub_ln1497_fu_446_p2[2], sub_ln1497_fu_446_p2[2], sub_ln1497_fu_446_p2[2], sub_ln1497_fu_446_p2[2], sub_ln1497_fu_446_p2[2], sub_ln1497_fu_446_p2[2], sub_ln1497_fu_446_p2[2], sub_ln1497_fu_446_p2[2], sub_ln1497_fu_446_p2[2], sub_ln1497_fu_446_p2[2], sub_ln1497_fu_446_p2[2], sub_ln1497_fu_446_p2[2], sub_ln1497_fu_446_p2[2], sub_ln1497_fu_446_p2[2], sub_ln1497_fu_446_p2[2], sub_ln1497_fu_446_p2[2], sub_ln1497_fu_446_p2[2], sub_ln1497_fu_446_p2[2], sub_ln1497_fu_446_p2[2], sub_ln1497_fu_446_p2 };
assign ret_V_24_fu_536_p2 = $signed(select_ln703_fu_526_p3) - $signed(op_11);
assign sub_ln1497_fu_446_p2 = $signed(1'h0) - $signed(ret_V_9_reg_717);
assign icmp_ln851_1_fu_201_p2 = _015_ ? 1'h1 : 1'h0;
assign icmp_ln851_2_fu_307_p2 = _016_ ? 1'h1 : 1'h0;
assign icmp_ln851_3_fu_564_p2 = _017_ ? 1'h1 : 1'h0;
assign icmp_ln851_fu_411_p2 = _018_ ? 1'h1 : 1'h0;
assign op_15_V_fu_470_p3 = ret_V_9_reg_717[1] ? trunc_ln1497_fu_462_p1 : trunc_ln1497_1_fu_466_p1;
assign ret_V_15_fu_584_p3 = ret_V_24_fu_536_p2[8] ? select_ln850_5_fu_576_p3 : { 1'h0, ret_V_24_fu_536_p2[7:6] };
assign ret_V_19_fu_221_p3 = op_3[31] ? select_ln850_fu_213_p3 : op_3[18:17];
assign ret_V_23_fu_632_p3 = ret_V_22_reg_739[6] ? select_ln850_4_fu_624_p3 : { tmp_1_reg_744[5], tmp_1_reg_744 };
assign ret_V_25_fu_359_p3 = op_3[31] ? select_ln850_6_fu_351_p3 : op_3[20:17];
assign ret_V_9_fu_327_p3 = op_11[7] ? select_ln850_1_fu_319_p3 : { 1'h0, op_11[6] };
assign select_ln69_fu_675_p3 = ret_V_21_reg_711 ? 2'h1 : 2'h2;
assign select_ln703_fu_526_p3 = ret_V_21_reg_711 ? 9'h1c0 : 9'h000;
assign select_ln850_1_fu_319_p3 = icmp_ln851_2_fu_307_p2 ? { 1'h1, op_11[6] } : ret_V_8_fu_313_p2;
assign select_ln850_3_fu_482_p3 = icmp_ln851_fu_411_p2 ? { 1'h1, ret_V_18_fu_383_p2[9:6] } : ret_V_2_fu_417_p2;
assign select_ln850_4_fu_624_p3 = op_6[0] ? add_ln691_fu_618_p2 : { tmp_1_reg_744[5], tmp_1_reg_744 };
assign select_ln850_5_fu_576_p3 = icmp_ln851_3_fu_564_p2 ? { 1'h1, ret_V_24_fu_536_p2[7:6] } : ret_V_14_fu_570_p2;
assign select_ln850_6_fu_351_p3 = icmp_ln851_1_fu_201_p2 ? op_3[20:17] : ret_V_16_fu_345_p2;
assign select_ln850_7_fu_490_p3 = ret_V_18_fu_383_p2[10] ? select_ln850_3_fu_482_p3 : { 1'h0, ret_V_18_fu_383_p2[9:6] };
assign select_ln850_fu_213_p3 = icmp_ln851_1_fu_201_p2 ? op_3[18:17] : ret_V_3_fu_207_p2;
assign ret_V_21_fu_279_p2 = ret_V_20_fu_245_p2[17] ^ and_ln353_fu_273_p2;
assign ap_CS_fsm_state1 = ap_CS_fsm[0];
assign ap_CS_fsm_state2 = ap_CS_fsm[1];
assign ap_CS_fsm_state3 = ap_CS_fsm[2];
assign ap_CS_fsm_state4 = ap_CS_fsm[3];
assign ap_done = op_30_ap_vld;
assign ap_ready = op_30_ap_vld;
assign conv_i482_fu_436_p1 = { 24'h000000, op_2 };
assign lhs_fu_367_p3 = { op_0, 6'h00 };
assign lshr_ln1497_fu_456_p2[3:0] = trunc_ln1497_fu_462_p1;
assign op_30 = { add_ln69_5_fu_690_p2[8], add_ln69_5_fu_690_p2[8], add_ln69_5_fu_690_p2[8], add_ln69_5_fu_690_p2[8], add_ln69_5_fu_690_p2[8], add_ln69_5_fu_690_p2[8], add_ln69_5_fu_690_p2[8], add_ln69_5_fu_690_p2[8], add_ln69_5_fu_690_p2[8], add_ln69_5_fu_690_p2[8], add_ln69_5_fu_690_p2[8], add_ln69_5_fu_690_p2[8], add_ln69_5_fu_690_p2[8], add_ln69_5_fu_690_p2[8], add_ln69_5_fu_690_p2[8], add_ln69_5_fu_690_p2[8], add_ln69_5_fu_690_p2[8], add_ln69_5_fu_690_p2[8], add_ln69_5_fu_690_p2[8], add_ln69_5_fu_690_p2[8], add_ln69_5_fu_690_p2[8], add_ln69_5_fu_690_p2[8], add_ln69_5_fu_690_p2[8], add_ln69_5_fu_690_p2 };
assign p_Result_1_fu_189_p1 = op_3;
assign p_Result_1_fu_189_p3 = op_3[31];
assign p_Result_2_fu_259_p3 = ret_V_20_fu_245_p2[32];
assign p_Result_3_fu_295_p1 = op_11;
assign p_Result_3_fu_295_p3 = op_11[7];
assign p_Result_4_fu_608_p3 = ret_V_22_reg_739[6];
assign p_Result_5_fu_552_p3 = ret_V_24_fu_536_p2[8];
assign p_Result_s_fu_399_p3 = ret_V_18_fu_383_p2[10];
assign ret_V_13_fu_542_p4 = ret_V_24_fu_536_p2[8:6];
assign ret_V_3_cast5_fu_335_p1 = op_3;
assign ret_V_3_cast5_fu_335_p4 = op_3[20:17];
assign ret_V_3_cast_fu_179_p1 = op_3;
assign ret_V_3_cast_fu_179_p4 = op_3[18:17];
assign ret_V_7_fu_285_p1 = op_11;
assign ret_V_7_fu_285_p4 = op_11[7:6];
assign ret_V_fu_389_p4 = ret_V_18_fu_383_p2[10:6];
assign rhs_1_fu_498_p3 = { select_ln850_7_fu_490_p3, 1'h0 };
assign rhs_fu_233_p3 = { op_4, 17'h00000 };
assign sext_ln1192_1_fu_478_p0 = op_6;
assign sext_ln1192_1_fu_478_p1 = { op_6[1], op_6[1], op_6[1], op_6[1], op_6[1], op_6 };
assign sext_ln1192_2_fu_506_p1 = { select_ln850_7_fu_490_p3[4], select_ln850_7_fu_490_p3, 1'h0 };
assign sext_ln1192_fu_375_p1 = { op_0[3], op_0, 6'h00 };
assign sext_ln1193_fu_592_p1 = { ret_V_19_reg_706[1], ret_V_19_reg_706[1], ret_V_19_reg_706 };
assign sext_ln1497_1_fu_452_p1 = { sub_ln1497_fu_446_p2[2], sub_ln1497_fu_446_p2[2], sub_ln1497_fu_446_p2[2], sub_ln1497_fu_446_p2[2], sub_ln1497_fu_446_p2[2], sub_ln1497_fu_446_p2[2], sub_ln1497_fu_446_p2[2], sub_ln1497_fu_446_p2[2], sub_ln1497_fu_446_p2[2], sub_ln1497_fu_446_p2[2], sub_ln1497_fu_446_p2[2], sub_ln1497_fu_446_p2[2], sub_ln1497_fu_446_p2[2], sub_ln1497_fu_446_p2[2], sub_ln1497_fu_446_p2[2], sub_ln1497_fu_446_p2[2], sub_ln1497_fu_446_p2[2], sub_ln1497_fu_446_p2[2], sub_ln1497_fu_446_p2[2], sub_ln1497_fu_446_p2[2], sub_ln1497_fu_446_p2[2], sub_ln1497_fu_446_p2[2], sub_ln1497_fu_446_p2[2], sub_ln1497_fu_446_p2[2], sub_ln1497_fu_446_p2[2], sub_ln1497_fu_446_p2[2], sub_ln1497_fu_446_p2[2], sub_ln1497_fu_446_p2[2], sub_ln1497_fu_446_p2[2], sub_ln1497_fu_446_p2 };
assign sext_ln1497_fu_426_p1 = { ret_V_9_reg_717[1], ret_V_9_reg_717 };
assign sext_ln27_fu_644_p1 = { op_12[7], op_12 };
assign sext_ln545_fu_423_p1 = { ret_V_9_reg_717[1], ret_V_9_reg_717[1], ret_V_9_reg_717[1], ret_V_9_reg_717[1], ret_V_9_reg_717[1], ret_V_9_reg_717[1], ret_V_9_reg_717[1], ret_V_9_reg_717[1], ret_V_9_reg_717[1], ret_V_9_reg_717[1], ret_V_9_reg_717[1], ret_V_9_reg_717[1], ret_V_9_reg_717[1], ret_V_9_reg_717[1], ret_V_9_reg_717[1], ret_V_9_reg_717[1], ret_V_9_reg_717[1], ret_V_9_reg_717[1], ret_V_9_reg_717[1], ret_V_9_reg_717[1], ret_V_9_reg_717[1], ret_V_9_reg_717[1], ret_V_9_reg_717[1], ret_V_9_reg_717[1], ret_V_9_reg_717[1], ret_V_9_reg_717[1], ret_V_9_reg_717[1], ret_V_9_reg_717[1], ret_V_9_reg_717[1], ret_V_9_reg_717[1], ret_V_9_reg_717 };
assign sext_ln69_1_fu_595_p1 = { ret_V_15_fu_584_p3[2], ret_V_15_fu_584_p3 };
assign sext_ln69_2_fu_666_p1 = { add_ln69_3_reg_749[3], add_ln69_3_reg_749[3], add_ln69_3_reg_749 };
assign sext_ln69_3_fu_687_p1 = { add_ln69_4_reg_759[5], add_ln69_4_reg_759[5], add_ln69_4_reg_759[5], add_ln69_4_reg_759 };
assign sext_ln69_fu_651_p1 = { ret_V_25_reg_724[3], ret_V_25_reg_724[3], ret_V_25_reg_724 };
assign sext_ln703_1_fu_229_p0 = op_3;
assign sext_ln703_1_fu_229_p1 = { op_3[31], op_3 };
assign sext_ln703_2_fu_533_p0 = op_11;
assign sext_ln703_2_fu_533_p1 = { op_11[7], op_11 };
assign sext_ln703_fu_379_p0 = op_1;
assign sext_ln703_fu_379_p1 = { op_1[7], op_1[7], op_1[7], op_1 };
assign sext_ln831_fu_640_p1 = { ret_V_23_fu_632_p3[6], ret_V_23_fu_632_p3[6], ret_V_23_fu_632_p3 };
assign sext_ln850_fu_605_p1 = { tmp_1_reg_744[5], tmp_1_reg_744 };
assign shl_ln1497_fu_440_p2[3:0] = trunc_ln1497_1_fu_466_p1;
assign tmp_4_fu_429_p3 = ret_V_9_reg_717[1];
assign tmp_fu_251_p3 = ret_V_20_fu_245_p2[17];
assign trunc_ln851_1_fu_197_p0 = op_3;
assign trunc_ln851_1_fu_197_p1 = op_3[16:0];
assign trunc_ln851_2_fu_303_p0 = op_11;
assign trunc_ln851_2_fu_303_p1 = op_11[5:0];
assign trunc_ln851_3_fu_615_p0 = op_6;
assign trunc_ln851_3_fu_615_p1 = op_6[0];
assign trunc_ln851_4_fu_560_p1 = ret_V_24_fu_536_p2[5:0];
assign trunc_ln851_fu_407_p0 = op_1;
assign trunc_ln851_fu_407_p1 = op_1[5:0];
assign zext_ln1192_fu_241_p1 = { 12'h000, op_4, 17'h00000 };
assign zext_ln27_fu_648_p1 = { 2'h0, op_15_V_reg_734 };
endmodule


// Product machine:
module top_A_times_top_B (ap_start, op_0, op_1, op_10, op_11, op_12, op_2, op_3, op_4, op_6, ap_clk, unsafe_signal);
input ap_start;
input [3:0] op_0;
input [7:0] op_1;
input [7:0] op_10;
input [7:0] op_11;
input [7:0] op_12;
input [7:0] op_2;
input [31:0] op_3;
input [3:0] op_4;
input [1:0] op_6;
input ap_clk;
output unsafe_signal;
reg _setup;
initial _setup = 1'b0;
always @ (posedge ap_clk) _setup <= 1'b1;
reg ap_start_internal;
always @ (posedge ap_clk) if (!_setup) ap_start_internal <= ap_start;
reg [3:0] op_0_internal;
always @ (posedge ap_clk) if (!_setup) op_0_internal <= op_0;
reg [7:0] op_1_internal;
always @ (posedge ap_clk) if (!_setup) op_1_internal <= op_1;
reg [7:0] op_10_internal;
always @ (posedge ap_clk) if (!_setup) op_10_internal <= op_10;
reg [7:0] op_11_internal;
always @ (posedge ap_clk) if (!_setup) op_11_internal <= op_11;
reg [7:0] op_12_internal;
always @ (posedge ap_clk) if (!_setup) op_12_internal <= op_12;
reg [7:0] op_2_internal;
always @ (posedge ap_clk) if (!_setup) op_2_internal <= op_2;
reg [31:0] op_3_internal;
always @ (posedge ap_clk) if (!_setup) op_3_internal <= op_3;
reg [3:0] op_4_internal;
always @ (posedge ap_clk) if (!_setup) op_4_internal <= op_4;
reg [1:0] op_6_internal;
always @ (posedge ap_clk) if (!_setup) op_6_internal <= op_6;
wire ap_done_A;
wire ap_done_B;
wire ap_done_eq;
assign ap_done_eq = ap_done_A == ap_done_B;
wire ap_idle_A;
wire ap_idle_B;
wire ap_idle_eq;
assign ap_idle_eq = ap_idle_A == ap_idle_B;
wire ap_ready_A;
wire ap_ready_B;
wire ap_ready_eq;
assign ap_ready_eq = ap_ready_A == ap_ready_B;
wire [31:0] op_30_A;
wire [31:0] op_30_B;
wire op_30_eq;
assign op_30_eq = op_30_A == op_30_B;
wire op_30_ap_vld_A;
wire op_30_ap_vld_B;
wire clk_enable_A;
wire clk_enable_B;
assign clk_enable_A = _setup & (~op_30_ap_vld_A | op_30_ap_vld_B);
assign clk_enable_B = _setup;
wire divergent;
assign divergent = ~(ap_done_eq & ap_idle_eq & ap_ready_eq & op_30_eq);
assign unsafe_signal = op_30_ap_vld_A & op_30_ap_vld_B & divergent;
top_A instance_A (
    .ap_clk(ap_clk),
    .clk_enable(clk_enable_A),
    .ap_start(ap_start_internal),
    .op_0(op_0_internal),
    .op_1(op_1_internal),
    .op_10(op_10_internal),
    .op_11(op_11_internal),
    .op_12(op_12_internal),
    .op_2(op_2_internal),
    .op_3(op_3_internal),
    .op_4(op_4_internal),
    .op_6(op_6_internal),
    .ap_done(ap_done_A),
    .ap_idle(ap_idle_A),
    .ap_ready(ap_ready_A),
    .op_30(op_30_A),
    .op_30_ap_vld(op_30_ap_vld_A)
);
top_B instance_B (
    .ap_clk(ap_clk),
    .clk_enable(clk_enable_B),
    .ap_start(ap_start_internal),
    .op_0(op_0_internal),
    .op_1(op_1_internal),
    .op_10(op_10_internal),
    .op_11(op_11_internal),
    .op_12(op_12_internal),
    .op_2(op_2_internal),
    .op_3(op_3_internal),
    .op_4(op_4_internal),
    .op_6(op_6_internal),
    .ap_done(ap_done_B),
    .ap_idle(ap_idle_B),
    .ap_ready(ap_ready_B),
    .op_30(op_30_B),
    .op_30_ap_vld(op_30_ap_vld_B)
);
endmodule
