// Processed by function `construct_kairos` in `verilog_tricks.py`.
// Machine A:
// Processed by function `add_clk_enable_signal` in `verilog_tricks.py`.
// Processed by function `remove_reset_signal` in `verilog_tricks.py`.
module top_A (
  ap_clk,
  ap_start,
  ap_done,
  ap_idle,
  ap_ready,
  op_0,
  op_3,
  op_4,
  op_5,
  op_6,
  op_7,
  op_9,
  op_10,
  op_11,
  op_12,
  op_13,
  op_15,
  op_16,
  op_17,
  op_18,
  op_19,
  op_33,
  op_33_ap_vld,
clk_enable
);
input clk_enable;


input ap_clk;
wire ap_rst;
assign ap_rst = op_33_ap_vld;
input ap_start;
input [7:0] op_0;
input [7:0] op_10;
input [3:0] op_11;
input [15:0] op_12;
input [1:0] op_13;
input [1:0] op_15;
input [31:0] op_16;
input [3:0] op_17;
input [7:0] op_18;
input [7:0] op_19;
input [7:0] op_3;
input op_4;
input [7:0] op_5;
input [3:0] op_6;
input [3:0] op_7;
input [1:0] op_9;
output ap_done;
output ap_idle;
output ap_ready;
output [31:0] op_33;
output op_33_ap_vld;


reg [31:0] add_ln691_1_reg_747;
reg [31:0] add_ln691_2_reg_769;
reg [31:0] add_ln691_4_reg_843;
reg [7:0] add_ln691_reg_725;
reg [8:0] add_ln69_1_reg_779;
reg [4:0] add_ln69_4_reg_816;
reg [31:0] add_ln69_reg_774;
reg [13:0] ap_CS_fsm = 14'h0001;
reg icmp_ln851_1_reg_714;
reg icmp_ln851_2_reg_794;
reg [31:0] op_31_V_reg_821;
reg [31:0] ret_V_11_cast_reg_762;
reg [8:0] ret_V_12_reg_704;
reg [33:0] ret_V_13_reg_735;
reg [33:0] ret_V_14_reg_757;
reg [31:0] ret_V_15_cast_reg_804;
reg [31:0] ret_V_16_reg_789;
reg [31:0] ret_V_18_cast_reg_836;
reg [31:0] ret_V_18_reg_811;
reg [33:0] ret_V_19_reg_831;
reg [31:0] ret_V_8_cast_reg_740;
reg [7:0] ret_V_reg_784;
reg [7:0] sext_ln850_reg_719;
reg [6:0] tmp_reg_709;
reg [32:0] _080_;
wire [31:0] _000_;
wire [31:0] _001_;
wire [31:0] _002_;
wire [7:0] _003_;
wire [8:0] _004_;
wire [4:0] _005_;
wire [31:0] _006_;
wire [13:0] _007_;
wire _008_;
wire _009_;
wire [31:0] _010_;
wire [31:0] _011_;
wire [8:0] _012_;
wire [33:0] _013_;
wire [33:0] _014_;
wire [31:0] _015_;
wire [31:0] _016_;
wire [32:0] _017_;
wire [31:0] _018_;
wire [31:0] _019_;
wire [33:0] _020_;
wire [31:0] _021_;
wire [4:0] _022_;
wire [7:0] _023_;
wire [6:0] _024_;
wire [1:0] _025_;
wire _026_;
wire _027_;
wire _028_;
wire _029_;
wire _030_;
wire _031_;
wire _032_;
wire _033_;
wire _034_;
wire _035_;
wire _036_;
wire _037_;
wire _038_;
wire _039_;
wire _040_;
wire _041_;
wire _042_;
wire _043_;
wire _044_;
wire _045_;
wire _046_;
wire _047_;
wire [31:0] add_ln691_1_fu_381_p2;
wire [31:0] add_ln691_2_fu_437_p2;
wire [31:0] add_ln691_3_fu_588_p2;
wire [31:0] add_ln691_4_fu_665_p2;
wire [7:0] add_ln691_fu_320_p2;
wire [8:0] add_ln69_1_fu_483_p2;
wire [31:0] add_ln69_3_fu_620_p2;
wire [4:0] add_ln69_4_fu_614_p2;
wire [31:0] add_ln69_fu_477_p2;
wire ap_CS_fsm_state1;
wire ap_CS_fsm_state10;
wire ap_CS_fsm_state11;
wire ap_CS_fsm_state12;
wire ap_CS_fsm_state13;
wire ap_CS_fsm_state14;
wire ap_CS_fsm_state2;
wire ap_CS_fsm_state3;
wire ap_CS_fsm_state4;
wire ap_CS_fsm_state5;
wire ap_CS_fsm_state6;
wire ap_CS_fsm_state7;
wire ap_CS_fsm_state8;
wire ap_CS_fsm_state9;
wire [13:0] ap_NS_fsm;
wire ap_clk;
wire ap_done;
wire ap_idle;
wire ap_ready;
wire ap_rst;
wire ap_start;
wire icmp_ln851_1_fu_311_p2;
wire icmp_ln851_2_fu_537_p2;
wire icmp_ln851_fu_251_p2;
wire [7:0] op_0;
wire [7:0] op_10;
wire [3:0] op_11;
wire [15:0] op_12;
wire [1:0] op_13;
wire [18:0] op_14_V_fu_543_p3;
wire [1:0] op_15;
wire [31:0] op_16;
wire [3:0] op_17;
wire [7:0] op_18;
wire [7:0] op_19;
wire [31:0] op_26_V_fu_510_p2;
wire [7:0] op_3;
wire [31:0] op_31_V_fu_628_p2;
wire [31:0] op_33;
wire op_33_ap_vld;
wire op_4;
wire op_4_read_read_fu_140_p2;
wire [7:0] op_5;
wire [3:0] op_6;
wire [3:0] op_7;
wire [1:0] op_9;
wire p_Result_1_fu_326_p3;
wire p_Result_2_fu_386_p3;
wire p_Result_3_fu_442_p3;
wire p_Result_4_fu_581_p3;
wire p_Result_5_fu_670_p3;
wire [13:0] p_Result_7_fu_529_p3;
wire p_Result_s_fu_239_p3;
wire [8:0] ret_V_12_fu_291_p2;
wire [33:0] ret_V_13_fu_365_p2;
wire [33:0] ret_V_14_fu_421_p2;
wire [31:0] ret_V_15_fu_458_p3;
wire [31:0] ret_V_16_fu_519_p2;
wire [46:0] ret_V_17_fu_565_p2;
wire [46:0] ret_V_17_reg_799;
wire [31:0] ret_V_18_fu_599_p3;
wire [33:0] ret_V_19_fu_649_p2;
wire [5:0] ret_V_1_fu_225_p4;
wire [31:0] ret_V_20_fu_686_p3;
wire [6:0] ret_V_2_fu_257_p2;
wire [7:0] ret_V_fu_501_p2;
wire [8:0] rhs_1_fu_283_p3;
wire [32:0] rhs_2_fu_409_p3;
wire [45:0] rhs_5_fu_554_p3;
wire [32:0] rhs_7_fu_638_p3;
wire [6:0] rhs_fu_489_p3;
wire [31:0] select_ln353_1_fu_402_p3;
wire [7:0] select_ln353_fu_346_p3;
wire [33:0] select_ln703_fu_333_p3;
wire [6:0] select_ln850_1_fu_275_p3;
wire [7:0] select_ln850_2_fu_341_p3;
wire [31:0] select_ln850_3_fu_452_p3;
wire [31:0] select_ln850_4_fu_593_p3;
wire [31:0] select_ln850_5_fu_680_p3;
wire [31:0] select_ln850_6_fu_397_p3;
wire [6:0] select_ln850_fu_267_p3;
wire [33:0] sext_ln1192_1_fu_361_p1;
wire [33:0] sext_ln1192_2_fu_417_p1;
wire [31:0] sext_ln1192_3_fu_515_p1;
wire [46:0] sext_ln1192_4_fu_561_p1;
wire [33:0] sext_ln1192_5_fu_645_p1;
wire [3:0] sext_ln1192_fu_263_p0;
wire [8:0] sext_ln1192_fu_263_p1;
wire [7:0] sext_ln1194_fu_497_p1;
wire [31:0] sext_ln69_1_fu_507_p1;
wire [31:0] sext_ln69_2_fu_693_p1;
wire [4:0] sext_ln69_3_fu_610_p1;
wire [31:0] sext_ln69_4_fu_625_p1;
wire [8:0] sext_ln69_fu_465_p1;
wire [46:0] sext_ln703_1_fu_550_p1;
wire [7:0] sext_ln703_2_fu_634_p0;
wire [33:0] sext_ln703_2_fu_634_p1;
wire [1:0] sext_ln703_fu_393_p0;
wire [33:0] sext_ln703_fu_393_p1;
wire [6:0] sext_ln835_fu_235_p1;
wire [7:0] sext_ln850_fu_317_p1;
wire [8:0] tmp_3_fu_353_p3;
wire [3:0] trunc_ln851_1_fu_307_p0;
wire [1:0] trunc_ln851_1_fu_307_p1;
wire [1:0] trunc_ln851_2_fu_449_p0;
wire trunc_ln851_2_fu_449_p1;
wire [2:0] trunc_ln851_3_fu_525_p1;
wire [7:0] trunc_ln851_4_fu_677_p0;
wire trunc_ln851_4_fu_677_p1;
wire [1:0] trunc_ln851_fu_247_p1;
wire [31:0] zext_ln69_1_fu_473_p1;
wire [4:0] zext_ln69_2_fu_606_p1;
wire [8:0] zext_ln69_fu_469_p1;


assign add_ln691_1_fu_381_p2 = ret_V_8_cast_reg_740 + 1'h1;
assign add_ln691_2_fu_437_p2 = ret_V_11_cast_reg_762 + 1'h1;
assign add_ln691_3_fu_588_p2 = ret_V_15_cast_reg_804 + 1'h1;
assign add_ln691_4_fu_665_p2 = ret_V_18_cast_reg_836 + 1'h1;
assign add_ln691_fu_320_p2 = $signed(tmp_reg_709) + $signed(2'h1);
assign add_ln69_1_fu_483_p2 = $signed(op_10) + $signed({ 1'h0, op_11 });
assign add_ln69_3_fu_620_p2 = ret_V_18_reg_811 + op_16;
assign add_ln69_4_fu_614_p2 = $signed(op_17) + $signed({ 1'h0, op_15 });
assign add_ln69_fu_477_p2 = ret_V_15_fu_458_p3 + op_12;
assign op_26_V_fu_510_p2 = $signed(add_ln69_1_reg_779) + $signed(add_ln69_reg_774);
assign op_31_V_fu_628_p2 = $signed(add_ln69_4_reg_816) + $signed(add_ln69_3_fu_620_p2);
assign op_33 = $signed(ret_V_20_fu_686_p3) + $signed(op_19);
assign ret_V_12_fu_291_p2 = $signed({ select_ln850_1_fu_275_p3, 2'h0 }) + $signed(op_7);
assign ret_V_13_fu_365_p2 = $signed({ select_ln353_fu_346_p3, 1'h0 }) + $signed(select_ln703_fu_333_p3);
assign ret_V_14_fu_421_p2 = $signed({ select_ln353_1_fu_402_p3, 1'h0 }) + $signed(op_9);
assign ret_V_16_fu_519_p2 = $signed(op_26_V_fu_510_p2) + $signed(op_13);
assign ret_V_17_fu_565_p2 = $signed({ ret_V_16_reg_789, 14'h0000 }) + $signed({ ret_V_reg_784, 11'h000 });
assign ret_V_19_fu_649_p2 = $signed({ op_31_V_reg_821, 1'h0 }) + $signed(op_18);
assign ret_V_2_fu_257_p2 = $signed(op_5[7:2]) + $signed(2'h1);
assign _026_ = op_4 & ap_CS_fsm[3];
assign _027_ = icmp_ln851_1_reg_714 & ap_CS_fsm[1];
assign _028_ = ap_CS_fsm[0] & _030_;
assign _029_ = ap_CS_fsm[0] & ap_start;
assign ret_V_fu_501_p2 = { op_6[3], op_6, 3'h0 } & op_3;
assign _030_ = ~ ap_start;
assign _031_ = ! op_5[1:0];
assign _032_ = | op_7[1:0];
assign _033_ = | { ret_V_fu_501_p2[2:0], 11'h000 };
always @(posedge ap_clk)
ret_V_reg_784[2:0] <= 3'h0;
always @(posedge ap_clk)
sext_ln850_reg_719 <= _023_;
always @(posedge ap_clk)
ret_V_19_reg_831 <= _020_;
always @(posedge ap_clk)
ret_V_18_cast_reg_836 <= _018_;
always @(posedge ap_clk)
_080_ <= _017_;
assign ret_V_17_reg_799[46:14] = _080_;
always @(posedge ap_clk)
ret_V_15_cast_reg_804 <= _015_;
always @(posedge ap_clk)
ret_V_13_reg_735 <= _013_;
always @(posedge ap_clk)
ret_V_8_cast_reg_740 <= _021_;
always @(posedge ap_clk)
ret_V_14_reg_757 <= _014_;
always @(posedge ap_clk)
ret_V_11_cast_reg_762 <= _011_;
always @(posedge ap_clk)
op_31_V_reg_821 <= _010_;
always @(posedge ap_clk)
ret_V_reg_784[7:3] <= _022_;
always @(posedge ap_clk)
ret_V_16_reg_789 <= _016_;
always @(posedge ap_clk)
icmp_ln851_2_reg_794 <= _009_;
always @(posedge ap_clk)
ret_V_12_reg_704 <= _012_;
always @(posedge ap_clk)
tmp_reg_709 <= _024_;
always @(posedge ap_clk)
icmp_ln851_1_reg_714 <= _008_;
always @(posedge ap_clk)
ret_V_18_reg_811 <= _019_;
always @(posedge ap_clk)
add_ln69_4_reg_816 <= _005_;
always @(posedge ap_clk)
add_ln69_reg_774 <= _006_;
always @(posedge ap_clk)
add_ln69_1_reg_779 <= _004_;
always @(posedge ap_clk)
add_ln691_reg_725 <= _003_;
always @(posedge ap_clk)
add_ln691_4_reg_843 <= _002_;
always @(posedge ap_clk)
add_ln691_2_reg_769 <= _001_;
always @(posedge ap_clk)
add_ln691_1_reg_747 <= _000_;
always @(posedge ap_clk)
ap_CS_fsm <= _007_;
assign _025_ = _029_ ? 2'h2 : 2'h1;
assign _034_ = ap_CS_fsm == 1'h1;
function [13:0] _104_;
input [13:0] a;
input [195:0] b;
input [13:0] s;
case (s)
14'b00000000000001:
_104_ = b[13:0];
14'b00000000000010:
_104_ = b[27:14];
14'b00000000000100:
_104_ = b[41:28];
14'b00000000001000:
_104_ = b[55:42];
14'b00000000010000:
_104_ = b[69:56];
14'b00000000100000:
_104_ = b[83:70];
14'b00000001000000:
_104_ = b[97:84];
14'b00000010000000:
_104_ = b[111:98];
14'b00000100000000:
_104_ = b[125:112];
14'b00001000000000:
_104_ = b[139:126];
14'b00010000000000:
_104_ = b[153:140];
14'b00100000000000:
_104_ = b[167:154];
14'b01000000000000:
_104_ = b[181:168];
14'b10000000000000:
_104_ = b[195:182];
14'b00000000000000:
_104_ = a;
default:
_104_ = 14'bx;
endcase
endfunction
assign ap_NS_fsm = _104_(14'hxxxx, { 12'h000, _025_, 182'h0004002001000800400200100080040020010008000001 }, { _034_, _047_, _046_, _045_, _044_, _043_, _042_, _041_, _040_, _039_, _038_, _037_, _036_, _035_ });
assign _035_ = ap_CS_fsm == 14'h2000;
assign _036_ = ap_CS_fsm == 13'h1000;
assign _037_ = ap_CS_fsm == 12'h800;
assign _038_ = ap_CS_fsm == 11'h400;
assign _039_ = ap_CS_fsm == 10'h200;
assign _040_ = ap_CS_fsm == 9'h100;
assign _041_ = ap_CS_fsm == 8'h80;
assign _042_ = ap_CS_fsm == 7'h40;
assign _043_ = ap_CS_fsm == 6'h20;
assign _044_ = ap_CS_fsm == 5'h10;
assign _045_ = ap_CS_fsm == 4'h8;
assign _046_ = ap_CS_fsm == 3'h4;
assign _047_ = ap_CS_fsm == 2'h2;
assign op_33_ap_vld = ap_CS_fsm[13] ? 1'h1 : 1'h0;
assign ap_idle = _028_ ? 1'h1 : 1'h0;
assign _023_ = ap_CS_fsm[1] ? { tmp_reg_709[6], tmp_reg_709 } : sext_ln850_reg_719;
assign _018_ = ap_CS_fsm[11] ? ret_V_19_fu_649_p2[32:1] : ret_V_18_cast_reg_836;
assign _020_ = ap_CS_fsm[11] ? ret_V_19_fu_649_p2 : ret_V_19_reg_831;
assign _015_ = ap_CS_fsm[8] ? ret_V_17_fu_565_p2[45:14] : ret_V_15_cast_reg_804;
assign _017_ = ap_CS_fsm[8] ? ret_V_17_fu_565_p2[46:14] : ret_V_17_reg_799[46:14];
assign _021_ = ap_CS_fsm[2] ? ret_V_13_fu_365_p2[32:1] : ret_V_8_cast_reg_740;
assign _013_ = ap_CS_fsm[2] ? ret_V_13_fu_365_p2 : ret_V_13_reg_735;
assign _011_ = ap_CS_fsm[4] ? ret_V_14_fu_421_p2[32:1] : ret_V_11_cast_reg_762;
assign _014_ = ap_CS_fsm[4] ? ret_V_14_fu_421_p2 : ret_V_14_reg_757;
assign _010_ = ap_CS_fsm[10] ? op_31_V_fu_628_p2 : op_31_V_reg_821;
assign _009_ = ap_CS_fsm[7] ? icmp_ln851_2_fu_537_p2 : icmp_ln851_2_reg_794;
assign _016_ = ap_CS_fsm[7] ? ret_V_16_fu_519_p2 : ret_V_16_reg_789;
assign _022_ = ap_CS_fsm[7] ? ret_V_fu_501_p2[7:3] : ret_V_reg_784[7:3];
assign _008_ = ap_CS_fsm[0] ? icmp_ln851_1_fu_311_p2 : icmp_ln851_1_reg_714;
assign _024_ = ap_CS_fsm[0] ? ret_V_12_fu_291_p2[8:2] : tmp_reg_709;
assign _012_ = ap_CS_fsm[0] ? ret_V_12_fu_291_p2 : ret_V_12_reg_704;
assign _005_ = ap_CS_fsm[9] ? add_ln69_4_fu_614_p2 : add_ln69_4_reg_816;
assign _019_ = ap_CS_fsm[9] ? ret_V_18_fu_599_p3 : ret_V_18_reg_811;
assign _004_ = ap_CS_fsm[6] ? add_ln69_1_fu_483_p2 : add_ln69_1_reg_779;
assign _006_ = ap_CS_fsm[6] ? add_ln69_fu_477_p2 : add_ln69_reg_774;
assign _003_ = _027_ ? add_ln691_fu_320_p2 : add_ln691_reg_725;
assign _002_ = ap_CS_fsm[12] ? add_ln691_4_fu_665_p2 : add_ln691_4_reg_843;
assign _001_ = ap_CS_fsm[5] ? add_ln691_2_fu_437_p2 : add_ln691_2_reg_769;
assign _000_ = _026_ ? add_ln691_1_fu_381_p2 : add_ln691_1_reg_747;
assign _007_ = ap_rst ? 14'h0001 : ap_NS_fsm;
assign icmp_ln851_1_fu_311_p2 = _032_ ? 1'h1 : 1'h0;
assign icmp_ln851_2_fu_537_p2 = _033_ ? 1'h1 : 1'h0;
assign icmp_ln851_fu_251_p2 = _031_ ? 1'h1 : 1'h0;
assign ret_V_15_fu_458_p3 = ret_V_14_reg_757[33] ? select_ln850_3_fu_452_p3 : ret_V_11_cast_reg_762;
assign ret_V_18_fu_599_p3 = ret_V_17_reg_799[46] ? select_ln850_4_fu_593_p3 : ret_V_15_cast_reg_804;
assign ret_V_20_fu_686_p3 = ret_V_19_reg_831[33] ? select_ln850_5_fu_680_p3 : ret_V_18_cast_reg_836;
assign select_ln353_1_fu_402_p3 = ret_V_13_reg_735[33] ? select_ln850_6_fu_397_p3 : ret_V_8_cast_reg_740;
assign select_ln353_fu_346_p3 = ret_V_12_reg_704[8] ? select_ln850_2_fu_341_p3 : sext_ln850_reg_719;
assign select_ln703_fu_333_p3 = op_4 ? 34'h3ffffffff : 34'h000000000;
assign select_ln850_1_fu_275_p3 = op_5[7] ? select_ln850_fu_267_p3 : { 2'h0, op_5[6:2] };
assign select_ln850_2_fu_341_p3 = icmp_ln851_1_reg_714 ? add_ln691_reg_725 : sext_ln850_reg_719;
assign select_ln850_3_fu_452_p3 = op_9[0] ? add_ln691_2_reg_769 : ret_V_11_cast_reg_762;
assign select_ln850_4_fu_593_p3 = icmp_ln851_2_reg_794 ? add_ln691_3_fu_588_p2 : ret_V_15_cast_reg_804;
assign select_ln850_5_fu_680_p3 = op_18[0] ? add_ln691_4_reg_843 : ret_V_18_cast_reg_836;
assign select_ln850_6_fu_397_p3 = op_4 ? add_ln691_1_reg_747 : ret_V_8_cast_reg_740;
assign select_ln850_fu_267_p3 = icmp_ln851_fu_251_p2 ? { 2'h3, op_5[6:2] } : ret_V_2_fu_257_p2;
assign ap_CS_fsm_state1 = ap_CS_fsm[0];
assign ap_CS_fsm_state10 = ap_CS_fsm[9];
assign ap_CS_fsm_state11 = ap_CS_fsm[10];
assign ap_CS_fsm_state12 = ap_CS_fsm[11];
assign ap_CS_fsm_state13 = ap_CS_fsm[12];
assign ap_CS_fsm_state14 = ap_CS_fsm[13];
assign ap_CS_fsm_state2 = ap_CS_fsm[1];
assign ap_CS_fsm_state3 = ap_CS_fsm[2];
assign ap_CS_fsm_state4 = ap_CS_fsm[3];
assign ap_CS_fsm_state5 = ap_CS_fsm[4];
assign ap_CS_fsm_state6 = ap_CS_fsm[5];
assign ap_CS_fsm_state7 = ap_CS_fsm[6];
assign ap_CS_fsm_state8 = ap_CS_fsm[7];
assign ap_CS_fsm_state9 = ap_CS_fsm[8];
assign ap_done = op_33_ap_vld;
assign ap_ready = op_33_ap_vld;
assign op_14_V_fu_543_p3 = { ret_V_reg_784, 11'h000 };
assign op_4_read_read_fu_140_p2 = op_4;
assign p_Result_1_fu_326_p3 = ret_V_12_reg_704[8];
assign p_Result_2_fu_386_p3 = ret_V_13_reg_735[33];
assign p_Result_3_fu_442_p3 = ret_V_14_reg_757[33];
assign p_Result_4_fu_581_p3 = ret_V_17_reg_799[46];
assign p_Result_5_fu_670_p3 = ret_V_19_reg_831[33];
assign p_Result_7_fu_529_p3 = { ret_V_fu_501_p2[2:0], 11'h000 };
assign p_Result_s_fu_239_p3 = op_5[7];
assign ret_V_1_fu_225_p4 = op_5[7:2];
assign rhs_1_fu_283_p3 = { select_ln850_1_fu_275_p3, 2'h0 };
assign rhs_2_fu_409_p3 = { select_ln353_1_fu_402_p3, 1'h0 };
assign rhs_5_fu_554_p3 = { ret_V_16_reg_789, 14'h0000 };
assign rhs_7_fu_638_p3 = { op_31_V_reg_821, 1'h0 };
assign rhs_fu_489_p3 = { op_6, 3'h0 };
assign sext_ln1192_1_fu_361_p1 = { select_ln353_fu_346_p3[7], select_ln353_fu_346_p3[7], select_ln353_fu_346_p3[7], select_ln353_fu_346_p3[7], select_ln353_fu_346_p3[7], select_ln353_fu_346_p3[7], select_ln353_fu_346_p3[7], select_ln353_fu_346_p3[7], select_ln353_fu_346_p3[7], select_ln353_fu_346_p3[7], select_ln353_fu_346_p3[7], select_ln353_fu_346_p3[7], select_ln353_fu_346_p3[7], select_ln353_fu_346_p3[7], select_ln353_fu_346_p3[7], select_ln353_fu_346_p3[7], select_ln353_fu_346_p3[7], select_ln353_fu_346_p3[7], select_ln353_fu_346_p3[7], select_ln353_fu_346_p3[7], select_ln353_fu_346_p3[7], select_ln353_fu_346_p3[7], select_ln353_fu_346_p3[7], select_ln353_fu_346_p3[7], select_ln353_fu_346_p3[7], select_ln353_fu_346_p3, 1'h0 };
assign sext_ln1192_2_fu_417_p1 = { select_ln353_1_fu_402_p3[31], select_ln353_1_fu_402_p3, 1'h0 };
assign sext_ln1192_3_fu_515_p1 = { op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13 };
assign sext_ln1192_4_fu_561_p1 = { ret_V_16_reg_789[31], ret_V_16_reg_789, 14'h0000 };
assign sext_ln1192_5_fu_645_p1 = { op_31_V_reg_821[31], op_31_V_reg_821, 1'h0 };
assign sext_ln1192_fu_263_p0 = op_7;
assign sext_ln1192_fu_263_p1 = { op_7[3], op_7[3], op_7[3], op_7[3], op_7[3], op_7 };
assign sext_ln1194_fu_497_p1 = { op_6[3], op_6, 3'h0 };
assign sext_ln69_1_fu_507_p1 = { add_ln69_1_reg_779[8], add_ln69_1_reg_779[8], add_ln69_1_reg_779[8], add_ln69_1_reg_779[8], add_ln69_1_reg_779[8], add_ln69_1_reg_779[8], add_ln69_1_reg_779[8], add_ln69_1_reg_779[8], add_ln69_1_reg_779[8], add_ln69_1_reg_779[8], add_ln69_1_reg_779[8], add_ln69_1_reg_779[8], add_ln69_1_reg_779[8], add_ln69_1_reg_779[8], add_ln69_1_reg_779[8], add_ln69_1_reg_779[8], add_ln69_1_reg_779[8], add_ln69_1_reg_779[8], add_ln69_1_reg_779[8], add_ln69_1_reg_779[8], add_ln69_1_reg_779[8], add_ln69_1_reg_779[8], add_ln69_1_reg_779[8], add_ln69_1_reg_779 };
assign sext_ln69_2_fu_693_p1 = { op_19[7], op_19[7], op_19[7], op_19[7], op_19[7], op_19[7], op_19[7], op_19[7], op_19[7], op_19[7], op_19[7], op_19[7], op_19[7], op_19[7], op_19[7], op_19[7], op_19[7], op_19[7], op_19[7], op_19[7], op_19[7], op_19[7], op_19[7], op_19[7], op_19 };
assign sext_ln69_3_fu_610_p1 = { op_17[3], op_17 };
assign sext_ln69_4_fu_625_p1 = { add_ln69_4_reg_816[4], add_ln69_4_reg_816[4], add_ln69_4_reg_816[4], add_ln69_4_reg_816[4], add_ln69_4_reg_816[4], add_ln69_4_reg_816[4], add_ln69_4_reg_816[4], add_ln69_4_reg_816[4], add_ln69_4_reg_816[4], add_ln69_4_reg_816[4], add_ln69_4_reg_816[4], add_ln69_4_reg_816[4], add_ln69_4_reg_816[4], add_ln69_4_reg_816[4], add_ln69_4_reg_816[4], add_ln69_4_reg_816[4], add_ln69_4_reg_816[4], add_ln69_4_reg_816[4], add_ln69_4_reg_816[4], add_ln69_4_reg_816[4], add_ln69_4_reg_816[4], add_ln69_4_reg_816[4], add_ln69_4_reg_816[4], add_ln69_4_reg_816[4], add_ln69_4_reg_816[4], add_ln69_4_reg_816[4], add_ln69_4_reg_816[4], add_ln69_4_reg_816 };
assign sext_ln69_fu_465_p1 = { op_10[7], op_10 };
assign sext_ln703_1_fu_550_p1 = { ret_V_reg_784[7], ret_V_reg_784[7], ret_V_reg_784[7], ret_V_reg_784[7], ret_V_reg_784[7], ret_V_reg_784[7], ret_V_reg_784[7], ret_V_reg_784[7], ret_V_reg_784[7], ret_V_reg_784[7], ret_V_reg_784[7], ret_V_reg_784[7], ret_V_reg_784[7], ret_V_reg_784[7], ret_V_reg_784[7], ret_V_reg_784[7], ret_V_reg_784[7], ret_V_reg_784[7], ret_V_reg_784[7], ret_V_reg_784[7], ret_V_reg_784[7], ret_V_reg_784[7], ret_V_reg_784[7], ret_V_reg_784[7], ret_V_reg_784[7], ret_V_reg_784[7], ret_V_reg_784[7], ret_V_reg_784[7], ret_V_reg_784, 11'h000 };
assign sext_ln703_2_fu_634_p0 = op_18;
assign sext_ln703_2_fu_634_p1 = { op_18[7], op_18[7], op_18[7], op_18[7], op_18[7], op_18[7], op_18[7], op_18[7], op_18[7], op_18[7], op_18[7], op_18[7], op_18[7], op_18[7], op_18[7], op_18[7], op_18[7], op_18[7], op_18[7], op_18[7], op_18[7], op_18[7], op_18[7], op_18[7], op_18[7], op_18[7], op_18 };
assign sext_ln703_fu_393_p0 = op_9;
assign sext_ln703_fu_393_p1 = { op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9 };
assign sext_ln835_fu_235_p1 = { op_5[7], op_5[7:2] };
assign sext_ln850_fu_317_p1 = { tmp_reg_709[6], tmp_reg_709 };
assign tmp_3_fu_353_p3 = { select_ln353_fu_346_p3, 1'h0 };
assign trunc_ln851_1_fu_307_p0 = op_7;
assign trunc_ln851_1_fu_307_p1 = op_7[1:0];
assign trunc_ln851_2_fu_449_p0 = op_9;
assign trunc_ln851_2_fu_449_p1 = op_9[0];
assign trunc_ln851_3_fu_525_p1 = ret_V_fu_501_p2[2:0];
assign trunc_ln851_4_fu_677_p0 = op_18;
assign trunc_ln851_4_fu_677_p1 = op_18[0];
assign trunc_ln851_fu_247_p1 = op_5[1:0];
assign zext_ln69_1_fu_473_p1 = { 16'h0000, op_12 };
assign zext_ln69_2_fu_606_p1 = { 3'h0, op_15 };
assign zext_ln69_fu_469_p1 = { 5'h00, op_11 };
endmodule


// Machine B:
// Processed by function `add_clk_enable_signal` in `verilog_tricks.py`.
// Processed by function `remove_reset_signal` in `verilog_tricks.py`.
module top_B (
  ap_clk,
  ap_start,
  ap_done,
  ap_idle,
  ap_ready,
  op_0,
  op_3,
  op_4,
  op_5,
  op_6,
  op_7,
  op_9,
  op_10,
  op_11,
  op_12,
  op_13,
  op_15,
  op_16,
  op_17,
  op_18,
  op_19,
  op_33,
  op_33_ap_vld,
clk_enable
);
input clk_enable;


input ap_clk;
wire ap_rst;
assign ap_rst = op_33_ap_vld;
input ap_start;
input [7:0] op_0;
input [7:0] op_10;
input [3:0] op_11;
input [15:0] op_12;
input [1:0] op_13;
input [1:0] op_15;
input [31:0] op_16;
input [3:0] op_17;
input [7:0] op_18;
input [7:0] op_19;
input [7:0] op_3;
input op_4;
input [7:0] op_5;
input [3:0] op_6;
input [3:0] op_7;
input [1:0] op_9;
output ap_done;
output ap_idle;
output ap_ready;
output [31:0] op_33;
output op_33_ap_vld;


reg [15:0] \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_4_U.ain_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_4_U.bin_s1 ;
reg \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_4_U.carry_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_4_U.sum_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_4_U.ain_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_4_U.bin_s1 ;
reg \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_4_U.carry_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_4_U.sum_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_4_U.ain_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_4_U.bin_s1 ;
reg \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_4_U.carry_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_4_U.sum_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.ain_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.bin_s1 ;
reg \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.carry_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.sum_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_4_U.ain_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_4_U.bin_s1 ;
reg \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_4_U.carry_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_4_U.sum_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.ain_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.bin_s1 ;
reg \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.carry_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.sum_s1 ;
reg [15:0] \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.ain_s1 ;
reg [15:0] \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.bin_s1 ;
reg \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.carry_s1 ;
reg [15:0] \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.sum_s1 ;
reg [15:0] \add_32ns_32s_32_2_1_U19.top_add_32ns_32s_32_2_1_Adder_8_U.ain_s1 ;
reg [15:0] \add_32ns_32s_32_2_1_U19.top_add_32ns_32s_32_2_1_Adder_8_U.bin_s1 ;
reg \add_32ns_32s_32_2_1_U19.top_add_32ns_32s_32_2_1_Adder_8_U.carry_s1 ;
reg [15:0] \add_32ns_32s_32_2_1_U19.top_add_32ns_32s_32_2_1_Adder_8_U.sum_s1 ;
reg [15:0] \add_32s_32ns_32_2_1_U10.top_add_32s_32ns_32_2_1_Adder_7_U.ain_s1 ;
reg [15:0] \add_32s_32ns_32_2_1_U10.top_add_32s_32ns_32_2_1_Adder_7_U.bin_s1 ;
reg \add_32s_32ns_32_2_1_U10.top_add_32s_32ns_32_2_1_Adder_7_U.carry_s1 ;
reg [15:0] \add_32s_32ns_32_2_1_U10.top_add_32s_32ns_32_2_1_Adder_7_U.sum_s1 ;
reg [15:0] \add_32s_32ns_32_2_1_U16.top_add_32s_32ns_32_2_1_Adder_7_U.ain_s1 ;
reg [15:0] \add_32s_32ns_32_2_1_U16.top_add_32s_32ns_32_2_1_Adder_7_U.bin_s1 ;
reg \add_32s_32ns_32_2_1_U16.top_add_32s_32ns_32_2_1_Adder_7_U.carry_s1 ;
reg [15:0] \add_32s_32ns_32_2_1_U16.top_add_32s_32ns_32_2_1_Adder_7_U.sum_s1 ;
reg [16:0] \add_34s_34ns_34_2_1_U4.top_add_34s_34ns_34_2_1_Adder_3_U.ain_s1 ;
reg [16:0] \add_34s_34ns_34_2_1_U4.top_add_34s_34ns_34_2_1_Adder_3_U.bin_s1 ;
reg \add_34s_34ns_34_2_1_U4.top_add_34s_34ns_34_2_1_Adder_3_U.carry_s1 ;
reg [16:0] \add_34s_34ns_34_2_1_U4.top_add_34s_34ns_34_2_1_Adder_3_U.sum_s1 ;
reg [16:0] \add_34s_34s_34_2_1_U17.top_add_34s_34s_34_2_1_Adder_5_U.ain_s1 ;
reg [16:0] \add_34s_34s_34_2_1_U17.top_add_34s_34s_34_2_1_Adder_5_U.bin_s1 ;
reg \add_34s_34s_34_2_1_U17.top_add_34s_34s_34_2_1_Adder_5_U.carry_s1 ;
reg [16:0] \add_34s_34s_34_2_1_U17.top_add_34s_34s_34_2_1_Adder_5_U.sum_s1 ;
reg [16:0] \add_34s_34s_34_2_1_U6.top_add_34s_34s_34_2_1_Adder_5_U.ain_s1 ;
reg [16:0] \add_34s_34s_34_2_1_U6.top_add_34s_34s_34_2_1_Adder_5_U.bin_s1 ;
reg \add_34s_34s_34_2_1_U6.top_add_34s_34s_34_2_1_Adder_5_U.carry_s1 ;
reg [16:0] \add_34s_34s_34_2_1_U6.top_add_34s_34s_34_2_1_Adder_5_U.sum_s1 ;
reg [23:0] \add_47s_47s_47_2_1_U12.top_add_47s_47s_47_2_1_Adder_9_U.ain_s1 ;
reg [23:0] \add_47s_47s_47_2_1_U12.top_add_47s_47s_47_2_1_Adder_9_U.bin_s1 ;
reg \add_47s_47s_47_2_1_U12.top_add_47s_47s_47_2_1_Adder_9_U.carry_s1 ;
reg [22:0] \add_47s_47s_47_2_1_U12.top_add_47s_47s_47_2_1_Adder_9_U.sum_s1 ;
reg [31:0] add_ln691_1_reg_769;
reg [31:0] add_ln691_2_reg_806;
reg [31:0] add_ln691_3_reg_888;
reg [31:0] add_ln691_4_reg_950;
reg [7:0] add_ln691_reg_732;
reg [8:0] add_ln69_1_reg_826;
reg [31:0] add_ln69_3_reg_903;
reg [4:0] add_ln69_4_reg_908;
reg [31:0] add_ln69_reg_821;
reg [35:0] ap_CS_fsm = 36'h000000001;
reg icmp_ln851_1_reg_721;
reg icmp_ln851_2_reg_871;
reg icmp_ln851_reg_701;
reg [31:0] op_26_V_reg_836;
reg [31:0] op_31_V_reg_918;
reg [31:0] ret_V_11_cast_reg_799;
reg [8:0] ret_V_12_reg_711;
reg [33:0] ret_V_13_reg_757;
reg [33:0] ret_V_14_reg_794;
reg [31:0] ret_V_15_cast_reg_881;
reg [31:0] ret_V_15_reg_811;
reg [31:0] ret_V_16_reg_851;
reg [46:0] ret_V_17_reg_876;
reg [31:0] ret_V_18_cast_reg_943;
reg [31:0] ret_V_18_reg_893;
reg [33:0] ret_V_19_reg_938;
reg [31:0] ret_V_20_reg_955;
reg [6:0] ret_V_2_reg_706;
reg [31:0] ret_V_8_cast_reg_762;
reg [7:0] ret_V_reg_846;
reg [31:0] select_ln353_1_reg_774;
reg [7:0] select_ln353_reg_747;
reg [33:0] select_ln703_reg_742;
reg [6:0] sext_ln835_reg_695;
reg [7:0] sext_ln850_reg_726;
reg [6:0] tmp_reg_716;
reg [2:0] trunc_ln851_3_reg_856;
wire [31:0] _000_;
wire [31:0] _001_;
wire [31:0] _002_;
wire [31:0] _003_;
wire [7:0] _004_;
wire [8:0] _005_;
wire [31:0] _006_;
wire [4:0] _007_;
wire [31:0] _008_;
wire [35:0] _009_;
wire _010_;
wire _011_;
wire _012_;
wire [31:0] _013_;
wire [31:0] _014_;
wire [31:0] _015_;
wire [8:0] _016_;
wire [33:0] _017_;
wire [33:0] _018_;
wire [31:0] _019_;
wire [31:0] _020_;
wire [31:0] _021_;
wire [46:0] _022_;
wire [31:0] _023_;
wire [31:0] _024_;
wire [33:0] _025_;
wire [31:0] _026_;
wire [6:0] _027_;
wire [31:0] _028_;
wire [4:0] _029_;
wire [31:0] _030_;
wire [7:0] _031_;
wire [33:0] _032_;
wire [6:0] _033_;
wire [7:0] _034_;
wire [6:0] _035_;
wire [1:0] _036_;
wire _037_;
wire _038_;
wire _039_;
wire _040_;
wire _041_;
wire _042_;
wire _043_;
wire [15:0] _044_;
wire [15:0] _045_;
wire _046_;
wire [15:0] _047_;
wire [16:0] _048_;
wire [16:0] _049_;
wire [15:0] _050_;
wire [15:0] _051_;
wire _052_;
wire [15:0] _053_;
wire [16:0] _054_;
wire [16:0] _055_;
wire [15:0] _056_;
wire [15:0] _057_;
wire _058_;
wire [15:0] _059_;
wire [16:0] _060_;
wire [16:0] _061_;
wire [15:0] _062_;
wire [15:0] _063_;
wire _064_;
wire [15:0] _065_;
wire [16:0] _066_;
wire [16:0] _067_;
wire [15:0] _068_;
wire [15:0] _069_;
wire _070_;
wire [15:0] _071_;
wire [16:0] _072_;
wire [16:0] _073_;
wire [15:0] _074_;
wire [15:0] _075_;
wire _076_;
wire [15:0] _077_;
wire [16:0] _078_;
wire [16:0] _079_;
wire [15:0] _080_;
wire [15:0] _081_;
wire _082_;
wire [15:0] _083_;
wire [16:0] _084_;
wire [16:0] _085_;
wire [15:0] _086_;
wire [15:0] _087_;
wire _088_;
wire [15:0] _089_;
wire [16:0] _090_;
wire [16:0] _091_;
wire [15:0] _092_;
wire [15:0] _093_;
wire _094_;
wire [15:0] _095_;
wire [16:0] _096_;
wire [16:0] _097_;
wire [15:0] _098_;
wire [15:0] _099_;
wire _100_;
wire [15:0] _101_;
wire [16:0] _102_;
wire [16:0] _103_;
wire [16:0] _104_;
wire [16:0] _105_;
wire _106_;
wire [16:0] _107_;
wire [17:0] _108_;
wire [17:0] _109_;
wire [16:0] _110_;
wire [16:0] _111_;
wire _112_;
wire [16:0] _113_;
wire [17:0] _114_;
wire [17:0] _115_;
wire [16:0] _116_;
wire [16:0] _117_;
wire _118_;
wire [16:0] _119_;
wire [17:0] _120_;
wire [17:0] _121_;
wire [23:0] _122_;
wire [23:0] _123_;
wire _124_;
wire [22:0] _125_;
wire [23:0] _126_;
wire [24:0] _127_;
wire _128_;
wire _129_;
wire _130_;
wire _131_;
wire _132_;
wire _133_;
wire _134_;
wire _135_;
wire _136_;
wire _137_;
wire _138_;
wire _139_;
wire _140_;
wire _141_;
wire _142_;
wire _143_;
wire _144_;
wire _145_;
wire _146_;
wire _147_;
wire _148_;
wire _149_;
wire _150_;
wire _151_;
wire _152_;
wire _153_;
wire _154_;
wire _155_;
wire _156_;
wire _157_;
wire _158_;
wire _159_;
wire _160_;
wire _161_;
wire _162_;
wire _163_;
wire _164_;
wire _165_;
wire \add_32ns_32ns_32_2_1_U13.ce ;
wire \add_32ns_32ns_32_2_1_U13.clk ;
wire [31:0] \add_32ns_32ns_32_2_1_U13.din0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U13.din1 ;
wire [31:0] \add_32ns_32ns_32_2_1_U13.dout ;
wire \add_32ns_32ns_32_2_1_U13.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_4_U.a ;
wire [31:0] \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_4_U.ain_s0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_4_U.b ;
wire [31:0] \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_4_U.bin_s0 ;
wire \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_4_U.ce ;
wire \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_4_U.clk ;
wire \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_4_U.facout_s1 ;
wire \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_4_U.facout_s2 ;
wire [15:0] \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_4_U.fas_s1 ;
wire [15:0] \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_4_U.fas_s2 ;
wire \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_4_U.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_4_U.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.b ;
wire \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.cin ;
wire \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.b ;
wire \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.cin ;
wire \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.s ;
wire \add_32ns_32ns_32_2_1_U14.ce ;
wire \add_32ns_32ns_32_2_1_U14.clk ;
wire [31:0] \add_32ns_32ns_32_2_1_U14.din0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U14.din1 ;
wire [31:0] \add_32ns_32ns_32_2_1_U14.dout ;
wire \add_32ns_32ns_32_2_1_U14.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_4_U.a ;
wire [31:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_4_U.ain_s0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_4_U.b ;
wire [31:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_4_U.bin_s0 ;
wire \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_4_U.ce ;
wire \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_4_U.clk ;
wire \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_4_U.facout_s1 ;
wire \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_4_U.facout_s2 ;
wire [15:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_4_U.fas_s1 ;
wire [15:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_4_U.fas_s2 ;
wire \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_4_U.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_4_U.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.b ;
wire \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.cin ;
wire \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.b ;
wire \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.cin ;
wire \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.s ;
wire \add_32ns_32ns_32_2_1_U18.ce ;
wire \add_32ns_32ns_32_2_1_U18.clk ;
wire [31:0] \add_32ns_32ns_32_2_1_U18.din0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U18.din1 ;
wire [31:0] \add_32ns_32ns_32_2_1_U18.dout ;
wire \add_32ns_32ns_32_2_1_U18.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_4_U.a ;
wire [31:0] \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_4_U.ain_s0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_4_U.b ;
wire [31:0] \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_4_U.bin_s0 ;
wire \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_4_U.ce ;
wire \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_4_U.clk ;
wire \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_4_U.facout_s1 ;
wire \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_4_U.facout_s2 ;
wire [15:0] \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_4_U.fas_s1 ;
wire [15:0] \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_4_U.fas_s2 ;
wire \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_4_U.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_4_U.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.b ;
wire \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.cin ;
wire \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.b ;
wire \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.cin ;
wire \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.s ;
wire \add_32ns_32ns_32_2_1_U5.ce ;
wire \add_32ns_32ns_32_2_1_U5.clk ;
wire [31:0] \add_32ns_32ns_32_2_1_U5.din0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U5.din1 ;
wire [31:0] \add_32ns_32ns_32_2_1_U5.dout ;
wire \add_32ns_32ns_32_2_1_U5.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.a ;
wire [31:0] \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.ain_s0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.b ;
wire [31:0] \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.bin_s0 ;
wire \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.ce ;
wire \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.clk ;
wire \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.facout_s1 ;
wire \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.facout_s2 ;
wire [15:0] \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.fas_s1 ;
wire [15:0] \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.fas_s2 ;
wire \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.b ;
wire \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.cin ;
wire \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.b ;
wire \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.cin ;
wire \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.s ;
wire \add_32ns_32ns_32_2_1_U7.ce ;
wire \add_32ns_32ns_32_2_1_U7.clk ;
wire [31:0] \add_32ns_32ns_32_2_1_U7.din0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U7.din1 ;
wire [31:0] \add_32ns_32ns_32_2_1_U7.dout ;
wire \add_32ns_32ns_32_2_1_U7.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_4_U.a ;
wire [31:0] \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_4_U.ain_s0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_4_U.b ;
wire [31:0] \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_4_U.bin_s0 ;
wire \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_4_U.ce ;
wire \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_4_U.clk ;
wire \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_4_U.facout_s1 ;
wire \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_4_U.facout_s2 ;
wire [15:0] \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_4_U.fas_s1 ;
wire [15:0] \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_4_U.fas_s2 ;
wire \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_4_U.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_4_U.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.b ;
wire \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.cin ;
wire \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.b ;
wire \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.cin ;
wire \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.s ;
wire \add_32ns_32ns_32_2_1_U8.ce ;
wire \add_32ns_32ns_32_2_1_U8.clk ;
wire [31:0] \add_32ns_32ns_32_2_1_U8.din0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U8.din1 ;
wire [31:0] \add_32ns_32ns_32_2_1_U8.dout ;
wire \add_32ns_32ns_32_2_1_U8.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.a ;
wire [31:0] \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.ain_s0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.b ;
wire [31:0] \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.bin_s0 ;
wire \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.ce ;
wire \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.clk ;
wire \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.facout_s1 ;
wire \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.facout_s2 ;
wire [15:0] \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.fas_s1 ;
wire [15:0] \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.fas_s2 ;
wire \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.b ;
wire \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.cin ;
wire \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.b ;
wire \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.cin ;
wire \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.s ;
wire \add_32ns_32s_32_2_1_U11.ce ;
wire \add_32ns_32s_32_2_1_U11.clk ;
wire [31:0] \add_32ns_32s_32_2_1_U11.din0 ;
wire [31:0] \add_32ns_32s_32_2_1_U11.din1 ;
wire [31:0] \add_32ns_32s_32_2_1_U11.dout ;
wire \add_32ns_32s_32_2_1_U11.reset ;
wire [31:0] \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.a ;
wire [31:0] \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.ain_s0 ;
wire [31:0] \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.b ;
wire [31:0] \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.bin_s0 ;
wire \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.ce ;
wire \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.clk ;
wire \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.facout_s1 ;
wire \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.facout_s2 ;
wire [15:0] \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.fas_s1 ;
wire [15:0] \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.fas_s2 ;
wire \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.reset ;
wire [31:0] \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.s ;
wire [15:0] \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.u1.a ;
wire [15:0] \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.u1.b ;
wire \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.u1.cin ;
wire \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.u1.cout ;
wire [15:0] \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.u1.s ;
wire [15:0] \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.u2.a ;
wire [15:0] \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.u2.b ;
wire \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.u2.cin ;
wire \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.u2.cout ;
wire [15:0] \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.u2.s ;
wire \add_32ns_32s_32_2_1_U19.ce ;
wire \add_32ns_32s_32_2_1_U19.clk ;
wire [31:0] \add_32ns_32s_32_2_1_U19.din0 ;
wire [31:0] \add_32ns_32s_32_2_1_U19.din1 ;
wire [31:0] \add_32ns_32s_32_2_1_U19.dout ;
wire \add_32ns_32s_32_2_1_U19.reset ;
wire [31:0] \add_32ns_32s_32_2_1_U19.top_add_32ns_32s_32_2_1_Adder_8_U.a ;
wire [31:0] \add_32ns_32s_32_2_1_U19.top_add_32ns_32s_32_2_1_Adder_8_U.ain_s0 ;
wire [31:0] \add_32ns_32s_32_2_1_U19.top_add_32ns_32s_32_2_1_Adder_8_U.b ;
wire [31:0] \add_32ns_32s_32_2_1_U19.top_add_32ns_32s_32_2_1_Adder_8_U.bin_s0 ;
wire \add_32ns_32s_32_2_1_U19.top_add_32ns_32s_32_2_1_Adder_8_U.ce ;
wire \add_32ns_32s_32_2_1_U19.top_add_32ns_32s_32_2_1_Adder_8_U.clk ;
wire \add_32ns_32s_32_2_1_U19.top_add_32ns_32s_32_2_1_Adder_8_U.facout_s1 ;
wire \add_32ns_32s_32_2_1_U19.top_add_32ns_32s_32_2_1_Adder_8_U.facout_s2 ;
wire [15:0] \add_32ns_32s_32_2_1_U19.top_add_32ns_32s_32_2_1_Adder_8_U.fas_s1 ;
wire [15:0] \add_32ns_32s_32_2_1_U19.top_add_32ns_32s_32_2_1_Adder_8_U.fas_s2 ;
wire \add_32ns_32s_32_2_1_U19.top_add_32ns_32s_32_2_1_Adder_8_U.reset ;
wire [31:0] \add_32ns_32s_32_2_1_U19.top_add_32ns_32s_32_2_1_Adder_8_U.s ;
wire [15:0] \add_32ns_32s_32_2_1_U19.top_add_32ns_32s_32_2_1_Adder_8_U.u1.a ;
wire [15:0] \add_32ns_32s_32_2_1_U19.top_add_32ns_32s_32_2_1_Adder_8_U.u1.b ;
wire \add_32ns_32s_32_2_1_U19.top_add_32ns_32s_32_2_1_Adder_8_U.u1.cin ;
wire \add_32ns_32s_32_2_1_U19.top_add_32ns_32s_32_2_1_Adder_8_U.u1.cout ;
wire [15:0] \add_32ns_32s_32_2_1_U19.top_add_32ns_32s_32_2_1_Adder_8_U.u1.s ;
wire [15:0] \add_32ns_32s_32_2_1_U19.top_add_32ns_32s_32_2_1_Adder_8_U.u2.a ;
wire [15:0] \add_32ns_32s_32_2_1_U19.top_add_32ns_32s_32_2_1_Adder_8_U.u2.b ;
wire \add_32ns_32s_32_2_1_U19.top_add_32ns_32s_32_2_1_Adder_8_U.u2.cin ;
wire \add_32ns_32s_32_2_1_U19.top_add_32ns_32s_32_2_1_Adder_8_U.u2.cout ;
wire [15:0] \add_32ns_32s_32_2_1_U19.top_add_32ns_32s_32_2_1_Adder_8_U.u2.s ;
wire \add_32s_32ns_32_2_1_U10.ce ;
wire \add_32s_32ns_32_2_1_U10.clk ;
wire [31:0] \add_32s_32ns_32_2_1_U10.din0 ;
wire [31:0] \add_32s_32ns_32_2_1_U10.din1 ;
wire [31:0] \add_32s_32ns_32_2_1_U10.dout ;
wire \add_32s_32ns_32_2_1_U10.reset ;
wire [31:0] \add_32s_32ns_32_2_1_U10.top_add_32s_32ns_32_2_1_Adder_7_U.a ;
wire [31:0] \add_32s_32ns_32_2_1_U10.top_add_32s_32ns_32_2_1_Adder_7_U.ain_s0 ;
wire [31:0] \add_32s_32ns_32_2_1_U10.top_add_32s_32ns_32_2_1_Adder_7_U.b ;
wire [31:0] \add_32s_32ns_32_2_1_U10.top_add_32s_32ns_32_2_1_Adder_7_U.bin_s0 ;
wire \add_32s_32ns_32_2_1_U10.top_add_32s_32ns_32_2_1_Adder_7_U.ce ;
wire \add_32s_32ns_32_2_1_U10.top_add_32s_32ns_32_2_1_Adder_7_U.clk ;
wire \add_32s_32ns_32_2_1_U10.top_add_32s_32ns_32_2_1_Adder_7_U.facout_s1 ;
wire \add_32s_32ns_32_2_1_U10.top_add_32s_32ns_32_2_1_Adder_7_U.facout_s2 ;
wire [15:0] \add_32s_32ns_32_2_1_U10.top_add_32s_32ns_32_2_1_Adder_7_U.fas_s1 ;
wire [15:0] \add_32s_32ns_32_2_1_U10.top_add_32s_32ns_32_2_1_Adder_7_U.fas_s2 ;
wire \add_32s_32ns_32_2_1_U10.top_add_32s_32ns_32_2_1_Adder_7_U.reset ;
wire [31:0] \add_32s_32ns_32_2_1_U10.top_add_32s_32ns_32_2_1_Adder_7_U.s ;
wire [15:0] \add_32s_32ns_32_2_1_U10.top_add_32s_32ns_32_2_1_Adder_7_U.u1.a ;
wire [15:0] \add_32s_32ns_32_2_1_U10.top_add_32s_32ns_32_2_1_Adder_7_U.u1.b ;
wire \add_32s_32ns_32_2_1_U10.top_add_32s_32ns_32_2_1_Adder_7_U.u1.cin ;
wire \add_32s_32ns_32_2_1_U10.top_add_32s_32ns_32_2_1_Adder_7_U.u1.cout ;
wire [15:0] \add_32s_32ns_32_2_1_U10.top_add_32s_32ns_32_2_1_Adder_7_U.u1.s ;
wire [15:0] \add_32s_32ns_32_2_1_U10.top_add_32s_32ns_32_2_1_Adder_7_U.u2.a ;
wire [15:0] \add_32s_32ns_32_2_1_U10.top_add_32s_32ns_32_2_1_Adder_7_U.u2.b ;
wire \add_32s_32ns_32_2_1_U10.top_add_32s_32ns_32_2_1_Adder_7_U.u2.cin ;
wire \add_32s_32ns_32_2_1_U10.top_add_32s_32ns_32_2_1_Adder_7_U.u2.cout ;
wire [15:0] \add_32s_32ns_32_2_1_U10.top_add_32s_32ns_32_2_1_Adder_7_U.u2.s ;
wire \add_32s_32ns_32_2_1_U16.ce ;
wire \add_32s_32ns_32_2_1_U16.clk ;
wire [31:0] \add_32s_32ns_32_2_1_U16.din0 ;
wire [31:0] \add_32s_32ns_32_2_1_U16.din1 ;
wire [31:0] \add_32s_32ns_32_2_1_U16.dout ;
wire \add_32s_32ns_32_2_1_U16.reset ;
wire [31:0] \add_32s_32ns_32_2_1_U16.top_add_32s_32ns_32_2_1_Adder_7_U.a ;
wire [31:0] \add_32s_32ns_32_2_1_U16.top_add_32s_32ns_32_2_1_Adder_7_U.ain_s0 ;
wire [31:0] \add_32s_32ns_32_2_1_U16.top_add_32s_32ns_32_2_1_Adder_7_U.b ;
wire [31:0] \add_32s_32ns_32_2_1_U16.top_add_32s_32ns_32_2_1_Adder_7_U.bin_s0 ;
wire \add_32s_32ns_32_2_1_U16.top_add_32s_32ns_32_2_1_Adder_7_U.ce ;
wire \add_32s_32ns_32_2_1_U16.top_add_32s_32ns_32_2_1_Adder_7_U.clk ;
wire \add_32s_32ns_32_2_1_U16.top_add_32s_32ns_32_2_1_Adder_7_U.facout_s1 ;
wire \add_32s_32ns_32_2_1_U16.top_add_32s_32ns_32_2_1_Adder_7_U.facout_s2 ;
wire [15:0] \add_32s_32ns_32_2_1_U16.top_add_32s_32ns_32_2_1_Adder_7_U.fas_s1 ;
wire [15:0] \add_32s_32ns_32_2_1_U16.top_add_32s_32ns_32_2_1_Adder_7_U.fas_s2 ;
wire \add_32s_32ns_32_2_1_U16.top_add_32s_32ns_32_2_1_Adder_7_U.reset ;
wire [31:0] \add_32s_32ns_32_2_1_U16.top_add_32s_32ns_32_2_1_Adder_7_U.s ;
wire [15:0] \add_32s_32ns_32_2_1_U16.top_add_32s_32ns_32_2_1_Adder_7_U.u1.a ;
wire [15:0] \add_32s_32ns_32_2_1_U16.top_add_32s_32ns_32_2_1_Adder_7_U.u1.b ;
wire \add_32s_32ns_32_2_1_U16.top_add_32s_32ns_32_2_1_Adder_7_U.u1.cin ;
wire \add_32s_32ns_32_2_1_U16.top_add_32s_32ns_32_2_1_Adder_7_U.u1.cout ;
wire [15:0] \add_32s_32ns_32_2_1_U16.top_add_32s_32ns_32_2_1_Adder_7_U.u1.s ;
wire [15:0] \add_32s_32ns_32_2_1_U16.top_add_32s_32ns_32_2_1_Adder_7_U.u2.a ;
wire [15:0] \add_32s_32ns_32_2_1_U16.top_add_32s_32ns_32_2_1_Adder_7_U.u2.b ;
wire \add_32s_32ns_32_2_1_U16.top_add_32s_32ns_32_2_1_Adder_7_U.u2.cin ;
wire \add_32s_32ns_32_2_1_U16.top_add_32s_32ns_32_2_1_Adder_7_U.u2.cout ;
wire [15:0] \add_32s_32ns_32_2_1_U16.top_add_32s_32ns_32_2_1_Adder_7_U.u2.s ;
wire \add_34s_34ns_34_2_1_U4.ce ;
wire \add_34s_34ns_34_2_1_U4.clk ;
wire [33:0] \add_34s_34ns_34_2_1_U4.din0 ;
wire [33:0] \add_34s_34ns_34_2_1_U4.din1 ;
wire [33:0] \add_34s_34ns_34_2_1_U4.dout ;
wire \add_34s_34ns_34_2_1_U4.reset ;
wire [33:0] \add_34s_34ns_34_2_1_U4.top_add_34s_34ns_34_2_1_Adder_3_U.a ;
wire [33:0] \add_34s_34ns_34_2_1_U4.top_add_34s_34ns_34_2_1_Adder_3_U.ain_s0 ;
wire [33:0] \add_34s_34ns_34_2_1_U4.top_add_34s_34ns_34_2_1_Adder_3_U.b ;
wire [33:0] \add_34s_34ns_34_2_1_U4.top_add_34s_34ns_34_2_1_Adder_3_U.bin_s0 ;
wire \add_34s_34ns_34_2_1_U4.top_add_34s_34ns_34_2_1_Adder_3_U.ce ;
wire \add_34s_34ns_34_2_1_U4.top_add_34s_34ns_34_2_1_Adder_3_U.clk ;
wire \add_34s_34ns_34_2_1_U4.top_add_34s_34ns_34_2_1_Adder_3_U.facout_s1 ;
wire \add_34s_34ns_34_2_1_U4.top_add_34s_34ns_34_2_1_Adder_3_U.facout_s2 ;
wire [16:0] \add_34s_34ns_34_2_1_U4.top_add_34s_34ns_34_2_1_Adder_3_U.fas_s1 ;
wire [16:0] \add_34s_34ns_34_2_1_U4.top_add_34s_34ns_34_2_1_Adder_3_U.fas_s2 ;
wire \add_34s_34ns_34_2_1_U4.top_add_34s_34ns_34_2_1_Adder_3_U.reset ;
wire [33:0] \add_34s_34ns_34_2_1_U4.top_add_34s_34ns_34_2_1_Adder_3_U.s ;
wire [16:0] \add_34s_34ns_34_2_1_U4.top_add_34s_34ns_34_2_1_Adder_3_U.u1.a ;
wire [16:0] \add_34s_34ns_34_2_1_U4.top_add_34s_34ns_34_2_1_Adder_3_U.u1.b ;
wire \add_34s_34ns_34_2_1_U4.top_add_34s_34ns_34_2_1_Adder_3_U.u1.cin ;
wire \add_34s_34ns_34_2_1_U4.top_add_34s_34ns_34_2_1_Adder_3_U.u1.cout ;
wire [16:0] \add_34s_34ns_34_2_1_U4.top_add_34s_34ns_34_2_1_Adder_3_U.u1.s ;
wire [16:0] \add_34s_34ns_34_2_1_U4.top_add_34s_34ns_34_2_1_Adder_3_U.u2.a ;
wire [16:0] \add_34s_34ns_34_2_1_U4.top_add_34s_34ns_34_2_1_Adder_3_U.u2.b ;
wire \add_34s_34ns_34_2_1_U4.top_add_34s_34ns_34_2_1_Adder_3_U.u2.cin ;
wire \add_34s_34ns_34_2_1_U4.top_add_34s_34ns_34_2_1_Adder_3_U.u2.cout ;
wire [16:0] \add_34s_34ns_34_2_1_U4.top_add_34s_34ns_34_2_1_Adder_3_U.u2.s ;
wire \add_34s_34s_34_2_1_U17.ce ;
wire \add_34s_34s_34_2_1_U17.clk ;
wire [33:0] \add_34s_34s_34_2_1_U17.din0 ;
wire [33:0] \add_34s_34s_34_2_1_U17.din1 ;
wire [33:0] \add_34s_34s_34_2_1_U17.dout ;
wire \add_34s_34s_34_2_1_U17.reset ;
wire [33:0] \add_34s_34s_34_2_1_U17.top_add_34s_34s_34_2_1_Adder_5_U.a ;
wire [33:0] \add_34s_34s_34_2_1_U17.top_add_34s_34s_34_2_1_Adder_5_U.ain_s0 ;
wire [33:0] \add_34s_34s_34_2_1_U17.top_add_34s_34s_34_2_1_Adder_5_U.b ;
wire [33:0] \add_34s_34s_34_2_1_U17.top_add_34s_34s_34_2_1_Adder_5_U.bin_s0 ;
wire \add_34s_34s_34_2_1_U17.top_add_34s_34s_34_2_1_Adder_5_U.ce ;
wire \add_34s_34s_34_2_1_U17.top_add_34s_34s_34_2_1_Adder_5_U.clk ;
wire \add_34s_34s_34_2_1_U17.top_add_34s_34s_34_2_1_Adder_5_U.facout_s1 ;
wire \add_34s_34s_34_2_1_U17.top_add_34s_34s_34_2_1_Adder_5_U.facout_s2 ;
wire [16:0] \add_34s_34s_34_2_1_U17.top_add_34s_34s_34_2_1_Adder_5_U.fas_s1 ;
wire [16:0] \add_34s_34s_34_2_1_U17.top_add_34s_34s_34_2_1_Adder_5_U.fas_s2 ;
wire \add_34s_34s_34_2_1_U17.top_add_34s_34s_34_2_1_Adder_5_U.reset ;
wire [33:0] \add_34s_34s_34_2_1_U17.top_add_34s_34s_34_2_1_Adder_5_U.s ;
wire [16:0] \add_34s_34s_34_2_1_U17.top_add_34s_34s_34_2_1_Adder_5_U.u1.a ;
wire [16:0] \add_34s_34s_34_2_1_U17.top_add_34s_34s_34_2_1_Adder_5_U.u1.b ;
wire \add_34s_34s_34_2_1_U17.top_add_34s_34s_34_2_1_Adder_5_U.u1.cin ;
wire \add_34s_34s_34_2_1_U17.top_add_34s_34s_34_2_1_Adder_5_U.u1.cout ;
wire [16:0] \add_34s_34s_34_2_1_U17.top_add_34s_34s_34_2_1_Adder_5_U.u1.s ;
wire [16:0] \add_34s_34s_34_2_1_U17.top_add_34s_34s_34_2_1_Adder_5_U.u2.a ;
wire [16:0] \add_34s_34s_34_2_1_U17.top_add_34s_34s_34_2_1_Adder_5_U.u2.b ;
wire \add_34s_34s_34_2_1_U17.top_add_34s_34s_34_2_1_Adder_5_U.u2.cin ;
wire \add_34s_34s_34_2_1_U17.top_add_34s_34s_34_2_1_Adder_5_U.u2.cout ;
wire [16:0] \add_34s_34s_34_2_1_U17.top_add_34s_34s_34_2_1_Adder_5_U.u2.s ;
wire \add_34s_34s_34_2_1_U6.ce ;
wire \add_34s_34s_34_2_1_U6.clk ;
wire [33:0] \add_34s_34s_34_2_1_U6.din0 ;
wire [33:0] \add_34s_34s_34_2_1_U6.din1 ;
wire [33:0] \add_34s_34s_34_2_1_U6.dout ;
wire \add_34s_34s_34_2_1_U6.reset ;
wire [33:0] \add_34s_34s_34_2_1_U6.top_add_34s_34s_34_2_1_Adder_5_U.a ;
wire [33:0] \add_34s_34s_34_2_1_U6.top_add_34s_34s_34_2_1_Adder_5_U.ain_s0 ;
wire [33:0] \add_34s_34s_34_2_1_U6.top_add_34s_34s_34_2_1_Adder_5_U.b ;
wire [33:0] \add_34s_34s_34_2_1_U6.top_add_34s_34s_34_2_1_Adder_5_U.bin_s0 ;
wire \add_34s_34s_34_2_1_U6.top_add_34s_34s_34_2_1_Adder_5_U.ce ;
wire \add_34s_34s_34_2_1_U6.top_add_34s_34s_34_2_1_Adder_5_U.clk ;
wire \add_34s_34s_34_2_1_U6.top_add_34s_34s_34_2_1_Adder_5_U.facout_s1 ;
wire \add_34s_34s_34_2_1_U6.top_add_34s_34s_34_2_1_Adder_5_U.facout_s2 ;
wire [16:0] \add_34s_34s_34_2_1_U6.top_add_34s_34s_34_2_1_Adder_5_U.fas_s1 ;
wire [16:0] \add_34s_34s_34_2_1_U6.top_add_34s_34s_34_2_1_Adder_5_U.fas_s2 ;
wire \add_34s_34s_34_2_1_U6.top_add_34s_34s_34_2_1_Adder_5_U.reset ;
wire [33:0] \add_34s_34s_34_2_1_U6.top_add_34s_34s_34_2_1_Adder_5_U.s ;
wire [16:0] \add_34s_34s_34_2_1_U6.top_add_34s_34s_34_2_1_Adder_5_U.u1.a ;
wire [16:0] \add_34s_34s_34_2_1_U6.top_add_34s_34s_34_2_1_Adder_5_U.u1.b ;
wire \add_34s_34s_34_2_1_U6.top_add_34s_34s_34_2_1_Adder_5_U.u1.cin ;
wire \add_34s_34s_34_2_1_U6.top_add_34s_34s_34_2_1_Adder_5_U.u1.cout ;
wire [16:0] \add_34s_34s_34_2_1_U6.top_add_34s_34s_34_2_1_Adder_5_U.u1.s ;
wire [16:0] \add_34s_34s_34_2_1_U6.top_add_34s_34s_34_2_1_Adder_5_U.u2.a ;
wire [16:0] \add_34s_34s_34_2_1_U6.top_add_34s_34s_34_2_1_Adder_5_U.u2.b ;
wire \add_34s_34s_34_2_1_U6.top_add_34s_34s_34_2_1_Adder_5_U.u2.cin ;
wire \add_34s_34s_34_2_1_U6.top_add_34s_34s_34_2_1_Adder_5_U.u2.cout ;
wire [16:0] \add_34s_34s_34_2_1_U6.top_add_34s_34s_34_2_1_Adder_5_U.u2.s ;
wire \add_47s_47s_47_2_1_U12.ce ;
wire \add_47s_47s_47_2_1_U12.clk ;
wire [46:0] \add_47s_47s_47_2_1_U12.din0 ;
wire [46:0] \add_47s_47s_47_2_1_U12.din1 ;
wire [46:0] \add_47s_47s_47_2_1_U12.dout ;
wire \add_47s_47s_47_2_1_U12.reset ;
wire [46:0] \add_47s_47s_47_2_1_U12.top_add_47s_47s_47_2_1_Adder_9_U.a ;
wire [46:0] \add_47s_47s_47_2_1_U12.top_add_47s_47s_47_2_1_Adder_9_U.ain_s0 ;
wire [46:0] \add_47s_47s_47_2_1_U12.top_add_47s_47s_47_2_1_Adder_9_U.b ;
wire [46:0] \add_47s_47s_47_2_1_U12.top_add_47s_47s_47_2_1_Adder_9_U.bin_s0 ;
wire \add_47s_47s_47_2_1_U12.top_add_47s_47s_47_2_1_Adder_9_U.ce ;
wire \add_47s_47s_47_2_1_U12.top_add_47s_47s_47_2_1_Adder_9_U.clk ;
wire \add_47s_47s_47_2_1_U12.top_add_47s_47s_47_2_1_Adder_9_U.facout_s1 ;
wire \add_47s_47s_47_2_1_U12.top_add_47s_47s_47_2_1_Adder_9_U.facout_s2 ;
wire [22:0] \add_47s_47s_47_2_1_U12.top_add_47s_47s_47_2_1_Adder_9_U.fas_s1 ;
wire [23:0] \add_47s_47s_47_2_1_U12.top_add_47s_47s_47_2_1_Adder_9_U.fas_s2 ;
wire \add_47s_47s_47_2_1_U12.top_add_47s_47s_47_2_1_Adder_9_U.reset ;
wire [46:0] \add_47s_47s_47_2_1_U12.top_add_47s_47s_47_2_1_Adder_9_U.s ;
wire [22:0] \add_47s_47s_47_2_1_U12.top_add_47s_47s_47_2_1_Adder_9_U.u1.a ;
wire [22:0] \add_47s_47s_47_2_1_U12.top_add_47s_47s_47_2_1_Adder_9_U.u1.b ;
wire \add_47s_47s_47_2_1_U12.top_add_47s_47s_47_2_1_Adder_9_U.u1.cin ;
wire \add_47s_47s_47_2_1_U12.top_add_47s_47s_47_2_1_Adder_9_U.u1.cout ;
wire [22:0] \add_47s_47s_47_2_1_U12.top_add_47s_47s_47_2_1_Adder_9_U.u1.s ;
wire [23:0] \add_47s_47s_47_2_1_U12.top_add_47s_47s_47_2_1_Adder_9_U.u2.a ;
wire [23:0] \add_47s_47s_47_2_1_U12.top_add_47s_47s_47_2_1_Adder_9_U.u2.b ;
wire \add_47s_47s_47_2_1_U12.top_add_47s_47s_47_2_1_Adder_9_U.u2.cin ;
wire \add_47s_47s_47_2_1_U12.top_add_47s_47s_47_2_1_Adder_9_U.u2.cout ;
wire [23:0] \add_47s_47s_47_2_1_U12.top_add_47s_47s_47_2_1_Adder_9_U.u2.s ;
wire [4:0] \add_5s_5ns_5_1_1_U15.din0 ;
wire [4:0] \add_5s_5ns_5_1_1_U15.din1 ;
wire [4:0] \add_5s_5ns_5_1_1_U15.dout ;
wire [4:0] \add_5s_5ns_5_1_1_U15.top_add_5s_5ns_5_1_1_Adder_10_U.a ;
wire [4:0] \add_5s_5ns_5_1_1_U15.top_add_5s_5ns_5_1_1_Adder_10_U.b ;
wire [4:0] \add_5s_5ns_5_1_1_U15.top_add_5s_5ns_5_1_1_Adder_10_U.s ;
wire [6:0] \add_7s_7ns_7_1_1_U1.din0 ;
wire [6:0] \add_7s_7ns_7_1_1_U1.din1 ;
wire [6:0] \add_7s_7ns_7_1_1_U1.dout ;
wire [6:0] \add_7s_7ns_7_1_1_U1.top_add_7s_7ns_7_1_1_Adder_0_U.a ;
wire [6:0] \add_7s_7ns_7_1_1_U1.top_add_7s_7ns_7_1_1_Adder_0_U.b ;
wire [6:0] \add_7s_7ns_7_1_1_U1.top_add_7s_7ns_7_1_1_Adder_0_U.s ;
wire [7:0] \add_8s_8ns_8_1_1_U3.din0 ;
wire [7:0] \add_8s_8ns_8_1_1_U3.din1 ;
wire [7:0] \add_8s_8ns_8_1_1_U3.dout ;
wire [7:0] \add_8s_8ns_8_1_1_U3.top_add_8s_8ns_8_1_1_Adder_2_U.a ;
wire [7:0] \add_8s_8ns_8_1_1_U3.top_add_8s_8ns_8_1_1_Adder_2_U.b ;
wire [7:0] \add_8s_8ns_8_1_1_U3.top_add_8s_8ns_8_1_1_Adder_2_U.s ;
wire [8:0] \add_9ns_9s_9_1_1_U2.din0 ;
wire [8:0] \add_9ns_9s_9_1_1_U2.din1 ;
wire [8:0] \add_9ns_9s_9_1_1_U2.dout ;
wire [8:0] \add_9ns_9s_9_1_1_U2.top_add_9ns_9s_9_1_1_Adder_1_U.a ;
wire [8:0] \add_9ns_9s_9_1_1_U2.top_add_9ns_9s_9_1_1_Adder_1_U.b ;
wire [8:0] \add_9ns_9s_9_1_1_U2.top_add_9ns_9s_9_1_1_Adder_1_U.s ;
wire [8:0] \add_9s_9ns_9_1_1_U9.din0 ;
wire [8:0] \add_9s_9ns_9_1_1_U9.din1 ;
wire [8:0] \add_9s_9ns_9_1_1_U9.dout ;
wire [8:0] \add_9s_9ns_9_1_1_U9.top_add_9s_9ns_9_1_1_Adder_6_U.a ;
wire [8:0] \add_9s_9ns_9_1_1_U9.top_add_9s_9ns_9_1_1_Adder_6_U.b ;
wire [8:0] \add_9s_9ns_9_1_1_U9.top_add_9s_9ns_9_1_1_Adder_6_U.s ;
wire [7:0] add_ln691_fu_315_p0;
wire [7:0] add_ln691_fu_315_p2;
wire [8:0] add_ln69_1_fu_474_p0;
wire [8:0] add_ln69_1_fu_474_p1;
wire [8:0] add_ln69_1_fu_474_p2;
wire [4:0] add_ln69_4_fu_607_p0;
wire [4:0] add_ln69_4_fu_607_p1;
wire [4:0] add_ln69_4_fu_607_p2;
wire ap_CS_fsm_state1;
wire ap_CS_fsm_state10;
wire ap_CS_fsm_state11;
wire ap_CS_fsm_state12;
wire ap_CS_fsm_state13;
wire ap_CS_fsm_state14;
wire ap_CS_fsm_state15;
wire ap_CS_fsm_state16;
wire ap_CS_fsm_state17;
wire ap_CS_fsm_state18;
wire ap_CS_fsm_state19;
wire ap_CS_fsm_state2;
wire ap_CS_fsm_state20;
wire ap_CS_fsm_state21;
wire ap_CS_fsm_state22;
wire ap_CS_fsm_state23;
wire ap_CS_fsm_state24;
wire ap_CS_fsm_state25;
wire ap_CS_fsm_state26;
wire ap_CS_fsm_state27;
wire ap_CS_fsm_state28;
wire ap_CS_fsm_state29;
wire ap_CS_fsm_state3;
wire ap_CS_fsm_state30;
wire ap_CS_fsm_state31;
wire ap_CS_fsm_state32;
wire ap_CS_fsm_state33;
wire ap_CS_fsm_state34;
wire ap_CS_fsm_state35;
wire ap_CS_fsm_state36;
wire ap_CS_fsm_state4;
wire ap_CS_fsm_state5;
wire ap_CS_fsm_state6;
wire ap_CS_fsm_state7;
wire ap_CS_fsm_state8;
wire ap_CS_fsm_state9;
wire [35:0] ap_NS_fsm;
wire ap_clk;
wire ap_done;
wire ap_idle;
wire ap_ready;
wire ap_rst;
wire ap_start;
wire [33:0] grp_fu_359_p0;
wire [33:0] grp_fu_359_p2;
wire [31:0] grp_fu_374_p2;
wire [33:0] grp_fu_413_p0;
wire [33:0] grp_fu_413_p1;
wire [33:0] grp_fu_413_p2;
wire [31:0] grp_fu_429_p2;
wire [31:0] grp_fu_461_p1;
wire [31:0] grp_fu_461_p2;
wire [31:0] grp_fu_483_p0;
wire [31:0] grp_fu_483_p2;
wire [31:0] grp_fu_492_p1;
wire [31:0] grp_fu_492_p2;
wire [46:0] grp_fu_541_p0;
wire [46:0] grp_fu_541_p1;
wire [46:0] grp_fu_541_p2;
wire [31:0] grp_fu_570_p2;
wire [31:0] grp_fu_594_p2;
wire [31:0] grp_fu_616_p0;
wire [31:0] grp_fu_616_p2;
wire [33:0] grp_fu_636_p0;
wire [33:0] grp_fu_636_p1;
wire [33:0] grp_fu_636_p2;
wire [31:0] grp_fu_652_p2;
wire [31:0] grp_fu_684_p1;
wire [31:0] grp_fu_684_p2;
wire icmp_ln851_1_fu_306_p2;
wire icmp_ln851_2_fu_554_p2;
wire icmp_ln851_fu_243_p2;
wire [7:0] op_0;
wire [7:0] op_10;
wire [3:0] op_11;
wire [15:0] op_12;
wire [1:0] op_13;
wire [18:0] op_14_V_fu_519_p3;
wire [1:0] op_15;
wire [31:0] op_16;
wire [3:0] op_17;
wire [7:0] op_18;
wire [7:0] op_19;
wire [7:0] op_3;
wire [31:0] op_33;
wire op_33_ap_vld;
wire op_4;
wire op_4_read_read_fu_140_p2;
wire [7:0] op_5;
wire [3:0] op_6;
wire [3:0] op_7;
wire [1:0] op_9;
wire p_Result_1_fu_321_p3;
wire p_Result_2_fu_379_p3;
wire p_Result_3_fu_434_p3;
wire p_Result_4_fu_575_p3;
wire p_Result_5_fu_657_p3;
wire [13:0] p_Result_7_fu_547_p3;
wire p_Result_s_fu_255_p3;
wire [8:0] ret_V_12_fu_286_p0;
wire [8:0] ret_V_12_fu_286_p1;
wire [8:0] ret_V_12_fu_286_p2;
wire [31:0] ret_V_15_fu_450_p3;
wire [31:0] ret_V_18_fu_587_p3;
wire [5:0] ret_V_1_fu_225_p4;
wire [31:0] ret_V_20_fu_673_p3;
wire [6:0] ret_V_2_fu_249_p0;
wire [6:0] ret_V_2_fu_249_p2;
wire [7:0] ret_V_fu_509_p2;
wire [32:0] rhs_2_fu_402_p3;
wire [45:0] rhs_5_fu_530_p3;
wire [32:0] rhs_7_fu_625_p3;
wire [6:0] rhs_fu_497_p3;
wire [31:0] select_ln353_1_fu_391_p3;
wire [7:0] select_ln353_fu_341_p3;
wire [33:0] select_ln703_fu_328_p3;
wire [6:0] select_ln850_1_fu_271_p3;
wire [7:0] select_ln850_2_fu_336_p3;
wire [31:0] select_ln850_3_fu_444_p3;
wire [31:0] select_ln850_4_fu_582_p3;
wire [31:0] select_ln850_5_fu_667_p3;
wire [31:0] select_ln850_6_fu_386_p3;
wire [6:0] select_ln850_fu_266_p3;
wire [3:0] sext_ln1192_fu_262_p0;
wire [7:0] sext_ln1194_fu_505_p1;
wire [7:0] sext_ln703_2_fu_621_p0;
wire [1:0] sext_ln703_fu_398_p0;
wire [6:0] sext_ln835_fu_235_p1;
wire [7:0] sext_ln850_fu_312_p1;
wire [8:0] tmp_3_fu_348_p3;
wire [3:0] trunc_ln851_1_fu_302_p0;
wire [1:0] trunc_ln851_1_fu_302_p1;
wire [1:0] trunc_ln851_2_fu_441_p0;
wire trunc_ln851_2_fu_441_p1;
wire [2:0] trunc_ln851_3_fu_515_p1;
wire [7:0] trunc_ln851_4_fu_664_p0;
wire trunc_ln851_4_fu_664_p1;
wire [1:0] trunc_ln851_fu_239_p1;


assign _037_ = ap_CS_fsm[7] & op_4;
assign _038_ = icmp_ln851_2_reg_871 & ap_CS_fsm[23];
assign _039_ = icmp_ln851_1_reg_721 & ap_CS_fsm[2];
assign _040_ = _042_ & ap_CS_fsm[0];
assign _041_ = ap_start & ap_CS_fsm[0];
assign ret_V_fu_509_p2 = { op_6[3], op_6, 3'h0 } & op_3;
assign _042_ = ~ ap_start;
assign _043_ = ! op_5[1:0];
always @(posedge \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_4_U.clk )
\add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_4_U.bin_s1  <= _045_;
always @(posedge \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_4_U.clk )
\add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_4_U.ain_s1  <= _044_;
always @(posedge \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_4_U.clk )
\add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_4_U.sum_s1  <= _047_;
always @(posedge \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_4_U.clk )
\add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_4_U.carry_s1  <= _046_;
assign _045_ = \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_4_U.ce  ? \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_4_U.b [31:16] : \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_4_U.bin_s1 ;
assign _044_ = \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_4_U.ce  ? \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_4_U.a [31:16] : \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_4_U.ain_s1 ;
assign _046_ = \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_4_U.ce  ? \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_4_U.facout_s1  : \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_4_U.carry_s1 ;
assign _047_ = \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_4_U.ce  ? \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_4_U.fas_s1  : \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_4_U.sum_s1 ;
assign _048_ = \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.a  + \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.b ;
assign { \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.cout , \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.s  } = _048_ + \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.cin ;
assign _049_ = \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.a  + \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.b ;
assign { \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.cout , \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.s  } = _049_ + \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.cin ;
always @(posedge \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_4_U.clk )
\add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_4_U.bin_s1  <= _051_;
always @(posedge \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_4_U.clk )
\add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_4_U.ain_s1  <= _050_;
always @(posedge \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_4_U.clk )
\add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_4_U.sum_s1  <= _053_;
always @(posedge \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_4_U.clk )
\add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_4_U.carry_s1  <= _052_;
assign _051_ = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_4_U.ce  ? \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_4_U.b [31:16] : \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_4_U.bin_s1 ;
assign _050_ = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_4_U.ce  ? \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_4_U.a [31:16] : \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_4_U.ain_s1 ;
assign _052_ = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_4_U.ce  ? \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_4_U.facout_s1  : \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_4_U.carry_s1 ;
assign _053_ = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_4_U.ce  ? \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_4_U.fas_s1  : \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_4_U.sum_s1 ;
assign _054_ = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.a  + \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.b ;
assign { \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.cout , \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.s  } = _054_ + \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.cin ;
assign _055_ = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.a  + \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.b ;
assign { \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.cout , \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.s  } = _055_ + \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.cin ;
always @(posedge \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_4_U.clk )
\add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_4_U.bin_s1  <= _057_;
always @(posedge \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_4_U.clk )
\add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_4_U.ain_s1  <= _056_;
always @(posedge \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_4_U.clk )
\add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_4_U.sum_s1  <= _059_;
always @(posedge \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_4_U.clk )
\add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_4_U.carry_s1  <= _058_;
assign _057_ = \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_4_U.ce  ? \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_4_U.b [31:16] : \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_4_U.bin_s1 ;
assign _056_ = \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_4_U.ce  ? \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_4_U.a [31:16] : \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_4_U.ain_s1 ;
assign _058_ = \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_4_U.ce  ? \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_4_U.facout_s1  : \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_4_U.carry_s1 ;
assign _059_ = \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_4_U.ce  ? \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_4_U.fas_s1  : \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_4_U.sum_s1 ;
assign _060_ = \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.a  + \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.b ;
assign { \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.cout , \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.s  } = _060_ + \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.cin ;
assign _061_ = \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.a  + \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.b ;
assign { \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.cout , \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.s  } = _061_ + \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.cin ;
always @(posedge \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.clk )
\add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.bin_s1  <= _063_;
always @(posedge \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.clk )
\add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.ain_s1  <= _062_;
always @(posedge \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.clk )
\add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.sum_s1  <= _065_;
always @(posedge \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.clk )
\add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.carry_s1  <= _064_;
assign _063_ = \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.ce  ? \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.b [31:16] : \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.bin_s1 ;
assign _062_ = \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.ce  ? \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.a [31:16] : \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.ain_s1 ;
assign _064_ = \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.ce  ? \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.facout_s1  : \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.carry_s1 ;
assign _065_ = \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.ce  ? \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.fas_s1  : \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.sum_s1 ;
assign _066_ = \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.a  + \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.b ;
assign { \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.cout , \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.s  } = _066_ + \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.cin ;
assign _067_ = \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.a  + \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.b ;
assign { \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.cout , \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.s  } = _067_ + \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.cin ;
always @(posedge \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_4_U.clk )
\add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_4_U.bin_s1  <= _069_;
always @(posedge \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_4_U.clk )
\add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_4_U.ain_s1  <= _068_;
always @(posedge \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_4_U.clk )
\add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_4_U.sum_s1  <= _071_;
always @(posedge \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_4_U.clk )
\add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_4_U.carry_s1  <= _070_;
assign _069_ = \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_4_U.ce  ? \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_4_U.b [31:16] : \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_4_U.bin_s1 ;
assign _068_ = \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_4_U.ce  ? \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_4_U.a [31:16] : \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_4_U.ain_s1 ;
assign _070_ = \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_4_U.ce  ? \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_4_U.facout_s1  : \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_4_U.carry_s1 ;
assign _071_ = \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_4_U.ce  ? \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_4_U.fas_s1  : \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_4_U.sum_s1 ;
assign _072_ = \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.a  + \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.b ;
assign { \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.cout , \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.s  } = _072_ + \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.cin ;
assign _073_ = \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.a  + \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.b ;
assign { \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.cout , \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.s  } = _073_ + \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.cin ;
always @(posedge \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.clk )
\add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.bin_s1  <= _075_;
always @(posedge \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.clk )
\add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.ain_s1  <= _074_;
always @(posedge \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.clk )
\add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.sum_s1  <= _077_;
always @(posedge \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.clk )
\add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.carry_s1  <= _076_;
assign _075_ = \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.ce  ? \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.b [31:16] : \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.bin_s1 ;
assign _074_ = \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.ce  ? \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.a [31:16] : \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.ain_s1 ;
assign _076_ = \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.ce  ? \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.facout_s1  : \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.carry_s1 ;
assign _077_ = \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.ce  ? \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.fas_s1  : \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.sum_s1 ;
assign _078_ = \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.a  + \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.b ;
assign { \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.cout , \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.s  } = _078_ + \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.cin ;
assign _079_ = \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.a  + \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.b ;
assign { \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.cout , \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.s  } = _079_ + \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.cin ;
always @(posedge \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.clk )
\add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.bin_s1  <= _081_;
always @(posedge \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.clk )
\add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.ain_s1  <= _080_;
always @(posedge \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.clk )
\add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.sum_s1  <= _083_;
always @(posedge \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.clk )
\add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.carry_s1  <= _082_;
assign _081_ = \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.ce  ? \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.b [31:16] : \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.bin_s1 ;
assign _080_ = \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.ce  ? \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.a [31:16] : \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.ain_s1 ;
assign _082_ = \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.ce  ? \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.facout_s1  : \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.carry_s1 ;
assign _083_ = \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.ce  ? \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.fas_s1  : \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.sum_s1 ;
assign _084_ = \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.u1.a  + \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.u1.b ;
assign { \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.u1.cout , \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.u1.s  } = _084_ + \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.u1.cin ;
assign _085_ = \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.u2.a  + \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.u2.b ;
assign { \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.u2.cout , \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.u2.s  } = _085_ + \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.u2.cin ;
always @(posedge \add_32ns_32s_32_2_1_U19.top_add_32ns_32s_32_2_1_Adder_8_U.clk )
\add_32ns_32s_32_2_1_U19.top_add_32ns_32s_32_2_1_Adder_8_U.bin_s1  <= _087_;
always @(posedge \add_32ns_32s_32_2_1_U19.top_add_32ns_32s_32_2_1_Adder_8_U.clk )
\add_32ns_32s_32_2_1_U19.top_add_32ns_32s_32_2_1_Adder_8_U.ain_s1  <= _086_;
always @(posedge \add_32ns_32s_32_2_1_U19.top_add_32ns_32s_32_2_1_Adder_8_U.clk )
\add_32ns_32s_32_2_1_U19.top_add_32ns_32s_32_2_1_Adder_8_U.sum_s1  <= _089_;
always @(posedge \add_32ns_32s_32_2_1_U19.top_add_32ns_32s_32_2_1_Adder_8_U.clk )
\add_32ns_32s_32_2_1_U19.top_add_32ns_32s_32_2_1_Adder_8_U.carry_s1  <= _088_;
assign _087_ = \add_32ns_32s_32_2_1_U19.top_add_32ns_32s_32_2_1_Adder_8_U.ce  ? \add_32ns_32s_32_2_1_U19.top_add_32ns_32s_32_2_1_Adder_8_U.b [31:16] : \add_32ns_32s_32_2_1_U19.top_add_32ns_32s_32_2_1_Adder_8_U.bin_s1 ;
assign _086_ = \add_32ns_32s_32_2_1_U19.top_add_32ns_32s_32_2_1_Adder_8_U.ce  ? \add_32ns_32s_32_2_1_U19.top_add_32ns_32s_32_2_1_Adder_8_U.a [31:16] : \add_32ns_32s_32_2_1_U19.top_add_32ns_32s_32_2_1_Adder_8_U.ain_s1 ;
assign _088_ = \add_32ns_32s_32_2_1_U19.top_add_32ns_32s_32_2_1_Adder_8_U.ce  ? \add_32ns_32s_32_2_1_U19.top_add_32ns_32s_32_2_1_Adder_8_U.facout_s1  : \add_32ns_32s_32_2_1_U19.top_add_32ns_32s_32_2_1_Adder_8_U.carry_s1 ;
assign _089_ = \add_32ns_32s_32_2_1_U19.top_add_32ns_32s_32_2_1_Adder_8_U.ce  ? \add_32ns_32s_32_2_1_U19.top_add_32ns_32s_32_2_1_Adder_8_U.fas_s1  : \add_32ns_32s_32_2_1_U19.top_add_32ns_32s_32_2_1_Adder_8_U.sum_s1 ;
assign _090_ = \add_32ns_32s_32_2_1_U19.top_add_32ns_32s_32_2_1_Adder_8_U.u1.a  + \add_32ns_32s_32_2_1_U19.top_add_32ns_32s_32_2_1_Adder_8_U.u1.b ;
assign { \add_32ns_32s_32_2_1_U19.top_add_32ns_32s_32_2_1_Adder_8_U.u1.cout , \add_32ns_32s_32_2_1_U19.top_add_32ns_32s_32_2_1_Adder_8_U.u1.s  } = _090_ + \add_32ns_32s_32_2_1_U19.top_add_32ns_32s_32_2_1_Adder_8_U.u1.cin ;
assign _091_ = \add_32ns_32s_32_2_1_U19.top_add_32ns_32s_32_2_1_Adder_8_U.u2.a  + \add_32ns_32s_32_2_1_U19.top_add_32ns_32s_32_2_1_Adder_8_U.u2.b ;
assign { \add_32ns_32s_32_2_1_U19.top_add_32ns_32s_32_2_1_Adder_8_U.u2.cout , \add_32ns_32s_32_2_1_U19.top_add_32ns_32s_32_2_1_Adder_8_U.u2.s  } = _091_ + \add_32ns_32s_32_2_1_U19.top_add_32ns_32s_32_2_1_Adder_8_U.u2.cin ;
always @(posedge \add_32s_32ns_32_2_1_U10.top_add_32s_32ns_32_2_1_Adder_7_U.clk )
\add_32s_32ns_32_2_1_U10.top_add_32s_32ns_32_2_1_Adder_7_U.bin_s1  <= _093_;
always @(posedge \add_32s_32ns_32_2_1_U10.top_add_32s_32ns_32_2_1_Adder_7_U.clk )
\add_32s_32ns_32_2_1_U10.top_add_32s_32ns_32_2_1_Adder_7_U.ain_s1  <= _092_;
always @(posedge \add_32s_32ns_32_2_1_U10.top_add_32s_32ns_32_2_1_Adder_7_U.clk )
\add_32s_32ns_32_2_1_U10.top_add_32s_32ns_32_2_1_Adder_7_U.sum_s1  <= _095_;
always @(posedge \add_32s_32ns_32_2_1_U10.top_add_32s_32ns_32_2_1_Adder_7_U.clk )
\add_32s_32ns_32_2_1_U10.top_add_32s_32ns_32_2_1_Adder_7_U.carry_s1  <= _094_;
assign _093_ = \add_32s_32ns_32_2_1_U10.top_add_32s_32ns_32_2_1_Adder_7_U.ce  ? \add_32s_32ns_32_2_1_U10.top_add_32s_32ns_32_2_1_Adder_7_U.b [31:16] : \add_32s_32ns_32_2_1_U10.top_add_32s_32ns_32_2_1_Adder_7_U.bin_s1 ;
assign _092_ = \add_32s_32ns_32_2_1_U10.top_add_32s_32ns_32_2_1_Adder_7_U.ce  ? \add_32s_32ns_32_2_1_U10.top_add_32s_32ns_32_2_1_Adder_7_U.a [31:16] : \add_32s_32ns_32_2_1_U10.top_add_32s_32ns_32_2_1_Adder_7_U.ain_s1 ;
assign _094_ = \add_32s_32ns_32_2_1_U10.top_add_32s_32ns_32_2_1_Adder_7_U.ce  ? \add_32s_32ns_32_2_1_U10.top_add_32s_32ns_32_2_1_Adder_7_U.facout_s1  : \add_32s_32ns_32_2_1_U10.top_add_32s_32ns_32_2_1_Adder_7_U.carry_s1 ;
assign _095_ = \add_32s_32ns_32_2_1_U10.top_add_32s_32ns_32_2_1_Adder_7_U.ce  ? \add_32s_32ns_32_2_1_U10.top_add_32s_32ns_32_2_1_Adder_7_U.fas_s1  : \add_32s_32ns_32_2_1_U10.top_add_32s_32ns_32_2_1_Adder_7_U.sum_s1 ;
assign _096_ = \add_32s_32ns_32_2_1_U10.top_add_32s_32ns_32_2_1_Adder_7_U.u1.a  + \add_32s_32ns_32_2_1_U10.top_add_32s_32ns_32_2_1_Adder_7_U.u1.b ;
assign { \add_32s_32ns_32_2_1_U10.top_add_32s_32ns_32_2_1_Adder_7_U.u1.cout , \add_32s_32ns_32_2_1_U10.top_add_32s_32ns_32_2_1_Adder_7_U.u1.s  } = _096_ + \add_32s_32ns_32_2_1_U10.top_add_32s_32ns_32_2_1_Adder_7_U.u1.cin ;
assign _097_ = \add_32s_32ns_32_2_1_U10.top_add_32s_32ns_32_2_1_Adder_7_U.u2.a  + \add_32s_32ns_32_2_1_U10.top_add_32s_32ns_32_2_1_Adder_7_U.u2.b ;
assign { \add_32s_32ns_32_2_1_U10.top_add_32s_32ns_32_2_1_Adder_7_U.u2.cout , \add_32s_32ns_32_2_1_U10.top_add_32s_32ns_32_2_1_Adder_7_U.u2.s  } = _097_ + \add_32s_32ns_32_2_1_U10.top_add_32s_32ns_32_2_1_Adder_7_U.u2.cin ;
always @(posedge \add_32s_32ns_32_2_1_U16.top_add_32s_32ns_32_2_1_Adder_7_U.clk )
\add_32s_32ns_32_2_1_U16.top_add_32s_32ns_32_2_1_Adder_7_U.bin_s1  <= _099_;
always @(posedge \add_32s_32ns_32_2_1_U16.top_add_32s_32ns_32_2_1_Adder_7_U.clk )
\add_32s_32ns_32_2_1_U16.top_add_32s_32ns_32_2_1_Adder_7_U.ain_s1  <= _098_;
always @(posedge \add_32s_32ns_32_2_1_U16.top_add_32s_32ns_32_2_1_Adder_7_U.clk )
\add_32s_32ns_32_2_1_U16.top_add_32s_32ns_32_2_1_Adder_7_U.sum_s1  <= _101_;
always @(posedge \add_32s_32ns_32_2_1_U16.top_add_32s_32ns_32_2_1_Adder_7_U.clk )
\add_32s_32ns_32_2_1_U16.top_add_32s_32ns_32_2_1_Adder_7_U.carry_s1  <= _100_;
assign _099_ = \add_32s_32ns_32_2_1_U16.top_add_32s_32ns_32_2_1_Adder_7_U.ce  ? \add_32s_32ns_32_2_1_U16.top_add_32s_32ns_32_2_1_Adder_7_U.b [31:16] : \add_32s_32ns_32_2_1_U16.top_add_32s_32ns_32_2_1_Adder_7_U.bin_s1 ;
assign _098_ = \add_32s_32ns_32_2_1_U16.top_add_32s_32ns_32_2_1_Adder_7_U.ce  ? \add_32s_32ns_32_2_1_U16.top_add_32s_32ns_32_2_1_Adder_7_U.a [31:16] : \add_32s_32ns_32_2_1_U16.top_add_32s_32ns_32_2_1_Adder_7_U.ain_s1 ;
assign _100_ = \add_32s_32ns_32_2_1_U16.top_add_32s_32ns_32_2_1_Adder_7_U.ce  ? \add_32s_32ns_32_2_1_U16.top_add_32s_32ns_32_2_1_Adder_7_U.facout_s1  : \add_32s_32ns_32_2_1_U16.top_add_32s_32ns_32_2_1_Adder_7_U.carry_s1 ;
assign _101_ = \add_32s_32ns_32_2_1_U16.top_add_32s_32ns_32_2_1_Adder_7_U.ce  ? \add_32s_32ns_32_2_1_U16.top_add_32s_32ns_32_2_1_Adder_7_U.fas_s1  : \add_32s_32ns_32_2_1_U16.top_add_32s_32ns_32_2_1_Adder_7_U.sum_s1 ;
assign _102_ = \add_32s_32ns_32_2_1_U16.top_add_32s_32ns_32_2_1_Adder_7_U.u1.a  + \add_32s_32ns_32_2_1_U16.top_add_32s_32ns_32_2_1_Adder_7_U.u1.b ;
assign { \add_32s_32ns_32_2_1_U16.top_add_32s_32ns_32_2_1_Adder_7_U.u1.cout , \add_32s_32ns_32_2_1_U16.top_add_32s_32ns_32_2_1_Adder_7_U.u1.s  } = _102_ + \add_32s_32ns_32_2_1_U16.top_add_32s_32ns_32_2_1_Adder_7_U.u1.cin ;
assign _103_ = \add_32s_32ns_32_2_1_U16.top_add_32s_32ns_32_2_1_Adder_7_U.u2.a  + \add_32s_32ns_32_2_1_U16.top_add_32s_32ns_32_2_1_Adder_7_U.u2.b ;
assign { \add_32s_32ns_32_2_1_U16.top_add_32s_32ns_32_2_1_Adder_7_U.u2.cout , \add_32s_32ns_32_2_1_U16.top_add_32s_32ns_32_2_1_Adder_7_U.u2.s  } = _103_ + \add_32s_32ns_32_2_1_U16.top_add_32s_32ns_32_2_1_Adder_7_U.u2.cin ;
always @(posedge \add_34s_34ns_34_2_1_U4.top_add_34s_34ns_34_2_1_Adder_3_U.clk )
\add_34s_34ns_34_2_1_U4.top_add_34s_34ns_34_2_1_Adder_3_U.bin_s1  <= _105_;
always @(posedge \add_34s_34ns_34_2_1_U4.top_add_34s_34ns_34_2_1_Adder_3_U.clk )
\add_34s_34ns_34_2_1_U4.top_add_34s_34ns_34_2_1_Adder_3_U.ain_s1  <= _104_;
always @(posedge \add_34s_34ns_34_2_1_U4.top_add_34s_34ns_34_2_1_Adder_3_U.clk )
\add_34s_34ns_34_2_1_U4.top_add_34s_34ns_34_2_1_Adder_3_U.sum_s1  <= _107_;
always @(posedge \add_34s_34ns_34_2_1_U4.top_add_34s_34ns_34_2_1_Adder_3_U.clk )
\add_34s_34ns_34_2_1_U4.top_add_34s_34ns_34_2_1_Adder_3_U.carry_s1  <= _106_;
assign _105_ = \add_34s_34ns_34_2_1_U4.top_add_34s_34ns_34_2_1_Adder_3_U.ce  ? \add_34s_34ns_34_2_1_U4.top_add_34s_34ns_34_2_1_Adder_3_U.b [33:17] : \add_34s_34ns_34_2_1_U4.top_add_34s_34ns_34_2_1_Adder_3_U.bin_s1 ;
assign _104_ = \add_34s_34ns_34_2_1_U4.top_add_34s_34ns_34_2_1_Adder_3_U.ce  ? \add_34s_34ns_34_2_1_U4.top_add_34s_34ns_34_2_1_Adder_3_U.a [33:17] : \add_34s_34ns_34_2_1_U4.top_add_34s_34ns_34_2_1_Adder_3_U.ain_s1 ;
assign _106_ = \add_34s_34ns_34_2_1_U4.top_add_34s_34ns_34_2_1_Adder_3_U.ce  ? \add_34s_34ns_34_2_1_U4.top_add_34s_34ns_34_2_1_Adder_3_U.facout_s1  : \add_34s_34ns_34_2_1_U4.top_add_34s_34ns_34_2_1_Adder_3_U.carry_s1 ;
assign _107_ = \add_34s_34ns_34_2_1_U4.top_add_34s_34ns_34_2_1_Adder_3_U.ce  ? \add_34s_34ns_34_2_1_U4.top_add_34s_34ns_34_2_1_Adder_3_U.fas_s1  : \add_34s_34ns_34_2_1_U4.top_add_34s_34ns_34_2_1_Adder_3_U.sum_s1 ;
assign _108_ = \add_34s_34ns_34_2_1_U4.top_add_34s_34ns_34_2_1_Adder_3_U.u1.a  + \add_34s_34ns_34_2_1_U4.top_add_34s_34ns_34_2_1_Adder_3_U.u1.b ;
assign { \add_34s_34ns_34_2_1_U4.top_add_34s_34ns_34_2_1_Adder_3_U.u1.cout , \add_34s_34ns_34_2_1_U4.top_add_34s_34ns_34_2_1_Adder_3_U.u1.s  } = _108_ + \add_34s_34ns_34_2_1_U4.top_add_34s_34ns_34_2_1_Adder_3_U.u1.cin ;
assign _109_ = \add_34s_34ns_34_2_1_U4.top_add_34s_34ns_34_2_1_Adder_3_U.u2.a  + \add_34s_34ns_34_2_1_U4.top_add_34s_34ns_34_2_1_Adder_3_U.u2.b ;
assign { \add_34s_34ns_34_2_1_U4.top_add_34s_34ns_34_2_1_Adder_3_U.u2.cout , \add_34s_34ns_34_2_1_U4.top_add_34s_34ns_34_2_1_Adder_3_U.u2.s  } = _109_ + \add_34s_34ns_34_2_1_U4.top_add_34s_34ns_34_2_1_Adder_3_U.u2.cin ;
always @(posedge \add_34s_34s_34_2_1_U17.top_add_34s_34s_34_2_1_Adder_5_U.clk )
\add_34s_34s_34_2_1_U17.top_add_34s_34s_34_2_1_Adder_5_U.bin_s1  <= _111_;
always @(posedge \add_34s_34s_34_2_1_U17.top_add_34s_34s_34_2_1_Adder_5_U.clk )
\add_34s_34s_34_2_1_U17.top_add_34s_34s_34_2_1_Adder_5_U.ain_s1  <= _110_;
always @(posedge \add_34s_34s_34_2_1_U17.top_add_34s_34s_34_2_1_Adder_5_U.clk )
\add_34s_34s_34_2_1_U17.top_add_34s_34s_34_2_1_Adder_5_U.sum_s1  <= _113_;
always @(posedge \add_34s_34s_34_2_1_U17.top_add_34s_34s_34_2_1_Adder_5_U.clk )
\add_34s_34s_34_2_1_U17.top_add_34s_34s_34_2_1_Adder_5_U.carry_s1  <= _112_;
assign _111_ = \add_34s_34s_34_2_1_U17.top_add_34s_34s_34_2_1_Adder_5_U.ce  ? \add_34s_34s_34_2_1_U17.top_add_34s_34s_34_2_1_Adder_5_U.b [33:17] : \add_34s_34s_34_2_1_U17.top_add_34s_34s_34_2_1_Adder_5_U.bin_s1 ;
assign _110_ = \add_34s_34s_34_2_1_U17.top_add_34s_34s_34_2_1_Adder_5_U.ce  ? \add_34s_34s_34_2_1_U17.top_add_34s_34s_34_2_1_Adder_5_U.a [33:17] : \add_34s_34s_34_2_1_U17.top_add_34s_34s_34_2_1_Adder_5_U.ain_s1 ;
assign _112_ = \add_34s_34s_34_2_1_U17.top_add_34s_34s_34_2_1_Adder_5_U.ce  ? \add_34s_34s_34_2_1_U17.top_add_34s_34s_34_2_1_Adder_5_U.facout_s1  : \add_34s_34s_34_2_1_U17.top_add_34s_34s_34_2_1_Adder_5_U.carry_s1 ;
assign _113_ = \add_34s_34s_34_2_1_U17.top_add_34s_34s_34_2_1_Adder_5_U.ce  ? \add_34s_34s_34_2_1_U17.top_add_34s_34s_34_2_1_Adder_5_U.fas_s1  : \add_34s_34s_34_2_1_U17.top_add_34s_34s_34_2_1_Adder_5_U.sum_s1 ;
assign _114_ = \add_34s_34s_34_2_1_U17.top_add_34s_34s_34_2_1_Adder_5_U.u1.a  + \add_34s_34s_34_2_1_U17.top_add_34s_34s_34_2_1_Adder_5_U.u1.b ;
assign { \add_34s_34s_34_2_1_U17.top_add_34s_34s_34_2_1_Adder_5_U.u1.cout , \add_34s_34s_34_2_1_U17.top_add_34s_34s_34_2_1_Adder_5_U.u1.s  } = _114_ + \add_34s_34s_34_2_1_U17.top_add_34s_34s_34_2_1_Adder_5_U.u1.cin ;
assign _115_ = \add_34s_34s_34_2_1_U17.top_add_34s_34s_34_2_1_Adder_5_U.u2.a  + \add_34s_34s_34_2_1_U17.top_add_34s_34s_34_2_1_Adder_5_U.u2.b ;
assign { \add_34s_34s_34_2_1_U17.top_add_34s_34s_34_2_1_Adder_5_U.u2.cout , \add_34s_34s_34_2_1_U17.top_add_34s_34s_34_2_1_Adder_5_U.u2.s  } = _115_ + \add_34s_34s_34_2_1_U17.top_add_34s_34s_34_2_1_Adder_5_U.u2.cin ;
always @(posedge \add_34s_34s_34_2_1_U6.top_add_34s_34s_34_2_1_Adder_5_U.clk )
\add_34s_34s_34_2_1_U6.top_add_34s_34s_34_2_1_Adder_5_U.bin_s1  <= _117_;
always @(posedge \add_34s_34s_34_2_1_U6.top_add_34s_34s_34_2_1_Adder_5_U.clk )
\add_34s_34s_34_2_1_U6.top_add_34s_34s_34_2_1_Adder_5_U.ain_s1  <= _116_;
always @(posedge \add_34s_34s_34_2_1_U6.top_add_34s_34s_34_2_1_Adder_5_U.clk )
\add_34s_34s_34_2_1_U6.top_add_34s_34s_34_2_1_Adder_5_U.sum_s1  <= _119_;
always @(posedge \add_34s_34s_34_2_1_U6.top_add_34s_34s_34_2_1_Adder_5_U.clk )
\add_34s_34s_34_2_1_U6.top_add_34s_34s_34_2_1_Adder_5_U.carry_s1  <= _118_;
assign _117_ = \add_34s_34s_34_2_1_U6.top_add_34s_34s_34_2_1_Adder_5_U.ce  ? \add_34s_34s_34_2_1_U6.top_add_34s_34s_34_2_1_Adder_5_U.b [33:17] : \add_34s_34s_34_2_1_U6.top_add_34s_34s_34_2_1_Adder_5_U.bin_s1 ;
assign _116_ = \add_34s_34s_34_2_1_U6.top_add_34s_34s_34_2_1_Adder_5_U.ce  ? \add_34s_34s_34_2_1_U6.top_add_34s_34s_34_2_1_Adder_5_U.a [33:17] : \add_34s_34s_34_2_1_U6.top_add_34s_34s_34_2_1_Adder_5_U.ain_s1 ;
assign _118_ = \add_34s_34s_34_2_1_U6.top_add_34s_34s_34_2_1_Adder_5_U.ce  ? \add_34s_34s_34_2_1_U6.top_add_34s_34s_34_2_1_Adder_5_U.facout_s1  : \add_34s_34s_34_2_1_U6.top_add_34s_34s_34_2_1_Adder_5_U.carry_s1 ;
assign _119_ = \add_34s_34s_34_2_1_U6.top_add_34s_34s_34_2_1_Adder_5_U.ce  ? \add_34s_34s_34_2_1_U6.top_add_34s_34s_34_2_1_Adder_5_U.fas_s1  : \add_34s_34s_34_2_1_U6.top_add_34s_34s_34_2_1_Adder_5_U.sum_s1 ;
assign _120_ = \add_34s_34s_34_2_1_U6.top_add_34s_34s_34_2_1_Adder_5_U.u1.a  + \add_34s_34s_34_2_1_U6.top_add_34s_34s_34_2_1_Adder_5_U.u1.b ;
assign { \add_34s_34s_34_2_1_U6.top_add_34s_34s_34_2_1_Adder_5_U.u1.cout , \add_34s_34s_34_2_1_U6.top_add_34s_34s_34_2_1_Adder_5_U.u1.s  } = _120_ + \add_34s_34s_34_2_1_U6.top_add_34s_34s_34_2_1_Adder_5_U.u1.cin ;
assign _121_ = \add_34s_34s_34_2_1_U6.top_add_34s_34s_34_2_1_Adder_5_U.u2.a  + \add_34s_34s_34_2_1_U6.top_add_34s_34s_34_2_1_Adder_5_U.u2.b ;
assign { \add_34s_34s_34_2_1_U6.top_add_34s_34s_34_2_1_Adder_5_U.u2.cout , \add_34s_34s_34_2_1_U6.top_add_34s_34s_34_2_1_Adder_5_U.u2.s  } = _121_ + \add_34s_34s_34_2_1_U6.top_add_34s_34s_34_2_1_Adder_5_U.u2.cin ;
always @(posedge \add_47s_47s_47_2_1_U12.top_add_47s_47s_47_2_1_Adder_9_U.clk )
\add_47s_47s_47_2_1_U12.top_add_47s_47s_47_2_1_Adder_9_U.bin_s1  <= _123_;
always @(posedge \add_47s_47s_47_2_1_U12.top_add_47s_47s_47_2_1_Adder_9_U.clk )
\add_47s_47s_47_2_1_U12.top_add_47s_47s_47_2_1_Adder_9_U.ain_s1  <= _122_;
always @(posedge \add_47s_47s_47_2_1_U12.top_add_47s_47s_47_2_1_Adder_9_U.clk )
\add_47s_47s_47_2_1_U12.top_add_47s_47s_47_2_1_Adder_9_U.sum_s1  <= _125_;
always @(posedge \add_47s_47s_47_2_1_U12.top_add_47s_47s_47_2_1_Adder_9_U.clk )
\add_47s_47s_47_2_1_U12.top_add_47s_47s_47_2_1_Adder_9_U.carry_s1  <= _124_;
assign _123_ = \add_47s_47s_47_2_1_U12.top_add_47s_47s_47_2_1_Adder_9_U.ce  ? \add_47s_47s_47_2_1_U12.top_add_47s_47s_47_2_1_Adder_9_U.b [46:23] : \add_47s_47s_47_2_1_U12.top_add_47s_47s_47_2_1_Adder_9_U.bin_s1 ;
assign _122_ = \add_47s_47s_47_2_1_U12.top_add_47s_47s_47_2_1_Adder_9_U.ce  ? \add_47s_47s_47_2_1_U12.top_add_47s_47s_47_2_1_Adder_9_U.a [46:23] : \add_47s_47s_47_2_1_U12.top_add_47s_47s_47_2_1_Adder_9_U.ain_s1 ;
assign _124_ = \add_47s_47s_47_2_1_U12.top_add_47s_47s_47_2_1_Adder_9_U.ce  ? \add_47s_47s_47_2_1_U12.top_add_47s_47s_47_2_1_Adder_9_U.facout_s1  : \add_47s_47s_47_2_1_U12.top_add_47s_47s_47_2_1_Adder_9_U.carry_s1 ;
assign _125_ = \add_47s_47s_47_2_1_U12.top_add_47s_47s_47_2_1_Adder_9_U.ce  ? \add_47s_47s_47_2_1_U12.top_add_47s_47s_47_2_1_Adder_9_U.fas_s1  : \add_47s_47s_47_2_1_U12.top_add_47s_47s_47_2_1_Adder_9_U.sum_s1 ;
assign _126_ = \add_47s_47s_47_2_1_U12.top_add_47s_47s_47_2_1_Adder_9_U.u1.a  + \add_47s_47s_47_2_1_U12.top_add_47s_47s_47_2_1_Adder_9_U.u1.b ;
assign { \add_47s_47s_47_2_1_U12.top_add_47s_47s_47_2_1_Adder_9_U.u1.cout , \add_47s_47s_47_2_1_U12.top_add_47s_47s_47_2_1_Adder_9_U.u1.s  } = _126_ + \add_47s_47s_47_2_1_U12.top_add_47s_47s_47_2_1_Adder_9_U.u1.cin ;
assign _127_ = \add_47s_47s_47_2_1_U12.top_add_47s_47s_47_2_1_Adder_9_U.u2.a  + \add_47s_47s_47_2_1_U12.top_add_47s_47s_47_2_1_Adder_9_U.u2.b ;
assign { \add_47s_47s_47_2_1_U12.top_add_47s_47s_47_2_1_Adder_9_U.u2.cout , \add_47s_47s_47_2_1_U12.top_add_47s_47s_47_2_1_Adder_9_U.u2.s  } = _127_ + \add_47s_47s_47_2_1_U12.top_add_47s_47s_47_2_1_Adder_9_U.u2.cin ;
assign \add_5s_5ns_5_1_1_U15.top_add_5s_5ns_5_1_1_Adder_10_U.s  = \add_5s_5ns_5_1_1_U15.top_add_5s_5ns_5_1_1_Adder_10_U.a  + \add_5s_5ns_5_1_1_U15.top_add_5s_5ns_5_1_1_Adder_10_U.b ;
assign \add_7s_7ns_7_1_1_U1.top_add_7s_7ns_7_1_1_Adder_0_U.s  = \add_7s_7ns_7_1_1_U1.top_add_7s_7ns_7_1_1_Adder_0_U.a  + \add_7s_7ns_7_1_1_U1.top_add_7s_7ns_7_1_1_Adder_0_U.b ;
assign \add_8s_8ns_8_1_1_U3.top_add_8s_8ns_8_1_1_Adder_2_U.s  = \add_8s_8ns_8_1_1_U3.top_add_8s_8ns_8_1_1_Adder_2_U.a  + \add_8s_8ns_8_1_1_U3.top_add_8s_8ns_8_1_1_Adder_2_U.b ;
assign \add_9ns_9s_9_1_1_U2.top_add_9ns_9s_9_1_1_Adder_1_U.s  = \add_9ns_9s_9_1_1_U2.top_add_9ns_9s_9_1_1_Adder_1_U.a  + \add_9ns_9s_9_1_1_U2.top_add_9ns_9s_9_1_1_Adder_1_U.b ;
assign \add_9s_9ns_9_1_1_U9.top_add_9s_9ns_9_1_1_Adder_6_U.s  = \add_9s_9ns_9_1_1_U9.top_add_9s_9ns_9_1_1_Adder_6_U.a  + \add_9s_9ns_9_1_1_U9.top_add_9s_9ns_9_1_1_Adder_6_U.b ;
assign _128_ = | op_7[1:0];
assign _129_ = | { trunc_ln851_3_reg_856, 11'h000 };
always @(posedge ap_clk)
ret_V_reg_846[2:0] <= 3'h0;
always @(posedge ap_clk)
trunc_ln851_3_reg_856 <= 3'h0;
always @(posedge ap_clk)
sext_ln850_reg_726 <= _034_;
always @(posedge ap_clk)
select_ln703_reg_742 <= _032_;
always @(posedge ap_clk)
select_ln353_reg_747 <= _031_;
always @(posedge ap_clk)
select_ln353_1_reg_774 <= _030_;
always @(posedge ap_clk)
ret_V_20_reg_955 <= _026_;
always @(posedge ap_clk)
ret_V_18_reg_893 <= _024_;
always @(posedge ap_clk)
ret_V_19_reg_938 <= _025_;
always @(posedge ap_clk)
ret_V_18_cast_reg_943 <= _023_;
always @(posedge ap_clk)
ret_V_reg_846[7:3] <= _029_;
always @(posedge ap_clk)
ret_V_16_reg_851 <= _021_;
always @(posedge ap_clk)
ret_V_15_reg_811 <= _020_;
always @(posedge ap_clk)
ret_V_17_reg_876 <= _022_;
always @(posedge ap_clk)
ret_V_15_cast_reg_881 <= _019_;
always @(posedge ap_clk)
ret_V_13_reg_757 <= _017_;
always @(posedge ap_clk)
ret_V_8_cast_reg_762 <= _028_;
always @(posedge ap_clk)
ret_V_14_reg_794 <= _018_;
always @(posedge ap_clk)
ret_V_11_cast_reg_799 <= _015_;
always @(posedge ap_clk)
op_31_V_reg_918 <= _014_;
always @(posedge ap_clk)
op_26_V_reg_836 <= _013_;
always @(posedge ap_clk)
sext_ln835_reg_695 <= _033_;
always @(posedge ap_clk)
icmp_ln851_reg_701 <= _012_;
always @(posedge ap_clk)
ret_V_2_reg_706 <= _027_;
always @(posedge ap_clk)
icmp_ln851_2_reg_871 <= _011_;
always @(posedge ap_clk)
ret_V_12_reg_711 <= _016_;
always @(posedge ap_clk)
tmp_reg_716 <= _035_;
always @(posedge ap_clk)
icmp_ln851_1_reg_721 <= _010_;
always @(posedge ap_clk)
add_ln69_3_reg_903 <= _006_;
always @(posedge ap_clk)
add_ln69_4_reg_908 <= _007_;
always @(posedge ap_clk)
add_ln69_reg_821 <= _008_;
always @(posedge ap_clk)
add_ln69_1_reg_826 <= _005_;
always @(posedge ap_clk)
add_ln691_reg_732 <= _004_;
always @(posedge ap_clk)
add_ln691_4_reg_950 <= _003_;
always @(posedge ap_clk)
add_ln691_3_reg_888 <= _002_;
always @(posedge ap_clk)
add_ln691_2_reg_806 <= _001_;
always @(posedge ap_clk)
add_ln691_1_reg_769 <= _000_;
always @(posedge ap_clk)
ap_CS_fsm <= _009_;
assign _036_ = _041_ ? 2'h2 : 2'h1;
assign _130_ = ap_CS_fsm == 1'h1;
function [35:0] _389_;
input [35:0] a;
input [1295:0] b;
input [35:0] s;
case (s)
36'b000000000000000000000000000000000001:
_389_ = b[35:0];
36'b000000000000000000000000000000000010:
_389_ = b[71:36];
36'b000000000000000000000000000000000100:
_389_ = b[107:72];
36'b000000000000000000000000000000001000:
_389_ = b[143:108];
36'b000000000000000000000000000000010000:
_389_ = b[179:144];
36'b000000000000000000000000000000100000:
_389_ = b[215:180];
36'b000000000000000000000000000001000000:
_389_ = b[251:216];
36'b000000000000000000000000000010000000:
_389_ = b[287:252];
36'b000000000000000000000000000100000000:
_389_ = b[323:288];
36'b000000000000000000000000001000000000:
_389_ = b[359:324];
36'b000000000000000000000000010000000000:
_389_ = b[395:360];
36'b000000000000000000000000100000000000:
_389_ = b[431:396];
36'b000000000000000000000001000000000000:
_389_ = b[467:432];
36'b000000000000000000000010000000000000:
_389_ = b[503:468];
36'b000000000000000000000100000000000000:
_389_ = b[539:504];
36'b000000000000000000001000000000000000:
_389_ = b[575:540];
36'b000000000000000000010000000000000000:
_389_ = b[611:576];
36'b000000000000000000100000000000000000:
_389_ = b[647:612];
36'b000000000000000001000000000000000000:
_389_ = b[683:648];
36'b000000000000000010000000000000000000:
_389_ = b[719:684];
36'b000000000000000100000000000000000000:
_389_ = b[755:720];
36'b000000000000001000000000000000000000:
_389_ = b[791:756];
36'b000000000000010000000000000000000000:
_389_ = b[827:792];
36'b000000000000100000000000000000000000:
_389_ = b[863:828];
36'b000000000001000000000000000000000000:
_389_ = b[899:864];
36'b000000000010000000000000000000000000:
_389_ = b[935:900];
36'b000000000100000000000000000000000000:
_389_ = b[971:936];
36'b000000001000000000000000000000000000:
_389_ = b[1007:972];
36'b000000010000000000000000000000000000:
_389_ = b[1043:1008];
36'b000000100000000000000000000000000000:
_389_ = b[1079:1044];
36'b000001000000000000000000000000000000:
_389_ = b[1115:1080];
36'b000010000000000000000000000000000000:
_389_ = b[1151:1116];
36'b000100000000000000000000000000000000:
_389_ = b[1187:1152];
36'b001000000000000000000000000000000000:
_389_ = b[1223:1188];
36'b010000000000000000000000000000000000:
_389_ = b[1259:1224];
36'b100000000000000000000000000000000000:
_389_ = b[1295:1260];
36'b000000000000000000000000000000000000:
_389_ = a;
default:
_389_ = 36'bx;
endcase
endfunction
assign ap_NS_fsm = _389_(36'hxxxxxxxxx, { 34'h000000000, _036_, 1260'h000000004000000008000000010000000020000000040000000080000000100000000200000000400000000800000001000000002000000004000000008000000010000000020000000040000000080000000100000000200000000400000000800000001000000002000000004000000008000000010000000020000000040000000080000000100000000200000000400000000800000000000000001 }, { _130_, _165_, _164_, _163_, _162_, _161_, _160_, _159_, _158_, _157_, _156_, _155_, _154_, _153_, _152_, _151_, _150_, _149_, _148_, _147_, _146_, _145_, _144_, _143_, _142_, _141_, _140_, _139_, _138_, _137_, _136_, _135_, _134_, _133_, _132_, _131_ });
assign _131_ = ap_CS_fsm == 36'h800000000;
assign _132_ = ap_CS_fsm == 35'h400000000;
assign _133_ = ap_CS_fsm == 34'h200000000;
assign _134_ = ap_CS_fsm == 33'h100000000;
assign _135_ = ap_CS_fsm == 32'd2147483648;
assign _136_ = ap_CS_fsm == 31'h40000000;
assign _137_ = ap_CS_fsm == 30'h20000000;
assign _138_ = ap_CS_fsm == 29'h10000000;
assign _139_ = ap_CS_fsm == 28'h8000000;
assign _140_ = ap_CS_fsm == 27'h4000000;
assign _141_ = ap_CS_fsm == 26'h2000000;
assign _142_ = ap_CS_fsm == 25'h1000000;
assign _143_ = ap_CS_fsm == 24'h800000;
assign _144_ = ap_CS_fsm == 23'h400000;
assign _145_ = ap_CS_fsm == 22'h200000;
assign _146_ = ap_CS_fsm == 21'h100000;
assign _147_ = ap_CS_fsm == 20'h80000;
assign _148_ = ap_CS_fsm == 19'h40000;
assign _149_ = ap_CS_fsm == 18'h20000;
assign _150_ = ap_CS_fsm == 17'h10000;
assign _151_ = ap_CS_fsm == 16'h8000;
assign _152_ = ap_CS_fsm == 15'h4000;
assign _153_ = ap_CS_fsm == 14'h2000;
assign _154_ = ap_CS_fsm == 13'h1000;
assign _155_ = ap_CS_fsm == 12'h800;
assign _156_ = ap_CS_fsm == 11'h400;
assign _157_ = ap_CS_fsm == 10'h200;
assign _158_ = ap_CS_fsm == 9'h100;
assign _159_ = ap_CS_fsm == 8'h80;
assign _160_ = ap_CS_fsm == 7'h40;
assign _161_ = ap_CS_fsm == 6'h20;
assign _162_ = ap_CS_fsm == 5'h10;
assign _163_ = ap_CS_fsm == 4'h8;
assign _164_ = ap_CS_fsm == 3'h4;
assign _165_ = ap_CS_fsm == 2'h2;
assign op_33_ap_vld = ap_CS_fsm[35] ? 1'h1 : 1'h0;
assign ap_idle = _040_ ? 1'h1 : 1'h0;
assign _034_ = ap_CS_fsm[2] ? { tmp_reg_716[6], tmp_reg_716 } : sext_ln850_reg_726;
assign _031_ = ap_CS_fsm[3] ? select_ln353_fu_341_p3 : select_ln353_reg_747;
assign _032_ = ap_CS_fsm[3] ? select_ln703_fu_328_p3 : select_ln703_reg_742;
assign _030_ = ap_CS_fsm[8] ? select_ln353_1_fu_391_p3 : select_ln353_1_reg_774;
assign _026_ = ap_CS_fsm[33] ? ret_V_20_fu_673_p3 : ret_V_20_reg_955;
assign _024_ = ap_CS_fsm[24] ? ret_V_18_fu_587_p3 : ret_V_18_reg_893;
assign _023_ = ap_CS_fsm[30] ? grp_fu_636_p2[32:1] : ret_V_18_cast_reg_943;
assign _025_ = ap_CS_fsm[30] ? grp_fu_636_p2 : ret_V_19_reg_938;
assign _021_ = ap_CS_fsm[19] ? grp_fu_492_p2 : ret_V_16_reg_851;
assign _029_ = ap_CS_fsm[19] ? ret_V_fu_509_p2[7:3] : ret_V_reg_846[7:3];
assign _020_ = ap_CS_fsm[13] ? ret_V_15_fu_450_p3 : ret_V_15_reg_811;
assign _019_ = ap_CS_fsm[21] ? grp_fu_541_p2[45:14] : ret_V_15_cast_reg_881;
assign _022_ = ap_CS_fsm[21] ? grp_fu_541_p2 : ret_V_17_reg_876;
assign _028_ = ap_CS_fsm[5] ? grp_fu_359_p2[32:1] : ret_V_8_cast_reg_762;
assign _017_ = ap_CS_fsm[5] ? grp_fu_359_p2 : ret_V_13_reg_757;
assign _015_ = ap_CS_fsm[10] ? grp_fu_413_p2[32:1] : ret_V_11_cast_reg_799;
assign _018_ = ap_CS_fsm[10] ? grp_fu_413_p2 : ret_V_14_reg_794;
assign _014_ = ap_CS_fsm[28] ? grp_fu_616_p2 : op_31_V_reg_918;
assign _013_ = ap_CS_fsm[17] ? grp_fu_483_p2 : op_26_V_reg_836;
assign _027_ = ap_CS_fsm[0] ? ret_V_2_fu_249_p2 : ret_V_2_reg_706;
assign _012_ = ap_CS_fsm[0] ? icmp_ln851_fu_243_p2 : icmp_ln851_reg_701;
assign _033_ = ap_CS_fsm[0] ? { op_5[7], op_5[7:2] } : sext_ln835_reg_695;
assign _011_ = ap_CS_fsm[20] ? icmp_ln851_2_fu_554_p2 : icmp_ln851_2_reg_871;
assign _010_ = ap_CS_fsm[1] ? icmp_ln851_1_fu_306_p2 : icmp_ln851_1_reg_721;
assign _035_ = ap_CS_fsm[1] ? ret_V_12_fu_286_p2[8:2] : tmp_reg_716;
assign _016_ = ap_CS_fsm[1] ? ret_V_12_fu_286_p2 : ret_V_12_reg_711;
assign _007_ = ap_CS_fsm[26] ? add_ln69_4_fu_607_p2 : add_ln69_4_reg_908;
assign _006_ = ap_CS_fsm[26] ? grp_fu_594_p2 : add_ln69_3_reg_903;
assign _005_ = ap_CS_fsm[15] ? add_ln69_1_fu_474_p2 : add_ln69_1_reg_826;
assign _008_ = ap_CS_fsm[15] ? grp_fu_461_p2 : add_ln69_reg_821;
assign _004_ = _039_ ? add_ln691_fu_315_p2 : add_ln691_reg_732;
assign _003_ = ap_CS_fsm[32] ? grp_fu_652_p2 : add_ln691_4_reg_950;
assign _002_ = _038_ ? grp_fu_570_p2 : add_ln691_3_reg_888;
assign _001_ = ap_CS_fsm[12] ? grp_fu_429_p2 : add_ln691_2_reg_806;
assign _000_ = _037_ ? grp_fu_374_p2 : add_ln691_1_reg_769;
assign _009_ = ap_rst ? 36'h000000001 : ap_NS_fsm;
assign icmp_ln851_1_fu_306_p2 = _128_ ? 1'h1 : 1'h0;
assign icmp_ln851_2_fu_554_p2 = _129_ ? 1'h1 : 1'h0;
assign icmp_ln851_fu_243_p2 = _043_ ? 1'h1 : 1'h0;
assign ret_V_15_fu_450_p3 = ret_V_14_reg_794[33] ? select_ln850_3_fu_444_p3 : ret_V_11_cast_reg_799;
assign ret_V_18_fu_587_p3 = ret_V_17_reg_876[46] ? select_ln850_4_fu_582_p3 : ret_V_15_cast_reg_881;
assign ret_V_20_fu_673_p3 = ret_V_19_reg_938[33] ? select_ln850_5_fu_667_p3 : ret_V_18_cast_reg_943;
assign select_ln353_1_fu_391_p3 = ret_V_13_reg_757[33] ? select_ln850_6_fu_386_p3 : ret_V_8_cast_reg_762;
assign select_ln353_fu_341_p3 = ret_V_12_reg_711[8] ? select_ln850_2_fu_336_p3 : sext_ln850_reg_726;
assign select_ln703_fu_328_p3 = op_4 ? 34'h3ffffffff : 34'h000000000;
assign select_ln850_1_fu_271_p3 = op_5[7] ? select_ln850_fu_266_p3 : sext_ln835_reg_695;
assign select_ln850_2_fu_336_p3 = icmp_ln851_1_reg_721 ? add_ln691_reg_732 : sext_ln850_reg_726;
assign select_ln850_3_fu_444_p3 = op_9[0] ? add_ln691_2_reg_806 : ret_V_11_cast_reg_799;
assign select_ln850_4_fu_582_p3 = icmp_ln851_2_reg_871 ? add_ln691_3_reg_888 : ret_V_15_cast_reg_881;
assign select_ln850_5_fu_667_p3 = op_18[0] ? add_ln691_4_reg_950 : ret_V_18_cast_reg_943;
assign select_ln850_6_fu_386_p3 = op_4 ? add_ln691_1_reg_769 : ret_V_8_cast_reg_762;
assign select_ln850_fu_266_p3 = icmp_ln851_reg_701 ? sext_ln835_reg_695 : ret_V_2_reg_706;
assign add_ln691_fu_315_p0 = { tmp_reg_716[6], tmp_reg_716 };
assign add_ln69_1_fu_474_p0 = { op_10[7], op_10 };
assign add_ln69_1_fu_474_p1 = { 5'h00, op_11 };
assign add_ln69_4_fu_607_p0 = { op_17[3], op_17 };
assign add_ln69_4_fu_607_p1 = { 3'h0, op_15 };
assign ap_CS_fsm_state1 = ap_CS_fsm[0];
assign ap_CS_fsm_state10 = ap_CS_fsm[9];
assign ap_CS_fsm_state11 = ap_CS_fsm[10];
assign ap_CS_fsm_state12 = ap_CS_fsm[11];
assign ap_CS_fsm_state13 = ap_CS_fsm[12];
assign ap_CS_fsm_state14 = ap_CS_fsm[13];
assign ap_CS_fsm_state15 = ap_CS_fsm[14];
assign ap_CS_fsm_state16 = ap_CS_fsm[15];
assign ap_CS_fsm_state17 = ap_CS_fsm[16];
assign ap_CS_fsm_state18 = ap_CS_fsm[17];
assign ap_CS_fsm_state19 = ap_CS_fsm[18];
assign ap_CS_fsm_state2 = ap_CS_fsm[1];
assign ap_CS_fsm_state20 = ap_CS_fsm[19];
assign ap_CS_fsm_state21 = ap_CS_fsm[20];
assign ap_CS_fsm_state22 = ap_CS_fsm[21];
assign ap_CS_fsm_state23 = ap_CS_fsm[22];
assign ap_CS_fsm_state24 = ap_CS_fsm[23];
assign ap_CS_fsm_state25 = ap_CS_fsm[24];
assign ap_CS_fsm_state26 = ap_CS_fsm[25];
assign ap_CS_fsm_state27 = ap_CS_fsm[26];
assign ap_CS_fsm_state28 = ap_CS_fsm[27];
assign ap_CS_fsm_state29 = ap_CS_fsm[28];
assign ap_CS_fsm_state3 = ap_CS_fsm[2];
assign ap_CS_fsm_state30 = ap_CS_fsm[29];
assign ap_CS_fsm_state31 = ap_CS_fsm[30];
assign ap_CS_fsm_state32 = ap_CS_fsm[31];
assign ap_CS_fsm_state33 = ap_CS_fsm[32];
assign ap_CS_fsm_state34 = ap_CS_fsm[33];
assign ap_CS_fsm_state35 = ap_CS_fsm[34];
assign ap_CS_fsm_state36 = ap_CS_fsm[35];
assign ap_CS_fsm_state4 = ap_CS_fsm[3];
assign ap_CS_fsm_state5 = ap_CS_fsm[4];
assign ap_CS_fsm_state6 = ap_CS_fsm[5];
assign ap_CS_fsm_state7 = ap_CS_fsm[6];
assign ap_CS_fsm_state8 = ap_CS_fsm[7];
assign ap_CS_fsm_state9 = ap_CS_fsm[8];
assign ap_done = op_33_ap_vld;
assign ap_ready = op_33_ap_vld;
assign grp_fu_359_p0 = { select_ln353_reg_747[7], select_ln353_reg_747[7], select_ln353_reg_747[7], select_ln353_reg_747[7], select_ln353_reg_747[7], select_ln353_reg_747[7], select_ln353_reg_747[7], select_ln353_reg_747[7], select_ln353_reg_747[7], select_ln353_reg_747[7], select_ln353_reg_747[7], select_ln353_reg_747[7], select_ln353_reg_747[7], select_ln353_reg_747[7], select_ln353_reg_747[7], select_ln353_reg_747[7], select_ln353_reg_747[7], select_ln353_reg_747[7], select_ln353_reg_747[7], select_ln353_reg_747[7], select_ln353_reg_747[7], select_ln353_reg_747[7], select_ln353_reg_747[7], select_ln353_reg_747[7], select_ln353_reg_747[7], select_ln353_reg_747, 1'h0 };
assign grp_fu_413_p0 = { select_ln353_1_reg_774[31], select_ln353_1_reg_774, 1'h0 };
assign grp_fu_413_p1 = { op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9 };
assign grp_fu_461_p1 = { 16'h0000, op_12 };
assign grp_fu_483_p0 = { add_ln69_1_reg_826[8], add_ln69_1_reg_826[8], add_ln69_1_reg_826[8], add_ln69_1_reg_826[8], add_ln69_1_reg_826[8], add_ln69_1_reg_826[8], add_ln69_1_reg_826[8], add_ln69_1_reg_826[8], add_ln69_1_reg_826[8], add_ln69_1_reg_826[8], add_ln69_1_reg_826[8], add_ln69_1_reg_826[8], add_ln69_1_reg_826[8], add_ln69_1_reg_826[8], add_ln69_1_reg_826[8], add_ln69_1_reg_826[8], add_ln69_1_reg_826[8], add_ln69_1_reg_826[8], add_ln69_1_reg_826[8], add_ln69_1_reg_826[8], add_ln69_1_reg_826[8], add_ln69_1_reg_826[8], add_ln69_1_reg_826[8], add_ln69_1_reg_826 };
assign grp_fu_492_p1 = { op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13 };
assign grp_fu_541_p0 = { ret_V_16_reg_851[31], ret_V_16_reg_851, 14'h0000 };
assign grp_fu_541_p1 = { ret_V_reg_846[7], ret_V_reg_846[7], ret_V_reg_846[7], ret_V_reg_846[7], ret_V_reg_846[7], ret_V_reg_846[7], ret_V_reg_846[7], ret_V_reg_846[7], ret_V_reg_846[7], ret_V_reg_846[7], ret_V_reg_846[7], ret_V_reg_846[7], ret_V_reg_846[7], ret_V_reg_846[7], ret_V_reg_846[7], ret_V_reg_846[7], ret_V_reg_846[7], ret_V_reg_846[7], ret_V_reg_846[7], ret_V_reg_846[7], ret_V_reg_846[7], ret_V_reg_846[7], ret_V_reg_846[7], ret_V_reg_846[7], ret_V_reg_846[7], ret_V_reg_846[7], ret_V_reg_846[7], ret_V_reg_846[7], ret_V_reg_846, 11'h000 };
assign grp_fu_616_p0 = { add_ln69_4_reg_908[4], add_ln69_4_reg_908[4], add_ln69_4_reg_908[4], add_ln69_4_reg_908[4], add_ln69_4_reg_908[4], add_ln69_4_reg_908[4], add_ln69_4_reg_908[4], add_ln69_4_reg_908[4], add_ln69_4_reg_908[4], add_ln69_4_reg_908[4], add_ln69_4_reg_908[4], add_ln69_4_reg_908[4], add_ln69_4_reg_908[4], add_ln69_4_reg_908[4], add_ln69_4_reg_908[4], add_ln69_4_reg_908[4], add_ln69_4_reg_908[4], add_ln69_4_reg_908[4], add_ln69_4_reg_908[4], add_ln69_4_reg_908[4], add_ln69_4_reg_908[4], add_ln69_4_reg_908[4], add_ln69_4_reg_908[4], add_ln69_4_reg_908[4], add_ln69_4_reg_908[4], add_ln69_4_reg_908[4], add_ln69_4_reg_908[4], add_ln69_4_reg_908 };
assign grp_fu_636_p0 = { op_31_V_reg_918[31], op_31_V_reg_918, 1'h0 };
assign grp_fu_636_p1 = { op_18[7], op_18[7], op_18[7], op_18[7], op_18[7], op_18[7], op_18[7], op_18[7], op_18[7], op_18[7], op_18[7], op_18[7], op_18[7], op_18[7], op_18[7], op_18[7], op_18[7], op_18[7], op_18[7], op_18[7], op_18[7], op_18[7], op_18[7], op_18[7], op_18[7], op_18[7], op_18 };
assign grp_fu_684_p1 = { op_19[7], op_19[7], op_19[7], op_19[7], op_19[7], op_19[7], op_19[7], op_19[7], op_19[7], op_19[7], op_19[7], op_19[7], op_19[7], op_19[7], op_19[7], op_19[7], op_19[7], op_19[7], op_19[7], op_19[7], op_19[7], op_19[7], op_19[7], op_19[7], op_19 };
assign op_14_V_fu_519_p3 = { ret_V_reg_846, 11'h000 };
assign op_33 = grp_fu_684_p2;
assign op_4_read_read_fu_140_p2 = op_4;
assign p_Result_1_fu_321_p3 = ret_V_12_reg_711[8];
assign p_Result_2_fu_379_p3 = ret_V_13_reg_757[33];
assign p_Result_3_fu_434_p3 = ret_V_14_reg_794[33];
assign p_Result_4_fu_575_p3 = ret_V_17_reg_876[46];
assign p_Result_5_fu_657_p3 = ret_V_19_reg_938[33];
assign p_Result_7_fu_547_p3 = { trunc_ln851_3_reg_856, 11'h000 };
assign p_Result_s_fu_255_p3 = op_5[7];
assign ret_V_12_fu_286_p0 = { select_ln850_1_fu_271_p3, 2'h0 };
assign ret_V_12_fu_286_p1 = { op_7[3], op_7[3], op_7[3], op_7[3], op_7[3], op_7 };
assign ret_V_1_fu_225_p4 = op_5[7:2];
assign ret_V_2_fu_249_p0 = { op_5[7], op_5[7:2] };
assign rhs_2_fu_402_p3 = { select_ln353_1_reg_774, 1'h0 };
assign rhs_5_fu_530_p3 = { ret_V_16_reg_851, 14'h0000 };
assign rhs_7_fu_625_p3 = { op_31_V_reg_918, 1'h0 };
assign rhs_fu_497_p3 = { op_6, 3'h0 };
assign sext_ln1192_fu_262_p0 = op_7;
assign sext_ln1194_fu_505_p1 = { op_6[3], op_6, 3'h0 };
assign sext_ln703_2_fu_621_p0 = op_18;
assign sext_ln703_fu_398_p0 = op_9;
assign sext_ln835_fu_235_p1 = { op_5[7], op_5[7:2] };
assign sext_ln850_fu_312_p1 = { tmp_reg_716[6], tmp_reg_716 };
assign tmp_3_fu_348_p3 = { select_ln353_reg_747, 1'h0 };
assign trunc_ln851_1_fu_302_p0 = op_7;
assign trunc_ln851_1_fu_302_p1 = op_7[1:0];
assign trunc_ln851_2_fu_441_p0 = op_9;
assign trunc_ln851_2_fu_441_p1 = op_9[0];
assign trunc_ln851_3_fu_515_p1 = ret_V_fu_509_p2[2:0];
assign trunc_ln851_4_fu_664_p0 = op_18;
assign trunc_ln851_4_fu_664_p1 = op_18[0];
assign trunc_ln851_fu_239_p1 = op_5[1:0];
assign \add_9s_9ns_9_1_1_U9.top_add_9s_9ns_9_1_1_Adder_6_U.a  = \add_9s_9ns_9_1_1_U9.din0 ;
assign \add_9s_9ns_9_1_1_U9.top_add_9s_9ns_9_1_1_Adder_6_U.b  = \add_9s_9ns_9_1_1_U9.din1 ;
assign \add_9s_9ns_9_1_1_U9.dout  = \add_9s_9ns_9_1_1_U9.top_add_9s_9ns_9_1_1_Adder_6_U.s ;
assign \add_9s_9ns_9_1_1_U9.din0  = { op_10[7], op_10 };
assign \add_9s_9ns_9_1_1_U9.din1  = { 5'h00, op_11 };
assign add_ln69_1_fu_474_p2 = \add_9s_9ns_9_1_1_U9.dout ;
assign \add_9ns_9s_9_1_1_U2.top_add_9ns_9s_9_1_1_Adder_1_U.a  = \add_9ns_9s_9_1_1_U2.din0 ;
assign \add_9ns_9s_9_1_1_U2.top_add_9ns_9s_9_1_1_Adder_1_U.b  = \add_9ns_9s_9_1_1_U2.din1 ;
assign \add_9ns_9s_9_1_1_U2.dout  = \add_9ns_9s_9_1_1_U2.top_add_9ns_9s_9_1_1_Adder_1_U.s ;
assign \add_9ns_9s_9_1_1_U2.din0  = { select_ln850_1_fu_271_p3, 2'h0 };
assign \add_9ns_9s_9_1_1_U2.din1  = { op_7[3], op_7[3], op_7[3], op_7[3], op_7[3], op_7 };
assign ret_V_12_fu_286_p2 = \add_9ns_9s_9_1_1_U2.dout ;
assign \add_8s_8ns_8_1_1_U3.top_add_8s_8ns_8_1_1_Adder_2_U.a  = \add_8s_8ns_8_1_1_U3.din0 ;
assign \add_8s_8ns_8_1_1_U3.top_add_8s_8ns_8_1_1_Adder_2_U.b  = \add_8s_8ns_8_1_1_U3.din1 ;
assign \add_8s_8ns_8_1_1_U3.dout  = \add_8s_8ns_8_1_1_U3.top_add_8s_8ns_8_1_1_Adder_2_U.s ;
assign \add_8s_8ns_8_1_1_U3.din0  = { tmp_reg_716[6], tmp_reg_716 };
assign \add_8s_8ns_8_1_1_U3.din1  = 8'h01;
assign add_ln691_fu_315_p2 = \add_8s_8ns_8_1_1_U3.dout ;
assign \add_7s_7ns_7_1_1_U1.top_add_7s_7ns_7_1_1_Adder_0_U.a  = \add_7s_7ns_7_1_1_U1.din0 ;
assign \add_7s_7ns_7_1_1_U1.top_add_7s_7ns_7_1_1_Adder_0_U.b  = \add_7s_7ns_7_1_1_U1.din1 ;
assign \add_7s_7ns_7_1_1_U1.dout  = \add_7s_7ns_7_1_1_U1.top_add_7s_7ns_7_1_1_Adder_0_U.s ;
assign \add_7s_7ns_7_1_1_U1.din0  = { op_5[7], op_5[7:2] };
assign \add_7s_7ns_7_1_1_U1.din1  = 7'h01;
assign ret_V_2_fu_249_p2 = \add_7s_7ns_7_1_1_U1.dout ;
assign \add_5s_5ns_5_1_1_U15.top_add_5s_5ns_5_1_1_Adder_10_U.a  = \add_5s_5ns_5_1_1_U15.din0 ;
assign \add_5s_5ns_5_1_1_U15.top_add_5s_5ns_5_1_1_Adder_10_U.b  = \add_5s_5ns_5_1_1_U15.din1 ;
assign \add_5s_5ns_5_1_1_U15.dout  = \add_5s_5ns_5_1_1_U15.top_add_5s_5ns_5_1_1_Adder_10_U.s ;
assign \add_5s_5ns_5_1_1_U15.din0  = { op_17[3], op_17 };
assign \add_5s_5ns_5_1_1_U15.din1  = { 3'h0, op_15 };
assign add_ln69_4_fu_607_p2 = \add_5s_5ns_5_1_1_U15.dout ;
assign \add_47s_47s_47_2_1_U12.top_add_47s_47s_47_2_1_Adder_9_U.ain_s0  = \add_47s_47s_47_2_1_U12.top_add_47s_47s_47_2_1_Adder_9_U.a ;
assign \add_47s_47s_47_2_1_U12.top_add_47s_47s_47_2_1_Adder_9_U.bin_s0  = \add_47s_47s_47_2_1_U12.top_add_47s_47s_47_2_1_Adder_9_U.b ;
assign \add_47s_47s_47_2_1_U12.top_add_47s_47s_47_2_1_Adder_9_U.s  = { \add_47s_47s_47_2_1_U12.top_add_47s_47s_47_2_1_Adder_9_U.fas_s2 , \add_47s_47s_47_2_1_U12.top_add_47s_47s_47_2_1_Adder_9_U.sum_s1  };
assign \add_47s_47s_47_2_1_U12.top_add_47s_47s_47_2_1_Adder_9_U.u2.a  = \add_47s_47s_47_2_1_U12.top_add_47s_47s_47_2_1_Adder_9_U.ain_s1 ;
assign \add_47s_47s_47_2_1_U12.top_add_47s_47s_47_2_1_Adder_9_U.u2.b  = \add_47s_47s_47_2_1_U12.top_add_47s_47s_47_2_1_Adder_9_U.bin_s1 ;
assign \add_47s_47s_47_2_1_U12.top_add_47s_47s_47_2_1_Adder_9_U.u2.cin  = \add_47s_47s_47_2_1_U12.top_add_47s_47s_47_2_1_Adder_9_U.carry_s1 ;
assign \add_47s_47s_47_2_1_U12.top_add_47s_47s_47_2_1_Adder_9_U.facout_s2  = \add_47s_47s_47_2_1_U12.top_add_47s_47s_47_2_1_Adder_9_U.u2.cout ;
assign \add_47s_47s_47_2_1_U12.top_add_47s_47s_47_2_1_Adder_9_U.fas_s2  = \add_47s_47s_47_2_1_U12.top_add_47s_47s_47_2_1_Adder_9_U.u2.s ;
assign \add_47s_47s_47_2_1_U12.top_add_47s_47s_47_2_1_Adder_9_U.u1.a  = \add_47s_47s_47_2_1_U12.top_add_47s_47s_47_2_1_Adder_9_U.a [22:0];
assign \add_47s_47s_47_2_1_U12.top_add_47s_47s_47_2_1_Adder_9_U.u1.b  = \add_47s_47s_47_2_1_U12.top_add_47s_47s_47_2_1_Adder_9_U.b [22:0];
assign \add_47s_47s_47_2_1_U12.top_add_47s_47s_47_2_1_Adder_9_U.u1.cin  = 1'h0;
assign \add_47s_47s_47_2_1_U12.top_add_47s_47s_47_2_1_Adder_9_U.facout_s1  = \add_47s_47s_47_2_1_U12.top_add_47s_47s_47_2_1_Adder_9_U.u1.cout ;
assign \add_47s_47s_47_2_1_U12.top_add_47s_47s_47_2_1_Adder_9_U.fas_s1  = \add_47s_47s_47_2_1_U12.top_add_47s_47s_47_2_1_Adder_9_U.u1.s ;
assign \add_47s_47s_47_2_1_U12.top_add_47s_47s_47_2_1_Adder_9_U.a  = \add_47s_47s_47_2_1_U12.din0 ;
assign \add_47s_47s_47_2_1_U12.top_add_47s_47s_47_2_1_Adder_9_U.b  = \add_47s_47s_47_2_1_U12.din1 ;
assign \add_47s_47s_47_2_1_U12.top_add_47s_47s_47_2_1_Adder_9_U.ce  = \add_47s_47s_47_2_1_U12.ce ;
assign \add_47s_47s_47_2_1_U12.top_add_47s_47s_47_2_1_Adder_9_U.clk  = \add_47s_47s_47_2_1_U12.clk ;
assign \add_47s_47s_47_2_1_U12.top_add_47s_47s_47_2_1_Adder_9_U.reset  = \add_47s_47s_47_2_1_U12.reset ;
assign \add_47s_47s_47_2_1_U12.dout  = \add_47s_47s_47_2_1_U12.top_add_47s_47s_47_2_1_Adder_9_U.s ;
assign \add_47s_47s_47_2_1_U12.ce  = 1'h1;
assign \add_47s_47s_47_2_1_U12.clk  = ap_clk;
assign \add_47s_47s_47_2_1_U12.din0  = { ret_V_16_reg_851[31], ret_V_16_reg_851, 14'h0000 };
assign \add_47s_47s_47_2_1_U12.din1  = { ret_V_reg_846[7], ret_V_reg_846[7], ret_V_reg_846[7], ret_V_reg_846[7], ret_V_reg_846[7], ret_V_reg_846[7], ret_V_reg_846[7], ret_V_reg_846[7], ret_V_reg_846[7], ret_V_reg_846[7], ret_V_reg_846[7], ret_V_reg_846[7], ret_V_reg_846[7], ret_V_reg_846[7], ret_V_reg_846[7], ret_V_reg_846[7], ret_V_reg_846[7], ret_V_reg_846[7], ret_V_reg_846[7], ret_V_reg_846[7], ret_V_reg_846[7], ret_V_reg_846[7], ret_V_reg_846[7], ret_V_reg_846[7], ret_V_reg_846[7], ret_V_reg_846[7], ret_V_reg_846[7], ret_V_reg_846[7], ret_V_reg_846, 11'h000 };
assign grp_fu_541_p2 = \add_47s_47s_47_2_1_U12.dout ;
assign \add_47s_47s_47_2_1_U12.reset  = ap_rst;
assign \add_34s_34s_34_2_1_U6.top_add_34s_34s_34_2_1_Adder_5_U.ain_s0  = \add_34s_34s_34_2_1_U6.top_add_34s_34s_34_2_1_Adder_5_U.a ;
assign \add_34s_34s_34_2_1_U6.top_add_34s_34s_34_2_1_Adder_5_U.bin_s0  = \add_34s_34s_34_2_1_U6.top_add_34s_34s_34_2_1_Adder_5_U.b ;
assign \add_34s_34s_34_2_1_U6.top_add_34s_34s_34_2_1_Adder_5_U.s  = { \add_34s_34s_34_2_1_U6.top_add_34s_34s_34_2_1_Adder_5_U.fas_s2 , \add_34s_34s_34_2_1_U6.top_add_34s_34s_34_2_1_Adder_5_U.sum_s1  };
assign \add_34s_34s_34_2_1_U6.top_add_34s_34s_34_2_1_Adder_5_U.u2.a  = \add_34s_34s_34_2_1_U6.top_add_34s_34s_34_2_1_Adder_5_U.ain_s1 ;
assign \add_34s_34s_34_2_1_U6.top_add_34s_34s_34_2_1_Adder_5_U.u2.b  = \add_34s_34s_34_2_1_U6.top_add_34s_34s_34_2_1_Adder_5_U.bin_s1 ;
assign \add_34s_34s_34_2_1_U6.top_add_34s_34s_34_2_1_Adder_5_U.u2.cin  = \add_34s_34s_34_2_1_U6.top_add_34s_34s_34_2_1_Adder_5_U.carry_s1 ;
assign \add_34s_34s_34_2_1_U6.top_add_34s_34s_34_2_1_Adder_5_U.facout_s2  = \add_34s_34s_34_2_1_U6.top_add_34s_34s_34_2_1_Adder_5_U.u2.cout ;
assign \add_34s_34s_34_2_1_U6.top_add_34s_34s_34_2_1_Adder_5_U.fas_s2  = \add_34s_34s_34_2_1_U6.top_add_34s_34s_34_2_1_Adder_5_U.u2.s ;
assign \add_34s_34s_34_2_1_U6.top_add_34s_34s_34_2_1_Adder_5_U.u1.a  = \add_34s_34s_34_2_1_U6.top_add_34s_34s_34_2_1_Adder_5_U.a [16:0];
assign \add_34s_34s_34_2_1_U6.top_add_34s_34s_34_2_1_Adder_5_U.u1.b  = \add_34s_34s_34_2_1_U6.top_add_34s_34s_34_2_1_Adder_5_U.b [16:0];
assign \add_34s_34s_34_2_1_U6.top_add_34s_34s_34_2_1_Adder_5_U.u1.cin  = 1'h0;
assign \add_34s_34s_34_2_1_U6.top_add_34s_34s_34_2_1_Adder_5_U.facout_s1  = \add_34s_34s_34_2_1_U6.top_add_34s_34s_34_2_1_Adder_5_U.u1.cout ;
assign \add_34s_34s_34_2_1_U6.top_add_34s_34s_34_2_1_Adder_5_U.fas_s1  = \add_34s_34s_34_2_1_U6.top_add_34s_34s_34_2_1_Adder_5_U.u1.s ;
assign \add_34s_34s_34_2_1_U6.top_add_34s_34s_34_2_1_Adder_5_U.a  = \add_34s_34s_34_2_1_U6.din0 ;
assign \add_34s_34s_34_2_1_U6.top_add_34s_34s_34_2_1_Adder_5_U.b  = \add_34s_34s_34_2_1_U6.din1 ;
assign \add_34s_34s_34_2_1_U6.top_add_34s_34s_34_2_1_Adder_5_U.ce  = \add_34s_34s_34_2_1_U6.ce ;
assign \add_34s_34s_34_2_1_U6.top_add_34s_34s_34_2_1_Adder_5_U.clk  = \add_34s_34s_34_2_1_U6.clk ;
assign \add_34s_34s_34_2_1_U6.top_add_34s_34s_34_2_1_Adder_5_U.reset  = \add_34s_34s_34_2_1_U6.reset ;
assign \add_34s_34s_34_2_1_U6.dout  = \add_34s_34s_34_2_1_U6.top_add_34s_34s_34_2_1_Adder_5_U.s ;
assign \add_34s_34s_34_2_1_U6.ce  = 1'h1;
assign \add_34s_34s_34_2_1_U6.clk  = ap_clk;
assign \add_34s_34s_34_2_1_U6.din0  = { select_ln353_1_reg_774[31], select_ln353_1_reg_774, 1'h0 };
assign \add_34s_34s_34_2_1_U6.din1  = { op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9 };
assign grp_fu_413_p2 = \add_34s_34s_34_2_1_U6.dout ;
assign \add_34s_34s_34_2_1_U6.reset  = ap_rst;
assign \add_34s_34s_34_2_1_U17.top_add_34s_34s_34_2_1_Adder_5_U.ain_s0  = \add_34s_34s_34_2_1_U17.top_add_34s_34s_34_2_1_Adder_5_U.a ;
assign \add_34s_34s_34_2_1_U17.top_add_34s_34s_34_2_1_Adder_5_U.bin_s0  = \add_34s_34s_34_2_1_U17.top_add_34s_34s_34_2_1_Adder_5_U.b ;
assign \add_34s_34s_34_2_1_U17.top_add_34s_34s_34_2_1_Adder_5_U.s  = { \add_34s_34s_34_2_1_U17.top_add_34s_34s_34_2_1_Adder_5_U.fas_s2 , \add_34s_34s_34_2_1_U17.top_add_34s_34s_34_2_1_Adder_5_U.sum_s1  };
assign \add_34s_34s_34_2_1_U17.top_add_34s_34s_34_2_1_Adder_5_U.u2.a  = \add_34s_34s_34_2_1_U17.top_add_34s_34s_34_2_1_Adder_5_U.ain_s1 ;
assign \add_34s_34s_34_2_1_U17.top_add_34s_34s_34_2_1_Adder_5_U.u2.b  = \add_34s_34s_34_2_1_U17.top_add_34s_34s_34_2_1_Adder_5_U.bin_s1 ;
assign \add_34s_34s_34_2_1_U17.top_add_34s_34s_34_2_1_Adder_5_U.u2.cin  = \add_34s_34s_34_2_1_U17.top_add_34s_34s_34_2_1_Adder_5_U.carry_s1 ;
assign \add_34s_34s_34_2_1_U17.top_add_34s_34s_34_2_1_Adder_5_U.facout_s2  = \add_34s_34s_34_2_1_U17.top_add_34s_34s_34_2_1_Adder_5_U.u2.cout ;
assign \add_34s_34s_34_2_1_U17.top_add_34s_34s_34_2_1_Adder_5_U.fas_s2  = \add_34s_34s_34_2_1_U17.top_add_34s_34s_34_2_1_Adder_5_U.u2.s ;
assign \add_34s_34s_34_2_1_U17.top_add_34s_34s_34_2_1_Adder_5_U.u1.a  = \add_34s_34s_34_2_1_U17.top_add_34s_34s_34_2_1_Adder_5_U.a [16:0];
assign \add_34s_34s_34_2_1_U17.top_add_34s_34s_34_2_1_Adder_5_U.u1.b  = \add_34s_34s_34_2_1_U17.top_add_34s_34s_34_2_1_Adder_5_U.b [16:0];
assign \add_34s_34s_34_2_1_U17.top_add_34s_34s_34_2_1_Adder_5_U.u1.cin  = 1'h0;
assign \add_34s_34s_34_2_1_U17.top_add_34s_34s_34_2_1_Adder_5_U.facout_s1  = \add_34s_34s_34_2_1_U17.top_add_34s_34s_34_2_1_Adder_5_U.u1.cout ;
assign \add_34s_34s_34_2_1_U17.top_add_34s_34s_34_2_1_Adder_5_U.fas_s1  = \add_34s_34s_34_2_1_U17.top_add_34s_34s_34_2_1_Adder_5_U.u1.s ;
assign \add_34s_34s_34_2_1_U17.top_add_34s_34s_34_2_1_Adder_5_U.a  = \add_34s_34s_34_2_1_U17.din0 ;
assign \add_34s_34s_34_2_1_U17.top_add_34s_34s_34_2_1_Adder_5_U.b  = \add_34s_34s_34_2_1_U17.din1 ;
assign \add_34s_34s_34_2_1_U17.top_add_34s_34s_34_2_1_Adder_5_U.ce  = \add_34s_34s_34_2_1_U17.ce ;
assign \add_34s_34s_34_2_1_U17.top_add_34s_34s_34_2_1_Adder_5_U.clk  = \add_34s_34s_34_2_1_U17.clk ;
assign \add_34s_34s_34_2_1_U17.top_add_34s_34s_34_2_1_Adder_5_U.reset  = \add_34s_34s_34_2_1_U17.reset ;
assign \add_34s_34s_34_2_1_U17.dout  = \add_34s_34s_34_2_1_U17.top_add_34s_34s_34_2_1_Adder_5_U.s ;
assign \add_34s_34s_34_2_1_U17.ce  = 1'h1;
assign \add_34s_34s_34_2_1_U17.clk  = ap_clk;
assign \add_34s_34s_34_2_1_U17.din0  = { op_31_V_reg_918[31], op_31_V_reg_918, 1'h0 };
assign \add_34s_34s_34_2_1_U17.din1  = { op_18[7], op_18[7], op_18[7], op_18[7], op_18[7], op_18[7], op_18[7], op_18[7], op_18[7], op_18[7], op_18[7], op_18[7], op_18[7], op_18[7], op_18[7], op_18[7], op_18[7], op_18[7], op_18[7], op_18[7], op_18[7], op_18[7], op_18[7], op_18[7], op_18[7], op_18[7], op_18 };
assign grp_fu_636_p2 = \add_34s_34s_34_2_1_U17.dout ;
assign \add_34s_34s_34_2_1_U17.reset  = ap_rst;
assign \add_34s_34ns_34_2_1_U4.top_add_34s_34ns_34_2_1_Adder_3_U.ain_s0  = \add_34s_34ns_34_2_1_U4.top_add_34s_34ns_34_2_1_Adder_3_U.a ;
assign \add_34s_34ns_34_2_1_U4.top_add_34s_34ns_34_2_1_Adder_3_U.bin_s0  = \add_34s_34ns_34_2_1_U4.top_add_34s_34ns_34_2_1_Adder_3_U.b ;
assign \add_34s_34ns_34_2_1_U4.top_add_34s_34ns_34_2_1_Adder_3_U.s  = { \add_34s_34ns_34_2_1_U4.top_add_34s_34ns_34_2_1_Adder_3_U.fas_s2 , \add_34s_34ns_34_2_1_U4.top_add_34s_34ns_34_2_1_Adder_3_U.sum_s1  };
assign \add_34s_34ns_34_2_1_U4.top_add_34s_34ns_34_2_1_Adder_3_U.u2.a  = \add_34s_34ns_34_2_1_U4.top_add_34s_34ns_34_2_1_Adder_3_U.ain_s1 ;
assign \add_34s_34ns_34_2_1_U4.top_add_34s_34ns_34_2_1_Adder_3_U.u2.b  = \add_34s_34ns_34_2_1_U4.top_add_34s_34ns_34_2_1_Adder_3_U.bin_s1 ;
assign \add_34s_34ns_34_2_1_U4.top_add_34s_34ns_34_2_1_Adder_3_U.u2.cin  = \add_34s_34ns_34_2_1_U4.top_add_34s_34ns_34_2_1_Adder_3_U.carry_s1 ;
assign \add_34s_34ns_34_2_1_U4.top_add_34s_34ns_34_2_1_Adder_3_U.facout_s2  = \add_34s_34ns_34_2_1_U4.top_add_34s_34ns_34_2_1_Adder_3_U.u2.cout ;
assign \add_34s_34ns_34_2_1_U4.top_add_34s_34ns_34_2_1_Adder_3_U.fas_s2  = \add_34s_34ns_34_2_1_U4.top_add_34s_34ns_34_2_1_Adder_3_U.u2.s ;
assign \add_34s_34ns_34_2_1_U4.top_add_34s_34ns_34_2_1_Adder_3_U.u1.a  = \add_34s_34ns_34_2_1_U4.top_add_34s_34ns_34_2_1_Adder_3_U.a [16:0];
assign \add_34s_34ns_34_2_1_U4.top_add_34s_34ns_34_2_1_Adder_3_U.u1.b  = \add_34s_34ns_34_2_1_U4.top_add_34s_34ns_34_2_1_Adder_3_U.b [16:0];
assign \add_34s_34ns_34_2_1_U4.top_add_34s_34ns_34_2_1_Adder_3_U.u1.cin  = 1'h0;
assign \add_34s_34ns_34_2_1_U4.top_add_34s_34ns_34_2_1_Adder_3_U.facout_s1  = \add_34s_34ns_34_2_1_U4.top_add_34s_34ns_34_2_1_Adder_3_U.u1.cout ;
assign \add_34s_34ns_34_2_1_U4.top_add_34s_34ns_34_2_1_Adder_3_U.fas_s1  = \add_34s_34ns_34_2_1_U4.top_add_34s_34ns_34_2_1_Adder_3_U.u1.s ;
assign \add_34s_34ns_34_2_1_U4.top_add_34s_34ns_34_2_1_Adder_3_U.a  = \add_34s_34ns_34_2_1_U4.din0 ;
assign \add_34s_34ns_34_2_1_U4.top_add_34s_34ns_34_2_1_Adder_3_U.b  = \add_34s_34ns_34_2_1_U4.din1 ;
assign \add_34s_34ns_34_2_1_U4.top_add_34s_34ns_34_2_1_Adder_3_U.ce  = \add_34s_34ns_34_2_1_U4.ce ;
assign \add_34s_34ns_34_2_1_U4.top_add_34s_34ns_34_2_1_Adder_3_U.clk  = \add_34s_34ns_34_2_1_U4.clk ;
assign \add_34s_34ns_34_2_1_U4.top_add_34s_34ns_34_2_1_Adder_3_U.reset  = \add_34s_34ns_34_2_1_U4.reset ;
assign \add_34s_34ns_34_2_1_U4.dout  = \add_34s_34ns_34_2_1_U4.top_add_34s_34ns_34_2_1_Adder_3_U.s ;
assign \add_34s_34ns_34_2_1_U4.ce  = 1'h1;
assign \add_34s_34ns_34_2_1_U4.clk  = ap_clk;
assign \add_34s_34ns_34_2_1_U4.din0  = { select_ln353_reg_747[7], select_ln353_reg_747[7], select_ln353_reg_747[7], select_ln353_reg_747[7], select_ln353_reg_747[7], select_ln353_reg_747[7], select_ln353_reg_747[7], select_ln353_reg_747[7], select_ln353_reg_747[7], select_ln353_reg_747[7], select_ln353_reg_747[7], select_ln353_reg_747[7], select_ln353_reg_747[7], select_ln353_reg_747[7], select_ln353_reg_747[7], select_ln353_reg_747[7], select_ln353_reg_747[7], select_ln353_reg_747[7], select_ln353_reg_747[7], select_ln353_reg_747[7], select_ln353_reg_747[7], select_ln353_reg_747[7], select_ln353_reg_747[7], select_ln353_reg_747[7], select_ln353_reg_747[7], select_ln353_reg_747, 1'h0 };
assign \add_34s_34ns_34_2_1_U4.din1  = select_ln703_reg_742;
assign grp_fu_359_p2 = \add_34s_34ns_34_2_1_U4.dout ;
assign \add_34s_34ns_34_2_1_U4.reset  = ap_rst;
assign \add_32s_32ns_32_2_1_U16.top_add_32s_32ns_32_2_1_Adder_7_U.ain_s0  = \add_32s_32ns_32_2_1_U16.top_add_32s_32ns_32_2_1_Adder_7_U.a ;
assign \add_32s_32ns_32_2_1_U16.top_add_32s_32ns_32_2_1_Adder_7_U.bin_s0  = \add_32s_32ns_32_2_1_U16.top_add_32s_32ns_32_2_1_Adder_7_U.b ;
assign \add_32s_32ns_32_2_1_U16.top_add_32s_32ns_32_2_1_Adder_7_U.s  = { \add_32s_32ns_32_2_1_U16.top_add_32s_32ns_32_2_1_Adder_7_U.fas_s2 , \add_32s_32ns_32_2_1_U16.top_add_32s_32ns_32_2_1_Adder_7_U.sum_s1  };
assign \add_32s_32ns_32_2_1_U16.top_add_32s_32ns_32_2_1_Adder_7_U.u2.a  = \add_32s_32ns_32_2_1_U16.top_add_32s_32ns_32_2_1_Adder_7_U.ain_s1 ;
assign \add_32s_32ns_32_2_1_U16.top_add_32s_32ns_32_2_1_Adder_7_U.u2.b  = \add_32s_32ns_32_2_1_U16.top_add_32s_32ns_32_2_1_Adder_7_U.bin_s1 ;
assign \add_32s_32ns_32_2_1_U16.top_add_32s_32ns_32_2_1_Adder_7_U.u2.cin  = \add_32s_32ns_32_2_1_U16.top_add_32s_32ns_32_2_1_Adder_7_U.carry_s1 ;
assign \add_32s_32ns_32_2_1_U16.top_add_32s_32ns_32_2_1_Adder_7_U.facout_s2  = \add_32s_32ns_32_2_1_U16.top_add_32s_32ns_32_2_1_Adder_7_U.u2.cout ;
assign \add_32s_32ns_32_2_1_U16.top_add_32s_32ns_32_2_1_Adder_7_U.fas_s2  = \add_32s_32ns_32_2_1_U16.top_add_32s_32ns_32_2_1_Adder_7_U.u2.s ;
assign \add_32s_32ns_32_2_1_U16.top_add_32s_32ns_32_2_1_Adder_7_U.u1.a  = \add_32s_32ns_32_2_1_U16.top_add_32s_32ns_32_2_1_Adder_7_U.a [15:0];
assign \add_32s_32ns_32_2_1_U16.top_add_32s_32ns_32_2_1_Adder_7_U.u1.b  = \add_32s_32ns_32_2_1_U16.top_add_32s_32ns_32_2_1_Adder_7_U.b [15:0];
assign \add_32s_32ns_32_2_1_U16.top_add_32s_32ns_32_2_1_Adder_7_U.u1.cin  = 1'h0;
assign \add_32s_32ns_32_2_1_U16.top_add_32s_32ns_32_2_1_Adder_7_U.facout_s1  = \add_32s_32ns_32_2_1_U16.top_add_32s_32ns_32_2_1_Adder_7_U.u1.cout ;
assign \add_32s_32ns_32_2_1_U16.top_add_32s_32ns_32_2_1_Adder_7_U.fas_s1  = \add_32s_32ns_32_2_1_U16.top_add_32s_32ns_32_2_1_Adder_7_U.u1.s ;
assign \add_32s_32ns_32_2_1_U16.top_add_32s_32ns_32_2_1_Adder_7_U.a  = \add_32s_32ns_32_2_1_U16.din0 ;
assign \add_32s_32ns_32_2_1_U16.top_add_32s_32ns_32_2_1_Adder_7_U.b  = \add_32s_32ns_32_2_1_U16.din1 ;
assign \add_32s_32ns_32_2_1_U16.top_add_32s_32ns_32_2_1_Adder_7_U.ce  = \add_32s_32ns_32_2_1_U16.ce ;
assign \add_32s_32ns_32_2_1_U16.top_add_32s_32ns_32_2_1_Adder_7_U.clk  = \add_32s_32ns_32_2_1_U16.clk ;
assign \add_32s_32ns_32_2_1_U16.top_add_32s_32ns_32_2_1_Adder_7_U.reset  = \add_32s_32ns_32_2_1_U16.reset ;
assign \add_32s_32ns_32_2_1_U16.dout  = \add_32s_32ns_32_2_1_U16.top_add_32s_32ns_32_2_1_Adder_7_U.s ;
assign \add_32s_32ns_32_2_1_U16.ce  = 1'h1;
assign \add_32s_32ns_32_2_1_U16.clk  = ap_clk;
assign \add_32s_32ns_32_2_1_U16.din0  = { add_ln69_4_reg_908[4], add_ln69_4_reg_908[4], add_ln69_4_reg_908[4], add_ln69_4_reg_908[4], add_ln69_4_reg_908[4], add_ln69_4_reg_908[4], add_ln69_4_reg_908[4], add_ln69_4_reg_908[4], add_ln69_4_reg_908[4], add_ln69_4_reg_908[4], add_ln69_4_reg_908[4], add_ln69_4_reg_908[4], add_ln69_4_reg_908[4], add_ln69_4_reg_908[4], add_ln69_4_reg_908[4], add_ln69_4_reg_908[4], add_ln69_4_reg_908[4], add_ln69_4_reg_908[4], add_ln69_4_reg_908[4], add_ln69_4_reg_908[4], add_ln69_4_reg_908[4], add_ln69_4_reg_908[4], add_ln69_4_reg_908[4], add_ln69_4_reg_908[4], add_ln69_4_reg_908[4], add_ln69_4_reg_908[4], add_ln69_4_reg_908[4], add_ln69_4_reg_908 };
assign \add_32s_32ns_32_2_1_U16.din1  = add_ln69_3_reg_903;
assign grp_fu_616_p2 = \add_32s_32ns_32_2_1_U16.dout ;
assign \add_32s_32ns_32_2_1_U16.reset  = ap_rst;
assign \add_32s_32ns_32_2_1_U10.top_add_32s_32ns_32_2_1_Adder_7_U.ain_s0  = \add_32s_32ns_32_2_1_U10.top_add_32s_32ns_32_2_1_Adder_7_U.a ;
assign \add_32s_32ns_32_2_1_U10.top_add_32s_32ns_32_2_1_Adder_7_U.bin_s0  = \add_32s_32ns_32_2_1_U10.top_add_32s_32ns_32_2_1_Adder_7_U.b ;
assign \add_32s_32ns_32_2_1_U10.top_add_32s_32ns_32_2_1_Adder_7_U.s  = { \add_32s_32ns_32_2_1_U10.top_add_32s_32ns_32_2_1_Adder_7_U.fas_s2 , \add_32s_32ns_32_2_1_U10.top_add_32s_32ns_32_2_1_Adder_7_U.sum_s1  };
assign \add_32s_32ns_32_2_1_U10.top_add_32s_32ns_32_2_1_Adder_7_U.u2.a  = \add_32s_32ns_32_2_1_U10.top_add_32s_32ns_32_2_1_Adder_7_U.ain_s1 ;
assign \add_32s_32ns_32_2_1_U10.top_add_32s_32ns_32_2_1_Adder_7_U.u2.b  = \add_32s_32ns_32_2_1_U10.top_add_32s_32ns_32_2_1_Adder_7_U.bin_s1 ;
assign \add_32s_32ns_32_2_1_U10.top_add_32s_32ns_32_2_1_Adder_7_U.u2.cin  = \add_32s_32ns_32_2_1_U10.top_add_32s_32ns_32_2_1_Adder_7_U.carry_s1 ;
assign \add_32s_32ns_32_2_1_U10.top_add_32s_32ns_32_2_1_Adder_7_U.facout_s2  = \add_32s_32ns_32_2_1_U10.top_add_32s_32ns_32_2_1_Adder_7_U.u2.cout ;
assign \add_32s_32ns_32_2_1_U10.top_add_32s_32ns_32_2_1_Adder_7_U.fas_s2  = \add_32s_32ns_32_2_1_U10.top_add_32s_32ns_32_2_1_Adder_7_U.u2.s ;
assign \add_32s_32ns_32_2_1_U10.top_add_32s_32ns_32_2_1_Adder_7_U.u1.a  = \add_32s_32ns_32_2_1_U10.top_add_32s_32ns_32_2_1_Adder_7_U.a [15:0];
assign \add_32s_32ns_32_2_1_U10.top_add_32s_32ns_32_2_1_Adder_7_U.u1.b  = \add_32s_32ns_32_2_1_U10.top_add_32s_32ns_32_2_1_Adder_7_U.b [15:0];
assign \add_32s_32ns_32_2_1_U10.top_add_32s_32ns_32_2_1_Adder_7_U.u1.cin  = 1'h0;
assign \add_32s_32ns_32_2_1_U10.top_add_32s_32ns_32_2_1_Adder_7_U.facout_s1  = \add_32s_32ns_32_2_1_U10.top_add_32s_32ns_32_2_1_Adder_7_U.u1.cout ;
assign \add_32s_32ns_32_2_1_U10.top_add_32s_32ns_32_2_1_Adder_7_U.fas_s1  = \add_32s_32ns_32_2_1_U10.top_add_32s_32ns_32_2_1_Adder_7_U.u1.s ;
assign \add_32s_32ns_32_2_1_U10.top_add_32s_32ns_32_2_1_Adder_7_U.a  = \add_32s_32ns_32_2_1_U10.din0 ;
assign \add_32s_32ns_32_2_1_U10.top_add_32s_32ns_32_2_1_Adder_7_U.b  = \add_32s_32ns_32_2_1_U10.din1 ;
assign \add_32s_32ns_32_2_1_U10.top_add_32s_32ns_32_2_1_Adder_7_U.ce  = \add_32s_32ns_32_2_1_U10.ce ;
assign \add_32s_32ns_32_2_1_U10.top_add_32s_32ns_32_2_1_Adder_7_U.clk  = \add_32s_32ns_32_2_1_U10.clk ;
assign \add_32s_32ns_32_2_1_U10.top_add_32s_32ns_32_2_1_Adder_7_U.reset  = \add_32s_32ns_32_2_1_U10.reset ;
assign \add_32s_32ns_32_2_1_U10.dout  = \add_32s_32ns_32_2_1_U10.top_add_32s_32ns_32_2_1_Adder_7_U.s ;
assign \add_32s_32ns_32_2_1_U10.ce  = 1'h1;
assign \add_32s_32ns_32_2_1_U10.clk  = ap_clk;
assign \add_32s_32ns_32_2_1_U10.din0  = { add_ln69_1_reg_826[8], add_ln69_1_reg_826[8], add_ln69_1_reg_826[8], add_ln69_1_reg_826[8], add_ln69_1_reg_826[8], add_ln69_1_reg_826[8], add_ln69_1_reg_826[8], add_ln69_1_reg_826[8], add_ln69_1_reg_826[8], add_ln69_1_reg_826[8], add_ln69_1_reg_826[8], add_ln69_1_reg_826[8], add_ln69_1_reg_826[8], add_ln69_1_reg_826[8], add_ln69_1_reg_826[8], add_ln69_1_reg_826[8], add_ln69_1_reg_826[8], add_ln69_1_reg_826[8], add_ln69_1_reg_826[8], add_ln69_1_reg_826[8], add_ln69_1_reg_826[8], add_ln69_1_reg_826[8], add_ln69_1_reg_826[8], add_ln69_1_reg_826 };
assign \add_32s_32ns_32_2_1_U10.din1  = add_ln69_reg_821;
assign grp_fu_483_p2 = \add_32s_32ns_32_2_1_U10.dout ;
assign \add_32s_32ns_32_2_1_U10.reset  = ap_rst;
assign \add_32ns_32s_32_2_1_U19.top_add_32ns_32s_32_2_1_Adder_8_U.ain_s0  = \add_32ns_32s_32_2_1_U19.top_add_32ns_32s_32_2_1_Adder_8_U.a ;
assign \add_32ns_32s_32_2_1_U19.top_add_32ns_32s_32_2_1_Adder_8_U.bin_s0  = \add_32ns_32s_32_2_1_U19.top_add_32ns_32s_32_2_1_Adder_8_U.b ;
assign \add_32ns_32s_32_2_1_U19.top_add_32ns_32s_32_2_1_Adder_8_U.s  = { \add_32ns_32s_32_2_1_U19.top_add_32ns_32s_32_2_1_Adder_8_U.fas_s2 , \add_32ns_32s_32_2_1_U19.top_add_32ns_32s_32_2_1_Adder_8_U.sum_s1  };
assign \add_32ns_32s_32_2_1_U19.top_add_32ns_32s_32_2_1_Adder_8_U.u2.a  = \add_32ns_32s_32_2_1_U19.top_add_32ns_32s_32_2_1_Adder_8_U.ain_s1 ;
assign \add_32ns_32s_32_2_1_U19.top_add_32ns_32s_32_2_1_Adder_8_U.u2.b  = \add_32ns_32s_32_2_1_U19.top_add_32ns_32s_32_2_1_Adder_8_U.bin_s1 ;
assign \add_32ns_32s_32_2_1_U19.top_add_32ns_32s_32_2_1_Adder_8_U.u2.cin  = \add_32ns_32s_32_2_1_U19.top_add_32ns_32s_32_2_1_Adder_8_U.carry_s1 ;
assign \add_32ns_32s_32_2_1_U19.top_add_32ns_32s_32_2_1_Adder_8_U.facout_s2  = \add_32ns_32s_32_2_1_U19.top_add_32ns_32s_32_2_1_Adder_8_U.u2.cout ;
assign \add_32ns_32s_32_2_1_U19.top_add_32ns_32s_32_2_1_Adder_8_U.fas_s2  = \add_32ns_32s_32_2_1_U19.top_add_32ns_32s_32_2_1_Adder_8_U.u2.s ;
assign \add_32ns_32s_32_2_1_U19.top_add_32ns_32s_32_2_1_Adder_8_U.u1.a  = \add_32ns_32s_32_2_1_U19.top_add_32ns_32s_32_2_1_Adder_8_U.a [15:0];
assign \add_32ns_32s_32_2_1_U19.top_add_32ns_32s_32_2_1_Adder_8_U.u1.b  = \add_32ns_32s_32_2_1_U19.top_add_32ns_32s_32_2_1_Adder_8_U.b [15:0];
assign \add_32ns_32s_32_2_1_U19.top_add_32ns_32s_32_2_1_Adder_8_U.u1.cin  = 1'h0;
assign \add_32ns_32s_32_2_1_U19.top_add_32ns_32s_32_2_1_Adder_8_U.facout_s1  = \add_32ns_32s_32_2_1_U19.top_add_32ns_32s_32_2_1_Adder_8_U.u1.cout ;
assign \add_32ns_32s_32_2_1_U19.top_add_32ns_32s_32_2_1_Adder_8_U.fas_s1  = \add_32ns_32s_32_2_1_U19.top_add_32ns_32s_32_2_1_Adder_8_U.u1.s ;
assign \add_32ns_32s_32_2_1_U19.top_add_32ns_32s_32_2_1_Adder_8_U.a  = \add_32ns_32s_32_2_1_U19.din0 ;
assign \add_32ns_32s_32_2_1_U19.top_add_32ns_32s_32_2_1_Adder_8_U.b  = \add_32ns_32s_32_2_1_U19.din1 ;
assign \add_32ns_32s_32_2_1_U19.top_add_32ns_32s_32_2_1_Adder_8_U.ce  = \add_32ns_32s_32_2_1_U19.ce ;
assign \add_32ns_32s_32_2_1_U19.top_add_32ns_32s_32_2_1_Adder_8_U.clk  = \add_32ns_32s_32_2_1_U19.clk ;
assign \add_32ns_32s_32_2_1_U19.top_add_32ns_32s_32_2_1_Adder_8_U.reset  = \add_32ns_32s_32_2_1_U19.reset ;
assign \add_32ns_32s_32_2_1_U19.dout  = \add_32ns_32s_32_2_1_U19.top_add_32ns_32s_32_2_1_Adder_8_U.s ;
assign \add_32ns_32s_32_2_1_U19.ce  = 1'h1;
assign \add_32ns_32s_32_2_1_U19.clk  = ap_clk;
assign \add_32ns_32s_32_2_1_U19.din0  = ret_V_20_reg_955;
assign \add_32ns_32s_32_2_1_U19.din1  = { op_19[7], op_19[7], op_19[7], op_19[7], op_19[7], op_19[7], op_19[7], op_19[7], op_19[7], op_19[7], op_19[7], op_19[7], op_19[7], op_19[7], op_19[7], op_19[7], op_19[7], op_19[7], op_19[7], op_19[7], op_19[7], op_19[7], op_19[7], op_19[7], op_19 };
assign grp_fu_684_p2 = \add_32ns_32s_32_2_1_U19.dout ;
assign \add_32ns_32s_32_2_1_U19.reset  = ap_rst;
assign \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.ain_s0  = \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.a ;
assign \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.bin_s0  = \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.b ;
assign \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.s  = { \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.fas_s2 , \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.sum_s1  };
assign \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.u2.a  = \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.ain_s1 ;
assign \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.u2.b  = \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.bin_s1 ;
assign \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.u2.cin  = \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.carry_s1 ;
assign \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.facout_s2  = \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.u2.cout ;
assign \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.fas_s2  = \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.u2.s ;
assign \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.u1.a  = \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.a [15:0];
assign \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.u1.b  = \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.b [15:0];
assign \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.u1.cin  = 1'h0;
assign \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.facout_s1  = \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.u1.cout ;
assign \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.fas_s1  = \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.u1.s ;
assign \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.a  = \add_32ns_32s_32_2_1_U11.din0 ;
assign \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.b  = \add_32ns_32s_32_2_1_U11.din1 ;
assign \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.ce  = \add_32ns_32s_32_2_1_U11.ce ;
assign \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.clk  = \add_32ns_32s_32_2_1_U11.clk ;
assign \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.reset  = \add_32ns_32s_32_2_1_U11.reset ;
assign \add_32ns_32s_32_2_1_U11.dout  = \add_32ns_32s_32_2_1_U11.top_add_32ns_32s_32_2_1_Adder_8_U.s ;
assign \add_32ns_32s_32_2_1_U11.ce  = 1'h1;
assign \add_32ns_32s_32_2_1_U11.clk  = ap_clk;
assign \add_32ns_32s_32_2_1_U11.din0  = op_26_V_reg_836;
assign \add_32ns_32s_32_2_1_U11.din1  = { op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13[1], op_13 };
assign grp_fu_492_p2 = \add_32ns_32s_32_2_1_U11.dout ;
assign \add_32ns_32s_32_2_1_U11.reset  = ap_rst;
assign \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.ain_s0  = \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.a ;
assign \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.bin_s0  = \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.b ;
assign \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.s  = { \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.fas_s2 , \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.sum_s1  };
assign \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.a  = \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.ain_s1 ;
assign \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.b  = \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.bin_s1 ;
assign \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.cin  = \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.carry_s1 ;
assign \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.facout_s2  = \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.cout ;
assign \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.fas_s2  = \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.s ;
assign \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.a  = \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.a [15:0];
assign \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.b  = \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.b [15:0];
assign \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.cin  = 1'h0;
assign \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.facout_s1  = \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.cout ;
assign \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.fas_s1  = \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.s ;
assign \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.a  = \add_32ns_32ns_32_2_1_U8.din0 ;
assign \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.b  = \add_32ns_32ns_32_2_1_U8.din1 ;
assign \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.ce  = \add_32ns_32ns_32_2_1_U8.ce ;
assign \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.clk  = \add_32ns_32ns_32_2_1_U8.clk ;
assign \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.reset  = \add_32ns_32ns_32_2_1_U8.reset ;
assign \add_32ns_32ns_32_2_1_U8.dout  = \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_4_U.s ;
assign \add_32ns_32ns_32_2_1_U8.ce  = 1'h1;
assign \add_32ns_32ns_32_2_1_U8.clk  = ap_clk;
assign \add_32ns_32ns_32_2_1_U8.din0  = ret_V_15_reg_811;
assign \add_32ns_32ns_32_2_1_U8.din1  = { 16'h0000, op_12 };
assign grp_fu_461_p2 = \add_32ns_32ns_32_2_1_U8.dout ;
assign \add_32ns_32ns_32_2_1_U8.reset  = ap_rst;
assign \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_4_U.ain_s0  = \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_4_U.a ;
assign \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_4_U.bin_s0  = \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_4_U.b ;
assign \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_4_U.s  = { \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_4_U.fas_s2 , \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_4_U.sum_s1  };
assign \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.a  = \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_4_U.ain_s1 ;
assign \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.b  = \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_4_U.bin_s1 ;
assign \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.cin  = \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_4_U.carry_s1 ;
assign \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_4_U.facout_s2  = \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.cout ;
assign \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_4_U.fas_s2  = \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.s ;
assign \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.a  = \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_4_U.a [15:0];
assign \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.b  = \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_4_U.b [15:0];
assign \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.cin  = 1'h0;
assign \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_4_U.facout_s1  = \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.cout ;
assign \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_4_U.fas_s1  = \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.s ;
assign \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_4_U.a  = \add_32ns_32ns_32_2_1_U7.din0 ;
assign \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_4_U.b  = \add_32ns_32ns_32_2_1_U7.din1 ;
assign \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_4_U.ce  = \add_32ns_32ns_32_2_1_U7.ce ;
assign \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_4_U.clk  = \add_32ns_32ns_32_2_1_U7.clk ;
assign \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_4_U.reset  = \add_32ns_32ns_32_2_1_U7.reset ;
assign \add_32ns_32ns_32_2_1_U7.dout  = \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_4_U.s ;
assign \add_32ns_32ns_32_2_1_U7.ce  = 1'h1;
assign \add_32ns_32ns_32_2_1_U7.clk  = ap_clk;
assign \add_32ns_32ns_32_2_1_U7.din0  = ret_V_11_cast_reg_799;
assign \add_32ns_32ns_32_2_1_U7.din1  = 32'd1;
assign grp_fu_429_p2 = \add_32ns_32ns_32_2_1_U7.dout ;
assign \add_32ns_32ns_32_2_1_U7.reset  = ap_rst;
assign \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.ain_s0  = \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.a ;
assign \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.bin_s0  = \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.b ;
assign \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.s  = { \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.fas_s2 , \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.sum_s1  };
assign \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.a  = \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.ain_s1 ;
assign \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.b  = \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.bin_s1 ;
assign \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.cin  = \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.carry_s1 ;
assign \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.facout_s2  = \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.cout ;
assign \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.fas_s2  = \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.s ;
assign \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.a  = \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.a [15:0];
assign \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.b  = \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.b [15:0];
assign \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.cin  = 1'h0;
assign \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.facout_s1  = \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.cout ;
assign \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.fas_s1  = \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.s ;
assign \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.a  = \add_32ns_32ns_32_2_1_U5.din0 ;
assign \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.b  = \add_32ns_32ns_32_2_1_U5.din1 ;
assign \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.ce  = \add_32ns_32ns_32_2_1_U5.ce ;
assign \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.clk  = \add_32ns_32ns_32_2_1_U5.clk ;
assign \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.reset  = \add_32ns_32ns_32_2_1_U5.reset ;
assign \add_32ns_32ns_32_2_1_U5.dout  = \add_32ns_32ns_32_2_1_U5.top_add_32ns_32ns_32_2_1_Adder_4_U.s ;
assign \add_32ns_32ns_32_2_1_U5.ce  = 1'h1;
assign \add_32ns_32ns_32_2_1_U5.clk  = ap_clk;
assign \add_32ns_32ns_32_2_1_U5.din0  = ret_V_8_cast_reg_762;
assign \add_32ns_32ns_32_2_1_U5.din1  = 32'd1;
assign grp_fu_374_p2 = \add_32ns_32ns_32_2_1_U5.dout ;
assign \add_32ns_32ns_32_2_1_U5.reset  = ap_rst;
assign \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_4_U.ain_s0  = \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_4_U.a ;
assign \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_4_U.bin_s0  = \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_4_U.b ;
assign \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_4_U.s  = { \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_4_U.fas_s2 , \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_4_U.sum_s1  };
assign \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.a  = \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_4_U.ain_s1 ;
assign \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.b  = \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_4_U.bin_s1 ;
assign \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.cin  = \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_4_U.carry_s1 ;
assign \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_4_U.facout_s2  = \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.cout ;
assign \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_4_U.fas_s2  = \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.s ;
assign \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.a  = \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_4_U.a [15:0];
assign \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.b  = \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_4_U.b [15:0];
assign \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.cin  = 1'h0;
assign \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_4_U.facout_s1  = \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.cout ;
assign \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_4_U.fas_s1  = \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.s ;
assign \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_4_U.a  = \add_32ns_32ns_32_2_1_U18.din0 ;
assign \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_4_U.b  = \add_32ns_32ns_32_2_1_U18.din1 ;
assign \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_4_U.ce  = \add_32ns_32ns_32_2_1_U18.ce ;
assign \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_4_U.clk  = \add_32ns_32ns_32_2_1_U18.clk ;
assign \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_4_U.reset  = \add_32ns_32ns_32_2_1_U18.reset ;
assign \add_32ns_32ns_32_2_1_U18.dout  = \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_4_U.s ;
assign \add_32ns_32ns_32_2_1_U18.ce  = 1'h1;
assign \add_32ns_32ns_32_2_1_U18.clk  = ap_clk;
assign \add_32ns_32ns_32_2_1_U18.din0  = ret_V_18_cast_reg_943;
assign \add_32ns_32ns_32_2_1_U18.din1  = 32'd1;
assign grp_fu_652_p2 = \add_32ns_32ns_32_2_1_U18.dout ;
assign \add_32ns_32ns_32_2_1_U18.reset  = ap_rst;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_4_U.ain_s0  = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_4_U.a ;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_4_U.bin_s0  = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_4_U.b ;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_4_U.s  = { \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_4_U.fas_s2 , \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_4_U.sum_s1  };
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.a  = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_4_U.ain_s1 ;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.b  = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_4_U.bin_s1 ;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.cin  = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_4_U.carry_s1 ;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_4_U.facout_s2  = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.cout ;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_4_U.fas_s2  = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.s ;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.a  = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_4_U.a [15:0];
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.b  = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_4_U.b [15:0];
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.cin  = 1'h0;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_4_U.facout_s1  = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.cout ;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_4_U.fas_s1  = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.s ;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_4_U.a  = \add_32ns_32ns_32_2_1_U14.din0 ;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_4_U.b  = \add_32ns_32ns_32_2_1_U14.din1 ;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_4_U.ce  = \add_32ns_32ns_32_2_1_U14.ce ;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_4_U.clk  = \add_32ns_32ns_32_2_1_U14.clk ;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_4_U.reset  = \add_32ns_32ns_32_2_1_U14.reset ;
assign \add_32ns_32ns_32_2_1_U14.dout  = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_4_U.s ;
assign \add_32ns_32ns_32_2_1_U14.ce  = 1'h1;
assign \add_32ns_32ns_32_2_1_U14.clk  = ap_clk;
assign \add_32ns_32ns_32_2_1_U14.din0  = ret_V_18_reg_893;
assign \add_32ns_32ns_32_2_1_U14.din1  = op_16;
assign grp_fu_594_p2 = \add_32ns_32ns_32_2_1_U14.dout ;
assign \add_32ns_32ns_32_2_1_U14.reset  = ap_rst;
assign \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_4_U.ain_s0  = \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_4_U.a ;
assign \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_4_U.bin_s0  = \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_4_U.b ;
assign \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_4_U.s  = { \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_4_U.fas_s2 , \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_4_U.sum_s1  };
assign \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.a  = \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_4_U.ain_s1 ;
assign \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.b  = \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_4_U.bin_s1 ;
assign \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.cin  = \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_4_U.carry_s1 ;
assign \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_4_U.facout_s2  = \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.cout ;
assign \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_4_U.fas_s2  = \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_4_U.u2.s ;
assign \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.a  = \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_4_U.a [15:0];
assign \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.b  = \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_4_U.b [15:0];
assign \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.cin  = 1'h0;
assign \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_4_U.facout_s1  = \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.cout ;
assign \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_4_U.fas_s1  = \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_4_U.u1.s ;
assign \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_4_U.a  = \add_32ns_32ns_32_2_1_U13.din0 ;
assign \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_4_U.b  = \add_32ns_32ns_32_2_1_U13.din1 ;
assign \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_4_U.ce  = \add_32ns_32ns_32_2_1_U13.ce ;
assign \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_4_U.clk  = \add_32ns_32ns_32_2_1_U13.clk ;
assign \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_4_U.reset  = \add_32ns_32ns_32_2_1_U13.reset ;
assign \add_32ns_32ns_32_2_1_U13.dout  = \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_4_U.s ;
assign \add_32ns_32ns_32_2_1_U13.ce  = 1'h1;
assign \add_32ns_32ns_32_2_1_U13.clk  = ap_clk;
assign \add_32ns_32ns_32_2_1_U13.din0  = ret_V_15_cast_reg_881;
assign \add_32ns_32ns_32_2_1_U13.din1  = 32'd1;
assign grp_fu_570_p2 = \add_32ns_32ns_32_2_1_U13.dout ;
assign \add_32ns_32ns_32_2_1_U13.reset  = ap_rst;
endmodule


// Product machine:
module top_A_times_top_B (ap_start, op_0, op_10, op_11, op_12, op_13, op_15, op_16, op_17, op_18, op_19, op_3, op_4, op_5, op_6, op_7, op_9, ap_clk, unsafe_signal);
input ap_start;
input [7:0] op_0;
input [7:0] op_10;
input [3:0] op_11;
input [15:0] op_12;
input [1:0] op_13;
input [1:0] op_15;
input [31:0] op_16;
input [3:0] op_17;
input [7:0] op_18;
input [7:0] op_19;
input [7:0] op_3;
input op_4;
input [7:0] op_5;
input [3:0] op_6;
input [3:0] op_7;
input [1:0] op_9;
input ap_clk;
output unsafe_signal;
reg _setup;
initial _setup = 1'b0;
always @ (posedge ap_clk) _setup <= 1'b1;
reg ap_start_internal;
always @ (posedge ap_clk) if (!_setup) ap_start_internal <= ap_start;
reg [7:0] op_0_internal;
always @ (posedge ap_clk) if (!_setup) op_0_internal <= op_0;
reg [7:0] op_10_internal;
always @ (posedge ap_clk) if (!_setup) op_10_internal <= op_10;
reg [3:0] op_11_internal;
always @ (posedge ap_clk) if (!_setup) op_11_internal <= op_11;
reg [15:0] op_12_internal;
always @ (posedge ap_clk) if (!_setup) op_12_internal <= op_12;
reg [1:0] op_13_internal;
always @ (posedge ap_clk) if (!_setup) op_13_internal <= op_13;
reg [1:0] op_15_internal;
always @ (posedge ap_clk) if (!_setup) op_15_internal <= op_15;
reg [31:0] op_16_internal;
always @ (posedge ap_clk) if (!_setup) op_16_internal <= op_16;
reg [3:0] op_17_internal;
always @ (posedge ap_clk) if (!_setup) op_17_internal <= op_17;
reg [7:0] op_18_internal;
always @ (posedge ap_clk) if (!_setup) op_18_internal <= op_18;
reg [7:0] op_19_internal;
always @ (posedge ap_clk) if (!_setup) op_19_internal <= op_19;
reg [7:0] op_3_internal;
always @ (posedge ap_clk) if (!_setup) op_3_internal <= op_3;
reg op_4_internal;
always @ (posedge ap_clk) if (!_setup) op_4_internal <= op_4;
reg [7:0] op_5_internal;
always @ (posedge ap_clk) if (!_setup) op_5_internal <= op_5;
reg [3:0] op_6_internal;
always @ (posedge ap_clk) if (!_setup) op_6_internal <= op_6;
reg [3:0] op_7_internal;
always @ (posedge ap_clk) if (!_setup) op_7_internal <= op_7;
reg [1:0] op_9_internal;
always @ (posedge ap_clk) if (!_setup) op_9_internal <= op_9;
wire ap_done_A;
wire ap_done_B;
wire ap_done_eq;
assign ap_done_eq = ap_done_A == ap_done_B;
wire ap_idle_A;
wire ap_idle_B;
wire ap_idle_eq;
assign ap_idle_eq = ap_idle_A == ap_idle_B;
wire ap_ready_A;
wire ap_ready_B;
wire ap_ready_eq;
assign ap_ready_eq = ap_ready_A == ap_ready_B;
wire [31:0] op_33_A;
wire [31:0] op_33_B;
wire op_33_eq;
assign op_33_eq = op_33_A == op_33_B;
wire op_33_ap_vld_A;
wire op_33_ap_vld_B;
wire clk_enable_A;
wire clk_enable_B;
assign clk_enable_A = _setup & (~op_33_ap_vld_A | op_33_ap_vld_B);
assign clk_enable_B = _setup;
wire divergent;
assign divergent = ~(ap_done_eq & ap_idle_eq & ap_ready_eq & op_33_eq);
assign unsafe_signal = op_33_ap_vld_A & op_33_ap_vld_B & divergent;
top_A instance_A (
    .ap_clk(ap_clk),
    .clk_enable(clk_enable_A),
    .ap_start(ap_start_internal),
    .op_0(op_0_internal),
    .op_10(op_10_internal),
    .op_11(op_11_internal),
    .op_12(op_12_internal),
    .op_13(op_13_internal),
    .op_15(op_15_internal),
    .op_16(op_16_internal),
    .op_17(op_17_internal),
    .op_18(op_18_internal),
    .op_19(op_19_internal),
    .op_3(op_3_internal),
    .op_4(op_4_internal),
    .op_5(op_5_internal),
    .op_6(op_6_internal),
    .op_7(op_7_internal),
    .op_9(op_9_internal),
    .ap_done(ap_done_A),
    .ap_idle(ap_idle_A),
    .ap_ready(ap_ready_A),
    .op_33(op_33_A),
    .op_33_ap_vld(op_33_ap_vld_A)
);
top_B instance_B (
    .ap_clk(ap_clk),
    .clk_enable(clk_enable_B),
    .ap_start(ap_start_internal),
    .op_0(op_0_internal),
    .op_10(op_10_internal),
    .op_11(op_11_internal),
    .op_12(op_12_internal),
    .op_13(op_13_internal),
    .op_15(op_15_internal),
    .op_16(op_16_internal),
    .op_17(op_17_internal),
    .op_18(op_18_internal),
    .op_19(op_19_internal),
    .op_3(op_3_internal),
    .op_4(op_4_internal),
    .op_5(op_5_internal),
    .op_6(op_6_internal),
    .op_7(op_7_internal),
    .op_9(op_9_internal),
    .ap_done(ap_done_B),
    .ap_idle(ap_idle_B),
    .ap_ready(ap_ready_B),
    .op_33(op_33_B),
    .op_33_ap_vld(op_33_ap_vld_B)
);
endmodule
