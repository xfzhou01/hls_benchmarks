// Processed by function `construct_kairos` in `verilog_tricks.py`.
// Machine A:
// Processed by function `add_clk_enable_signal` in `verilog_tricks.py`.
// Processed by function `remove_reset_signal` in `verilog_tricks.py`.
module top_A (
  ap_clk,
  ap_start,
  ap_done,
  ap_idle,
  ap_ready,
  op_0,
  op_1,
  op_7,
  op_8,
  op_9,
  op_19,
  op_27,
  op_27_ap_vld,
clk_enable
);
input clk_enable;


input ap_clk;
wire ap_rst;
assign ap_rst = op_27_ap_vld;
input ap_start;
input [3:0] op_0;
input [3:0] op_1;
input [15:0] op_19;
input [31:0] op_7;
input [3:0] op_8;
input [31:0] op_9;
output ap_done;
output ap_idle;
output ap_ready;
output [31:0] op_27;
output op_27_ap_vld;


reg [31:0] add_ln691_2_reg_1415;
reg [4:0] add_ln69_1_reg_1374;
reg [1:0] add_ln731_1_reg_1295;
reg and_ln785_1_reg_1250;
reg [7:0] ap_CS_fsm = 8'h01;
reg icmp_ln768_2_reg_1364;
reg icmp_ln786_2_reg_1311;
reg icmp_ln790_reg_1316;
reg icmp_ln850_reg_1354;
reg icmp_ln851_1_reg_1338;
reg icmp_ln851_2_reg_1399;
reg lhs_V_3_reg_1279;
reg newsignbit_reg_1240;
reg op_16_V_reg_1379;
reg [31:0] op_18_V_reg_1389;
reg [31:0] op_23_V_reg_1384;
reg [31:0] op_25_V_reg_1394;
reg op_2_V_reg_1268;
reg [3:0] op_4_V_reg_1255;
reg overflow_3_reg_1305;
reg p_Result_19_reg_1290;
reg p_Result_20_reg_1300;
reg [19:0] r_V_reg_1348;
reg [3:0] ret_V_11_reg_1273;
reg [31:0] ret_V_12_reg_1343;
reg [62:0] ret_V_15_reg_1326;
reg [31:0] ret_V_16_reg_1369;
reg [31:0] ret_V_18_cast_reg_1409;
reg [31:0] ret_V_7_cast_reg_1331;
reg [3:0] ret_V_reg_1321;
reg select_ln340_reg_1245;
reg [4:0] sext_ln1346_reg_1285;
reg [10:0] trunc_ln731_1_reg_1359;
reg [32:0] _142_;
wire [31:0] _000_;
wire [4:0] _001_;
wire [1:0] _002_;
wire _003_;
wire [7:0] _004_;
wire _005_;
wire _006_;
wire _007_;
wire _008_;
wire _009_;
wire _010_;
wire _011_;
wire _012_;
wire _013_;
wire [10:0] _014_;
wire [31:0] _015_;
wire [31:0] _016_;
wire _017_;
wire [3:0] _018_;
wire _019_;
wire _020_;
wire _021_;
wire [19:0] _022_;
wire [3:0] _023_;
wire [31:0] _024_;
wire [62:0] _025_;
wire [31:0] _026_;
wire [31:0] _027_;
wire [32:0] _028_;
wire [31:0] _029_;
wire [3:0] _030_;
wire _031_;
wire [4:0] _032_;
wire [10:0] _033_;
wire [1:0] _034_;
wire _035_;
wire _036_;
wire _037_;
wire _038_;
wire _039_;
wire _040_;
wire _041_;
wire _042_;
wire _043_;
wire _044_;
wire _045_;
wire _046_;
wire _047_;
wire _048_;
wire _049_;
wire _050_;
wire _051_;
wire _052_;
wire _053_;
wire _054_;
wire _055_;
wire _056_;
wire _057_;
wire _058_;
wire _059_;
wire _060_;
wire _061_;
wire [31:0] add_ln691_1_fu_960_p2;
wire [31:0] add_ln691_2_fu_1137_p2;
wire [31:0] add_ln691_3_fu_1212_p2;
wire [3:0] add_ln691_fu_745_p2;
wire [4:0] add_ln69_1_fu_982_p2;
wire [31:0] add_ln69_fu_1026_p2;
wire [1:0] add_ln731_1_fu_621_p2;
wire [10:0] add_ln731_fu_1042_p2;
wire and_ln340_1_fu_489_p2;
wire and_ln340_2_fu_541_p2;
wire and_ln340_fu_313_p2;
wire and_ln353_fu_1002_p2;
wire and_ln785_1_fu_351_p2;
wire and_ln785_3_fu_527_p2;
wire and_ln785_4_fu_547_p2;
wire and_ln785_fu_345_p2;
wire and_ln786_fu_509_p2;
wire ap_CS_fsm_state1;
wire ap_CS_fsm_state2;
wire ap_CS_fsm_state3;
wire ap_CS_fsm_state4;
wire ap_CS_fsm_state5;
wire ap_CS_fsm_state6;
wire ap_CS_fsm_state7;
wire ap_CS_fsm_state8;
wire [7:0] ap_NS_fsm;
wire ap_clk;
wire ap_done;
wire ap_idle;
wire ap_ready;
wire ap_rst;
wire ap_start;
wire icmp_ln1498_fu_879_p2;
wire icmp_ln768_1_fu_399_p2;
wire icmp_ln768_2_fu_939_p2;
wire icmp_ln768_3_fu_645_p2;
wire icmp_ln768_fu_237_p2;
wire icmp_ln786_1_fu_429_p2;
wire icmp_ln786_2_fu_669_p2;
wire icmp_ln786_fu_267_p2;
wire icmp_ln790_fu_687_p2;
wire icmp_ln850_fu_905_p2;
wire icmp_ln851_1_fu_850_p2;
wire icmp_ln851_2_fu_1101_p2;
wire icmp_ln851_3_fu_1206_p2;
wire icmp_ln851_fu_739_p2;
wire lhs_V_3_fu_585_p2;
wire [61:0] lhs_V_4_fu_814_p3;
wire [15:0] \mul_16ns_4s_20_1_1_U1.din0 ;
wire [3:0] \mul_16ns_4s_20_1_1_U1.din1 ;
wire [19:0] \mul_16ns_4s_20_1_1_U1.dout ;
wire [15:0] \mul_16ns_4s_20_1_1_U1.top_mul_16ns_4s_20_1_1_Multiplier_0_U.a ;
wire [3:0] \mul_16ns_4s_20_1_1_U1.top_mul_16ns_4s_20_1_1_Multiplier_0_U.b ;
wire [19:0] \mul_16ns_4s_20_1_1_U1.top_mul_16ns_4s_20_1_1_Multiplier_0_U.p ;
wire newsignbit_fu_215_p1;
wire [3:0] op_0;
wire [3:0] op_1;
wire [31:0] op_12_V_fu_806_p3;
wire [4:0] op_15_V_fu_948_p2;
wire [3:0] op_16_V_fu_1021_p1;
wire op_16_V_fu_1021_p2;
wire [31:0] op_18_V_fu_1068_p3;
wire [15:0] op_19;
wire [31:0] op_23_V_fu_1033_p2;
wire [31:0] op_25_V_fu_1091_p2;
wire [31:0] op_27;
wire op_27_ap_vld;
wire op_2_V_fu_573_p3;
wire [3:0] op_4_V_fu_565_p3;
wire [31:0] op_7;
wire [3:0] op_8;
wire [31:0] op_9;
wire or_ln340_1_fu_441_p2;
wire or_ln340_fu_279_p2;
wire or_ln384_fu_801_p2;
wire or_ln785_1_fu_405_p2;
wire or_ln785_2_fu_339_p2;
wire or_ln785_3_fu_651_p2;
wire or_ln785_4_fu_521_p2;
wire or_ln785_5_fu_553_p2;
wire or_ln785_fu_243_p2;
wire or_ln786_1_fu_435_p2;
wire or_ln786_fu_273_p2;
wire or_ln788_1_fu_784_p2;
wire or_ln788_fu_779_p2;
wire overflow_1_fu_417_p2;
wire overflow_2_fu_1063_p2;
wire overflow_3_fu_663_p2;
wire overflow_fu_255_p2;
wire p_Result_10_fu_953_p3;
wire p_Result_11_fu_1143_p3;
wire p_Result_12_fu_1194_p3;
wire p_Result_13_fu_207_p3;
wire p_Result_14_fu_219_p3;
wire [3:0] p_Result_15_fu_357_p1;
wire p_Result_15_fu_357_p3;
wire p_Result_16_fu_375_p2;
wire [3:0] p_Result_17_fu_381_p1;
wire p_Result_17_fu_381_p3;
wire p_Result_18_fu_1055_p3;
wire p_Result_19_fu_605_p3;
wire [3:0] p_Result_1_fu_389_p1;
wire [2:0] p_Result_1_fu_389_p4;
wire p_Result_20_fu_627_p3;
wire p_Result_3_fu_995_p3;
wire [21:0] p_Result_4_fu_929_p4;
wire p_Result_6_fu_727_p3;
wire [30:0] p_Result_8_fu_679_p3;
wire [3:0] p_Result_s_16_fu_473_p4;
wire [3:0] p_Result_s_fu_227_p4;
wire [31:0] p_Val2_11_fu_767_p3;
wire p_Val2_1_fu_261_p2;
wire [3:0] p_Val2_2_fu_369_p0;
wire [3:0] p_Val2_2_fu_369_p2;
wire [2:0] p_Val2_3_fu_467_p2;
wire [31:0] p_Val2_7_fu_1047_p3;
wire [15:0] r_V_fu_895_p0;
wire [19:0] r_V_fu_895_p00;
wire [19:0] r_V_fu_895_p2;
wire [32:0] ret_1_fu_919_p2;
wire [4:0] ret_2_fu_599_p2;
wire [3:0] ret_V_11_fu_578_p2;
wire [3:0] ret_V_11_fu_578_p3;
wire [31:0] ret_V_12_fu_863_p2;
wire ret_V_13_fu_1007_p2;
wire [4:0] ret_V_14_fu_707_p2;
wire [62:0] ret_V_15_fu_830_p2;
wire [31:0] ret_V_16_fu_971_p3;
wire [31:0] ret_V_17_fu_1083_p2;
wire [31:0] ret_V_18_cast_fu_1127_p4;
wire [53:0] ret_V_18_fu_1121_p2;
wire [53:0] ret_V_18_reg_1404;
wire [46:0] ret_V_19_fu_1178_p2;
wire [31:0] ret_V_20_cast_fu_1184_p4;
wire [3:0] ret_V_fu_759_p3;
wire [4:0] ret_fu_201_p2;
wire [2:0] rhs_1_fu_696_p3;
wire [52:0] rhs_4_fu_1110_p3;
wire [45:0] rhs_5_fu_1166_p3;
wire sel_tmp18_fu_559_p2;
wire [31:0] select_ln1192_1_fu_1076_p3;
wire [31:0] select_ln1192_fu_856_p3;
wire [3:0] select_ln340_1_fu_495_p3;
wire select_ln340_fu_319_p3;
wire [31:0] select_ln353_fu_1159_p3;
wire select_ln365_fu_299_p3;
wire [31:0] select_ln384_fu_794_p3;
wire [3:0] select_ln785_fu_533_p3;
wire [31:0] select_ln850_1_fu_965_p3;
wire [31:0] select_ln850_2_fu_1154_p3;
wire [31:0] select_ln850_3_fu_1218_p3;
wire [3:0] select_ln850_fu_751_p3;
wire [3:0] select_ln874_fu_1013_p3;
wire [15:0] sext_ln1118_fu_888_p1;
wire [53:0] sext_ln1192_1_fu_1117_p1;
wire [46:0] sext_ln1192_2_fu_1174_p1;
wire [62:0] sext_ln1192_fu_822_p1;
wire [4:0] sext_ln1193_fu_693_p1;
wire [3:0] sext_ln1346_fu_595_p0;
wire [4:0] sext_ln1346_fu_595_p1;
wire [3:0] sext_ln1347_fu_197_p0;
wire [4:0] sext_ln1347_fu_197_p1;
wire [4:0] sext_ln215_fu_193_p1;
wire [31:0] sext_ln69_fu_1030_p1;
wire [15:0] sext_ln703_1_fu_1150_p0;
wire [46:0] sext_ln703_1_fu_1150_p1;
wire [62:0] sext_ln703_fu_826_p1;
wire [5:0] sext_ln727_fu_869_p1;
wire [10:0] sext_ln731_fu_1039_p1;
wire [4:0] sext_ln831_fu_945_p1;
wire [3:0] sext_ln850_fu_723_p1;
wire [3:0] shl_ln_fu_872_p1;
wire [5:0] shl_ln_fu_872_p3;
wire [2:0] tmp_2_fu_713_p4;
wire [2:0] tmp_3_fu_635_p4;
wire [3:0] tmp_5_fu_447_p1;
wire tmp_5_fu_447_p3;
wire tmp_7_fu_988_p3;
wire tmp_fu_285_p3;
wire [10:0] trunc_ln731_1_fu_925_p1;
wire [3:0] trunc_ln731_2_fu_613_p0;
wire [1:0] trunc_ln731_2_fu_613_p1;
wire [3:0] trunc_ln731_fu_365_p0;
wire trunc_ln731_fu_365_p1;
wire trunc_ln790_fu_675_p1;
wire [1:0] trunc_ln851_1_fu_735_p1;
wire [29:0] trunc_ln851_2_fu_846_p1;
wire [20:0] trunc_ln851_3_fu_1097_p1;
wire [15:0] trunc_ln851_4_fu_1202_p0;
wire [13:0] trunc_ln851_4_fu_1202_p1;
wire [1:0] trunc_ln851_fu_901_p1;
wire underflow_2_fu_789_p2;
wire xor_ln340_1_fu_483_p2;
wire xor_ln340_fu_307_p2;
wire xor_ln365_1_fu_455_p2;
wire xor_ln365_2_fu_461_p2;
wire xor_ln365_fu_293_p2;
wire xor_ln785_1_fu_411_p2;
wire xor_ln785_2_fu_657_p2;
wire xor_ln785_3_fu_333_p2;
wire xor_ln785_4_fu_515_p2;
wire xor_ln785_fu_249_p2;
wire xor_ln786_1_fu_774_p2;
wire xor_ln786_3_fu_327_p2;
wire xor_ln786_4_fu_503_p2;
wire xor_ln786_fu_423_p2;
wire [4:0] zext_ln1193_fu_703_p1;
wire [4:0] zext_ln1346_fu_591_p1;
wire [32:0] zext_ln215_1_fu_915_p1;
wire [32:0] zext_ln215_fu_911_p1;
wire [31:0] zext_ln69_1_fu_1088_p1;
wire [4:0] zext_ln69_fu_978_p1;
wire [53:0] zext_ln703_fu_1107_p1;
wire [1:0] zext_ln731_fu_617_p1;


assign add_ln691_1_fu_960_p2 = ret_V_7_cast_reg_1331 + 1'h1;
assign add_ln691_2_fu_1137_p2 = ret_V_18_fu_1121_p2[52:21] + 1'h1;
assign add_ln691_3_fu_1212_p2 = ret_V_19_fu_1178_p2[45:14] + 1'h1;
assign add_ln691_fu_745_p2 = $signed(ret_V_14_fu_707_p2[4:2]) + $signed(2'h1);
assign add_ln69_1_fu_982_p2 = op_15_V_fu_948_p2 + icmp_ln1498_fu_879_p2;
assign add_ln69_fu_1026_p2 = ret_V_12_reg_1343 + ret_V_16_reg_1369;
assign add_ln731_1_fu_621_p2 = op_8[1:0] + lhs_V_3_fu_585_p2;
assign add_ln731_fu_1042_p2 = $signed(trunc_ln731_1_reg_1359) + $signed(ret_V_11_reg_1273);
assign op_23_V_fu_1033_p2 = $signed(add_ln69_1_reg_1374) + $signed(add_ln69_fu_1026_p2);
assign op_25_V_fu_1091_p2 = ret_V_17_fu_1083_p2 + lhs_V_3_reg_1279;
assign ret_1_fu_919_p2 = op_9 + { ret_V_11_reg_1273[3], ret_V_11_reg_1273[3], ret_V_11_reg_1273[3], ret_V_11_reg_1273[3], ret_V_11_reg_1273[3], ret_V_11_reg_1273[3], ret_V_11_reg_1273[3], ret_V_11_reg_1273[3], ret_V_11_reg_1273[3], ret_V_11_reg_1273[3], ret_V_11_reg_1273[3], ret_V_11_reg_1273[3], ret_V_11_reg_1273 };
assign ret_2_fu_599_p2 = $signed(op_8) + $signed({ 1'h0, lhs_V_3_fu_585_p2 });
assign ret_V_12_fu_863_p2 = select_ln1192_fu_856_p3 + op_9;
assign ret_V_15_fu_830_p2 = $signed({ op_7, 30'h00000000 }) + $signed(op_12_V_fu_806_p3);
assign ret_V_17_fu_1083_p2 = op_23_V_reg_1384 + select_ln1192_1_fu_1076_p3;
assign ret_V_18_fu_1121_p2 = $signed({ op_25_V_reg_1394, 21'h000000 }) + $signed({ 1'h0, op_18_V_reg_1389 });
assign ret_V_19_fu_1178_p2 = $signed({ select_ln353_fu_1159_p3, 14'h0000 }) + $signed(op_19);
assign _035_ = ap_CS_fsm[6] & icmp_ln851_2_reg_1399;
assign _036_ = ap_CS_fsm[0] & _038_;
assign _037_ = ap_CS_fsm[0] & ap_start;
assign and_ln340_1_fu_489_p2 = xor_ln340_1_fu_483_p2 & or_ln786_1_fu_435_p2;
assign and_ln340_2_fu_541_p2 = or_ln786_1_fu_435_p2 & or_ln340_1_fu_441_p2;
assign and_ln340_fu_313_p2 = xor_ln340_fu_307_p2 & or_ln786_fu_273_p2;
assign and_ln353_fu_1002_p2 = r_V_reg_1348[19] & icmp_ln850_reg_1354;
assign and_ln785_1_fu_351_p2 = ret_fu_201_p2[0] & and_ln785_fu_345_p2;
assign and_ln785_3_fu_527_p2 = or_ln785_4_fu_521_p2 & and_ln786_fu_509_p2;
assign and_ln785_4_fu_547_p2 = xor_ln785_1_fu_411_p2 & and_ln786_fu_509_p2;
assign and_ln785_fu_345_p2 = xor_ln786_3_fu_327_p2 & or_ln785_2_fu_339_p2;
assign and_ln786_fu_509_p2 = xor_ln786_4_fu_503_p2 & p_Result_16_fu_375_p2;
assign overflow_1_fu_417_p2 = xor_ln785_1_fu_411_p2 & or_ln785_1_fu_405_p2;
assign overflow_3_fu_663_p2 = xor_ln785_2_fu_657_p2 & or_ln785_3_fu_651_p2;
assign overflow_fu_255_p2 = xor_ln785_fu_249_p2 & or_ln785_fu_243_p2;
assign sel_tmp18_fu_559_p2 = xor_ln365_2_fu_461_p2 & or_ln785_5_fu_553_p2;
assign underflow_2_fu_789_p2 = p_Result_19_reg_1290 & or_ln788_1_fu_784_p2;
assign lhs_V_3_fu_585_p2 = ~ op_2_V_fu_573_p3;
assign xor_ln786_fu_423_p2 = ~ p_Result_16_fu_375_p2;
assign xor_ln785_1_fu_411_p2 = ~ op_1[3];
assign xor_ln340_1_fu_483_p2 = ~ or_ln340_1_fu_441_p2;
assign p_Val2_1_fu_261_p2 = ~ ret_fu_201_p2[0];
assign xor_ln785_fu_249_p2 = ~ ret_fu_201_p2[4];
assign xor_ln340_fu_307_p2 = ~ or_ln340_fu_279_p2;
assign xor_ln785_3_fu_333_p2 = ~ or_ln785_fu_243_p2;
assign xor_ln786_3_fu_327_p2 = ~ icmp_ln786_fu_267_p2;
assign xor_ln786_4_fu_503_p2 = ~ icmp_ln786_1_fu_429_p2;
assign xor_ln785_4_fu_515_p2 = ~ or_ln785_1_fu_405_p2;
assign xor_ln786_1_fu_774_p2 = ~ p_Result_20_reg_1300;
assign xor_ln365_2_fu_461_p2 = ~ xor_ln365_1_fu_455_p2;
assign xor_ln785_2_fu_657_p2 = ~ ret_2_fu_599_p2[4];
assign _038_ = ~ ap_start;
assign _039_ = { op_4_V_reg_1255[3], op_4_V_reg_1255[3], op_4_V_reg_1255 } == { op_8, 2'h0 };
assign _040_ = ! { add_ln731_1_fu_621_p2[0], 30'h00000000 };
assign \mul_16ns_4s_20_1_1_U1.top_mul_16ns_4s_20_1_1_Multiplier_0_U.p  = $signed({ 1'h0, \mul_16ns_4s_20_1_1_U1.top_mul_16ns_4s_20_1_1_Multiplier_0_U.a  }) * $signed(\mul_16ns_4s_20_1_1_U1.top_mul_16ns_4s_20_1_1_Multiplier_0_U.b );
assign _041_ = | op_1[3:1];
assign _042_ = | ret_1_fu_919_p2[32:11];
assign _043_ = | ret_2_fu_599_p2[4:2];
assign _044_ = | ret_fu_201_p2[4:1];
assign _045_ = op_1[3:1] != 3'h7;
assign _046_ = ret_2_fu_599_p2[4:2] != 3'h7;
assign _047_ = ret_fu_201_p2[4:1] != 4'hf;
assign _048_ = | r_V_fu_895_p2[1:0];
assign _049_ = | op_12_V_fu_806_p3[29:0];
assign _050_ = | op_18_V_fu_1068_p3[20:0];
assign _051_ = | op_19[13:0];
assign _052_ = | ret_V_14_fu_707_p2[1:0];
assign _053_ = select_ln874_fu_1013_p3 != op_8;
assign or_ln340_1_fu_441_p2 = op_1[3] | overflow_1_fu_417_p2;
assign or_ln340_fu_279_p2 = ret_fu_201_p2[4] | overflow_fu_255_p2;
assign or_ln384_fu_801_p2 = underflow_2_fu_789_p2 | overflow_3_reg_1305;
assign or_ln785_1_fu_405_p2 = p_Result_16_fu_375_p2 | icmp_ln768_1_fu_399_p2;
assign or_ln785_2_fu_339_p2 = xor_ln785_3_fu_333_p2 | ret_fu_201_p2[4];
assign or_ln785_3_fu_651_p2 = add_ln731_1_fu_621_p2[1] | icmp_ln768_3_fu_645_p2;
assign or_ln785_4_fu_521_p2 = xor_ln785_4_fu_515_p2 | op_1[3];
assign or_ln785_5_fu_553_p2 = and_ln785_4_fu_547_p2 | and_ln340_2_fu_541_p2;
assign or_ln785_fu_243_p2 = ret_fu_201_p2[0] | icmp_ln768_fu_237_p2;
assign or_ln786_1_fu_435_p2 = xor_ln786_fu_423_p2 | icmp_ln786_1_fu_429_p2;
assign or_ln786_fu_273_p2 = p_Val2_1_fu_261_p2 | icmp_ln786_fu_267_p2;
assign or_ln788_1_fu_784_p2 = or_ln788_fu_779_p2 | icmp_ln786_2_reg_1311;
assign or_ln788_fu_779_p2 = xor_ln786_1_fu_774_p2 | icmp_ln790_reg_1316;
assign overflow_2_fu_1063_p2 = add_ln731_fu_1042_p2[10] | icmp_ln768_2_reg_1364;
always @(posedge ap_clk)
op_18_V_reg_1389[20:0] <= 21'h000000;
always @(posedge ap_clk)
_142_ <= _028_;
assign ret_V_18_reg_1404[53:21] = _142_;
always @(posedge ap_clk)
ret_V_18_cast_reg_1409 <= _027_;
always @(posedge ap_clk)
op_16_V_reg_1379 <= _013_;
always @(posedge ap_clk)
op_23_V_reg_1384 <= _015_;
always @(posedge ap_clk)
op_18_V_reg_1389[31:21] <= _014_;
always @(posedge ap_clk)
op_25_V_reg_1394 <= _016_;
always @(posedge ap_clk)
icmp_ln851_2_reg_1399 <= _010_;
always @(posedge ap_clk)
ret_V_reg_1321 <= _030_;
always @(posedge ap_clk)
ret_V_15_reg_1326 <= _025_;
always @(posedge ap_clk)
ret_V_7_cast_reg_1331 <= _029_;
always @(posedge ap_clk)
icmp_ln851_1_reg_1338 <= _009_;
always @(posedge ap_clk)
newsignbit_reg_1240 <= _012_;
always @(posedge ap_clk)
select_ln340_reg_1245 <= _031_;
always @(posedge ap_clk)
and_ln785_1_reg_1250 <= _003_;
always @(posedge ap_clk)
op_4_V_reg_1255 <= _018_;
always @(posedge ap_clk)
op_2_V_reg_1268 <= _017_;
always @(posedge ap_clk)
ret_V_11_reg_1273 <= _023_;
always @(posedge ap_clk)
lhs_V_3_reg_1279 <= _011_;
always @(posedge ap_clk)
sext_ln1346_reg_1285 <= _032_;
always @(posedge ap_clk)
p_Result_19_reg_1290 <= _020_;
always @(posedge ap_clk)
add_ln731_1_reg_1295 <= _002_;
always @(posedge ap_clk)
p_Result_20_reg_1300 <= _021_;
always @(posedge ap_clk)
overflow_3_reg_1305 <= _019_;
always @(posedge ap_clk)
icmp_ln786_2_reg_1311 <= _006_;
always @(posedge ap_clk)
icmp_ln790_reg_1316 <= _007_;
always @(posedge ap_clk)
ret_V_12_reg_1343 <= _024_;
always @(posedge ap_clk)
r_V_reg_1348 <= _022_;
always @(posedge ap_clk)
icmp_ln850_reg_1354 <= _008_;
always @(posedge ap_clk)
trunc_ln731_1_reg_1359 <= _033_;
always @(posedge ap_clk)
icmp_ln768_2_reg_1364 <= _005_;
always @(posedge ap_clk)
ret_V_16_reg_1369 <= _026_;
always @(posedge ap_clk)
add_ln69_1_reg_1374 <= _001_;
always @(posedge ap_clk)
add_ln691_2_reg_1415 <= _000_;
always @(posedge ap_clk)
ap_CS_fsm <= _004_;
assign _034_ = _037_ ? 2'h2 : 2'h1;
assign _054_ = ap_CS_fsm == 1'h1;
function [7:0] _178_;
input [7:0] a;
input [63:0] b;
input [7:0] s;
case (s)
8'b00000001:
_178_ = b[7:0];
8'b00000010:
_178_ = b[15:8];
8'b00000100:
_178_ = b[23:16];
8'b00001000:
_178_ = b[31:24];
8'b00010000:
_178_ = b[39:32];
8'b00100000:
_178_ = b[47:40];
8'b01000000:
_178_ = b[55:48];
8'b10000000:
_178_ = b[63:56];
8'b00000000:
_178_ = a;
default:
_178_ = 8'bx;
endcase
endfunction
assign ap_NS_fsm = _178_(8'hxx, { 6'h00, _034_, 56'h04081020408001 }, { _054_, _061_, _060_, _059_, _058_, _057_, _056_, _055_ });
assign _055_ = ap_CS_fsm == 8'h80;
assign _056_ = ap_CS_fsm == 7'h40;
assign _057_ = ap_CS_fsm == 6'h20;
assign _058_ = ap_CS_fsm == 5'h10;
assign _059_ = ap_CS_fsm == 4'h8;
assign _060_ = ap_CS_fsm == 3'h4;
assign _061_ = ap_CS_fsm == 2'h2;
assign op_27_ap_vld = ap_CS_fsm[7] ? 1'h1 : 1'h0;
assign ap_idle = _036_ ? 1'h1 : 1'h0;
assign _027_ = ap_CS_fsm[6] ? ret_V_18_fu_1121_p2[52:21] : ret_V_18_cast_reg_1409;
assign _028_ = ap_CS_fsm[6] ? ret_V_18_fu_1121_p2[53:21] : ret_V_18_reg_1404[53:21];
assign _015_ = ap_CS_fsm[4] ? op_23_V_fu_1033_p2 : op_23_V_reg_1384;
assign _013_ = ap_CS_fsm[4] ? op_16_V_fu_1021_p2 : op_16_V_reg_1379;
assign _010_ = ap_CS_fsm[5] ? icmp_ln851_2_fu_1101_p2 : icmp_ln851_2_reg_1399;
assign _016_ = ap_CS_fsm[5] ? op_25_V_fu_1091_p2 : op_25_V_reg_1394;
assign _014_ = ap_CS_fsm[5] ? op_18_V_fu_1068_p3[31:21] : op_18_V_reg_1389[31:21];
assign _009_ = ap_CS_fsm[2] ? icmp_ln851_1_fu_850_p2 : icmp_ln851_1_reg_1338;
assign _029_ = ap_CS_fsm[2] ? ret_V_15_fu_830_p2[61:30] : ret_V_7_cast_reg_1331;
assign _025_ = ap_CS_fsm[2] ? ret_V_15_fu_830_p2 : ret_V_15_reg_1326;
assign _030_ = ap_CS_fsm[2] ? ret_V_fu_759_p3 : ret_V_reg_1321;
assign _018_ = ap_CS_fsm[0] ? op_4_V_fu_565_p3 : op_4_V_reg_1255;
assign _003_ = ap_CS_fsm[0] ? and_ln785_1_fu_351_p2 : and_ln785_1_reg_1250;
assign _031_ = ap_CS_fsm[0] ? select_ln340_fu_319_p3 : select_ln340_reg_1245;
assign _012_ = ap_CS_fsm[0] ? ret_fu_201_p2[0] : newsignbit_reg_1240;
assign _007_ = ap_CS_fsm[1] ? icmp_ln790_fu_687_p2 : icmp_ln790_reg_1316;
assign _006_ = ap_CS_fsm[1] ? icmp_ln786_2_fu_669_p2 : icmp_ln786_2_reg_1311;
assign _019_ = ap_CS_fsm[1] ? overflow_3_fu_663_p2 : overflow_3_reg_1305;
assign _021_ = ap_CS_fsm[1] ? add_ln731_1_fu_621_p2[1] : p_Result_20_reg_1300;
assign _002_ = ap_CS_fsm[1] ? add_ln731_1_fu_621_p2 : add_ln731_1_reg_1295;
assign _020_ = ap_CS_fsm[1] ? ret_2_fu_599_p2[4] : p_Result_19_reg_1290;
assign _032_ = ap_CS_fsm[1] ? { op_8[3], op_8 } : sext_ln1346_reg_1285;
assign _011_ = ap_CS_fsm[1] ? lhs_V_3_fu_585_p2 : lhs_V_3_reg_1279;
assign _023_ = ap_CS_fsm[1] ? ret_V_11_fu_578_p3 : ret_V_11_reg_1273;
assign _017_ = ap_CS_fsm[1] ? op_2_V_fu_573_p3 : op_2_V_reg_1268;
assign _001_ = ap_CS_fsm[3] ? add_ln69_1_fu_982_p2 : add_ln69_1_reg_1374;
assign _026_ = ap_CS_fsm[3] ? ret_V_16_fu_971_p3 : ret_V_16_reg_1369;
assign _005_ = ap_CS_fsm[3] ? icmp_ln768_2_fu_939_p2 : icmp_ln768_2_reg_1364;
assign _033_ = ap_CS_fsm[3] ? op_9[10:0] : trunc_ln731_1_reg_1359;
assign _008_ = ap_CS_fsm[3] ? icmp_ln850_fu_905_p2 : icmp_ln850_reg_1354;
assign _022_ = ap_CS_fsm[3] ? r_V_fu_895_p2 : r_V_reg_1348;
assign _024_ = ap_CS_fsm[3] ? ret_V_12_fu_863_p2 : ret_V_12_reg_1343;
assign _000_ = _035_ ? add_ln691_2_fu_1137_p2 : add_ln691_2_reg_1415;
assign _004_ = ap_rst ? 8'h01 : ap_NS_fsm;
assign op_15_V_fu_948_p2 = $signed(sext_ln1346_reg_1285) - $signed(ret_V_reg_1321);
assign ret_V_14_fu_707_p2 = $signed(op_4_V_reg_1255) - $signed({ 1'h0, lhs_V_3_reg_1279, 2'h0 });
assign ret_fu_201_p2 = $signed(op_0) - $signed(op_1);
assign icmp_ln1498_fu_879_p2 = _039_ ? 1'h1 : 1'h0;
assign icmp_ln768_1_fu_399_p2 = _041_ ? 1'h1 : 1'h0;
assign icmp_ln768_2_fu_939_p2 = _042_ ? 1'h1 : 1'h0;
assign icmp_ln768_3_fu_645_p2 = _043_ ? 1'h1 : 1'h0;
assign icmp_ln768_fu_237_p2 = _044_ ? 1'h1 : 1'h0;
assign icmp_ln786_1_fu_429_p2 = _045_ ? 1'h1 : 1'h0;
assign icmp_ln786_2_fu_669_p2 = _046_ ? 1'h1 : 1'h0;
assign icmp_ln786_fu_267_p2 = _047_ ? 1'h1 : 1'h0;
assign icmp_ln790_fu_687_p2 = _040_ ? 1'h1 : 1'h0;
assign icmp_ln850_fu_905_p2 = _048_ ? 1'h1 : 1'h0;
assign icmp_ln851_1_fu_850_p2 = _049_ ? 1'h1 : 1'h0;
assign icmp_ln851_2_fu_1101_p2 = _050_ ? 1'h1 : 1'h0;
assign icmp_ln851_3_fu_1206_p2 = _051_ ? 1'h1 : 1'h0;
assign icmp_ln851_fu_739_p2 = _052_ ? 1'h1 : 1'h0;
assign op_12_V_fu_806_p3 = or_ln384_fu_801_p2 ? select_ln384_fu_794_p3 : { add_ln731_1_reg_1295, 30'h00000000 };
assign op_16_V_fu_1021_p2 = _053_ ? 1'h1 : 1'h0;
assign op_18_V_fu_1068_p3 = overflow_2_fu_1063_p2 ? 32'd0 : { add_ln731_fu_1042_p2, 21'h000000 };
assign op_27 = ret_V_19_fu_1178_p2[46] ? select_ln850_3_fu_1218_p3 : ret_V_19_fu_1178_p2[45:14];
assign op_2_V_fu_573_p3 = and_ln785_1_reg_1250 ? newsignbit_reg_1240 : select_ln340_reg_1245;
assign op_4_V_fu_565_p3 = sel_tmp18_fu_559_p2 ? { op_1[0], 3'h0 } : select_ln785_fu_533_p3;
assign p_Result_16_fu_375_p2 = op_1[0] ? 1'h1 : 1'h0;
assign ret_V_11_fu_578_p3 = op_2_V_fu_573_p3 ? 4'hf : op_1;
assign ret_V_16_fu_971_p3 = ret_V_15_reg_1326[62] ? select_ln850_1_fu_965_p3 : ret_V_7_cast_reg_1331;
assign ret_V_fu_759_p3 = ret_V_14_fu_707_p2[4] ? select_ln850_fu_751_p3 : { 2'h0, ret_V_14_fu_707_p2[3:2] };
assign select_ln1192_1_fu_1076_p3 = op_16_V_reg_1379 ? 32'd4294967295 : 32'd0;
assign select_ln1192_fu_856_p3 = op_2_V_reg_1268 ? 32'd4294967295 : 32'd0;
assign select_ln340_1_fu_495_p3 = and_ln340_1_fu_489_p2 ? { op_1[0], 3'h0 } : { op_1[1], 3'h7 };
assign select_ln340_fu_319_p3 = and_ln340_fu_313_p2 ? ret_fu_201_p2[0] : select_ln365_fu_299_p3;
assign select_ln353_fu_1159_p3 = ret_V_18_reg_1404[53] ? select_ln850_2_fu_1154_p3 : ret_V_18_cast_reg_1409;
assign select_ln365_fu_299_p3 = xor_ln365_fu_293_p2 ? ret_fu_201_p2[1] : ret_fu_201_p2[0];
assign select_ln384_fu_794_p3 = overflow_3_reg_1305 ? 32'd2147483647 : 32'd2147483649;
assign select_ln785_fu_533_p3 = and_ln785_3_fu_527_p2 ? { op_1[0], 3'h0 } : select_ln340_1_fu_495_p3;
assign select_ln850_1_fu_965_p3 = icmp_ln851_1_reg_1338 ? add_ln691_1_fu_960_p2 : ret_V_7_cast_reg_1331;
assign select_ln850_2_fu_1154_p3 = icmp_ln851_2_reg_1399 ? add_ln691_2_reg_1415 : ret_V_18_cast_reg_1409;
assign select_ln850_3_fu_1218_p3 = icmp_ln851_3_fu_1206_p2 ? add_ln691_3_fu_1212_p2 : ret_V_19_fu_1178_p2[45:14];
assign select_ln850_fu_751_p3 = icmp_ln851_fu_739_p2 ? add_ln691_fu_745_p2 : { 2'h3, ret_V_14_fu_707_p2[3:2] };
assign select_ln874_fu_1013_p3 = ret_V_13_fu_1007_p2 ? 4'hf : 4'h0;
assign ret_V_13_fu_1007_p2 = r_V_reg_1348[2] ^ and_ln353_fu_1002_p2;
assign xor_ln365_1_fu_455_p2 = op_1[0] ^ op_1[1];
assign xor_ln365_fu_293_p2 = ret_fu_201_p2[1] ^ ret_fu_201_p2[0];
assign ap_CS_fsm_state1 = ap_CS_fsm[0];
assign ap_CS_fsm_state2 = ap_CS_fsm[1];
assign ap_CS_fsm_state3 = ap_CS_fsm[2];
assign ap_CS_fsm_state4 = ap_CS_fsm[3];
assign ap_CS_fsm_state5 = ap_CS_fsm[4];
assign ap_CS_fsm_state6 = ap_CS_fsm[5];
assign ap_CS_fsm_state7 = ap_CS_fsm[6];
assign ap_CS_fsm_state8 = ap_CS_fsm[7];
assign ap_done = op_27_ap_vld;
assign ap_ready = op_27_ap_vld;
assign lhs_V_4_fu_814_p3 = { op_7, 30'h00000000 };
assign newsignbit_fu_215_p1 = ret_fu_201_p2[0];
assign op_16_V_fu_1021_p1 = op_8;
assign p_Result_10_fu_953_p3 = ret_V_15_reg_1326[62];
assign p_Result_11_fu_1143_p3 = ret_V_18_reg_1404[53];
assign p_Result_12_fu_1194_p3 = ret_V_19_fu_1178_p2[46];
assign p_Result_13_fu_207_p3 = ret_fu_201_p2[4];
assign p_Result_14_fu_219_p3 = ret_fu_201_p2[1];
assign p_Result_15_fu_357_p1 = op_1;
assign p_Result_15_fu_357_p3 = op_1[3];
assign p_Result_17_fu_381_p1 = op_1;
assign p_Result_17_fu_381_p3 = op_1[1];
assign p_Result_18_fu_1055_p3 = add_ln731_fu_1042_p2[10];
assign p_Result_19_fu_605_p3 = ret_2_fu_599_p2[4];
assign p_Result_1_fu_389_p1 = op_1;
assign p_Result_1_fu_389_p4 = op_1[3:1];
assign p_Result_20_fu_627_p3 = add_ln731_1_fu_621_p2[1];
assign p_Result_3_fu_995_p3 = r_V_reg_1348[19];
assign p_Result_4_fu_929_p4 = ret_1_fu_919_p2[32:11];
assign p_Result_6_fu_727_p3 = ret_V_14_fu_707_p2[4];
assign p_Result_8_fu_679_p3 = { add_ln731_1_fu_621_p2[0], 30'h00000000 };
assign p_Result_s_16_fu_473_p4 = { op_1[1], 3'h7 };
assign p_Result_s_fu_227_p4 = ret_fu_201_p2[4:1];
assign p_Val2_11_fu_767_p3 = { add_ln731_1_reg_1295, 30'h00000000 };
assign p_Val2_2_fu_369_p0 = op_1;
assign p_Val2_2_fu_369_p2 = { op_1[0], 3'h0 };
assign p_Val2_3_fu_467_p2 = 3'h7;
assign p_Val2_7_fu_1047_p3 = { add_ln731_fu_1042_p2, 21'h000000 };
assign r_V_fu_895_p0 = { ret_V_11_reg_1273[3], ret_V_11_reg_1273[3], ret_V_11_reg_1273[3], ret_V_11_reg_1273[3], ret_V_11_reg_1273[3], ret_V_11_reg_1273[3], ret_V_11_reg_1273[3], ret_V_11_reg_1273[3], ret_V_11_reg_1273[3], ret_V_11_reg_1273[3], ret_V_11_reg_1273[3], ret_V_11_reg_1273[3], ret_V_11_reg_1273 };
assign r_V_fu_895_p00 = { 4'h0, ret_V_11_reg_1273[3], ret_V_11_reg_1273[3], ret_V_11_reg_1273[3], ret_V_11_reg_1273[3], ret_V_11_reg_1273[3], ret_V_11_reg_1273[3], ret_V_11_reg_1273[3], ret_V_11_reg_1273[3], ret_V_11_reg_1273[3], ret_V_11_reg_1273[3], ret_V_11_reg_1273[3], ret_V_11_reg_1273[3], ret_V_11_reg_1273 };
assign ret_V_11_fu_578_p2 = op_1;
assign ret_V_18_cast_fu_1127_p4 = ret_V_18_fu_1121_p2[52:21];
assign ret_V_20_cast_fu_1184_p4 = ret_V_19_fu_1178_p2[45:14];
assign rhs_1_fu_696_p3 = { lhs_V_3_reg_1279, 2'h0 };
assign rhs_4_fu_1110_p3 = { op_25_V_reg_1394, 21'h000000 };
assign rhs_5_fu_1166_p3 = { select_ln353_fu_1159_p3, 14'h0000 };
assign sext_ln1118_fu_888_p1 = { ret_V_11_reg_1273[3], ret_V_11_reg_1273[3], ret_V_11_reg_1273[3], ret_V_11_reg_1273[3], ret_V_11_reg_1273[3], ret_V_11_reg_1273[3], ret_V_11_reg_1273[3], ret_V_11_reg_1273[3], ret_V_11_reg_1273[3], ret_V_11_reg_1273[3], ret_V_11_reg_1273[3], ret_V_11_reg_1273[3], ret_V_11_reg_1273 };
assign sext_ln1192_1_fu_1117_p1 = { op_25_V_reg_1394[31], op_25_V_reg_1394, 21'h000000 };
assign sext_ln1192_2_fu_1174_p1 = { select_ln353_fu_1159_p3[31], select_ln353_fu_1159_p3, 14'h0000 };
assign sext_ln1192_fu_822_p1 = { op_7[31], op_7, 30'h00000000 };
assign sext_ln1193_fu_693_p1 = { op_4_V_reg_1255[3], op_4_V_reg_1255 };
assign sext_ln1346_fu_595_p0 = op_8;
assign sext_ln1346_fu_595_p1 = { op_8[3], op_8 };
assign sext_ln1347_fu_197_p0 = op_1;
assign sext_ln1347_fu_197_p1 = { op_1[3], op_1 };
assign sext_ln215_fu_193_p1 = { op_0[3], op_0 };
assign sext_ln69_fu_1030_p1 = { add_ln69_1_reg_1374[4], add_ln69_1_reg_1374[4], add_ln69_1_reg_1374[4], add_ln69_1_reg_1374[4], add_ln69_1_reg_1374[4], add_ln69_1_reg_1374[4], add_ln69_1_reg_1374[4], add_ln69_1_reg_1374[4], add_ln69_1_reg_1374[4], add_ln69_1_reg_1374[4], add_ln69_1_reg_1374[4], add_ln69_1_reg_1374[4], add_ln69_1_reg_1374[4], add_ln69_1_reg_1374[4], add_ln69_1_reg_1374[4], add_ln69_1_reg_1374[4], add_ln69_1_reg_1374[4], add_ln69_1_reg_1374[4], add_ln69_1_reg_1374[4], add_ln69_1_reg_1374[4], add_ln69_1_reg_1374[4], add_ln69_1_reg_1374[4], add_ln69_1_reg_1374[4], add_ln69_1_reg_1374[4], add_ln69_1_reg_1374[4], add_ln69_1_reg_1374[4], add_ln69_1_reg_1374[4], add_ln69_1_reg_1374 };
assign sext_ln703_1_fu_1150_p0 = op_19;
assign sext_ln703_1_fu_1150_p1 = { op_19[15], op_19[15], op_19[15], op_19[15], op_19[15], op_19[15], op_19[15], op_19[15], op_19[15], op_19[15], op_19[15], op_19[15], op_19[15], op_19[15], op_19[15], op_19[15], op_19[15], op_19[15], op_19[15], op_19[15], op_19[15], op_19[15], op_19[15], op_19[15], op_19[15], op_19[15], op_19[15], op_19[15], op_19[15], op_19[15], op_19[15], op_19 };
assign sext_ln703_fu_826_p1 = { op_12_V_fu_806_p3[31], op_12_V_fu_806_p3[31], op_12_V_fu_806_p3[31], op_12_V_fu_806_p3[31], op_12_V_fu_806_p3[31], op_12_V_fu_806_p3[31], op_12_V_fu_806_p3[31], op_12_V_fu_806_p3[31], op_12_V_fu_806_p3[31], op_12_V_fu_806_p3[31], op_12_V_fu_806_p3[31], op_12_V_fu_806_p3[31], op_12_V_fu_806_p3[31], op_12_V_fu_806_p3[31], op_12_V_fu_806_p3[31], op_12_V_fu_806_p3[31], op_12_V_fu_806_p3[31], op_12_V_fu_806_p3[31], op_12_V_fu_806_p3[31], op_12_V_fu_806_p3[31], op_12_V_fu_806_p3[31], op_12_V_fu_806_p3[31], op_12_V_fu_806_p3[31], op_12_V_fu_806_p3[31], op_12_V_fu_806_p3[31], op_12_V_fu_806_p3[31], op_12_V_fu_806_p3[31], op_12_V_fu_806_p3[31], op_12_V_fu_806_p3[31], op_12_V_fu_806_p3[31], op_12_V_fu_806_p3[31], op_12_V_fu_806_p3 };
assign sext_ln727_fu_869_p1 = { op_4_V_reg_1255[3], op_4_V_reg_1255[3], op_4_V_reg_1255 };
assign sext_ln731_fu_1039_p1 = { ret_V_11_reg_1273[3], ret_V_11_reg_1273[3], ret_V_11_reg_1273[3], ret_V_11_reg_1273[3], ret_V_11_reg_1273[3], ret_V_11_reg_1273[3], ret_V_11_reg_1273[3], ret_V_11_reg_1273 };
assign sext_ln831_fu_945_p1 = { ret_V_reg_1321[3], ret_V_reg_1321 };
assign sext_ln850_fu_723_p1 = { ret_V_14_fu_707_p2[4], ret_V_14_fu_707_p2[4:2] };
assign shl_ln_fu_872_p1 = op_8;
assign shl_ln_fu_872_p3 = { op_8, 2'h0 };
assign tmp_2_fu_713_p4 = ret_V_14_fu_707_p2[4:2];
assign tmp_3_fu_635_p4 = ret_2_fu_599_p2[4:2];
assign tmp_5_fu_447_p1 = op_1;
assign tmp_5_fu_447_p3 = op_1[1];
assign tmp_7_fu_988_p3 = r_V_reg_1348[2];
assign tmp_fu_285_p3 = ret_fu_201_p2[1];
assign trunc_ln731_1_fu_925_p1 = op_9[10:0];
assign trunc_ln731_2_fu_613_p0 = op_8;
assign trunc_ln731_2_fu_613_p1 = op_8[1:0];
assign trunc_ln731_fu_365_p0 = op_1;
assign trunc_ln731_fu_365_p1 = op_1[0];
assign trunc_ln790_fu_675_p1 = add_ln731_1_fu_621_p2[0];
assign trunc_ln851_1_fu_735_p1 = ret_V_14_fu_707_p2[1:0];
assign trunc_ln851_2_fu_846_p1 = op_12_V_fu_806_p3[29:0];
assign trunc_ln851_3_fu_1097_p1 = op_18_V_fu_1068_p3[20:0];
assign trunc_ln851_4_fu_1202_p0 = op_19;
assign trunc_ln851_4_fu_1202_p1 = op_19[13:0];
assign trunc_ln851_fu_901_p1 = r_V_fu_895_p2[1:0];
assign zext_ln1193_fu_703_p1 = { 2'h0, lhs_V_3_reg_1279, 2'h0 };
assign zext_ln1346_fu_591_p1 = { 4'h0, lhs_V_3_fu_585_p2 };
assign zext_ln215_1_fu_915_p1 = { 1'h0, op_9 };
assign zext_ln215_fu_911_p1 = { 17'h00000, ret_V_11_reg_1273[3], ret_V_11_reg_1273[3], ret_V_11_reg_1273[3], ret_V_11_reg_1273[3], ret_V_11_reg_1273[3], ret_V_11_reg_1273[3], ret_V_11_reg_1273[3], ret_V_11_reg_1273[3], ret_V_11_reg_1273[3], ret_V_11_reg_1273[3], ret_V_11_reg_1273[3], ret_V_11_reg_1273[3], ret_V_11_reg_1273 };
assign zext_ln69_1_fu_1088_p1 = { 31'h00000000, lhs_V_3_reg_1279 };
assign zext_ln69_fu_978_p1 = { 4'h0, icmp_ln1498_fu_879_p2 };
assign zext_ln703_fu_1107_p1 = { 22'h000000, op_18_V_reg_1389 };
assign zext_ln731_fu_617_p1 = { 1'h0, lhs_V_3_fu_585_p2 };
assign \mul_16ns_4s_20_1_1_U1.top_mul_16ns_4s_20_1_1_Multiplier_0_U.a  = \mul_16ns_4s_20_1_1_U1.din0 ;
assign \mul_16ns_4s_20_1_1_U1.top_mul_16ns_4s_20_1_1_Multiplier_0_U.b  = \mul_16ns_4s_20_1_1_U1.din1 ;
assign \mul_16ns_4s_20_1_1_U1.dout  = \mul_16ns_4s_20_1_1_U1.top_mul_16ns_4s_20_1_1_Multiplier_0_U.p ;
assign \mul_16ns_4s_20_1_1_U1.din0  = { ret_V_11_reg_1273[3], ret_V_11_reg_1273[3], ret_V_11_reg_1273[3], ret_V_11_reg_1273[3], ret_V_11_reg_1273[3], ret_V_11_reg_1273[3], ret_V_11_reg_1273[3], ret_V_11_reg_1273[3], ret_V_11_reg_1273[3], ret_V_11_reg_1273[3], ret_V_11_reg_1273[3], ret_V_11_reg_1273[3], ret_V_11_reg_1273 };
assign \mul_16ns_4s_20_1_1_U1.din1  = op_4_V_reg_1255;
assign r_V_fu_895_p2 = \mul_16ns_4s_20_1_1_U1.dout ;
endmodule


// Machine B:
// Processed by function `add_clk_enable_signal` in `verilog_tricks.py`.
// Processed by function `remove_reset_signal` in `verilog_tricks.py`.
module top_B (
  ap_clk,
  ap_start,
  ap_done,
  ap_idle,
  ap_ready,
  op_0,
  op_1,
  op_7,
  op_8,
  op_9,
  op_19,
  op_27,
  op_27_ap_vld,
clk_enable
);
input clk_enable;


input ap_clk;
wire ap_rst;
assign ap_rst = op_27_ap_vld;
input ap_start;
input [3:0] op_0;
input [3:0] op_1;
input [15:0] op_19;
input [31:0] op_7;
input [3:0] op_8;
input [31:0] op_9;
output ap_done;
output ap_idle;
output ap_ready;
output [31:0] op_27;
output op_27_ap_vld;


reg [5:0] \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_8_U.ain_s1 ;
reg [5:0] \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_8_U.bin_s1 ;
reg \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_8_U.carry_s1 ;
reg [4:0] \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_8_U.sum_s1 ;
reg \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_2_U.ain_s1 ;
reg \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_2_U.bin_s1 ;
reg \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_2_U.carry_s1 ;
reg \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_2_U.sum_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s1 ;
reg \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.carry_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.sum_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s1 ;
reg \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.carry_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.sum_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s1 ;
reg \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.carry_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.sum_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s1 ;
reg \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_6_U.carry_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_6_U.sum_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s1 ;
reg \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_6_U.carry_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_6_U.sum_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s1 ;
reg \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.carry_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.sum_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s1 ;
reg \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.carry_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.sum_s1 ;
reg [15:0] \add_32s_32ns_32_2_1_U15.top_add_32s_32ns_32_2_1_Adder_10_U.ain_s1 ;
reg [15:0] \add_32s_32ns_32_2_1_U15.top_add_32s_32ns_32_2_1_Adder_10_U.bin_s1 ;
reg \add_32s_32ns_32_2_1_U15.top_add_32s_32ns_32_2_1_Adder_10_U.carry_s1 ;
reg [15:0] \add_32s_32ns_32_2_1_U15.top_add_32s_32ns_32_2_1_Adder_10_U.sum_s1 ;
reg [16:0] \add_33ns_33ns_33_2_1_U10.top_add_33ns_33ns_33_2_1_Adder_7_U.ain_s1 ;
reg [16:0] \add_33ns_33ns_33_2_1_U10.top_add_33ns_33ns_33_2_1_Adder_7_U.bin_s1 ;
reg \add_33ns_33ns_33_2_1_U10.top_add_33ns_33ns_33_2_1_Adder_7_U.carry_s1 ;
reg [15:0] \add_33ns_33ns_33_2_1_U10.top_add_33ns_33ns_33_2_1_Adder_7_U.sum_s1 ;
reg [23:0] \add_47s_47s_47_2_1_U20.top_add_47s_47s_47_2_1_Adder_12_U.ain_s1 ;
reg [23:0] \add_47s_47s_47_2_1_U20.top_add_47s_47s_47_2_1_Adder_12_U.bin_s1 ;
reg \add_47s_47s_47_2_1_U20.top_add_47s_47s_47_2_1_Adder_12_U.carry_s1 ;
reg [22:0] \add_47s_47s_47_2_1_U20.top_add_47s_47s_47_2_1_Adder_12_U.sum_s1 ;
reg [1:0] \add_4s_4ns_4_2_1_U6.top_add_4s_4ns_4_2_1_Adder_4_U.ain_s1 ;
reg [1:0] \add_4s_4ns_4_2_1_U6.top_add_4s_4ns_4_2_1_Adder_4_U.bin_s1 ;
reg \add_4s_4ns_4_2_1_U6.top_add_4s_4ns_4_2_1_Adder_4_U.carry_s1 ;
reg [1:0] \add_4s_4ns_4_2_1_U6.top_add_4s_4ns_4_2_1_Adder_4_U.sum_s1 ;
reg [26:0] \add_54s_54ns_54_2_1_U18.top_add_54s_54ns_54_2_1_Adder_11_U.ain_s1 ;
reg [26:0] \add_54s_54ns_54_2_1_U18.top_add_54s_54ns_54_2_1_Adder_11_U.bin_s1 ;
reg \add_54s_54ns_54_2_1_U18.top_add_54s_54ns_54_2_1_Adder_11_U.carry_s1 ;
reg [26:0] \add_54s_54ns_54_2_1_U18.top_add_54s_54ns_54_2_1_Adder_11_U.sum_s1 ;
reg [2:0] \add_5ns_5ns_5_2_1_U14.top_add_5ns_5ns_5_2_1_Adder_9_U.ain_s1 ;
reg [2:0] \add_5ns_5ns_5_2_1_U14.top_add_5ns_5ns_5_2_1_Adder_9_U.bin_s1 ;
reg \add_5ns_5ns_5_2_1_U14.top_add_5ns_5ns_5_2_1_Adder_9_U.carry_s1 ;
reg [1:0] \add_5ns_5ns_5_2_1_U14.top_add_5ns_5ns_5_2_1_Adder_9_U.sum_s1 ;
reg [2:0] \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.ain_s1 ;
reg [2:0] \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.bin_s1 ;
reg \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.carry_s1 ;
reg [1:0] \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.sum_s1 ;
reg [31:0] \add_63s_63s_63_2_1_U7.top_add_63s_63s_63_2_1_Adder_5_U.ain_s1 ;
reg [31:0] \add_63s_63s_63_2_1_U7.top_add_63s_63s_63_2_1_Adder_5_U.bin_s1 ;
reg \add_63s_63s_63_2_1_U7.top_add_63s_63s_63_2_1_Adder_5_U.carry_s1 ;
reg [30:0] \add_63s_63s_63_2_1_U7.top_add_63s_63s_63_2_1_Adder_5_U.sum_s1 ;
reg [31:0] add_ln691_1_reg_1552;
reg [31:0] add_ln691_2_reg_1691;
reg [31:0] add_ln691_3_reg_1728;
reg [3:0] add_ln691_reg_1495;
reg [4:0] add_ln69_1_reg_1614;
reg [31:0] add_ln69_reg_1609;
reg [1:0] add_ln731_1_reg_1358;
reg [10:0] add_ln731_reg_1562;
reg and_ln340_reg_1229;
reg and_ln785_1_reg_1234;
reg and_ln786_reg_1304;
reg [36:0] ap_CS_fsm = 37'h0000000001;
reg icmp_ln1498_reg_1423;
reg icmp_ln768_1_reg_1171;
reg icmp_ln768_2_reg_1594;
reg icmp_ln768_3_reg_1369;
reg icmp_ln768_reg_1212;
reg icmp_ln786_1_reg_1176;
reg icmp_ln786_2_reg_1374;
reg icmp_ln786_reg_1217;
reg icmp_ln790_reg_1397;
reg icmp_ln850_reg_1604;
reg icmp_ln851_1_reg_1490;
reg icmp_ln851_2_reg_1674;
reg icmp_ln851_3_reg_1711;
reg icmp_ln851_reg_1475;
reg lhs_V_3_reg_1278;
reg [15:0] \mul_16ns_4s_20_7_1_U5.top_mul_16ns_4s_20_7_1_Mul_DSP_0_U.a_reg0 ;
reg [3:0] \mul_16ns_4s_20_7_1_U5.top_mul_16ns_4s_20_7_1_Mul_DSP_0_U.b_reg0 ;
reg [19:0] \mul_16ns_4s_20_7_1_U5.top_mul_16ns_4s_20_7_1_Mul_DSP_0_U.buff0 ;
reg [19:0] \mul_16ns_4s_20_7_1_U5.top_mul_16ns_4s_20_7_1_Mul_DSP_0_U.buff1 ;
reg [19:0] \mul_16ns_4s_20_7_1_U5.top_mul_16ns_4s_20_7_1_Mul_DSP_0_U.buff2 ;
reg [19:0] \mul_16ns_4s_20_7_1_U5.top_mul_16ns_4s_20_7_1_Mul_DSP_0_U.buff3 ;
reg [19:0] \mul_16ns_4s_20_7_1_U5.top_mul_16ns_4s_20_7_1_Mul_DSP_0_U.buff4 ;
reg newsignbit_reg_1195;
reg [31:0] op_12_V_reg_1458;
reg [4:0] op_15_V_reg_1573;
reg op_16_V_reg_1619;
reg [31:0] op_18_V_reg_1649;
reg [31:0] op_23_V_reg_1629;
reg [31:0] op_25_V_reg_1654;
reg op_2_V_reg_1244;
reg [3:0] op_4_V_reg_1384;
reg or_ln340_1_reg_1298;
reg or_ln384_reg_1418;
reg or_ln785_1_reg_1266;
reg or_ln785_reg_1223;
reg or_ln786_1_reg_1292;
reg overflow_3_reg_1391;
reg p_Result_13_reg_1188;
reg p_Result_15_reg_1164;
reg p_Result_16_reg_1259;
reg p_Result_19_reg_1336;
reg p_Result_20_reg_1363;
reg [21:0] p_Result_4_reg_1568;
reg [3:0] p_Result_s_reg_1206;
reg [3:0] p_Val2_2_reg_1251;
reg [19:0] r_V_reg_1583;
reg [3:0] ret_V_11_reg_1402;
reg [31:0] ret_V_12_reg_1557;
reg [4:0] ret_V_14_reg_1443;
reg [62:0] ret_V_15_reg_1500;
reg [31:0] ret_V_16_reg_1578;
reg [31:0] ret_V_17_reg_1639;
reg [31:0] ret_V_18_cast_reg_1684;
reg [53:0] ret_V_18_reg_1679;
reg [46:0] ret_V_19_reg_1716;
reg [31:0] ret_V_20_cast_reg_1721;
reg [31:0] ret_V_7_cast_reg_1505;
reg [3:0] ret_V_reg_1517;
reg [4:0] ret_reg_1182;
reg sel_tmp18_reg_1331;
reg [31:0] select_ln1192_1_reg_1634;
reg [31:0] select_ln1192_reg_1512;
reg [3:0] select_ln340_1_reg_1326;
reg select_ln340_reg_1239;
reg [31:0] select_ln353_reg_1696;
reg [3:0] select_ln785_reg_1353;
reg [15:0] sext_ln1118_reg_1433;
reg [4:0] sext_ln1346_reg_1315;
reg [3:0] sext_ln850_reg_1468;
reg [2:0] \sub_5s_5ns_5_2_1_U4.top_sub_5s_5ns_5_2_1_Adder_3_U.ain_s1 ;
reg [2:0] \sub_5s_5ns_5_2_1_U4.top_sub_5s_5ns_5_2_1_Adder_3_U.bin_s1 ;
reg \sub_5s_5ns_5_2_1_U4.top_sub_5s_5ns_5_2_1_Adder_3_U.carry_s1 ;
reg [1:0] \sub_5s_5ns_5_2_1_U4.top_sub_5s_5ns_5_2_1_Adder_3_U.sum_s1 ;
reg [2:0] \sub_5s_5s_5_2_1_U1.top_sub_5s_5s_5_2_1_Adder_0_U.ain_s1 ;
reg [2:0] \sub_5s_5s_5_2_1_U1.top_sub_5s_5s_5_2_1_Adder_0_U.bin_s1 ;
reg \sub_5s_5s_5_2_1_U1.top_sub_5s_5s_5_2_1_Adder_0_U.carry_s1 ;
reg [1:0] \sub_5s_5s_5_2_1_U1.top_sub_5s_5s_5_2_1_Adder_0_U.sum_s1 ;
reg [2:0] \sub_5s_5s_5_2_1_U12.top_sub_5s_5s_5_2_1_Adder_0_U.ain_s1 ;
reg [2:0] \sub_5s_5s_5_2_1_U12.top_sub_5s_5s_5_2_1_Adder_0_U.bin_s1 ;
reg \sub_5s_5s_5_2_1_U12.top_sub_5s_5s_5_2_1_Adder_0_U.carry_s1 ;
reg [1:0] \sub_5s_5s_5_2_1_U12.top_sub_5s_5s_5_2_1_Adder_0_U.sum_s1 ;
reg [2:0] tmp_2_reg_1448;
reg [2:0] tmp_3_reg_1347;
reg [1:0] trunc_ln731_2_reg_1321;
reg trunc_ln790_reg_1379;
reg [1:0] trunc_ln851_1_reg_1453;
reg [29:0] trunc_ln851_2_reg_1463;
reg [20:0] trunc_ln851_3_reg_1659;
reg [1:0] trunc_ln851_reg_1589;
reg xor_ln785_1_reg_1272;
wire [31:0] _000_;
wire [31:0] _001_;
wire [31:0] _002_;
wire [3:0] _003_;
wire [4:0] _004_;
wire [31:0] _005_;
wire [1:0] _006_;
wire [10:0] _007_;
wire _008_;
wire _009_;
wire _010_;
wire [36:0] _011_;
wire _012_;
wire _013_;
wire _014_;
wire _015_;
wire _016_;
wire _017_;
wire _018_;
wire _019_;
wire _020_;
wire _021_;
wire _022_;
wire _023_;
wire _024_;
wire _025_;
wire _026_;
wire _027_;
wire [31:0] _028_;
wire [4:0] _029_;
wire _030_;
wire [10:0] _031_;
wire [31:0] _032_;
wire [31:0] _033_;
wire _034_;
wire [3:0] _035_;
wire _036_;
wire _037_;
wire _038_;
wire _039_;
wire _040_;
wire _041_;
wire _042_;
wire _043_;
wire _044_;
wire _045_;
wire _046_;
wire [21:0] _047_;
wire [3:0] _048_;
wire _049_;
wire [19:0] _050_;
wire [3:0] _051_;
wire [31:0] _052_;
wire [4:0] _053_;
wire [62:0] _054_;
wire [31:0] _055_;
wire [31:0] _056_;
wire [31:0] _057_;
wire [53:0] _058_;
wire [46:0] _059_;
wire [31:0] _060_;
wire [31:0] _061_;
wire [3:0] _062_;
wire [4:0] _063_;
wire _064_;
wire [31:0] _065_;
wire [31:0] _066_;
wire [3:0] _067_;
wire _068_;
wire [31:0] _069_;
wire [3:0] _070_;
wire [15:0] _071_;
wire [4:0] _072_;
wire [3:0] _073_;
wire [2:0] _074_;
wire [2:0] _075_;
wire [1:0] _076_;
wire _077_;
wire [1:0] _078_;
wire [29:0] _079_;
wire [1:0] _080_;
wire _081_;
wire [1:0] _082_;
wire _083_;
wire _084_;
wire _085_;
wire _086_;
wire _087_;
wire _088_;
wire _089_;
wire _090_;
wire _091_;
wire _092_;
wire _093_;
wire _094_;
wire [5:0] _095_;
wire [5:0] _096_;
wire _097_;
wire [4:0] _098_;
wire [5:0] _099_;
wire [6:0] _100_;
wire _101_;
wire _102_;
wire _103_;
wire _104_;
wire [1:0] _105_;
wire [1:0] _106_;
wire [15:0] _107_;
wire [15:0] _108_;
wire _109_;
wire [15:0] _110_;
wire [16:0] _111_;
wire [16:0] _112_;
wire [15:0] _113_;
wire [15:0] _114_;
wire _115_;
wire [15:0] _116_;
wire [16:0] _117_;
wire [16:0] _118_;
wire [15:0] _119_;
wire [15:0] _120_;
wire _121_;
wire [15:0] _122_;
wire [16:0] _123_;
wire [16:0] _124_;
wire [15:0] _125_;
wire [15:0] _126_;
wire _127_;
wire [15:0] _128_;
wire [16:0] _129_;
wire [16:0] _130_;
wire [15:0] _131_;
wire [15:0] _132_;
wire _133_;
wire [15:0] _134_;
wire [16:0] _135_;
wire [16:0] _136_;
wire [15:0] _137_;
wire [15:0] _138_;
wire _139_;
wire [15:0] _140_;
wire [16:0] _141_;
wire [16:0] _142_;
wire [15:0] _143_;
wire [15:0] _144_;
wire _145_;
wire [15:0] _146_;
wire [16:0] _147_;
wire [16:0] _148_;
wire [15:0] _149_;
wire [15:0] _150_;
wire _151_;
wire [15:0] _152_;
wire [16:0] _153_;
wire [16:0] _154_;
wire [16:0] _155_;
wire [16:0] _156_;
wire _157_;
wire [15:0] _158_;
wire [16:0] _159_;
wire [17:0] _160_;
wire [23:0] _161_;
wire [23:0] _162_;
wire _163_;
wire [22:0] _164_;
wire [23:0] _165_;
wire [24:0] _166_;
wire [1:0] _167_;
wire [1:0] _168_;
wire _169_;
wire [1:0] _170_;
wire [2:0] _171_;
wire [2:0] _172_;
wire [26:0] _173_;
wire [26:0] _174_;
wire _175_;
wire [26:0] _176_;
wire [27:0] _177_;
wire [27:0] _178_;
wire [2:0] _179_;
wire [2:0] _180_;
wire _181_;
wire [1:0] _182_;
wire [2:0] _183_;
wire [3:0] _184_;
wire [2:0] _185_;
wire [2:0] _186_;
wire _187_;
wire [1:0] _188_;
wire [2:0] _189_;
wire [3:0] _190_;
wire [31:0] _191_;
wire [31:0] _192_;
wire _193_;
wire [30:0] _194_;
wire [31:0] _195_;
wire [32:0] _196_;
wire [15:0] _197_;
wire [3:0] _198_;
wire [19:0] _199_;
wire [19:0] _200_;
wire [19:0] _201_;
wire [19:0] _202_;
wire [19:0] _203_;
wire [2:0] _204_;
wire [2:0] _205_;
wire _206_;
wire [1:0] _207_;
wire [2:0] _208_;
wire [3:0] _209_;
wire [2:0] _210_;
wire [2:0] _211_;
wire _212_;
wire [1:0] _213_;
wire [2:0] _214_;
wire [3:0] _215_;
wire [2:0] _216_;
wire [2:0] _217_;
wire _218_;
wire [1:0] _219_;
wire [2:0] _220_;
wire [3:0] _221_;
wire _222_;
wire _223_;
wire _224_;
wire _225_;
wire _226_;
wire _227_;
wire _228_;
wire _229_;
wire _230_;
wire _231_;
wire _232_;
wire _233_;
wire _234_;
wire _235_;
wire _236_;
wire _237_;
wire _238_;
wire _239_;
wire _240_;
wire _241_;
wire _242_;
wire _243_;
wire _244_;
wire _245_;
wire _246_;
wire _247_;
wire _248_;
wire _249_;
wire _250_;
wire _251_;
wire _252_;
wire _253_;
wire _254_;
wire _255_;
wire _256_;
wire _257_;
wire _258_;
wire _259_;
wire _260_;
wire _261_;
wire _262_;
wire _263_;
wire _264_;
wire _265_;
wire _266_;
wire _267_;
wire _268_;
wire _269_;
wire _270_;
wire _271_;
wire \add_11ns_11s_11_2_1_U11.ce ;
wire \add_11ns_11s_11_2_1_U11.clk ;
wire [10:0] \add_11ns_11s_11_2_1_U11.din0 ;
wire [10:0] \add_11ns_11s_11_2_1_U11.din1 ;
wire [10:0] \add_11ns_11s_11_2_1_U11.dout ;
wire \add_11ns_11s_11_2_1_U11.reset ;
wire [10:0] \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_8_U.a ;
wire [10:0] \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_8_U.ain_s0 ;
wire [10:0] \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_8_U.b ;
wire [10:0] \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_8_U.bin_s0 ;
wire \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_8_U.ce ;
wire \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_8_U.clk ;
wire \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_8_U.facout_s1 ;
wire \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_8_U.facout_s2 ;
wire [4:0] \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_8_U.fas_s1 ;
wire [5:0] \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_8_U.fas_s2 ;
wire \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_8_U.reset ;
wire [10:0] \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_8_U.s ;
wire [4:0] \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_8_U.u1.a ;
wire [4:0] \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_8_U.u1.b ;
wire \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_8_U.u1.cin ;
wire \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_8_U.u1.cout ;
wire [4:0] \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_8_U.u1.s ;
wire [5:0] \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_8_U.u2.a ;
wire [5:0] \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_8_U.u2.b ;
wire \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_8_U.u2.cin ;
wire \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_8_U.u2.cout ;
wire [5:0] \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_8_U.u2.s ;
wire \add_2ns_2ns_2_2_1_U3.ce ;
wire \add_2ns_2ns_2_2_1_U3.clk ;
wire [1:0] \add_2ns_2ns_2_2_1_U3.din0 ;
wire [1:0] \add_2ns_2ns_2_2_1_U3.din1 ;
wire [1:0] \add_2ns_2ns_2_2_1_U3.dout ;
wire \add_2ns_2ns_2_2_1_U3.reset ;
wire [1:0] \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_2_U.a ;
wire [1:0] \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_2_U.ain_s0 ;
wire [1:0] \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_2_U.b ;
wire [1:0] \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_2_U.bin_s0 ;
wire \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_2_U.ce ;
wire \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_2_U.clk ;
wire \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_2_U.facout_s1 ;
wire \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_2_U.facout_s2 ;
wire \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_2_U.fas_s1 ;
wire \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_2_U.fas_s2 ;
wire \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_2_U.reset ;
wire [1:0] \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_2_U.s ;
wire \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_2_U.u1.a ;
wire \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_2_U.u1.b ;
wire \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_2_U.u1.cin ;
wire \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_2_U.u1.cout ;
wire \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_2_U.u1.s ;
wire \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_2_U.u2.a ;
wire \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_2_U.u2.b ;
wire \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_2_U.u2.cin ;
wire \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_2_U.u2.cout ;
wire \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_2_U.u2.s ;
wire \add_32ns_32ns_32_2_1_U13.ce ;
wire \add_32ns_32ns_32_2_1_U13.clk ;
wire [31:0] \add_32ns_32ns_32_2_1_U13.din0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U13.din1 ;
wire [31:0] \add_32ns_32ns_32_2_1_U13.dout ;
wire \add_32ns_32ns_32_2_1_U13.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.a ;
wire [31:0] \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.b ;
wire [31:0] \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s0 ;
wire \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.ce ;
wire \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.clk ;
wire \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s1 ;
wire \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s2 ;
wire [15:0] \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s1 ;
wire [15:0] \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s2 ;
wire \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.b ;
wire \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cin ;
wire \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.b ;
wire \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cin ;
wire \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.s ;
wire \add_32ns_32ns_32_2_1_U16.ce ;
wire \add_32ns_32ns_32_2_1_U16.clk ;
wire [31:0] \add_32ns_32ns_32_2_1_U16.din0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U16.din1 ;
wire [31:0] \add_32ns_32ns_32_2_1_U16.dout ;
wire \add_32ns_32ns_32_2_1_U16.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.a ;
wire [31:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.b ;
wire [31:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s0 ;
wire \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.ce ;
wire \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.clk ;
wire \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s1 ;
wire \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s2 ;
wire [15:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s1 ;
wire [15:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s2 ;
wire \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.b ;
wire \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cin ;
wire \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.b ;
wire \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cin ;
wire \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.s ;
wire \add_32ns_32ns_32_2_1_U17.ce ;
wire \add_32ns_32ns_32_2_1_U17.clk ;
wire [31:0] \add_32ns_32ns_32_2_1_U17.din0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U17.din1 ;
wire [31:0] \add_32ns_32ns_32_2_1_U17.dout ;
wire \add_32ns_32ns_32_2_1_U17.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.a ;
wire [31:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.b ;
wire [31:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s0 ;
wire \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.ce ;
wire \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.clk ;
wire \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s1 ;
wire \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s2 ;
wire [15:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s1 ;
wire [15:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s2 ;
wire \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.b ;
wire \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cin ;
wire \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.b ;
wire \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cin ;
wire \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.s ;
wire \add_32ns_32ns_32_2_1_U19.ce ;
wire \add_32ns_32ns_32_2_1_U19.clk ;
wire [31:0] \add_32ns_32ns_32_2_1_U19.din0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U19.din1 ;
wire [31:0] \add_32ns_32ns_32_2_1_U19.dout ;
wire \add_32ns_32ns_32_2_1_U19.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_6_U.a ;
wire [31:0] \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_6_U.b ;
wire [31:0] \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s0 ;
wire \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_6_U.ce ;
wire \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_6_U.clk ;
wire \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s1 ;
wire \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s2 ;
wire [15:0] \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s1 ;
wire [15:0] \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s2 ;
wire \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_6_U.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_6_U.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.b ;
wire \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cin ;
wire \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.b ;
wire \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cin ;
wire \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.s ;
wire \add_32ns_32ns_32_2_1_U21.ce ;
wire \add_32ns_32ns_32_2_1_U21.clk ;
wire [31:0] \add_32ns_32ns_32_2_1_U21.din0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U21.din1 ;
wire [31:0] \add_32ns_32ns_32_2_1_U21.dout ;
wire \add_32ns_32ns_32_2_1_U21.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_6_U.a ;
wire [31:0] \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_6_U.b ;
wire [31:0] \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s0 ;
wire \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_6_U.ce ;
wire \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_6_U.clk ;
wire \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s1 ;
wire \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s2 ;
wire [15:0] \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s1 ;
wire [15:0] \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s2 ;
wire \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_6_U.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_6_U.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.b ;
wire \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cin ;
wire \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.b ;
wire \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cin ;
wire \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.s ;
wire \add_32ns_32ns_32_2_1_U8.ce ;
wire \add_32ns_32ns_32_2_1_U8.clk ;
wire [31:0] \add_32ns_32ns_32_2_1_U8.din0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U8.din1 ;
wire [31:0] \add_32ns_32ns_32_2_1_U8.dout ;
wire \add_32ns_32ns_32_2_1_U8.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.a ;
wire [31:0] \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.b ;
wire [31:0] \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s0 ;
wire \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.ce ;
wire \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.clk ;
wire \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s1 ;
wire \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s2 ;
wire [15:0] \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s1 ;
wire [15:0] \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s2 ;
wire \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.b ;
wire \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cin ;
wire \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.b ;
wire \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cin ;
wire \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.s ;
wire \add_32ns_32ns_32_2_1_U9.ce ;
wire \add_32ns_32ns_32_2_1_U9.clk ;
wire [31:0] \add_32ns_32ns_32_2_1_U9.din0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U9.din1 ;
wire [31:0] \add_32ns_32ns_32_2_1_U9.dout ;
wire \add_32ns_32ns_32_2_1_U9.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.a ;
wire [31:0] \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.b ;
wire [31:0] \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s0 ;
wire \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.ce ;
wire \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.clk ;
wire \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s1 ;
wire \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s2 ;
wire [15:0] \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s1 ;
wire [15:0] \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s2 ;
wire \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.b ;
wire \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cin ;
wire \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.b ;
wire \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cin ;
wire \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.s ;
wire \add_32s_32ns_32_2_1_U15.ce ;
wire \add_32s_32ns_32_2_1_U15.clk ;
wire [31:0] \add_32s_32ns_32_2_1_U15.din0 ;
wire [31:0] \add_32s_32ns_32_2_1_U15.din1 ;
wire [31:0] \add_32s_32ns_32_2_1_U15.dout ;
wire \add_32s_32ns_32_2_1_U15.reset ;
wire [31:0] \add_32s_32ns_32_2_1_U15.top_add_32s_32ns_32_2_1_Adder_10_U.a ;
wire [31:0] \add_32s_32ns_32_2_1_U15.top_add_32s_32ns_32_2_1_Adder_10_U.ain_s0 ;
wire [31:0] \add_32s_32ns_32_2_1_U15.top_add_32s_32ns_32_2_1_Adder_10_U.b ;
wire [31:0] \add_32s_32ns_32_2_1_U15.top_add_32s_32ns_32_2_1_Adder_10_U.bin_s0 ;
wire \add_32s_32ns_32_2_1_U15.top_add_32s_32ns_32_2_1_Adder_10_U.ce ;
wire \add_32s_32ns_32_2_1_U15.top_add_32s_32ns_32_2_1_Adder_10_U.clk ;
wire \add_32s_32ns_32_2_1_U15.top_add_32s_32ns_32_2_1_Adder_10_U.facout_s1 ;
wire \add_32s_32ns_32_2_1_U15.top_add_32s_32ns_32_2_1_Adder_10_U.facout_s2 ;
wire [15:0] \add_32s_32ns_32_2_1_U15.top_add_32s_32ns_32_2_1_Adder_10_U.fas_s1 ;
wire [15:0] \add_32s_32ns_32_2_1_U15.top_add_32s_32ns_32_2_1_Adder_10_U.fas_s2 ;
wire \add_32s_32ns_32_2_1_U15.top_add_32s_32ns_32_2_1_Adder_10_U.reset ;
wire [31:0] \add_32s_32ns_32_2_1_U15.top_add_32s_32ns_32_2_1_Adder_10_U.s ;
wire [15:0] \add_32s_32ns_32_2_1_U15.top_add_32s_32ns_32_2_1_Adder_10_U.u1.a ;
wire [15:0] \add_32s_32ns_32_2_1_U15.top_add_32s_32ns_32_2_1_Adder_10_U.u1.b ;
wire \add_32s_32ns_32_2_1_U15.top_add_32s_32ns_32_2_1_Adder_10_U.u1.cin ;
wire \add_32s_32ns_32_2_1_U15.top_add_32s_32ns_32_2_1_Adder_10_U.u1.cout ;
wire [15:0] \add_32s_32ns_32_2_1_U15.top_add_32s_32ns_32_2_1_Adder_10_U.u1.s ;
wire [15:0] \add_32s_32ns_32_2_1_U15.top_add_32s_32ns_32_2_1_Adder_10_U.u2.a ;
wire [15:0] \add_32s_32ns_32_2_1_U15.top_add_32s_32ns_32_2_1_Adder_10_U.u2.b ;
wire \add_32s_32ns_32_2_1_U15.top_add_32s_32ns_32_2_1_Adder_10_U.u2.cin ;
wire \add_32s_32ns_32_2_1_U15.top_add_32s_32ns_32_2_1_Adder_10_U.u2.cout ;
wire [15:0] \add_32s_32ns_32_2_1_U15.top_add_32s_32ns_32_2_1_Adder_10_U.u2.s ;
wire \add_33ns_33ns_33_2_1_U10.ce ;
wire \add_33ns_33ns_33_2_1_U10.clk ;
wire [32:0] \add_33ns_33ns_33_2_1_U10.din0 ;
wire [32:0] \add_33ns_33ns_33_2_1_U10.din1 ;
wire [32:0] \add_33ns_33ns_33_2_1_U10.dout ;
wire \add_33ns_33ns_33_2_1_U10.reset ;
wire [32:0] \add_33ns_33ns_33_2_1_U10.top_add_33ns_33ns_33_2_1_Adder_7_U.a ;
wire [32:0] \add_33ns_33ns_33_2_1_U10.top_add_33ns_33ns_33_2_1_Adder_7_U.ain_s0 ;
wire [32:0] \add_33ns_33ns_33_2_1_U10.top_add_33ns_33ns_33_2_1_Adder_7_U.b ;
wire [32:0] \add_33ns_33ns_33_2_1_U10.top_add_33ns_33ns_33_2_1_Adder_7_U.bin_s0 ;
wire \add_33ns_33ns_33_2_1_U10.top_add_33ns_33ns_33_2_1_Adder_7_U.ce ;
wire \add_33ns_33ns_33_2_1_U10.top_add_33ns_33ns_33_2_1_Adder_7_U.clk ;
wire \add_33ns_33ns_33_2_1_U10.top_add_33ns_33ns_33_2_1_Adder_7_U.facout_s1 ;
wire \add_33ns_33ns_33_2_1_U10.top_add_33ns_33ns_33_2_1_Adder_7_U.facout_s2 ;
wire [15:0] \add_33ns_33ns_33_2_1_U10.top_add_33ns_33ns_33_2_1_Adder_7_U.fas_s1 ;
wire [16:0] \add_33ns_33ns_33_2_1_U10.top_add_33ns_33ns_33_2_1_Adder_7_U.fas_s2 ;
wire \add_33ns_33ns_33_2_1_U10.top_add_33ns_33ns_33_2_1_Adder_7_U.reset ;
wire [32:0] \add_33ns_33ns_33_2_1_U10.top_add_33ns_33ns_33_2_1_Adder_7_U.s ;
wire [15:0] \add_33ns_33ns_33_2_1_U10.top_add_33ns_33ns_33_2_1_Adder_7_U.u1.a ;
wire [15:0] \add_33ns_33ns_33_2_1_U10.top_add_33ns_33ns_33_2_1_Adder_7_U.u1.b ;
wire \add_33ns_33ns_33_2_1_U10.top_add_33ns_33ns_33_2_1_Adder_7_U.u1.cin ;
wire \add_33ns_33ns_33_2_1_U10.top_add_33ns_33ns_33_2_1_Adder_7_U.u1.cout ;
wire [15:0] \add_33ns_33ns_33_2_1_U10.top_add_33ns_33ns_33_2_1_Adder_7_U.u1.s ;
wire [16:0] \add_33ns_33ns_33_2_1_U10.top_add_33ns_33ns_33_2_1_Adder_7_U.u2.a ;
wire [16:0] \add_33ns_33ns_33_2_1_U10.top_add_33ns_33ns_33_2_1_Adder_7_U.u2.b ;
wire \add_33ns_33ns_33_2_1_U10.top_add_33ns_33ns_33_2_1_Adder_7_U.u2.cin ;
wire \add_33ns_33ns_33_2_1_U10.top_add_33ns_33ns_33_2_1_Adder_7_U.u2.cout ;
wire [16:0] \add_33ns_33ns_33_2_1_U10.top_add_33ns_33ns_33_2_1_Adder_7_U.u2.s ;
wire \add_47s_47s_47_2_1_U20.ce ;
wire \add_47s_47s_47_2_1_U20.clk ;
wire [46:0] \add_47s_47s_47_2_1_U20.din0 ;
wire [46:0] \add_47s_47s_47_2_1_U20.din1 ;
wire [46:0] \add_47s_47s_47_2_1_U20.dout ;
wire \add_47s_47s_47_2_1_U20.reset ;
wire [46:0] \add_47s_47s_47_2_1_U20.top_add_47s_47s_47_2_1_Adder_12_U.a ;
wire [46:0] \add_47s_47s_47_2_1_U20.top_add_47s_47s_47_2_1_Adder_12_U.ain_s0 ;
wire [46:0] \add_47s_47s_47_2_1_U20.top_add_47s_47s_47_2_1_Adder_12_U.b ;
wire [46:0] \add_47s_47s_47_2_1_U20.top_add_47s_47s_47_2_1_Adder_12_U.bin_s0 ;
wire \add_47s_47s_47_2_1_U20.top_add_47s_47s_47_2_1_Adder_12_U.ce ;
wire \add_47s_47s_47_2_1_U20.top_add_47s_47s_47_2_1_Adder_12_U.clk ;
wire \add_47s_47s_47_2_1_U20.top_add_47s_47s_47_2_1_Adder_12_U.facout_s1 ;
wire \add_47s_47s_47_2_1_U20.top_add_47s_47s_47_2_1_Adder_12_U.facout_s2 ;
wire [22:0] \add_47s_47s_47_2_1_U20.top_add_47s_47s_47_2_1_Adder_12_U.fas_s1 ;
wire [23:0] \add_47s_47s_47_2_1_U20.top_add_47s_47s_47_2_1_Adder_12_U.fas_s2 ;
wire \add_47s_47s_47_2_1_U20.top_add_47s_47s_47_2_1_Adder_12_U.reset ;
wire [46:0] \add_47s_47s_47_2_1_U20.top_add_47s_47s_47_2_1_Adder_12_U.s ;
wire [22:0] \add_47s_47s_47_2_1_U20.top_add_47s_47s_47_2_1_Adder_12_U.u1.a ;
wire [22:0] \add_47s_47s_47_2_1_U20.top_add_47s_47s_47_2_1_Adder_12_U.u1.b ;
wire \add_47s_47s_47_2_1_U20.top_add_47s_47s_47_2_1_Adder_12_U.u1.cin ;
wire \add_47s_47s_47_2_1_U20.top_add_47s_47s_47_2_1_Adder_12_U.u1.cout ;
wire [22:0] \add_47s_47s_47_2_1_U20.top_add_47s_47s_47_2_1_Adder_12_U.u1.s ;
wire [23:0] \add_47s_47s_47_2_1_U20.top_add_47s_47s_47_2_1_Adder_12_U.u2.a ;
wire [23:0] \add_47s_47s_47_2_1_U20.top_add_47s_47s_47_2_1_Adder_12_U.u2.b ;
wire \add_47s_47s_47_2_1_U20.top_add_47s_47s_47_2_1_Adder_12_U.u2.cin ;
wire \add_47s_47s_47_2_1_U20.top_add_47s_47s_47_2_1_Adder_12_U.u2.cout ;
wire [23:0] \add_47s_47s_47_2_1_U20.top_add_47s_47s_47_2_1_Adder_12_U.u2.s ;
wire \add_4s_4ns_4_2_1_U6.ce ;
wire \add_4s_4ns_4_2_1_U6.clk ;
wire [3:0] \add_4s_4ns_4_2_1_U6.din0 ;
wire [3:0] \add_4s_4ns_4_2_1_U6.din1 ;
wire [3:0] \add_4s_4ns_4_2_1_U6.dout ;
wire \add_4s_4ns_4_2_1_U6.reset ;
wire [3:0] \add_4s_4ns_4_2_1_U6.top_add_4s_4ns_4_2_1_Adder_4_U.a ;
wire [3:0] \add_4s_4ns_4_2_1_U6.top_add_4s_4ns_4_2_1_Adder_4_U.ain_s0 ;
wire [3:0] \add_4s_4ns_4_2_1_U6.top_add_4s_4ns_4_2_1_Adder_4_U.b ;
wire [3:0] \add_4s_4ns_4_2_1_U6.top_add_4s_4ns_4_2_1_Adder_4_U.bin_s0 ;
wire \add_4s_4ns_4_2_1_U6.top_add_4s_4ns_4_2_1_Adder_4_U.ce ;
wire \add_4s_4ns_4_2_1_U6.top_add_4s_4ns_4_2_1_Adder_4_U.clk ;
wire \add_4s_4ns_4_2_1_U6.top_add_4s_4ns_4_2_1_Adder_4_U.facout_s1 ;
wire \add_4s_4ns_4_2_1_U6.top_add_4s_4ns_4_2_1_Adder_4_U.facout_s2 ;
wire [1:0] \add_4s_4ns_4_2_1_U6.top_add_4s_4ns_4_2_1_Adder_4_U.fas_s1 ;
wire [1:0] \add_4s_4ns_4_2_1_U6.top_add_4s_4ns_4_2_1_Adder_4_U.fas_s2 ;
wire \add_4s_4ns_4_2_1_U6.top_add_4s_4ns_4_2_1_Adder_4_U.reset ;
wire [3:0] \add_4s_4ns_4_2_1_U6.top_add_4s_4ns_4_2_1_Adder_4_U.s ;
wire [1:0] \add_4s_4ns_4_2_1_U6.top_add_4s_4ns_4_2_1_Adder_4_U.u1.a ;
wire [1:0] \add_4s_4ns_4_2_1_U6.top_add_4s_4ns_4_2_1_Adder_4_U.u1.b ;
wire \add_4s_4ns_4_2_1_U6.top_add_4s_4ns_4_2_1_Adder_4_U.u1.cin ;
wire \add_4s_4ns_4_2_1_U6.top_add_4s_4ns_4_2_1_Adder_4_U.u1.cout ;
wire [1:0] \add_4s_4ns_4_2_1_U6.top_add_4s_4ns_4_2_1_Adder_4_U.u1.s ;
wire [1:0] \add_4s_4ns_4_2_1_U6.top_add_4s_4ns_4_2_1_Adder_4_U.u2.a ;
wire [1:0] \add_4s_4ns_4_2_1_U6.top_add_4s_4ns_4_2_1_Adder_4_U.u2.b ;
wire \add_4s_4ns_4_2_1_U6.top_add_4s_4ns_4_2_1_Adder_4_U.u2.cin ;
wire \add_4s_4ns_4_2_1_U6.top_add_4s_4ns_4_2_1_Adder_4_U.u2.cout ;
wire [1:0] \add_4s_4ns_4_2_1_U6.top_add_4s_4ns_4_2_1_Adder_4_U.u2.s ;
wire \add_54s_54ns_54_2_1_U18.ce ;
wire \add_54s_54ns_54_2_1_U18.clk ;
wire [53:0] \add_54s_54ns_54_2_1_U18.din0 ;
wire [53:0] \add_54s_54ns_54_2_1_U18.din1 ;
wire [53:0] \add_54s_54ns_54_2_1_U18.dout ;
wire \add_54s_54ns_54_2_1_U18.reset ;
wire [53:0] \add_54s_54ns_54_2_1_U18.top_add_54s_54ns_54_2_1_Adder_11_U.a ;
wire [53:0] \add_54s_54ns_54_2_1_U18.top_add_54s_54ns_54_2_1_Adder_11_U.ain_s0 ;
wire [53:0] \add_54s_54ns_54_2_1_U18.top_add_54s_54ns_54_2_1_Adder_11_U.b ;
wire [53:0] \add_54s_54ns_54_2_1_U18.top_add_54s_54ns_54_2_1_Adder_11_U.bin_s0 ;
wire \add_54s_54ns_54_2_1_U18.top_add_54s_54ns_54_2_1_Adder_11_U.ce ;
wire \add_54s_54ns_54_2_1_U18.top_add_54s_54ns_54_2_1_Adder_11_U.clk ;
wire \add_54s_54ns_54_2_1_U18.top_add_54s_54ns_54_2_1_Adder_11_U.facout_s1 ;
wire \add_54s_54ns_54_2_1_U18.top_add_54s_54ns_54_2_1_Adder_11_U.facout_s2 ;
wire [26:0] \add_54s_54ns_54_2_1_U18.top_add_54s_54ns_54_2_1_Adder_11_U.fas_s1 ;
wire [26:0] \add_54s_54ns_54_2_1_U18.top_add_54s_54ns_54_2_1_Adder_11_U.fas_s2 ;
wire \add_54s_54ns_54_2_1_U18.top_add_54s_54ns_54_2_1_Adder_11_U.reset ;
wire [53:0] \add_54s_54ns_54_2_1_U18.top_add_54s_54ns_54_2_1_Adder_11_U.s ;
wire [26:0] \add_54s_54ns_54_2_1_U18.top_add_54s_54ns_54_2_1_Adder_11_U.u1.a ;
wire [26:0] \add_54s_54ns_54_2_1_U18.top_add_54s_54ns_54_2_1_Adder_11_U.u1.b ;
wire \add_54s_54ns_54_2_1_U18.top_add_54s_54ns_54_2_1_Adder_11_U.u1.cin ;
wire \add_54s_54ns_54_2_1_U18.top_add_54s_54ns_54_2_1_Adder_11_U.u1.cout ;
wire [26:0] \add_54s_54ns_54_2_1_U18.top_add_54s_54ns_54_2_1_Adder_11_U.u1.s ;
wire [26:0] \add_54s_54ns_54_2_1_U18.top_add_54s_54ns_54_2_1_Adder_11_U.u2.a ;
wire [26:0] \add_54s_54ns_54_2_1_U18.top_add_54s_54ns_54_2_1_Adder_11_U.u2.b ;
wire \add_54s_54ns_54_2_1_U18.top_add_54s_54ns_54_2_1_Adder_11_U.u2.cin ;
wire \add_54s_54ns_54_2_1_U18.top_add_54s_54ns_54_2_1_Adder_11_U.u2.cout ;
wire [26:0] \add_54s_54ns_54_2_1_U18.top_add_54s_54ns_54_2_1_Adder_11_U.u2.s ;
wire \add_5ns_5ns_5_2_1_U14.ce ;
wire \add_5ns_5ns_5_2_1_U14.clk ;
wire [4:0] \add_5ns_5ns_5_2_1_U14.din0 ;
wire [4:0] \add_5ns_5ns_5_2_1_U14.din1 ;
wire [4:0] \add_5ns_5ns_5_2_1_U14.dout ;
wire \add_5ns_5ns_5_2_1_U14.reset ;
wire [4:0] \add_5ns_5ns_5_2_1_U14.top_add_5ns_5ns_5_2_1_Adder_9_U.a ;
wire [4:0] \add_5ns_5ns_5_2_1_U14.top_add_5ns_5ns_5_2_1_Adder_9_U.ain_s0 ;
wire [4:0] \add_5ns_5ns_5_2_1_U14.top_add_5ns_5ns_5_2_1_Adder_9_U.b ;
wire [4:0] \add_5ns_5ns_5_2_1_U14.top_add_5ns_5ns_5_2_1_Adder_9_U.bin_s0 ;
wire \add_5ns_5ns_5_2_1_U14.top_add_5ns_5ns_5_2_1_Adder_9_U.ce ;
wire \add_5ns_5ns_5_2_1_U14.top_add_5ns_5ns_5_2_1_Adder_9_U.clk ;
wire \add_5ns_5ns_5_2_1_U14.top_add_5ns_5ns_5_2_1_Adder_9_U.facout_s1 ;
wire \add_5ns_5ns_5_2_1_U14.top_add_5ns_5ns_5_2_1_Adder_9_U.facout_s2 ;
wire [1:0] \add_5ns_5ns_5_2_1_U14.top_add_5ns_5ns_5_2_1_Adder_9_U.fas_s1 ;
wire [2:0] \add_5ns_5ns_5_2_1_U14.top_add_5ns_5ns_5_2_1_Adder_9_U.fas_s2 ;
wire \add_5ns_5ns_5_2_1_U14.top_add_5ns_5ns_5_2_1_Adder_9_U.reset ;
wire [4:0] \add_5ns_5ns_5_2_1_U14.top_add_5ns_5ns_5_2_1_Adder_9_U.s ;
wire [1:0] \add_5ns_5ns_5_2_1_U14.top_add_5ns_5ns_5_2_1_Adder_9_U.u1.a ;
wire [1:0] \add_5ns_5ns_5_2_1_U14.top_add_5ns_5ns_5_2_1_Adder_9_U.u1.b ;
wire \add_5ns_5ns_5_2_1_U14.top_add_5ns_5ns_5_2_1_Adder_9_U.u1.cin ;
wire \add_5ns_5ns_5_2_1_U14.top_add_5ns_5ns_5_2_1_Adder_9_U.u1.cout ;
wire [1:0] \add_5ns_5ns_5_2_1_U14.top_add_5ns_5ns_5_2_1_Adder_9_U.u1.s ;
wire [2:0] \add_5ns_5ns_5_2_1_U14.top_add_5ns_5ns_5_2_1_Adder_9_U.u2.a ;
wire [2:0] \add_5ns_5ns_5_2_1_U14.top_add_5ns_5ns_5_2_1_Adder_9_U.u2.b ;
wire \add_5ns_5ns_5_2_1_U14.top_add_5ns_5ns_5_2_1_Adder_9_U.u2.cin ;
wire \add_5ns_5ns_5_2_1_U14.top_add_5ns_5ns_5_2_1_Adder_9_U.u2.cout ;
wire [2:0] \add_5ns_5ns_5_2_1_U14.top_add_5ns_5ns_5_2_1_Adder_9_U.u2.s ;
wire \add_5s_5ns_5_2_1_U2.ce ;
wire \add_5s_5ns_5_2_1_U2.clk ;
wire [4:0] \add_5s_5ns_5_2_1_U2.din0 ;
wire [4:0] \add_5s_5ns_5_2_1_U2.din1 ;
wire [4:0] \add_5s_5ns_5_2_1_U2.dout ;
wire \add_5s_5ns_5_2_1_U2.reset ;
wire [4:0] \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.a ;
wire [4:0] \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.ain_s0 ;
wire [4:0] \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.b ;
wire [4:0] \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.bin_s0 ;
wire \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.ce ;
wire \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.clk ;
wire \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.facout_s1 ;
wire \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.facout_s2 ;
wire [1:0] \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.fas_s1 ;
wire [2:0] \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.fas_s2 ;
wire \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.reset ;
wire [4:0] \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.s ;
wire [1:0] \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.u1.a ;
wire [1:0] \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.u1.b ;
wire \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.u1.cin ;
wire \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.u1.cout ;
wire [1:0] \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.u1.s ;
wire [2:0] \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.u2.a ;
wire [2:0] \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.u2.b ;
wire \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.u2.cin ;
wire \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.u2.cout ;
wire [2:0] \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.u2.s ;
wire \add_63s_63s_63_2_1_U7.ce ;
wire \add_63s_63s_63_2_1_U7.clk ;
wire [62:0] \add_63s_63s_63_2_1_U7.din0 ;
wire [62:0] \add_63s_63s_63_2_1_U7.din1 ;
wire [62:0] \add_63s_63s_63_2_1_U7.dout ;
wire \add_63s_63s_63_2_1_U7.reset ;
wire [62:0] \add_63s_63s_63_2_1_U7.top_add_63s_63s_63_2_1_Adder_5_U.a ;
wire [62:0] \add_63s_63s_63_2_1_U7.top_add_63s_63s_63_2_1_Adder_5_U.ain_s0 ;
wire [62:0] \add_63s_63s_63_2_1_U7.top_add_63s_63s_63_2_1_Adder_5_U.b ;
wire [62:0] \add_63s_63s_63_2_1_U7.top_add_63s_63s_63_2_1_Adder_5_U.bin_s0 ;
wire \add_63s_63s_63_2_1_U7.top_add_63s_63s_63_2_1_Adder_5_U.ce ;
wire \add_63s_63s_63_2_1_U7.top_add_63s_63s_63_2_1_Adder_5_U.clk ;
wire \add_63s_63s_63_2_1_U7.top_add_63s_63s_63_2_1_Adder_5_U.facout_s1 ;
wire \add_63s_63s_63_2_1_U7.top_add_63s_63s_63_2_1_Adder_5_U.facout_s2 ;
wire [30:0] \add_63s_63s_63_2_1_U7.top_add_63s_63s_63_2_1_Adder_5_U.fas_s1 ;
wire [31:0] \add_63s_63s_63_2_1_U7.top_add_63s_63s_63_2_1_Adder_5_U.fas_s2 ;
wire \add_63s_63s_63_2_1_U7.top_add_63s_63s_63_2_1_Adder_5_U.reset ;
wire [62:0] \add_63s_63s_63_2_1_U7.top_add_63s_63s_63_2_1_Adder_5_U.s ;
wire [30:0] \add_63s_63s_63_2_1_U7.top_add_63s_63s_63_2_1_Adder_5_U.u1.a ;
wire [30:0] \add_63s_63s_63_2_1_U7.top_add_63s_63s_63_2_1_Adder_5_U.u1.b ;
wire \add_63s_63s_63_2_1_U7.top_add_63s_63s_63_2_1_Adder_5_U.u1.cin ;
wire \add_63s_63s_63_2_1_U7.top_add_63s_63s_63_2_1_Adder_5_U.u1.cout ;
wire [30:0] \add_63s_63s_63_2_1_U7.top_add_63s_63s_63_2_1_Adder_5_U.u1.s ;
wire [31:0] \add_63s_63s_63_2_1_U7.top_add_63s_63s_63_2_1_Adder_5_U.u2.a ;
wire [31:0] \add_63s_63s_63_2_1_U7.top_add_63s_63s_63_2_1_Adder_5_U.u2.b ;
wire \add_63s_63s_63_2_1_U7.top_add_63s_63s_63_2_1_Adder_5_U.u2.cin ;
wire \add_63s_63s_63_2_1_U7.top_add_63s_63s_63_2_1_Adder_5_U.u2.cout ;
wire [31:0] \add_63s_63s_63_2_1_U7.top_add_63s_63s_63_2_1_Adder_5_U.u2.s ;
wire and_ln340_1_fu_493_p2;
wire and_ln340_2_fu_505_p2;
wire and_ln340_fu_304_p2;
wire and_ln353_fu_938_p2;
wire and_ln785_1_fu_331_p2;
wire and_ln785_3_fu_561_p2;
wire and_ln785_4_fu_509_p2;
wire and_ln785_fu_325_p2;
wire and_ln786_fu_422_p2;
wire ap_CS_fsm_state1;
wire ap_CS_fsm_state10;
wire ap_CS_fsm_state11;
wire ap_CS_fsm_state12;
wire ap_CS_fsm_state13;
wire ap_CS_fsm_state14;
wire ap_CS_fsm_state15;
wire ap_CS_fsm_state16;
wire ap_CS_fsm_state17;
wire ap_CS_fsm_state18;
wire ap_CS_fsm_state19;
wire ap_CS_fsm_state2;
wire ap_CS_fsm_state20;
wire ap_CS_fsm_state21;
wire ap_CS_fsm_state22;
wire ap_CS_fsm_state23;
wire ap_CS_fsm_state24;
wire ap_CS_fsm_state25;
wire ap_CS_fsm_state26;
wire ap_CS_fsm_state27;
wire ap_CS_fsm_state28;
wire ap_CS_fsm_state29;
wire ap_CS_fsm_state3;
wire ap_CS_fsm_state30;
wire ap_CS_fsm_state31;
wire ap_CS_fsm_state32;
wire ap_CS_fsm_state33;
wire ap_CS_fsm_state34;
wire ap_CS_fsm_state35;
wire ap_CS_fsm_state36;
wire ap_CS_fsm_state37;
wire ap_CS_fsm_state4;
wire ap_CS_fsm_state5;
wire ap_CS_fsm_state6;
wire ap_CS_fsm_state7;
wire ap_CS_fsm_state8;
wire ap_CS_fsm_state9;
wire [36:0] ap_NS_fsm;
wire ap_clk;
wire ap_done;
wire ap_idle;
wire ap_ready;
wire ap_rst;
wire ap_start;
wire [53:0] grp_fu_1034_p0;
wire [53:0] grp_fu_1034_p1;
wire [53:0] grp_fu_1034_p2;
wire [31:0] grp_fu_1055_p2;
wire [46:0] grp_fu_1094_p0;
wire [46:0] grp_fu_1094_p1;
wire [46:0] grp_fu_1094_p2;
wire [31:0] grp_fu_1120_p2;
wire [4:0] grp_fu_201_p0;
wire [4:0] grp_fu_201_p1;
wire [4:0] grp_fu_201_p2;
wire [4:0] grp_fu_434_p0;
wire [4:0] grp_fu_434_p1;
wire [4:0] grp_fu_434_p2;
wire [1:0] grp_fu_536_p1;
wire [1:0] grp_fu_536_p2;
wire [4:0] grp_fu_647_p0;
wire [4:0] grp_fu_647_p1;
wire [4:0] grp_fu_647_p2;
wire [15:0] grp_fu_704_p0;
wire [19:0] grp_fu_704_p00;
wire [19:0] grp_fu_704_p2;
wire [3:0] grp_fu_757_p0;
wire [3:0] grp_fu_757_p2;
wire [62:0] grp_fu_778_p0;
wire [62:0] grp_fu_778_p1;
wire [62:0] grp_fu_778_p2;
wire [31:0] grp_fu_825_p2;
wire [31:0] grp_fu_830_p2;
wire [32:0] grp_fu_842_p0;
wire [32:0] grp_fu_842_p1;
wire [32:0] grp_fu_842_p2;
wire [10:0] grp_fu_855_p0;
wire [10:0] grp_fu_855_p1;
wire [10:0] grp_fu_855_p2;
wire [4:0] grp_fu_864_p1;
wire [4:0] grp_fu_864_p2;
wire [31:0] grp_fu_910_p2;
wire [4:0] grp_fu_914_p1;
wire [4:0] grp_fu_914_p2;
wire [31:0] grp_fu_965_p0;
wire [31:0] grp_fu_965_p2;
wire [31:0] grp_fu_977_p2;
wire [31:0] grp_fu_984_p1;
wire [31:0] grp_fu_984_p2;
wire icmp_ln1498_fu_688_p2;
wire icmp_ln768_1_fu_225_p2;
wire icmp_ln768_2_fu_902_p2;
wire icmp_ln768_3_fu_580_p2;
wire icmp_ln768_fu_259_p2;
wire icmp_ln786_1_fu_231_p2;
wire icmp_ln786_2_fu_585_p2;
wire icmp_ln786_fu_264_p2;
wire icmp_ln790_fu_621_p2;
wire icmp_ln850_fu_919_p2;
wire icmp_ln851_1_fu_784_p2;
wire icmp_ln851_2_fu_1040_p2;
wire icmp_ln851_3_fu_1104_p2;
wire icmp_ln851_fu_752_p2;
wire lhs_V_3_fu_393_p2;
wire [61:0] lhs_V_4_fu_763_p3;
wire \mul_16ns_4s_20_7_1_U5.ce ;
wire \mul_16ns_4s_20_7_1_U5.clk ;
wire [15:0] \mul_16ns_4s_20_7_1_U5.din0 ;
wire [3:0] \mul_16ns_4s_20_7_1_U5.din1 ;
wire [19:0] \mul_16ns_4s_20_7_1_U5.dout ;
wire \mul_16ns_4s_20_7_1_U5.reset ;
wire [15:0] \mul_16ns_4s_20_7_1_U5.top_mul_16ns_4s_20_7_1_Mul_DSP_0_U.a ;
wire [3:0] \mul_16ns_4s_20_7_1_U5.top_mul_16ns_4s_20_7_1_Mul_DSP_0_U.b ;
wire \mul_16ns_4s_20_7_1_U5.top_mul_16ns_4s_20_7_1_Mul_DSP_0_U.ce ;
wire \mul_16ns_4s_20_7_1_U5.top_mul_16ns_4s_20_7_1_Mul_DSP_0_U.clk ;
wire [19:0] \mul_16ns_4s_20_7_1_U5.top_mul_16ns_4s_20_7_1_Mul_DSP_0_U.p ;
wire [19:0] \mul_16ns_4s_20_7_1_U5.top_mul_16ns_4s_20_7_1_Mul_DSP_0_U.tmp_product ;
wire newsignbit_fu_245_p1;
wire [3:0] op_0;
wire [3:0] op_1;
wire [31:0] op_12_V_fu_738_p3;
wire [3:0] op_16_V_fu_957_p1;
wire op_16_V_fu_957_p2;
wire [31:0] op_18_V_fu_1008_p3;
wire [15:0] op_19;
wire [31:0] op_27;
wire op_27_ap_vld;
wire op_2_V_fu_368_p3;
wire [3:0] op_4_V_fu_594_p3;
wire [31:0] op_7;
wire [3:0] op_8;
wire [31:0] op_9;
wire or_ln340_1_fu_412_p2;
wire or_ln340_fu_293_p2;
wire or_ln384_fu_673_p2;
wire or_ln785_1_fu_384_p2;
wire or_ln785_2_fu_320_p2;
wire or_ln785_3_fu_599_p2;
wire or_ln785_4_fu_556_p2;
wire or_ln785_5_fu_513_p2;
wire or_ln785_fu_269_p2;
wire or_ln786_1_fu_407_p2;
wire or_ln786_fu_288_p2;
wire or_ln788_1_fu_663_p2;
wire or_ln788_fu_658_p2;
wire overflow_1_fu_398_p2;
wire overflow_2_fu_1003_p2;
wire overflow_3_fu_608_p2;
wire overflow_fu_278_p2;
wire p_Result_10_fu_879_p3;
wire p_Result_11_fu_1060_p3;
wire p_Result_12_fu_1125_p3;
wire p_Result_14_fu_336_p3;
wire [3:0] p_Result_15_fu_207_p1;
wire p_Result_16_fu_378_p2;
wire [3:0] p_Result_17_fu_447_p1;
wire p_Result_17_fu_447_p3;
wire p_Result_18_fu_996_p3;
wire [3:0] p_Result_1_fu_215_p1;
wire [2:0] p_Result_1_fu_215_p4;
wire p_Result_3_fu_931_p3;
wire p_Result_6_fu_806_p3;
wire [30:0] p_Result_8_fu_614_p3;
wire [3:0] p_Result_s_16_fu_478_p4;
wire [31:0] p_Val2_11_fu_724_p3;
wire p_Val2_1_fu_283_p2;
wire [3:0] p_Val2_2_fu_373_p0;
wire [3:0] p_Val2_2_fu_373_p2;
wire [2:0] p_Val2_3_fu_473_p2;
wire [31:0] p_Val2_7_fu_989_p3;
wire [3:0] ret_V_11_fu_627_p2;
wire [3:0] ret_V_11_fu_627_p3;
wire ret_V_13_fu_943_p2;
wire [31:0] ret_V_16_fu_891_p3;
wire [3:0] ret_V_fu_818_p3;
wire [2:0] rhs_1_fu_636_p3;
wire [52:0] rhs_4_fu_1023_p3;
wire [45:0] rhs_5_fu_1083_p3;
wire sel_tmp18_fu_519_p2;
wire [31:0] select_ln1192_1_fu_970_p3;
wire [31:0] select_ln1192_fu_799_p3;
wire [3:0] select_ln340_1_fu_498_p3;
wire select_ln340_fu_362_p3;
wire [31:0] select_ln353_fu_1072_p3;
wire select_ln365_fu_355_p3;
wire [31:0] select_ln384_fu_731_p3;
wire [3:0] select_ln785_fu_566_p3;
wire [31:0] select_ln850_1_fu_886_p3;
wire [31:0] select_ln850_2_fu_1067_p3;
wire [31:0] select_ln850_3_fu_1132_p3;
wire [3:0] select_ln850_fu_813_p3;
wire [3:0] select_ln874_fu_949_p3;
wire [15:0] sext_ln1118_fu_697_p1;
wire [3:0] sext_ln1346_fu_430_p0;
wire [4:0] sext_ln1346_fu_430_p1;
wire [3:0] sext_ln1347_fu_197_p0;
wire [15:0] sext_ln703_1_fu_1079_p0;
wire [5:0] sext_ln727_fu_678_p1;
wire [3:0] sext_ln850_fu_749_p1;
wire [3:0] shl_ln_fu_681_p1;
wire [5:0] shl_ln_fu_681_p3;
wire \sub_5s_5ns_5_2_1_U4.ce ;
wire \sub_5s_5ns_5_2_1_U4.clk ;
wire [4:0] \sub_5s_5ns_5_2_1_U4.din0 ;
wire [4:0] \sub_5s_5ns_5_2_1_U4.din1 ;
wire [4:0] \sub_5s_5ns_5_2_1_U4.dout ;
wire \sub_5s_5ns_5_2_1_U4.reset ;
wire [4:0] \sub_5s_5ns_5_2_1_U4.top_sub_5s_5ns_5_2_1_Adder_3_U.a ;
wire [4:0] \sub_5s_5ns_5_2_1_U4.top_sub_5s_5ns_5_2_1_Adder_3_U.ain_s0 ;
wire [4:0] \sub_5s_5ns_5_2_1_U4.top_sub_5s_5ns_5_2_1_Adder_3_U.b ;
wire [4:0] \sub_5s_5ns_5_2_1_U4.top_sub_5s_5ns_5_2_1_Adder_3_U.bin_s0 ;
wire \sub_5s_5ns_5_2_1_U4.top_sub_5s_5ns_5_2_1_Adder_3_U.ce ;
wire \sub_5s_5ns_5_2_1_U4.top_sub_5s_5ns_5_2_1_Adder_3_U.clk ;
wire \sub_5s_5ns_5_2_1_U4.top_sub_5s_5ns_5_2_1_Adder_3_U.facout_s1 ;
wire \sub_5s_5ns_5_2_1_U4.top_sub_5s_5ns_5_2_1_Adder_3_U.facout_s2 ;
wire [1:0] \sub_5s_5ns_5_2_1_U4.top_sub_5s_5ns_5_2_1_Adder_3_U.fas_s1 ;
wire [2:0] \sub_5s_5ns_5_2_1_U4.top_sub_5s_5ns_5_2_1_Adder_3_U.fas_s2 ;
wire \sub_5s_5ns_5_2_1_U4.top_sub_5s_5ns_5_2_1_Adder_3_U.reset ;
wire [4:0] \sub_5s_5ns_5_2_1_U4.top_sub_5s_5ns_5_2_1_Adder_3_U.s ;
wire [1:0] \sub_5s_5ns_5_2_1_U4.top_sub_5s_5ns_5_2_1_Adder_3_U.u1.a ;
wire [1:0] \sub_5s_5ns_5_2_1_U4.top_sub_5s_5ns_5_2_1_Adder_3_U.u1.b ;
wire \sub_5s_5ns_5_2_1_U4.top_sub_5s_5ns_5_2_1_Adder_3_U.u1.cin ;
wire \sub_5s_5ns_5_2_1_U4.top_sub_5s_5ns_5_2_1_Adder_3_U.u1.cout ;
wire [1:0] \sub_5s_5ns_5_2_1_U4.top_sub_5s_5ns_5_2_1_Adder_3_U.u1.s ;
wire [2:0] \sub_5s_5ns_5_2_1_U4.top_sub_5s_5ns_5_2_1_Adder_3_U.u2.a ;
wire [2:0] \sub_5s_5ns_5_2_1_U4.top_sub_5s_5ns_5_2_1_Adder_3_U.u2.b ;
wire \sub_5s_5ns_5_2_1_U4.top_sub_5s_5ns_5_2_1_Adder_3_U.u2.cin ;
wire \sub_5s_5ns_5_2_1_U4.top_sub_5s_5ns_5_2_1_Adder_3_U.u2.cout ;
wire [2:0] \sub_5s_5ns_5_2_1_U4.top_sub_5s_5ns_5_2_1_Adder_3_U.u2.s ;
wire \sub_5s_5s_5_2_1_U1.ce ;
wire \sub_5s_5s_5_2_1_U1.clk ;
wire [4:0] \sub_5s_5s_5_2_1_U1.din0 ;
wire [4:0] \sub_5s_5s_5_2_1_U1.din1 ;
wire [4:0] \sub_5s_5s_5_2_1_U1.dout ;
wire \sub_5s_5s_5_2_1_U1.reset ;
wire [4:0] \sub_5s_5s_5_2_1_U1.top_sub_5s_5s_5_2_1_Adder_0_U.a ;
wire [4:0] \sub_5s_5s_5_2_1_U1.top_sub_5s_5s_5_2_1_Adder_0_U.ain_s0 ;
wire [4:0] \sub_5s_5s_5_2_1_U1.top_sub_5s_5s_5_2_1_Adder_0_U.b ;
wire [4:0] \sub_5s_5s_5_2_1_U1.top_sub_5s_5s_5_2_1_Adder_0_U.bin_s0 ;
wire \sub_5s_5s_5_2_1_U1.top_sub_5s_5s_5_2_1_Adder_0_U.ce ;
wire \sub_5s_5s_5_2_1_U1.top_sub_5s_5s_5_2_1_Adder_0_U.clk ;
wire \sub_5s_5s_5_2_1_U1.top_sub_5s_5s_5_2_1_Adder_0_U.facout_s1 ;
wire \sub_5s_5s_5_2_1_U1.top_sub_5s_5s_5_2_1_Adder_0_U.facout_s2 ;
wire [1:0] \sub_5s_5s_5_2_1_U1.top_sub_5s_5s_5_2_1_Adder_0_U.fas_s1 ;
wire [2:0] \sub_5s_5s_5_2_1_U1.top_sub_5s_5s_5_2_1_Adder_0_U.fas_s2 ;
wire \sub_5s_5s_5_2_1_U1.top_sub_5s_5s_5_2_1_Adder_0_U.reset ;
wire [4:0] \sub_5s_5s_5_2_1_U1.top_sub_5s_5s_5_2_1_Adder_0_U.s ;
wire [1:0] \sub_5s_5s_5_2_1_U1.top_sub_5s_5s_5_2_1_Adder_0_U.u1.a ;
wire [1:0] \sub_5s_5s_5_2_1_U1.top_sub_5s_5s_5_2_1_Adder_0_U.u1.b ;
wire \sub_5s_5s_5_2_1_U1.top_sub_5s_5s_5_2_1_Adder_0_U.u1.cin ;
wire \sub_5s_5s_5_2_1_U1.top_sub_5s_5s_5_2_1_Adder_0_U.u1.cout ;
wire [1:0] \sub_5s_5s_5_2_1_U1.top_sub_5s_5s_5_2_1_Adder_0_U.u1.s ;
wire [2:0] \sub_5s_5s_5_2_1_U1.top_sub_5s_5s_5_2_1_Adder_0_U.u2.a ;
wire [2:0] \sub_5s_5s_5_2_1_U1.top_sub_5s_5s_5_2_1_Adder_0_U.u2.b ;
wire \sub_5s_5s_5_2_1_U1.top_sub_5s_5s_5_2_1_Adder_0_U.u2.cin ;
wire \sub_5s_5s_5_2_1_U1.top_sub_5s_5s_5_2_1_Adder_0_U.u2.cout ;
wire [2:0] \sub_5s_5s_5_2_1_U1.top_sub_5s_5s_5_2_1_Adder_0_U.u2.s ;
wire \sub_5s_5s_5_2_1_U12.ce ;
wire \sub_5s_5s_5_2_1_U12.clk ;
wire [4:0] \sub_5s_5s_5_2_1_U12.din0 ;
wire [4:0] \sub_5s_5s_5_2_1_U12.din1 ;
wire [4:0] \sub_5s_5s_5_2_1_U12.dout ;
wire \sub_5s_5s_5_2_1_U12.reset ;
wire [4:0] \sub_5s_5s_5_2_1_U12.top_sub_5s_5s_5_2_1_Adder_0_U.a ;
wire [4:0] \sub_5s_5s_5_2_1_U12.top_sub_5s_5s_5_2_1_Adder_0_U.ain_s0 ;
wire [4:0] \sub_5s_5s_5_2_1_U12.top_sub_5s_5s_5_2_1_Adder_0_U.b ;
wire [4:0] \sub_5s_5s_5_2_1_U12.top_sub_5s_5s_5_2_1_Adder_0_U.bin_s0 ;
wire \sub_5s_5s_5_2_1_U12.top_sub_5s_5s_5_2_1_Adder_0_U.ce ;
wire \sub_5s_5s_5_2_1_U12.top_sub_5s_5s_5_2_1_Adder_0_U.clk ;
wire \sub_5s_5s_5_2_1_U12.top_sub_5s_5s_5_2_1_Adder_0_U.facout_s1 ;
wire \sub_5s_5s_5_2_1_U12.top_sub_5s_5s_5_2_1_Adder_0_U.facout_s2 ;
wire [1:0] \sub_5s_5s_5_2_1_U12.top_sub_5s_5s_5_2_1_Adder_0_U.fas_s1 ;
wire [2:0] \sub_5s_5s_5_2_1_U12.top_sub_5s_5s_5_2_1_Adder_0_U.fas_s2 ;
wire \sub_5s_5s_5_2_1_U12.top_sub_5s_5s_5_2_1_Adder_0_U.reset ;
wire [4:0] \sub_5s_5s_5_2_1_U12.top_sub_5s_5s_5_2_1_Adder_0_U.s ;
wire [1:0] \sub_5s_5s_5_2_1_U12.top_sub_5s_5s_5_2_1_Adder_0_U.u1.a ;
wire [1:0] \sub_5s_5s_5_2_1_U12.top_sub_5s_5s_5_2_1_Adder_0_U.u1.b ;
wire \sub_5s_5s_5_2_1_U12.top_sub_5s_5s_5_2_1_Adder_0_U.u1.cin ;
wire \sub_5s_5s_5_2_1_U12.top_sub_5s_5s_5_2_1_Adder_0_U.u1.cout ;
wire [1:0] \sub_5s_5s_5_2_1_U12.top_sub_5s_5s_5_2_1_Adder_0_U.u1.s ;
wire [2:0] \sub_5s_5s_5_2_1_U12.top_sub_5s_5s_5_2_1_Adder_0_U.u2.a ;
wire [2:0] \sub_5s_5s_5_2_1_U12.top_sub_5s_5s_5_2_1_Adder_0_U.u2.b ;
wire \sub_5s_5s_5_2_1_U12.top_sub_5s_5s_5_2_1_Adder_0_U.u2.cin ;
wire \sub_5s_5s_5_2_1_U12.top_sub_5s_5s_5_2_1_Adder_0_U.u2.cout ;
wire [2:0] \sub_5s_5s_5_2_1_U12.top_sub_5s_5s_5_2_1_Adder_0_U.u2.s ;
wire [3:0] tmp_5_fu_454_p1;
wire tmp_5_fu_454_p3;
wire tmp_7_fu_924_p3;
wire tmp_fu_343_p3;
wire [3:0] trunc_ln731_2_fu_440_p0;
wire [1:0] trunc_ln731_2_fu_440_p1;
wire [3:0] trunc_ln731_fu_444_p0;
wire trunc_ln731_fu_444_p1;
wire trunc_ln790_fu_590_p1;
wire [1:0] trunc_ln851_1_fu_720_p1;
wire [29:0] trunc_ln851_2_fu_745_p1;
wire [20:0] trunc_ln851_3_fu_1016_p1;
wire [15:0] trunc_ln851_4_fu_1100_p0;
wire [13:0] trunc_ln851_4_fu_1100_p1;
wire [1:0] trunc_ln851_fu_898_p1;
wire underflow_2_fu_668_p2;
wire xor_ln340_1_fu_488_p2;
wire xor_ln340_fu_298_p2;
wire xor_ln365_1_fu_461_p2;
wire xor_ln365_2_fu_467_p2;
wire xor_ln365_fu_350_p2;
wire xor_ln785_1_fu_388_p2;
wire xor_ln785_2_fu_603_p2;
wire xor_ln785_3_fu_315_p2;
wire xor_ln785_4_fu_551_p2;
wire xor_ln785_fu_273_p2;
wire xor_ln786_1_fu_653_p2;
wire xor_ln786_3_fu_310_p2;
wire xor_ln786_4_fu_417_p2;
wire xor_ln786_fu_402_p2;


assign _083_ = icmp_ln851_1_reg_1490 & ap_CS_fsm[17];
assign _084_ = icmp_ln851_2_reg_1674 & ap_CS_fsm[30];
assign _085_ = icmp_ln851_3_reg_1711 & ap_CS_fsm[35];
assign _086_ = ap_CS_fsm[5] & _090_;
assign _087_ = ap_CS_fsm[10] & _091_;
assign _088_ = _092_ & ap_CS_fsm[0];
assign _089_ = ap_start & ap_CS_fsm[0];
assign and_ln340_1_fu_493_p2 = xor_ln340_1_fu_488_p2 & or_ln786_1_reg_1292;
assign and_ln340_2_fu_505_p2 = or_ln786_1_reg_1292 & or_ln340_1_reg_1298;
assign and_ln340_fu_304_p2 = xor_ln340_fu_298_p2 & or_ln786_fu_288_p2;
assign and_ln353_fu_938_p2 = r_V_reg_1583[19] & icmp_ln850_reg_1604;
assign and_ln785_1_fu_331_p2 = newsignbit_reg_1195 & and_ln785_fu_325_p2;
assign and_ln785_3_fu_561_p2 = or_ln785_4_fu_556_p2 & and_ln786_reg_1304;
assign and_ln785_4_fu_509_p2 = xor_ln785_1_reg_1272 & and_ln786_reg_1304;
assign and_ln785_fu_325_p2 = xor_ln786_3_fu_310_p2 & or_ln785_2_fu_320_p2;
assign and_ln786_fu_422_p2 = xor_ln786_4_fu_417_p2 & p_Result_16_reg_1259;
assign overflow_1_fu_398_p2 = xor_ln785_1_reg_1272 & or_ln785_1_reg_1266;
assign overflow_3_fu_608_p2 = xor_ln785_2_fu_603_p2 & or_ln785_3_fu_599_p2;
assign overflow_fu_278_p2 = xor_ln785_fu_273_p2 & or_ln785_reg_1223;
assign sel_tmp18_fu_519_p2 = xor_ln365_2_fu_467_p2 & or_ln785_5_fu_513_p2;
assign underflow_2_fu_668_p2 = p_Result_19_reg_1336 & or_ln788_1_fu_663_p2;
assign xor_ln340_1_fu_488_p2 = ~ or_ln340_1_reg_1298;
assign p_Val2_1_fu_283_p2 = ~ newsignbit_reg_1195;
assign xor_ln785_fu_273_p2 = ~ p_Result_13_reg_1188;
assign xor_ln340_fu_298_p2 = ~ or_ln340_fu_293_p2;
assign xor_ln785_3_fu_315_p2 = ~ or_ln785_reg_1223;
assign xor_ln786_3_fu_310_p2 = ~ icmp_ln786_reg_1217;
assign xor_ln785_4_fu_551_p2 = ~ or_ln785_1_reg_1266;
assign xor_ln786_4_fu_417_p2 = ~ icmp_ln786_1_reg_1176;
assign lhs_V_3_fu_393_p2 = ~ op_2_V_reg_1244;
assign xor_ln786_1_fu_653_p2 = ~ p_Result_20_reg_1363;
assign xor_ln786_fu_402_p2 = ~ p_Result_16_reg_1259;
assign xor_ln785_2_fu_603_p2 = ~ p_Result_19_reg_1336;
assign xor_ln365_2_fu_467_p2 = ~ xor_ln365_1_fu_461_p2;
assign xor_ln785_1_fu_388_p2 = ~ p_Result_15_reg_1164;
assign p_Val2_3_fu_473_p2 = ~ p_Val2_2_reg_1251[2:0];
assign _090_ = ~ and_ln785_1_reg_1234;
assign _091_ = ~ sel_tmp18_reg_1331;
assign _092_ = ~ ap_start;
assign _093_ = { op_4_V_reg_1384[3], op_4_V_reg_1384[3], op_4_V_reg_1384 } == { op_8, 2'h0 };
assign _094_ = ! { trunc_ln790_reg_1379, 30'h00000000 };
always @(posedge \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_8_U.clk )
\add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_8_U.bin_s1  <= _096_;
always @(posedge \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_8_U.clk )
\add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_8_U.ain_s1  <= _095_;
always @(posedge \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_8_U.clk )
\add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_8_U.sum_s1  <= _098_;
always @(posedge \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_8_U.clk )
\add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_8_U.carry_s1  <= _097_;
assign _096_ = \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_8_U.ce  ? \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_8_U.b [10:5] : \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_8_U.bin_s1 ;
assign _095_ = \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_8_U.ce  ? \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_8_U.a [10:5] : \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_8_U.ain_s1 ;
assign _097_ = \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_8_U.ce  ? \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_8_U.facout_s1  : \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_8_U.carry_s1 ;
assign _098_ = \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_8_U.ce  ? \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_8_U.fas_s1  : \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_8_U.sum_s1 ;
assign _099_ = \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_8_U.u1.a  + \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_8_U.u1.b ;
assign { \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_8_U.u1.cout , \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_8_U.u1.s  } = _099_ + \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_8_U.u1.cin ;
assign _100_ = \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_8_U.u2.a  + \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_8_U.u2.b ;
assign { \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_8_U.u2.cout , \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_8_U.u2.s  } = _100_ + \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_8_U.u2.cin ;
always @(posedge \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_2_U.clk )
\add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_2_U.bin_s1  <= _102_;
always @(posedge \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_2_U.clk )
\add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_2_U.ain_s1  <= _101_;
always @(posedge \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_2_U.clk )
\add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_2_U.sum_s1  <= _104_;
always @(posedge \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_2_U.clk )
\add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_2_U.carry_s1  <= _103_;
assign _102_ = \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_2_U.ce  ? \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_2_U.b [1] : \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_2_U.bin_s1 ;
assign _101_ = \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_2_U.ce  ? \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_2_U.a [1] : \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_2_U.ain_s1 ;
assign _103_ = \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_2_U.ce  ? \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_2_U.facout_s1  : \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_2_U.carry_s1 ;
assign _104_ = \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_2_U.ce  ? \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_2_U.fas_s1  : \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_2_U.sum_s1 ;
assign _105_ = \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_2_U.u1.a  + \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_2_U.u1.b ;
assign { \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_2_U.u1.cout , \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_2_U.u1.s  } = _105_ + \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_2_U.u1.cin ;
assign _106_ = \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_2_U.u2.a  + \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_2_U.u2.b ;
assign { \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_2_U.u2.cout , \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_2_U.u2.s  } = _106_ + \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_2_U.u2.cin ;
always @(posedge \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.clk )
\add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s1  <= _108_;
always @(posedge \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.clk )
\add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s1  <= _107_;
always @(posedge \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.clk )
\add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.sum_s1  <= _110_;
always @(posedge \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.clk )
\add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.carry_s1  <= _109_;
assign _108_ = \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  ? \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.b [31:16] : \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s1 ;
assign _107_ = \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  ? \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.a [31:16] : \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s1 ;
assign _109_ = \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  ? \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s1  : \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.carry_s1 ;
assign _110_ = \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  ? \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s1  : \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.sum_s1 ;
assign _111_ = \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.a  + \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.b ;
assign { \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cout , \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.s  } = _111_ + \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cin ;
assign _112_ = \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.a  + \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.b ;
assign { \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cout , \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.s  } = _112_ + \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cin ;
always @(posedge \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.clk )
\add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s1  <= _114_;
always @(posedge \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.clk )
\add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s1  <= _113_;
always @(posedge \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.clk )
\add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.sum_s1  <= _116_;
always @(posedge \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.clk )
\add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.carry_s1  <= _115_;
assign _114_ = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  ? \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.b [31:16] : \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s1 ;
assign _113_ = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  ? \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.a [31:16] : \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s1 ;
assign _115_ = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  ? \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s1  : \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.carry_s1 ;
assign _116_ = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  ? \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s1  : \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.sum_s1 ;
assign _117_ = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.a  + \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.b ;
assign { \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cout , \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.s  } = _117_ + \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cin ;
assign _118_ = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.a  + \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.b ;
assign { \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cout , \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.s  } = _118_ + \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cin ;
always @(posedge \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.clk )
\add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s1  <= _120_;
always @(posedge \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.clk )
\add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s1  <= _119_;
always @(posedge \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.clk )
\add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.sum_s1  <= _122_;
always @(posedge \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.clk )
\add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.carry_s1  <= _121_;
assign _120_ = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  ? \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.b [31:16] : \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s1 ;
assign _119_ = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  ? \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.a [31:16] : \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s1 ;
assign _121_ = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  ? \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s1  : \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.carry_s1 ;
assign _122_ = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  ? \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s1  : \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.sum_s1 ;
assign _123_ = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.a  + \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.b ;
assign { \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cout , \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.s  } = _123_ + \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cin ;
assign _124_ = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.a  + \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.b ;
assign { \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cout , \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.s  } = _124_ + \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cin ;
always @(posedge \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_6_U.clk )
\add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s1  <= _126_;
always @(posedge \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_6_U.clk )
\add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s1  <= _125_;
always @(posedge \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_6_U.clk )
\add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_6_U.sum_s1  <= _128_;
always @(posedge \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_6_U.clk )
\add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_6_U.carry_s1  <= _127_;
assign _126_ = \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  ? \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_6_U.b [31:16] : \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s1 ;
assign _125_ = \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  ? \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_6_U.a [31:16] : \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s1 ;
assign _127_ = \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  ? \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s1  : \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_6_U.carry_s1 ;
assign _128_ = \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  ? \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s1  : \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_6_U.sum_s1 ;
assign _129_ = \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.a  + \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.b ;
assign { \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cout , \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.s  } = _129_ + \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cin ;
assign _130_ = \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.a  + \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.b ;
assign { \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cout , \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.s  } = _130_ + \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cin ;
always @(posedge \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_6_U.clk )
\add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s1  <= _132_;
always @(posedge \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_6_U.clk )
\add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s1  <= _131_;
always @(posedge \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_6_U.clk )
\add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_6_U.sum_s1  <= _134_;
always @(posedge \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_6_U.clk )
\add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_6_U.carry_s1  <= _133_;
assign _132_ = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  ? \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_6_U.b [31:16] : \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s1 ;
assign _131_ = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  ? \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_6_U.a [31:16] : \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s1 ;
assign _133_ = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  ? \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s1  : \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_6_U.carry_s1 ;
assign _134_ = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  ? \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s1  : \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_6_U.sum_s1 ;
assign _135_ = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.a  + \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.b ;
assign { \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cout , \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.s  } = _135_ + \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cin ;
assign _136_ = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.a  + \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.b ;
assign { \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cout , \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.s  } = _136_ + \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cin ;
always @(posedge \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.clk )
\add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s1  <= _138_;
always @(posedge \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.clk )
\add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s1  <= _137_;
always @(posedge \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.clk )
\add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.sum_s1  <= _140_;
always @(posedge \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.clk )
\add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.carry_s1  <= _139_;
assign _138_ = \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  ? \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.b [31:16] : \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s1 ;
assign _137_ = \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  ? \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.a [31:16] : \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s1 ;
assign _139_ = \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  ? \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s1  : \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.carry_s1 ;
assign _140_ = \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  ? \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s1  : \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.sum_s1 ;
assign _141_ = \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.a  + \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.b ;
assign { \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cout , \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.s  } = _141_ + \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cin ;
assign _142_ = \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.a  + \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.b ;
assign { \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cout , \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.s  } = _142_ + \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cin ;
always @(posedge \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.clk )
\add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s1  <= _144_;
always @(posedge \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.clk )
\add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s1  <= _143_;
always @(posedge \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.clk )
\add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.sum_s1  <= _146_;
always @(posedge \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.clk )
\add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.carry_s1  <= _145_;
assign _144_ = \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  ? \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.b [31:16] : \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s1 ;
assign _143_ = \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  ? \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.a [31:16] : \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s1 ;
assign _145_ = \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  ? \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s1  : \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.carry_s1 ;
assign _146_ = \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  ? \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s1  : \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.sum_s1 ;
assign _147_ = \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.a  + \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.b ;
assign { \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cout , \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.s  } = _147_ + \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cin ;
assign _148_ = \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.a  + \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.b ;
assign { \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cout , \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.s  } = _148_ + \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cin ;
always @(posedge \add_32s_32ns_32_2_1_U15.top_add_32s_32ns_32_2_1_Adder_10_U.clk )
\add_32s_32ns_32_2_1_U15.top_add_32s_32ns_32_2_1_Adder_10_U.bin_s1  <= _150_;
always @(posedge \add_32s_32ns_32_2_1_U15.top_add_32s_32ns_32_2_1_Adder_10_U.clk )
\add_32s_32ns_32_2_1_U15.top_add_32s_32ns_32_2_1_Adder_10_U.ain_s1  <= _149_;
always @(posedge \add_32s_32ns_32_2_1_U15.top_add_32s_32ns_32_2_1_Adder_10_U.clk )
\add_32s_32ns_32_2_1_U15.top_add_32s_32ns_32_2_1_Adder_10_U.sum_s1  <= _152_;
always @(posedge \add_32s_32ns_32_2_1_U15.top_add_32s_32ns_32_2_1_Adder_10_U.clk )
\add_32s_32ns_32_2_1_U15.top_add_32s_32ns_32_2_1_Adder_10_U.carry_s1  <= _151_;
assign _150_ = \add_32s_32ns_32_2_1_U15.top_add_32s_32ns_32_2_1_Adder_10_U.ce  ? \add_32s_32ns_32_2_1_U15.top_add_32s_32ns_32_2_1_Adder_10_U.b [31:16] : \add_32s_32ns_32_2_1_U15.top_add_32s_32ns_32_2_1_Adder_10_U.bin_s1 ;
assign _149_ = \add_32s_32ns_32_2_1_U15.top_add_32s_32ns_32_2_1_Adder_10_U.ce  ? \add_32s_32ns_32_2_1_U15.top_add_32s_32ns_32_2_1_Adder_10_U.a [31:16] : \add_32s_32ns_32_2_1_U15.top_add_32s_32ns_32_2_1_Adder_10_U.ain_s1 ;
assign _151_ = \add_32s_32ns_32_2_1_U15.top_add_32s_32ns_32_2_1_Adder_10_U.ce  ? \add_32s_32ns_32_2_1_U15.top_add_32s_32ns_32_2_1_Adder_10_U.facout_s1  : \add_32s_32ns_32_2_1_U15.top_add_32s_32ns_32_2_1_Adder_10_U.carry_s1 ;
assign _152_ = \add_32s_32ns_32_2_1_U15.top_add_32s_32ns_32_2_1_Adder_10_U.ce  ? \add_32s_32ns_32_2_1_U15.top_add_32s_32ns_32_2_1_Adder_10_U.fas_s1  : \add_32s_32ns_32_2_1_U15.top_add_32s_32ns_32_2_1_Adder_10_U.sum_s1 ;
assign _153_ = \add_32s_32ns_32_2_1_U15.top_add_32s_32ns_32_2_1_Adder_10_U.u1.a  + \add_32s_32ns_32_2_1_U15.top_add_32s_32ns_32_2_1_Adder_10_U.u1.b ;
assign { \add_32s_32ns_32_2_1_U15.top_add_32s_32ns_32_2_1_Adder_10_U.u1.cout , \add_32s_32ns_32_2_1_U15.top_add_32s_32ns_32_2_1_Adder_10_U.u1.s  } = _153_ + \add_32s_32ns_32_2_1_U15.top_add_32s_32ns_32_2_1_Adder_10_U.u1.cin ;
assign _154_ = \add_32s_32ns_32_2_1_U15.top_add_32s_32ns_32_2_1_Adder_10_U.u2.a  + \add_32s_32ns_32_2_1_U15.top_add_32s_32ns_32_2_1_Adder_10_U.u2.b ;
assign { \add_32s_32ns_32_2_1_U15.top_add_32s_32ns_32_2_1_Adder_10_U.u2.cout , \add_32s_32ns_32_2_1_U15.top_add_32s_32ns_32_2_1_Adder_10_U.u2.s  } = _154_ + \add_32s_32ns_32_2_1_U15.top_add_32s_32ns_32_2_1_Adder_10_U.u2.cin ;
always @(posedge \add_33ns_33ns_33_2_1_U10.top_add_33ns_33ns_33_2_1_Adder_7_U.clk )
\add_33ns_33ns_33_2_1_U10.top_add_33ns_33ns_33_2_1_Adder_7_U.bin_s1  <= _156_;
always @(posedge \add_33ns_33ns_33_2_1_U10.top_add_33ns_33ns_33_2_1_Adder_7_U.clk )
\add_33ns_33ns_33_2_1_U10.top_add_33ns_33ns_33_2_1_Adder_7_U.ain_s1  <= _155_;
always @(posedge \add_33ns_33ns_33_2_1_U10.top_add_33ns_33ns_33_2_1_Adder_7_U.clk )
\add_33ns_33ns_33_2_1_U10.top_add_33ns_33ns_33_2_1_Adder_7_U.sum_s1  <= _158_;
always @(posedge \add_33ns_33ns_33_2_1_U10.top_add_33ns_33ns_33_2_1_Adder_7_U.clk )
\add_33ns_33ns_33_2_1_U10.top_add_33ns_33ns_33_2_1_Adder_7_U.carry_s1  <= _157_;
assign _156_ = \add_33ns_33ns_33_2_1_U10.top_add_33ns_33ns_33_2_1_Adder_7_U.ce  ? \add_33ns_33ns_33_2_1_U10.top_add_33ns_33ns_33_2_1_Adder_7_U.b [32:16] : \add_33ns_33ns_33_2_1_U10.top_add_33ns_33ns_33_2_1_Adder_7_U.bin_s1 ;
assign _155_ = \add_33ns_33ns_33_2_1_U10.top_add_33ns_33ns_33_2_1_Adder_7_U.ce  ? \add_33ns_33ns_33_2_1_U10.top_add_33ns_33ns_33_2_1_Adder_7_U.a [32:16] : \add_33ns_33ns_33_2_1_U10.top_add_33ns_33ns_33_2_1_Adder_7_U.ain_s1 ;
assign _157_ = \add_33ns_33ns_33_2_1_U10.top_add_33ns_33ns_33_2_1_Adder_7_U.ce  ? \add_33ns_33ns_33_2_1_U10.top_add_33ns_33ns_33_2_1_Adder_7_U.facout_s1  : \add_33ns_33ns_33_2_1_U10.top_add_33ns_33ns_33_2_1_Adder_7_U.carry_s1 ;
assign _158_ = \add_33ns_33ns_33_2_1_U10.top_add_33ns_33ns_33_2_1_Adder_7_U.ce  ? \add_33ns_33ns_33_2_1_U10.top_add_33ns_33ns_33_2_1_Adder_7_U.fas_s1  : \add_33ns_33ns_33_2_1_U10.top_add_33ns_33ns_33_2_1_Adder_7_U.sum_s1 ;
assign _159_ = \add_33ns_33ns_33_2_1_U10.top_add_33ns_33ns_33_2_1_Adder_7_U.u1.a  + \add_33ns_33ns_33_2_1_U10.top_add_33ns_33ns_33_2_1_Adder_7_U.u1.b ;
assign { \add_33ns_33ns_33_2_1_U10.top_add_33ns_33ns_33_2_1_Adder_7_U.u1.cout , \add_33ns_33ns_33_2_1_U10.top_add_33ns_33ns_33_2_1_Adder_7_U.u1.s  } = _159_ + \add_33ns_33ns_33_2_1_U10.top_add_33ns_33ns_33_2_1_Adder_7_U.u1.cin ;
assign _160_ = \add_33ns_33ns_33_2_1_U10.top_add_33ns_33ns_33_2_1_Adder_7_U.u2.a  + \add_33ns_33ns_33_2_1_U10.top_add_33ns_33ns_33_2_1_Adder_7_U.u2.b ;
assign { \add_33ns_33ns_33_2_1_U10.top_add_33ns_33ns_33_2_1_Adder_7_U.u2.cout , \add_33ns_33ns_33_2_1_U10.top_add_33ns_33ns_33_2_1_Adder_7_U.u2.s  } = _160_ + \add_33ns_33ns_33_2_1_U10.top_add_33ns_33ns_33_2_1_Adder_7_U.u2.cin ;
always @(posedge \add_47s_47s_47_2_1_U20.top_add_47s_47s_47_2_1_Adder_12_U.clk )
\add_47s_47s_47_2_1_U20.top_add_47s_47s_47_2_1_Adder_12_U.bin_s1  <= _162_;
always @(posedge \add_47s_47s_47_2_1_U20.top_add_47s_47s_47_2_1_Adder_12_U.clk )
\add_47s_47s_47_2_1_U20.top_add_47s_47s_47_2_1_Adder_12_U.ain_s1  <= _161_;
always @(posedge \add_47s_47s_47_2_1_U20.top_add_47s_47s_47_2_1_Adder_12_U.clk )
\add_47s_47s_47_2_1_U20.top_add_47s_47s_47_2_1_Adder_12_U.sum_s1  <= _164_;
always @(posedge \add_47s_47s_47_2_1_U20.top_add_47s_47s_47_2_1_Adder_12_U.clk )
\add_47s_47s_47_2_1_U20.top_add_47s_47s_47_2_1_Adder_12_U.carry_s1  <= _163_;
assign _162_ = \add_47s_47s_47_2_1_U20.top_add_47s_47s_47_2_1_Adder_12_U.ce  ? \add_47s_47s_47_2_1_U20.top_add_47s_47s_47_2_1_Adder_12_U.b [46:23] : \add_47s_47s_47_2_1_U20.top_add_47s_47s_47_2_1_Adder_12_U.bin_s1 ;
assign _161_ = \add_47s_47s_47_2_1_U20.top_add_47s_47s_47_2_1_Adder_12_U.ce  ? \add_47s_47s_47_2_1_U20.top_add_47s_47s_47_2_1_Adder_12_U.a [46:23] : \add_47s_47s_47_2_1_U20.top_add_47s_47s_47_2_1_Adder_12_U.ain_s1 ;
assign _163_ = \add_47s_47s_47_2_1_U20.top_add_47s_47s_47_2_1_Adder_12_U.ce  ? \add_47s_47s_47_2_1_U20.top_add_47s_47s_47_2_1_Adder_12_U.facout_s1  : \add_47s_47s_47_2_1_U20.top_add_47s_47s_47_2_1_Adder_12_U.carry_s1 ;
assign _164_ = \add_47s_47s_47_2_1_U20.top_add_47s_47s_47_2_1_Adder_12_U.ce  ? \add_47s_47s_47_2_1_U20.top_add_47s_47s_47_2_1_Adder_12_U.fas_s1  : \add_47s_47s_47_2_1_U20.top_add_47s_47s_47_2_1_Adder_12_U.sum_s1 ;
assign _165_ = \add_47s_47s_47_2_1_U20.top_add_47s_47s_47_2_1_Adder_12_U.u1.a  + \add_47s_47s_47_2_1_U20.top_add_47s_47s_47_2_1_Adder_12_U.u1.b ;
assign { \add_47s_47s_47_2_1_U20.top_add_47s_47s_47_2_1_Adder_12_U.u1.cout , \add_47s_47s_47_2_1_U20.top_add_47s_47s_47_2_1_Adder_12_U.u1.s  } = _165_ + \add_47s_47s_47_2_1_U20.top_add_47s_47s_47_2_1_Adder_12_U.u1.cin ;
assign _166_ = \add_47s_47s_47_2_1_U20.top_add_47s_47s_47_2_1_Adder_12_U.u2.a  + \add_47s_47s_47_2_1_U20.top_add_47s_47s_47_2_1_Adder_12_U.u2.b ;
assign { \add_47s_47s_47_2_1_U20.top_add_47s_47s_47_2_1_Adder_12_U.u2.cout , \add_47s_47s_47_2_1_U20.top_add_47s_47s_47_2_1_Adder_12_U.u2.s  } = _166_ + \add_47s_47s_47_2_1_U20.top_add_47s_47s_47_2_1_Adder_12_U.u2.cin ;
always @(posedge \add_4s_4ns_4_2_1_U6.top_add_4s_4ns_4_2_1_Adder_4_U.clk )
\add_4s_4ns_4_2_1_U6.top_add_4s_4ns_4_2_1_Adder_4_U.bin_s1  <= _168_;
always @(posedge \add_4s_4ns_4_2_1_U6.top_add_4s_4ns_4_2_1_Adder_4_U.clk )
\add_4s_4ns_4_2_1_U6.top_add_4s_4ns_4_2_1_Adder_4_U.ain_s1  <= _167_;
always @(posedge \add_4s_4ns_4_2_1_U6.top_add_4s_4ns_4_2_1_Adder_4_U.clk )
\add_4s_4ns_4_2_1_U6.top_add_4s_4ns_4_2_1_Adder_4_U.sum_s1  <= _170_;
always @(posedge \add_4s_4ns_4_2_1_U6.top_add_4s_4ns_4_2_1_Adder_4_U.clk )
\add_4s_4ns_4_2_1_U6.top_add_4s_4ns_4_2_1_Adder_4_U.carry_s1  <= _169_;
assign _168_ = \add_4s_4ns_4_2_1_U6.top_add_4s_4ns_4_2_1_Adder_4_U.ce  ? \add_4s_4ns_4_2_1_U6.top_add_4s_4ns_4_2_1_Adder_4_U.b [3:2] : \add_4s_4ns_4_2_1_U6.top_add_4s_4ns_4_2_1_Adder_4_U.bin_s1 ;
assign _167_ = \add_4s_4ns_4_2_1_U6.top_add_4s_4ns_4_2_1_Adder_4_U.ce  ? \add_4s_4ns_4_2_1_U6.top_add_4s_4ns_4_2_1_Adder_4_U.a [3:2] : \add_4s_4ns_4_2_1_U6.top_add_4s_4ns_4_2_1_Adder_4_U.ain_s1 ;
assign _169_ = \add_4s_4ns_4_2_1_U6.top_add_4s_4ns_4_2_1_Adder_4_U.ce  ? \add_4s_4ns_4_2_1_U6.top_add_4s_4ns_4_2_1_Adder_4_U.facout_s1  : \add_4s_4ns_4_2_1_U6.top_add_4s_4ns_4_2_1_Adder_4_U.carry_s1 ;
assign _170_ = \add_4s_4ns_4_2_1_U6.top_add_4s_4ns_4_2_1_Adder_4_U.ce  ? \add_4s_4ns_4_2_1_U6.top_add_4s_4ns_4_2_1_Adder_4_U.fas_s1  : \add_4s_4ns_4_2_1_U6.top_add_4s_4ns_4_2_1_Adder_4_U.sum_s1 ;
assign _171_ = \add_4s_4ns_4_2_1_U6.top_add_4s_4ns_4_2_1_Adder_4_U.u1.a  + \add_4s_4ns_4_2_1_U6.top_add_4s_4ns_4_2_1_Adder_4_U.u1.b ;
assign { \add_4s_4ns_4_2_1_U6.top_add_4s_4ns_4_2_1_Adder_4_U.u1.cout , \add_4s_4ns_4_2_1_U6.top_add_4s_4ns_4_2_1_Adder_4_U.u1.s  } = _171_ + \add_4s_4ns_4_2_1_U6.top_add_4s_4ns_4_2_1_Adder_4_U.u1.cin ;
assign _172_ = \add_4s_4ns_4_2_1_U6.top_add_4s_4ns_4_2_1_Adder_4_U.u2.a  + \add_4s_4ns_4_2_1_U6.top_add_4s_4ns_4_2_1_Adder_4_U.u2.b ;
assign { \add_4s_4ns_4_2_1_U6.top_add_4s_4ns_4_2_1_Adder_4_U.u2.cout , \add_4s_4ns_4_2_1_U6.top_add_4s_4ns_4_2_1_Adder_4_U.u2.s  } = _172_ + \add_4s_4ns_4_2_1_U6.top_add_4s_4ns_4_2_1_Adder_4_U.u2.cin ;
always @(posedge \add_54s_54ns_54_2_1_U18.top_add_54s_54ns_54_2_1_Adder_11_U.clk )
\add_54s_54ns_54_2_1_U18.top_add_54s_54ns_54_2_1_Adder_11_U.bin_s1  <= _174_;
always @(posedge \add_54s_54ns_54_2_1_U18.top_add_54s_54ns_54_2_1_Adder_11_U.clk )
\add_54s_54ns_54_2_1_U18.top_add_54s_54ns_54_2_1_Adder_11_U.ain_s1  <= _173_;
always @(posedge \add_54s_54ns_54_2_1_U18.top_add_54s_54ns_54_2_1_Adder_11_U.clk )
\add_54s_54ns_54_2_1_U18.top_add_54s_54ns_54_2_1_Adder_11_U.sum_s1  <= _176_;
always @(posedge \add_54s_54ns_54_2_1_U18.top_add_54s_54ns_54_2_1_Adder_11_U.clk )
\add_54s_54ns_54_2_1_U18.top_add_54s_54ns_54_2_1_Adder_11_U.carry_s1  <= _175_;
assign _174_ = \add_54s_54ns_54_2_1_U18.top_add_54s_54ns_54_2_1_Adder_11_U.ce  ? \add_54s_54ns_54_2_1_U18.top_add_54s_54ns_54_2_1_Adder_11_U.b [53:27] : \add_54s_54ns_54_2_1_U18.top_add_54s_54ns_54_2_1_Adder_11_U.bin_s1 ;
assign _173_ = \add_54s_54ns_54_2_1_U18.top_add_54s_54ns_54_2_1_Adder_11_U.ce  ? \add_54s_54ns_54_2_1_U18.top_add_54s_54ns_54_2_1_Adder_11_U.a [53:27] : \add_54s_54ns_54_2_1_U18.top_add_54s_54ns_54_2_1_Adder_11_U.ain_s1 ;
assign _175_ = \add_54s_54ns_54_2_1_U18.top_add_54s_54ns_54_2_1_Adder_11_U.ce  ? \add_54s_54ns_54_2_1_U18.top_add_54s_54ns_54_2_1_Adder_11_U.facout_s1  : \add_54s_54ns_54_2_1_U18.top_add_54s_54ns_54_2_1_Adder_11_U.carry_s1 ;
assign _176_ = \add_54s_54ns_54_2_1_U18.top_add_54s_54ns_54_2_1_Adder_11_U.ce  ? \add_54s_54ns_54_2_1_U18.top_add_54s_54ns_54_2_1_Adder_11_U.fas_s1  : \add_54s_54ns_54_2_1_U18.top_add_54s_54ns_54_2_1_Adder_11_U.sum_s1 ;
assign _177_ = \add_54s_54ns_54_2_1_U18.top_add_54s_54ns_54_2_1_Adder_11_U.u1.a  + \add_54s_54ns_54_2_1_U18.top_add_54s_54ns_54_2_1_Adder_11_U.u1.b ;
assign { \add_54s_54ns_54_2_1_U18.top_add_54s_54ns_54_2_1_Adder_11_U.u1.cout , \add_54s_54ns_54_2_1_U18.top_add_54s_54ns_54_2_1_Adder_11_U.u1.s  } = _177_ + \add_54s_54ns_54_2_1_U18.top_add_54s_54ns_54_2_1_Adder_11_U.u1.cin ;
assign _178_ = \add_54s_54ns_54_2_1_U18.top_add_54s_54ns_54_2_1_Adder_11_U.u2.a  + \add_54s_54ns_54_2_1_U18.top_add_54s_54ns_54_2_1_Adder_11_U.u2.b ;
assign { \add_54s_54ns_54_2_1_U18.top_add_54s_54ns_54_2_1_Adder_11_U.u2.cout , \add_54s_54ns_54_2_1_U18.top_add_54s_54ns_54_2_1_Adder_11_U.u2.s  } = _178_ + \add_54s_54ns_54_2_1_U18.top_add_54s_54ns_54_2_1_Adder_11_U.u2.cin ;
always @(posedge \add_5ns_5ns_5_2_1_U14.top_add_5ns_5ns_5_2_1_Adder_9_U.clk )
\add_5ns_5ns_5_2_1_U14.top_add_5ns_5ns_5_2_1_Adder_9_U.bin_s1  <= _180_;
always @(posedge \add_5ns_5ns_5_2_1_U14.top_add_5ns_5ns_5_2_1_Adder_9_U.clk )
\add_5ns_5ns_5_2_1_U14.top_add_5ns_5ns_5_2_1_Adder_9_U.ain_s1  <= _179_;
always @(posedge \add_5ns_5ns_5_2_1_U14.top_add_5ns_5ns_5_2_1_Adder_9_U.clk )
\add_5ns_5ns_5_2_1_U14.top_add_5ns_5ns_5_2_1_Adder_9_U.sum_s1  <= _182_;
always @(posedge \add_5ns_5ns_5_2_1_U14.top_add_5ns_5ns_5_2_1_Adder_9_U.clk )
\add_5ns_5ns_5_2_1_U14.top_add_5ns_5ns_5_2_1_Adder_9_U.carry_s1  <= _181_;
assign _180_ = \add_5ns_5ns_5_2_1_U14.top_add_5ns_5ns_5_2_1_Adder_9_U.ce  ? \add_5ns_5ns_5_2_1_U14.top_add_5ns_5ns_5_2_1_Adder_9_U.b [4:2] : \add_5ns_5ns_5_2_1_U14.top_add_5ns_5ns_5_2_1_Adder_9_U.bin_s1 ;
assign _179_ = \add_5ns_5ns_5_2_1_U14.top_add_5ns_5ns_5_2_1_Adder_9_U.ce  ? \add_5ns_5ns_5_2_1_U14.top_add_5ns_5ns_5_2_1_Adder_9_U.a [4:2] : \add_5ns_5ns_5_2_1_U14.top_add_5ns_5ns_5_2_1_Adder_9_U.ain_s1 ;
assign _181_ = \add_5ns_5ns_5_2_1_U14.top_add_5ns_5ns_5_2_1_Adder_9_U.ce  ? \add_5ns_5ns_5_2_1_U14.top_add_5ns_5ns_5_2_1_Adder_9_U.facout_s1  : \add_5ns_5ns_5_2_1_U14.top_add_5ns_5ns_5_2_1_Adder_9_U.carry_s1 ;
assign _182_ = \add_5ns_5ns_5_2_1_U14.top_add_5ns_5ns_5_2_1_Adder_9_U.ce  ? \add_5ns_5ns_5_2_1_U14.top_add_5ns_5ns_5_2_1_Adder_9_U.fas_s1  : \add_5ns_5ns_5_2_1_U14.top_add_5ns_5ns_5_2_1_Adder_9_U.sum_s1 ;
assign _183_ = \add_5ns_5ns_5_2_1_U14.top_add_5ns_5ns_5_2_1_Adder_9_U.u1.a  + \add_5ns_5ns_5_2_1_U14.top_add_5ns_5ns_5_2_1_Adder_9_U.u1.b ;
assign { \add_5ns_5ns_5_2_1_U14.top_add_5ns_5ns_5_2_1_Adder_9_U.u1.cout , \add_5ns_5ns_5_2_1_U14.top_add_5ns_5ns_5_2_1_Adder_9_U.u1.s  } = _183_ + \add_5ns_5ns_5_2_1_U14.top_add_5ns_5ns_5_2_1_Adder_9_U.u1.cin ;
assign _184_ = \add_5ns_5ns_5_2_1_U14.top_add_5ns_5ns_5_2_1_Adder_9_U.u2.a  + \add_5ns_5ns_5_2_1_U14.top_add_5ns_5ns_5_2_1_Adder_9_U.u2.b ;
assign { \add_5ns_5ns_5_2_1_U14.top_add_5ns_5ns_5_2_1_Adder_9_U.u2.cout , \add_5ns_5ns_5_2_1_U14.top_add_5ns_5ns_5_2_1_Adder_9_U.u2.s  } = _184_ + \add_5ns_5ns_5_2_1_U14.top_add_5ns_5ns_5_2_1_Adder_9_U.u2.cin ;
always @(posedge \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.clk )
\add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.bin_s1  <= _186_;
always @(posedge \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.clk )
\add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.ain_s1  <= _185_;
always @(posedge \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.clk )
\add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.sum_s1  <= _188_;
always @(posedge \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.clk )
\add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.carry_s1  <= _187_;
assign _186_ = \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.ce  ? \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.b [4:2] : \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.bin_s1 ;
assign _185_ = \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.ce  ? \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.a [4:2] : \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.ain_s1 ;
assign _187_ = \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.ce  ? \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.facout_s1  : \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.carry_s1 ;
assign _188_ = \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.ce  ? \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.fas_s1  : \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.sum_s1 ;
assign _189_ = \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.u1.a  + \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.u1.b ;
assign { \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.u1.cout , \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.u1.s  } = _189_ + \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.u1.cin ;
assign _190_ = \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.u2.a  + \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.u2.b ;
assign { \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.u2.cout , \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.u2.s  } = _190_ + \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.u2.cin ;
always @(posedge \add_63s_63s_63_2_1_U7.top_add_63s_63s_63_2_1_Adder_5_U.clk )
\add_63s_63s_63_2_1_U7.top_add_63s_63s_63_2_1_Adder_5_U.bin_s1  <= _192_;
always @(posedge \add_63s_63s_63_2_1_U7.top_add_63s_63s_63_2_1_Adder_5_U.clk )
\add_63s_63s_63_2_1_U7.top_add_63s_63s_63_2_1_Adder_5_U.ain_s1  <= _191_;
always @(posedge \add_63s_63s_63_2_1_U7.top_add_63s_63s_63_2_1_Adder_5_U.clk )
\add_63s_63s_63_2_1_U7.top_add_63s_63s_63_2_1_Adder_5_U.sum_s1  <= _194_;
always @(posedge \add_63s_63s_63_2_1_U7.top_add_63s_63s_63_2_1_Adder_5_U.clk )
\add_63s_63s_63_2_1_U7.top_add_63s_63s_63_2_1_Adder_5_U.carry_s1  <= _193_;
assign _192_ = \add_63s_63s_63_2_1_U7.top_add_63s_63s_63_2_1_Adder_5_U.ce  ? \add_63s_63s_63_2_1_U7.top_add_63s_63s_63_2_1_Adder_5_U.b [62:31] : \add_63s_63s_63_2_1_U7.top_add_63s_63s_63_2_1_Adder_5_U.bin_s1 ;
assign _191_ = \add_63s_63s_63_2_1_U7.top_add_63s_63s_63_2_1_Adder_5_U.ce  ? \add_63s_63s_63_2_1_U7.top_add_63s_63s_63_2_1_Adder_5_U.a [62:31] : \add_63s_63s_63_2_1_U7.top_add_63s_63s_63_2_1_Adder_5_U.ain_s1 ;
assign _193_ = \add_63s_63s_63_2_1_U7.top_add_63s_63s_63_2_1_Adder_5_U.ce  ? \add_63s_63s_63_2_1_U7.top_add_63s_63s_63_2_1_Adder_5_U.facout_s1  : \add_63s_63s_63_2_1_U7.top_add_63s_63s_63_2_1_Adder_5_U.carry_s1 ;
assign _194_ = \add_63s_63s_63_2_1_U7.top_add_63s_63s_63_2_1_Adder_5_U.ce  ? \add_63s_63s_63_2_1_U7.top_add_63s_63s_63_2_1_Adder_5_U.fas_s1  : \add_63s_63s_63_2_1_U7.top_add_63s_63s_63_2_1_Adder_5_U.sum_s1 ;
assign _195_ = \add_63s_63s_63_2_1_U7.top_add_63s_63s_63_2_1_Adder_5_U.u1.a  + \add_63s_63s_63_2_1_U7.top_add_63s_63s_63_2_1_Adder_5_U.u1.b ;
assign { \add_63s_63s_63_2_1_U7.top_add_63s_63s_63_2_1_Adder_5_U.u1.cout , \add_63s_63s_63_2_1_U7.top_add_63s_63s_63_2_1_Adder_5_U.u1.s  } = _195_ + \add_63s_63s_63_2_1_U7.top_add_63s_63s_63_2_1_Adder_5_U.u1.cin ;
assign _196_ = \add_63s_63s_63_2_1_U7.top_add_63s_63s_63_2_1_Adder_5_U.u2.a  + \add_63s_63s_63_2_1_U7.top_add_63s_63s_63_2_1_Adder_5_U.u2.b ;
assign { \add_63s_63s_63_2_1_U7.top_add_63s_63s_63_2_1_Adder_5_U.u2.cout , \add_63s_63s_63_2_1_U7.top_add_63s_63s_63_2_1_Adder_5_U.u2.s  } = _196_ + \add_63s_63s_63_2_1_U7.top_add_63s_63s_63_2_1_Adder_5_U.u2.cin ;
assign \mul_16ns_4s_20_7_1_U5.top_mul_16ns_4s_20_7_1_Mul_DSP_0_U.tmp_product  = $signed({ 1'h0, \mul_16ns_4s_20_7_1_U5.top_mul_16ns_4s_20_7_1_Mul_DSP_0_U.a_reg0  }) * $signed(\mul_16ns_4s_20_7_1_U5.top_mul_16ns_4s_20_7_1_Mul_DSP_0_U.b_reg0 );
always @(posedge \mul_16ns_4s_20_7_1_U5.top_mul_16ns_4s_20_7_1_Mul_DSP_0_U.clk )
\mul_16ns_4s_20_7_1_U5.top_mul_16ns_4s_20_7_1_Mul_DSP_0_U.a_reg0  <= _197_;
always @(posedge \mul_16ns_4s_20_7_1_U5.top_mul_16ns_4s_20_7_1_Mul_DSP_0_U.clk )
\mul_16ns_4s_20_7_1_U5.top_mul_16ns_4s_20_7_1_Mul_DSP_0_U.b_reg0  <= _198_;
always @(posedge \mul_16ns_4s_20_7_1_U5.top_mul_16ns_4s_20_7_1_Mul_DSP_0_U.clk )
\mul_16ns_4s_20_7_1_U5.top_mul_16ns_4s_20_7_1_Mul_DSP_0_U.buff0  <= _199_;
always @(posedge \mul_16ns_4s_20_7_1_U5.top_mul_16ns_4s_20_7_1_Mul_DSP_0_U.clk )
\mul_16ns_4s_20_7_1_U5.top_mul_16ns_4s_20_7_1_Mul_DSP_0_U.buff1  <= _200_;
always @(posedge \mul_16ns_4s_20_7_1_U5.top_mul_16ns_4s_20_7_1_Mul_DSP_0_U.clk )
\mul_16ns_4s_20_7_1_U5.top_mul_16ns_4s_20_7_1_Mul_DSP_0_U.buff2  <= _201_;
always @(posedge \mul_16ns_4s_20_7_1_U5.top_mul_16ns_4s_20_7_1_Mul_DSP_0_U.clk )
\mul_16ns_4s_20_7_1_U5.top_mul_16ns_4s_20_7_1_Mul_DSP_0_U.buff3  <= _202_;
always @(posedge \mul_16ns_4s_20_7_1_U5.top_mul_16ns_4s_20_7_1_Mul_DSP_0_U.clk )
\mul_16ns_4s_20_7_1_U5.top_mul_16ns_4s_20_7_1_Mul_DSP_0_U.buff4  <= _203_;
assign _203_ = \mul_16ns_4s_20_7_1_U5.top_mul_16ns_4s_20_7_1_Mul_DSP_0_U.ce  ? \mul_16ns_4s_20_7_1_U5.top_mul_16ns_4s_20_7_1_Mul_DSP_0_U.buff3  : \mul_16ns_4s_20_7_1_U5.top_mul_16ns_4s_20_7_1_Mul_DSP_0_U.buff4 ;
assign _202_ = \mul_16ns_4s_20_7_1_U5.top_mul_16ns_4s_20_7_1_Mul_DSP_0_U.ce  ? \mul_16ns_4s_20_7_1_U5.top_mul_16ns_4s_20_7_1_Mul_DSP_0_U.buff2  : \mul_16ns_4s_20_7_1_U5.top_mul_16ns_4s_20_7_1_Mul_DSP_0_U.buff3 ;
assign _201_ = \mul_16ns_4s_20_7_1_U5.top_mul_16ns_4s_20_7_1_Mul_DSP_0_U.ce  ? \mul_16ns_4s_20_7_1_U5.top_mul_16ns_4s_20_7_1_Mul_DSP_0_U.buff1  : \mul_16ns_4s_20_7_1_U5.top_mul_16ns_4s_20_7_1_Mul_DSP_0_U.buff2 ;
assign _200_ = \mul_16ns_4s_20_7_1_U5.top_mul_16ns_4s_20_7_1_Mul_DSP_0_U.ce  ? \mul_16ns_4s_20_7_1_U5.top_mul_16ns_4s_20_7_1_Mul_DSP_0_U.buff0  : \mul_16ns_4s_20_7_1_U5.top_mul_16ns_4s_20_7_1_Mul_DSP_0_U.buff1 ;
assign _199_ = \mul_16ns_4s_20_7_1_U5.top_mul_16ns_4s_20_7_1_Mul_DSP_0_U.ce  ? \mul_16ns_4s_20_7_1_U5.top_mul_16ns_4s_20_7_1_Mul_DSP_0_U.tmp_product  : \mul_16ns_4s_20_7_1_U5.top_mul_16ns_4s_20_7_1_Mul_DSP_0_U.buff0 ;
assign _198_ = \mul_16ns_4s_20_7_1_U5.top_mul_16ns_4s_20_7_1_Mul_DSP_0_U.ce  ? \mul_16ns_4s_20_7_1_U5.top_mul_16ns_4s_20_7_1_Mul_DSP_0_U.b  : \mul_16ns_4s_20_7_1_U5.top_mul_16ns_4s_20_7_1_Mul_DSP_0_U.b_reg0 ;
assign _197_ = \mul_16ns_4s_20_7_1_U5.top_mul_16ns_4s_20_7_1_Mul_DSP_0_U.ce  ? \mul_16ns_4s_20_7_1_U5.top_mul_16ns_4s_20_7_1_Mul_DSP_0_U.a  : \mul_16ns_4s_20_7_1_U5.top_mul_16ns_4s_20_7_1_Mul_DSP_0_U.a_reg0 ;
assign \sub_5s_5ns_5_2_1_U4.top_sub_5s_5ns_5_2_1_Adder_3_U.bin_s0  = ~ \sub_5s_5ns_5_2_1_U4.top_sub_5s_5ns_5_2_1_Adder_3_U.b ;
always @(posedge \sub_5s_5ns_5_2_1_U4.top_sub_5s_5ns_5_2_1_Adder_3_U.clk )
\sub_5s_5ns_5_2_1_U4.top_sub_5s_5ns_5_2_1_Adder_3_U.bin_s1  <= _205_;
always @(posedge \sub_5s_5ns_5_2_1_U4.top_sub_5s_5ns_5_2_1_Adder_3_U.clk )
\sub_5s_5ns_5_2_1_U4.top_sub_5s_5ns_5_2_1_Adder_3_U.ain_s1  <= _204_;
always @(posedge \sub_5s_5ns_5_2_1_U4.top_sub_5s_5ns_5_2_1_Adder_3_U.clk )
\sub_5s_5ns_5_2_1_U4.top_sub_5s_5ns_5_2_1_Adder_3_U.sum_s1  <= _207_;
always @(posedge \sub_5s_5ns_5_2_1_U4.top_sub_5s_5ns_5_2_1_Adder_3_U.clk )
\sub_5s_5ns_5_2_1_U4.top_sub_5s_5ns_5_2_1_Adder_3_U.carry_s1  <= _206_;
assign _205_ = \sub_5s_5ns_5_2_1_U4.top_sub_5s_5ns_5_2_1_Adder_3_U.ce  ? \sub_5s_5ns_5_2_1_U4.top_sub_5s_5ns_5_2_1_Adder_3_U.bin_s0 [4:2] : \sub_5s_5ns_5_2_1_U4.top_sub_5s_5ns_5_2_1_Adder_3_U.bin_s1 ;
assign _204_ = \sub_5s_5ns_5_2_1_U4.top_sub_5s_5ns_5_2_1_Adder_3_U.ce  ? \sub_5s_5ns_5_2_1_U4.top_sub_5s_5ns_5_2_1_Adder_3_U.a [4:2] : \sub_5s_5ns_5_2_1_U4.top_sub_5s_5ns_5_2_1_Adder_3_U.ain_s1 ;
assign _206_ = \sub_5s_5ns_5_2_1_U4.top_sub_5s_5ns_5_2_1_Adder_3_U.ce  ? \sub_5s_5ns_5_2_1_U4.top_sub_5s_5ns_5_2_1_Adder_3_U.facout_s1  : \sub_5s_5ns_5_2_1_U4.top_sub_5s_5ns_5_2_1_Adder_3_U.carry_s1 ;
assign _207_ = \sub_5s_5ns_5_2_1_U4.top_sub_5s_5ns_5_2_1_Adder_3_U.ce  ? \sub_5s_5ns_5_2_1_U4.top_sub_5s_5ns_5_2_1_Adder_3_U.fas_s1  : \sub_5s_5ns_5_2_1_U4.top_sub_5s_5ns_5_2_1_Adder_3_U.sum_s1 ;
assign _208_ = \sub_5s_5ns_5_2_1_U4.top_sub_5s_5ns_5_2_1_Adder_3_U.u1.a  + \sub_5s_5ns_5_2_1_U4.top_sub_5s_5ns_5_2_1_Adder_3_U.u1.b ;
assign { \sub_5s_5ns_5_2_1_U4.top_sub_5s_5ns_5_2_1_Adder_3_U.u1.cout , \sub_5s_5ns_5_2_1_U4.top_sub_5s_5ns_5_2_1_Adder_3_U.u1.s  } = _208_ + \sub_5s_5ns_5_2_1_U4.top_sub_5s_5ns_5_2_1_Adder_3_U.u1.cin ;
assign _209_ = \sub_5s_5ns_5_2_1_U4.top_sub_5s_5ns_5_2_1_Adder_3_U.u2.a  + \sub_5s_5ns_5_2_1_U4.top_sub_5s_5ns_5_2_1_Adder_3_U.u2.b ;
assign { \sub_5s_5ns_5_2_1_U4.top_sub_5s_5ns_5_2_1_Adder_3_U.u2.cout , \sub_5s_5ns_5_2_1_U4.top_sub_5s_5ns_5_2_1_Adder_3_U.u2.s  } = _209_ + \sub_5s_5ns_5_2_1_U4.top_sub_5s_5ns_5_2_1_Adder_3_U.u2.cin ;
assign \sub_5s_5s_5_2_1_U1.top_sub_5s_5s_5_2_1_Adder_0_U.bin_s0  = ~ \sub_5s_5s_5_2_1_U1.top_sub_5s_5s_5_2_1_Adder_0_U.b ;
always @(posedge \sub_5s_5s_5_2_1_U1.top_sub_5s_5s_5_2_1_Adder_0_U.clk )
\sub_5s_5s_5_2_1_U1.top_sub_5s_5s_5_2_1_Adder_0_U.bin_s1  <= _211_;
always @(posedge \sub_5s_5s_5_2_1_U1.top_sub_5s_5s_5_2_1_Adder_0_U.clk )
\sub_5s_5s_5_2_1_U1.top_sub_5s_5s_5_2_1_Adder_0_U.ain_s1  <= _210_;
always @(posedge \sub_5s_5s_5_2_1_U1.top_sub_5s_5s_5_2_1_Adder_0_U.clk )
\sub_5s_5s_5_2_1_U1.top_sub_5s_5s_5_2_1_Adder_0_U.sum_s1  <= _213_;
always @(posedge \sub_5s_5s_5_2_1_U1.top_sub_5s_5s_5_2_1_Adder_0_U.clk )
\sub_5s_5s_5_2_1_U1.top_sub_5s_5s_5_2_1_Adder_0_U.carry_s1  <= _212_;
assign _211_ = \sub_5s_5s_5_2_1_U1.top_sub_5s_5s_5_2_1_Adder_0_U.ce  ? \sub_5s_5s_5_2_1_U1.top_sub_5s_5s_5_2_1_Adder_0_U.bin_s0 [4:2] : \sub_5s_5s_5_2_1_U1.top_sub_5s_5s_5_2_1_Adder_0_U.bin_s1 ;
assign _210_ = \sub_5s_5s_5_2_1_U1.top_sub_5s_5s_5_2_1_Adder_0_U.ce  ? \sub_5s_5s_5_2_1_U1.top_sub_5s_5s_5_2_1_Adder_0_U.a [4:2] : \sub_5s_5s_5_2_1_U1.top_sub_5s_5s_5_2_1_Adder_0_U.ain_s1 ;
assign _212_ = \sub_5s_5s_5_2_1_U1.top_sub_5s_5s_5_2_1_Adder_0_U.ce  ? \sub_5s_5s_5_2_1_U1.top_sub_5s_5s_5_2_1_Adder_0_U.facout_s1  : \sub_5s_5s_5_2_1_U1.top_sub_5s_5s_5_2_1_Adder_0_U.carry_s1 ;
assign _213_ = \sub_5s_5s_5_2_1_U1.top_sub_5s_5s_5_2_1_Adder_0_U.ce  ? \sub_5s_5s_5_2_1_U1.top_sub_5s_5s_5_2_1_Adder_0_U.fas_s1  : \sub_5s_5s_5_2_1_U1.top_sub_5s_5s_5_2_1_Adder_0_U.sum_s1 ;
assign _214_ = \sub_5s_5s_5_2_1_U1.top_sub_5s_5s_5_2_1_Adder_0_U.u1.a  + \sub_5s_5s_5_2_1_U1.top_sub_5s_5s_5_2_1_Adder_0_U.u1.b ;
assign { \sub_5s_5s_5_2_1_U1.top_sub_5s_5s_5_2_1_Adder_0_U.u1.cout , \sub_5s_5s_5_2_1_U1.top_sub_5s_5s_5_2_1_Adder_0_U.u1.s  } = _214_ + \sub_5s_5s_5_2_1_U1.top_sub_5s_5s_5_2_1_Adder_0_U.u1.cin ;
assign _215_ = \sub_5s_5s_5_2_1_U1.top_sub_5s_5s_5_2_1_Adder_0_U.u2.a  + \sub_5s_5s_5_2_1_U1.top_sub_5s_5s_5_2_1_Adder_0_U.u2.b ;
assign { \sub_5s_5s_5_2_1_U1.top_sub_5s_5s_5_2_1_Adder_0_U.u2.cout , \sub_5s_5s_5_2_1_U1.top_sub_5s_5s_5_2_1_Adder_0_U.u2.s  } = _215_ + \sub_5s_5s_5_2_1_U1.top_sub_5s_5s_5_2_1_Adder_0_U.u2.cin ;
assign \sub_5s_5s_5_2_1_U12.top_sub_5s_5s_5_2_1_Adder_0_U.bin_s0  = ~ \sub_5s_5s_5_2_1_U12.top_sub_5s_5s_5_2_1_Adder_0_U.b ;
always @(posedge \sub_5s_5s_5_2_1_U12.top_sub_5s_5s_5_2_1_Adder_0_U.clk )
\sub_5s_5s_5_2_1_U12.top_sub_5s_5s_5_2_1_Adder_0_U.bin_s1  <= _217_;
always @(posedge \sub_5s_5s_5_2_1_U12.top_sub_5s_5s_5_2_1_Adder_0_U.clk )
\sub_5s_5s_5_2_1_U12.top_sub_5s_5s_5_2_1_Adder_0_U.ain_s1  <= _216_;
always @(posedge \sub_5s_5s_5_2_1_U12.top_sub_5s_5s_5_2_1_Adder_0_U.clk )
\sub_5s_5s_5_2_1_U12.top_sub_5s_5s_5_2_1_Adder_0_U.sum_s1  <= _219_;
always @(posedge \sub_5s_5s_5_2_1_U12.top_sub_5s_5s_5_2_1_Adder_0_U.clk )
\sub_5s_5s_5_2_1_U12.top_sub_5s_5s_5_2_1_Adder_0_U.carry_s1  <= _218_;
assign _217_ = \sub_5s_5s_5_2_1_U12.top_sub_5s_5s_5_2_1_Adder_0_U.ce  ? \sub_5s_5s_5_2_1_U12.top_sub_5s_5s_5_2_1_Adder_0_U.bin_s0 [4:2] : \sub_5s_5s_5_2_1_U12.top_sub_5s_5s_5_2_1_Adder_0_U.bin_s1 ;
assign _216_ = \sub_5s_5s_5_2_1_U12.top_sub_5s_5s_5_2_1_Adder_0_U.ce  ? \sub_5s_5s_5_2_1_U12.top_sub_5s_5s_5_2_1_Adder_0_U.a [4:2] : \sub_5s_5s_5_2_1_U12.top_sub_5s_5s_5_2_1_Adder_0_U.ain_s1 ;
assign _218_ = \sub_5s_5s_5_2_1_U12.top_sub_5s_5s_5_2_1_Adder_0_U.ce  ? \sub_5s_5s_5_2_1_U12.top_sub_5s_5s_5_2_1_Adder_0_U.facout_s1  : \sub_5s_5s_5_2_1_U12.top_sub_5s_5s_5_2_1_Adder_0_U.carry_s1 ;
assign _219_ = \sub_5s_5s_5_2_1_U12.top_sub_5s_5s_5_2_1_Adder_0_U.ce  ? \sub_5s_5s_5_2_1_U12.top_sub_5s_5s_5_2_1_Adder_0_U.fas_s1  : \sub_5s_5s_5_2_1_U12.top_sub_5s_5s_5_2_1_Adder_0_U.sum_s1 ;
assign _220_ = \sub_5s_5s_5_2_1_U12.top_sub_5s_5s_5_2_1_Adder_0_U.u1.a  + \sub_5s_5s_5_2_1_U12.top_sub_5s_5s_5_2_1_Adder_0_U.u1.b ;
assign { \sub_5s_5s_5_2_1_U12.top_sub_5s_5s_5_2_1_Adder_0_U.u1.cout , \sub_5s_5s_5_2_1_U12.top_sub_5s_5s_5_2_1_Adder_0_U.u1.s  } = _220_ + \sub_5s_5s_5_2_1_U12.top_sub_5s_5s_5_2_1_Adder_0_U.u1.cin ;
assign _221_ = \sub_5s_5s_5_2_1_U12.top_sub_5s_5s_5_2_1_Adder_0_U.u2.a  + \sub_5s_5s_5_2_1_U12.top_sub_5s_5s_5_2_1_Adder_0_U.u2.b ;
assign { \sub_5s_5s_5_2_1_U12.top_sub_5s_5s_5_2_1_Adder_0_U.u2.cout , \sub_5s_5s_5_2_1_U12.top_sub_5s_5s_5_2_1_Adder_0_U.u2.s  } = _221_ + \sub_5s_5s_5_2_1_U12.top_sub_5s_5s_5_2_1_Adder_0_U.u2.cin ;
assign _222_ = | op_1[3:1];
assign _223_ = | p_Result_4_reg_1568;
assign _224_ = | tmp_3_reg_1347;
assign _225_ = | p_Result_s_reg_1206;
assign _226_ = op_1[3:1] != 3'h7;
assign _227_ = tmp_3_reg_1347 != 3'h7;
assign _228_ = p_Result_s_reg_1206 != 4'hf;
assign _229_ = | trunc_ln851_reg_1589;
assign _230_ = | trunc_ln851_2_reg_1463;
assign _231_ = | trunc_ln851_3_reg_1659;
assign _232_ = | op_19[13:0];
assign _233_ = | trunc_ln851_1_reg_1453;
assign _234_ = select_ln874_fu_949_p3 != op_8;
assign or_ln340_1_fu_412_p2 = p_Result_15_reg_1164 | overflow_1_fu_398_p2;
assign or_ln340_fu_293_p2 = p_Result_13_reg_1188 | overflow_fu_278_p2;
assign or_ln384_fu_673_p2 = underflow_2_fu_668_p2 | overflow_3_reg_1391;
assign or_ln785_1_fu_384_p2 = p_Result_16_reg_1259 | icmp_ln768_1_reg_1171;
assign or_ln785_2_fu_320_p2 = xor_ln785_3_fu_315_p2 | p_Result_13_reg_1188;
assign or_ln785_3_fu_599_p2 = p_Result_20_reg_1363 | icmp_ln768_3_reg_1369;
assign or_ln785_4_fu_556_p2 = xor_ln785_4_fu_551_p2 | p_Result_15_reg_1164;
assign or_ln785_5_fu_513_p2 = and_ln785_4_fu_509_p2 | and_ln340_2_fu_505_p2;
assign or_ln785_fu_269_p2 = newsignbit_reg_1195 | icmp_ln768_reg_1212;
assign or_ln786_1_fu_407_p2 = xor_ln786_fu_402_p2 | icmp_ln786_1_reg_1176;
assign or_ln786_fu_288_p2 = p_Val2_1_fu_283_p2 | icmp_ln786_reg_1217;
assign or_ln788_1_fu_663_p2 = or_ln788_fu_658_p2 | icmp_ln786_2_reg_1374;
assign or_ln788_fu_658_p2 = xor_ln786_1_fu_653_p2 | icmp_ln790_reg_1397;
assign overflow_2_fu_1003_p2 = add_ln731_reg_1562[10] | icmp_ln768_2_reg_1594;
always @(posedge ap_clk)
p_Val2_2_reg_1251[2:0] <= 3'h0;
always @(posedge ap_clk)
op_18_V_reg_1649[20:0] <= 21'h000000;
always @(posedge ap_clk)
trunc_ln851_3_reg_1659 <= 21'h000000;
always @(posedge ap_clk)
select_ln785_reg_1353 <= _070_;
always @(posedge ap_clk)
select_ln353_reg_1696 <= _069_;
always @(posedge ap_clk)
select_ln340_reg_1239 <= _068_;
always @(posedge ap_clk)
select_ln1192_reg_1512 <= _066_;
always @(posedge ap_clk)
ret_V_reg_1517 <= _062_;
always @(posedge ap_clk)
ret_V_19_reg_1716 <= _059_;
always @(posedge ap_clk)
ret_V_20_cast_reg_1721 <= _060_;
always @(posedge ap_clk)
ret_V_18_reg_1679 <= _058_;
always @(posedge ap_clk)
ret_V_18_cast_reg_1684 <= _057_;
always @(posedge ap_clk)
ret_V_17_reg_1639 <= _056_;
always @(posedge ap_clk)
select_ln340_1_reg_1326 <= _067_;
always @(posedge ap_clk)
sel_tmp18_reg_1331 <= _064_;
always @(posedge ap_clk)
p_Result_19_reg_1336 <= _045_;
always @(posedge ap_clk)
tmp_3_reg_1347 <= _075_;
always @(posedge ap_clk)
or_ln785_reg_1223 <= _039_;
always @(posedge ap_clk)
ret_V_11_reg_1402 <= _051_;
always @(posedge ap_clk)
or_ln384_reg_1418 <= _037_;
always @(posedge ap_clk)
op_2_V_reg_1244 <= _034_;
always @(posedge ap_clk)
p_Val2_2_reg_1251[3] <= _049_;
always @(posedge ap_clk)
p_Result_16_reg_1259 <= _044_;
always @(posedge ap_clk)
op_23_V_reg_1629 <= _032_;
always @(posedge ap_clk)
select_ln1192_1_reg_1634 <= _065_;
always @(posedge ap_clk)
op_18_V_reg_1649[31:21] <= _031_;
always @(posedge ap_clk)
op_25_V_reg_1654 <= _033_;
always @(posedge ap_clk)
op_16_V_reg_1619 <= _030_;
always @(posedge ap_clk)
ret_reg_1182 <= _063_;
always @(posedge ap_clk)
p_Result_13_reg_1188 <= _042_;
always @(posedge ap_clk)
newsignbit_reg_1195 <= _027_;
always @(posedge ap_clk)
p_Result_s_reg_1206 <= _048_;
always @(posedge ap_clk)
or_ln785_1_reg_1266 <= _038_;
always @(posedge ap_clk)
xor_ln785_1_reg_1272 <= _081_;
always @(posedge ap_clk)
lhs_V_3_reg_1278 <= _026_;
always @(posedge ap_clk)
icmp_ln851_3_reg_1711 <= _024_;
always @(posedge ap_clk)
icmp_ln851_2_reg_1674 <= _023_;
always @(posedge ap_clk)
sext_ln850_reg_1468 <= _073_;
always @(posedge ap_clk)
icmp_ln851_reg_1475 <= _025_;
always @(posedge ap_clk)
icmp_ln851_1_reg_1490 <= _022_;
always @(posedge ap_clk)
op_4_V_reg_1384 <= _035_;
always @(posedge ap_clk)
overflow_3_reg_1391 <= _041_;
always @(posedge ap_clk)
icmp_ln790_reg_1397 <= _020_;
always @(posedge ap_clk)
icmp_ln768_reg_1212 <= _016_;
always @(posedge ap_clk)
icmp_ln786_reg_1217 <= _019_;
always @(posedge ap_clk)
r_V_reg_1583 <= _050_;
always @(posedge ap_clk)
trunc_ln851_reg_1589 <= _080_;
always @(posedge ap_clk)
icmp_ln768_2_reg_1594 <= _014_;
always @(posedge ap_clk)
p_Result_15_reg_1164 <= _043_;
always @(posedge ap_clk)
icmp_ln768_1_reg_1171 <= _013_;
always @(posedge ap_clk)
icmp_ln786_1_reg_1176 <= _017_;
always @(posedge ap_clk)
icmp_ln1498_reg_1423 <= _012_;
always @(posedge ap_clk)
sext_ln1118_reg_1433 <= _071_;
always @(posedge ap_clk)
ret_V_14_reg_1443 <= _053_;
always @(posedge ap_clk)
tmp_2_reg_1448 <= _074_;
always @(posedge ap_clk)
trunc_ln851_1_reg_1453 <= _078_;
always @(posedge ap_clk)
op_12_V_reg_1458 <= _028_;
always @(posedge ap_clk)
trunc_ln851_2_reg_1463 <= _079_;
always @(posedge ap_clk)
or_ln786_1_reg_1292 <= _040_;
always @(posedge ap_clk)
or_ln340_1_reg_1298 <= _036_;
always @(posedge ap_clk)
and_ln786_reg_1304 <= _010_;
always @(posedge ap_clk)
sext_ln1346_reg_1315 <= _072_;
always @(posedge ap_clk)
trunc_ln731_2_reg_1321 <= _076_;
always @(posedge ap_clk)
and_ln340_reg_1229 <= _008_;
always @(posedge ap_clk)
and_ln785_1_reg_1234 <= _009_;
always @(posedge ap_clk)
ret_V_12_reg_1557 <= _052_;
always @(posedge ap_clk)
add_ln731_reg_1562 <= _007_;
always @(posedge ap_clk)
p_Result_4_reg_1568 <= _047_;
always @(posedge ap_clk)
op_15_V_reg_1573 <= _029_;
always @(posedge ap_clk)
ret_V_16_reg_1578 <= _055_;
always @(posedge ap_clk)
add_ln731_1_reg_1358 <= _006_;
always @(posedge ap_clk)
p_Result_20_reg_1363 <= _046_;
always @(posedge ap_clk)
icmp_ln768_3_reg_1369 <= _015_;
always @(posedge ap_clk)
icmp_ln786_2_reg_1374 <= _018_;
always @(posedge ap_clk)
trunc_ln790_reg_1379 <= _077_;
always @(posedge ap_clk)
icmp_ln850_reg_1604 <= _021_;
always @(posedge ap_clk)
add_ln69_reg_1609 <= _005_;
always @(posedge ap_clk)
add_ln69_1_reg_1614 <= _004_;
always @(posedge ap_clk)
add_ln691_reg_1495 <= _003_;
always @(posedge ap_clk)
ret_V_15_reg_1500 <= _054_;
always @(posedge ap_clk)
ret_V_7_cast_reg_1505 <= _061_;
always @(posedge ap_clk)
add_ln691_3_reg_1728 <= _002_;
always @(posedge ap_clk)
add_ln691_2_reg_1691 <= _001_;
always @(posedge ap_clk)
add_ln691_1_reg_1552 <= _000_;
always @(posedge ap_clk)
ap_CS_fsm <= _011_;
assign _082_ = _089_ ? 2'h2 : 2'h1;
assign _235_ = ap_CS_fsm == 1'h1;
function [36:0] _685_;
input [36:0] a;
input [1368:0] b;
input [36:0] s;
case (s)
37'b0000000000000000000000000000000000001:
_685_ = b[36:0];
37'b0000000000000000000000000000000000010:
_685_ = b[73:37];
37'b0000000000000000000000000000000000100:
_685_ = b[110:74];
37'b0000000000000000000000000000000001000:
_685_ = b[147:111];
37'b0000000000000000000000000000000010000:
_685_ = b[184:148];
37'b0000000000000000000000000000000100000:
_685_ = b[221:185];
37'b0000000000000000000000000000001000000:
_685_ = b[258:222];
37'b0000000000000000000000000000010000000:
_685_ = b[295:259];
37'b0000000000000000000000000000100000000:
_685_ = b[332:296];
37'b0000000000000000000000000001000000000:
_685_ = b[369:333];
37'b0000000000000000000000000010000000000:
_685_ = b[406:370];
37'b0000000000000000000000000100000000000:
_685_ = b[443:407];
37'b0000000000000000000000001000000000000:
_685_ = b[480:444];
37'b0000000000000000000000010000000000000:
_685_ = b[517:481];
37'b0000000000000000000000100000000000000:
_685_ = b[554:518];
37'b0000000000000000000001000000000000000:
_685_ = b[591:555];
37'b0000000000000000000010000000000000000:
_685_ = b[628:592];
37'b0000000000000000000100000000000000000:
_685_ = b[665:629];
37'b0000000000000000001000000000000000000:
_685_ = b[702:666];
37'b0000000000000000010000000000000000000:
_685_ = b[739:703];
37'b0000000000000000100000000000000000000:
_685_ = b[776:740];
37'b0000000000000001000000000000000000000:
_685_ = b[813:777];
37'b0000000000000010000000000000000000000:
_685_ = b[850:814];
37'b0000000000000100000000000000000000000:
_685_ = b[887:851];
37'b0000000000001000000000000000000000000:
_685_ = b[924:888];
37'b0000000000010000000000000000000000000:
_685_ = b[961:925];
37'b0000000000100000000000000000000000000:
_685_ = b[998:962];
37'b0000000001000000000000000000000000000:
_685_ = b[1035:999];
37'b0000000010000000000000000000000000000:
_685_ = b[1072:1036];
37'b0000000100000000000000000000000000000:
_685_ = b[1109:1073];
37'b0000001000000000000000000000000000000:
_685_ = b[1146:1110];
37'b0000010000000000000000000000000000000:
_685_ = b[1183:1147];
37'b0000100000000000000000000000000000000:
_685_ = b[1220:1184];
37'b0001000000000000000000000000000000000:
_685_ = b[1257:1221];
37'b0010000000000000000000000000000000000:
_685_ = b[1294:1258];
37'b0100000000000000000000000000000000000:
_685_ = b[1331:1295];
37'b1000000000000000000000000000000000000:
_685_ = b[1368:1332];
37'b0000000000000000000000000000000000000:
_685_ = a;
default:
_685_ = 37'bx;
endcase
endfunction
assign ap_NS_fsm = _685_(37'hxxxxxxxxxx, { 35'h000000000, _082_, 1332'h000000002000000002000000002000000002000000002000000002000000002000000002000000002000000002000000002000000002000000002000000002000000002000000002000000002000000002000000002000000002000000002000000002000000002000000002000000002000000002000000002000000002000000002000000002000000002000000002000000002000000002000000002000000000000000001 }, { _235_, _271_, _270_, _269_, _268_, _267_, _266_, _265_, _264_, _263_, _262_, _261_, _260_, _259_, _258_, _257_, _256_, _255_, _254_, _253_, _252_, _251_, _250_, _249_, _248_, _247_, _246_, _245_, _244_, _243_, _242_, _241_, _240_, _239_, _238_, _237_, _236_ });
assign _236_ = ap_CS_fsm == 37'h1000000000;
assign _237_ = ap_CS_fsm == 36'h800000000;
assign _238_ = ap_CS_fsm == 35'h400000000;
assign _239_ = ap_CS_fsm == 34'h200000000;
assign _240_ = ap_CS_fsm == 33'h100000000;
assign _241_ = ap_CS_fsm == 32'd2147483648;
assign _242_ = ap_CS_fsm == 31'h40000000;
assign _243_ = ap_CS_fsm == 30'h20000000;
assign _244_ = ap_CS_fsm == 29'h10000000;
assign _245_ = ap_CS_fsm == 28'h8000000;
assign _246_ = ap_CS_fsm == 27'h4000000;
assign _247_ = ap_CS_fsm == 26'h2000000;
assign _248_ = ap_CS_fsm == 25'h1000000;
assign _249_ = ap_CS_fsm == 24'h800000;
assign _250_ = ap_CS_fsm == 23'h400000;
assign _251_ = ap_CS_fsm == 22'h200000;
assign _252_ = ap_CS_fsm == 21'h100000;
assign _253_ = ap_CS_fsm == 20'h80000;
assign _254_ = ap_CS_fsm == 19'h40000;
assign _255_ = ap_CS_fsm == 18'h20000;
assign _256_ = ap_CS_fsm == 17'h10000;
assign _257_ = ap_CS_fsm == 16'h8000;
assign _258_ = ap_CS_fsm == 15'h4000;
assign _259_ = ap_CS_fsm == 14'h2000;
assign _260_ = ap_CS_fsm == 13'h1000;
assign _261_ = ap_CS_fsm == 12'h800;
assign _262_ = ap_CS_fsm == 11'h400;
assign _263_ = ap_CS_fsm == 10'h200;
assign _264_ = ap_CS_fsm == 9'h100;
assign _265_ = ap_CS_fsm == 8'h80;
assign _266_ = ap_CS_fsm == 7'h40;
assign _267_ = ap_CS_fsm == 6'h20;
assign _268_ = ap_CS_fsm == 5'h10;
assign _269_ = ap_CS_fsm == 4'h8;
assign _270_ = ap_CS_fsm == 3'h4;
assign _271_ = ap_CS_fsm == 2'h2;
assign op_27_ap_vld = ap_CS_fsm[36] ? 1'h1 : 1'h0;
assign ap_idle = _088_ ? 1'h1 : 1'h0;
assign _070_ = _087_ ? select_ln785_fu_566_p3 : select_ln785_reg_1353;
assign _069_ = ap_CS_fsm[31] ? select_ln353_fu_1072_p3 : select_ln353_reg_1696;
assign _068_ = _086_ ? select_ln340_fu_362_p3 : select_ln340_reg_1239;
assign _062_ = ap_CS_fsm[16] ? ret_V_fu_818_p3 : ret_V_reg_1517;
assign _066_ = ap_CS_fsm[16] ? select_ln1192_fu_799_p3 : select_ln1192_reg_1512;
assign _060_ = ap_CS_fsm[33] ? grp_fu_1094_p2[45:14] : ret_V_20_cast_reg_1721;
assign _059_ = ap_CS_fsm[33] ? grp_fu_1094_p2 : ret_V_19_reg_1716;
assign _057_ = ap_CS_fsm[28] ? grp_fu_1034_p2[52:21] : ret_V_18_cast_reg_1684;
assign _058_ = ap_CS_fsm[28] ? grp_fu_1034_p2 : ret_V_18_reg_1679;
assign _056_ = ap_CS_fsm[24] ? grp_fu_977_p2 : ret_V_17_reg_1639;
assign _075_ = ap_CS_fsm[9] ? grp_fu_434_p2[4:2] : tmp_3_reg_1347;
assign _045_ = ap_CS_fsm[9] ? grp_fu_434_p2[4] : p_Result_19_reg_1336;
assign _064_ = ap_CS_fsm[9] ? sel_tmp18_fu_519_p2 : sel_tmp18_reg_1331;
assign _067_ = ap_CS_fsm[9] ? select_ln340_1_fu_498_p3 : select_ln340_1_reg_1326;
assign _039_ = ap_CS_fsm[3] ? or_ln785_fu_269_p2 : or_ln785_reg_1223;
assign _037_ = ap_CS_fsm[12] ? or_ln384_fu_673_p2 : or_ln384_reg_1418;
assign _051_ = ap_CS_fsm[12] ? ret_V_11_fu_627_p3 : ret_V_11_reg_1402;
assign _044_ = ap_CS_fsm[6] ? p_Result_16_fu_378_p2 : p_Result_16_reg_1259;
assign _049_ = ap_CS_fsm[6] ? op_1[0] : p_Val2_2_reg_1251[3];
assign _034_ = ap_CS_fsm[6] ? op_2_V_fu_368_p3 : op_2_V_reg_1244;
assign _065_ = ap_CS_fsm[22] ? select_ln1192_1_fu_970_p3 : select_ln1192_1_reg_1634;
assign _032_ = ap_CS_fsm[22] ? grp_fu_965_p2 : op_23_V_reg_1629;
assign _033_ = ap_CS_fsm[26] ? grp_fu_984_p2 : op_25_V_reg_1654;
assign _031_ = ap_CS_fsm[26] ? op_18_V_fu_1008_p3[31:21] : op_18_V_reg_1649[31:21];
assign _030_ = ap_CS_fsm[21] ? op_16_V_fu_957_p2 : op_16_V_reg_1619;
assign _048_ = ap_CS_fsm[1] ? grp_fu_201_p2[4:1] : p_Result_s_reg_1206;
assign _027_ = ap_CS_fsm[1] ? grp_fu_201_p2[0] : newsignbit_reg_1195;
assign _042_ = ap_CS_fsm[1] ? grp_fu_201_p2[4] : p_Result_13_reg_1188;
assign _063_ = ap_CS_fsm[1] ? grp_fu_201_p2 : ret_reg_1182;
assign _026_ = ap_CS_fsm[7] ? lhs_V_3_fu_393_p2 : lhs_V_3_reg_1278;
assign _081_ = ap_CS_fsm[7] ? xor_ln785_1_fu_388_p2 : xor_ln785_1_reg_1272;
assign _038_ = ap_CS_fsm[7] ? or_ln785_1_fu_384_p2 : or_ln785_1_reg_1266;
assign _024_ = ap_CS_fsm[32] ? icmp_ln851_3_fu_1104_p2 : icmp_ln851_3_reg_1711;
assign _023_ = ap_CS_fsm[27] ? icmp_ln851_2_fu_1040_p2 : icmp_ln851_2_reg_1674;
assign _022_ = ap_CS_fsm[14] ? icmp_ln851_1_fu_784_p2 : icmp_ln851_1_reg_1490;
assign _025_ = ap_CS_fsm[14] ? icmp_ln851_fu_752_p2 : icmp_ln851_reg_1475;
assign _073_ = ap_CS_fsm[14] ? { tmp_2_reg_1448[2], tmp_2_reg_1448 } : sext_ln850_reg_1468;
assign _020_ = ap_CS_fsm[11] ? icmp_ln790_fu_621_p2 : icmp_ln790_reg_1397;
assign _041_ = ap_CS_fsm[11] ? overflow_3_fu_608_p2 : overflow_3_reg_1391;
assign _035_ = ap_CS_fsm[11] ? op_4_V_fu_594_p3 : op_4_V_reg_1384;
assign _019_ = ap_CS_fsm[2] ? icmp_ln786_fu_264_p2 : icmp_ln786_reg_1217;
assign _016_ = ap_CS_fsm[2] ? icmp_ln768_fu_259_p2 : icmp_ln768_reg_1212;
assign _014_ = ap_CS_fsm[19] ? icmp_ln768_2_fu_902_p2 : icmp_ln768_2_reg_1594;
assign _080_ = ap_CS_fsm[19] ? grp_fu_704_p2[1:0] : trunc_ln851_reg_1589;
assign _050_ = ap_CS_fsm[19] ? grp_fu_704_p2 : r_V_reg_1583;
assign _017_ = ap_CS_fsm[0] ? icmp_ln786_1_fu_231_p2 : icmp_ln786_1_reg_1176;
assign _013_ = ap_CS_fsm[0] ? icmp_ln768_1_fu_225_p2 : icmp_ln768_1_reg_1171;
assign _043_ = ap_CS_fsm[0] ? op_1[3] : p_Result_15_reg_1164;
assign _079_ = ap_CS_fsm[13] ? op_12_V_fu_738_p3[29:0] : trunc_ln851_2_reg_1463;
assign _028_ = ap_CS_fsm[13] ? op_12_V_fu_738_p3 : op_12_V_reg_1458;
assign _078_ = ap_CS_fsm[13] ? grp_fu_647_p2[1:0] : trunc_ln851_1_reg_1453;
assign _074_ = ap_CS_fsm[13] ? grp_fu_647_p2[4:2] : tmp_2_reg_1448;
assign _053_ = ap_CS_fsm[13] ? grp_fu_647_p2 : ret_V_14_reg_1443;
assign _071_ = ap_CS_fsm[13] ? { ret_V_11_reg_1402[3], ret_V_11_reg_1402[3], ret_V_11_reg_1402[3], ret_V_11_reg_1402[3], ret_V_11_reg_1402[3], ret_V_11_reg_1402[3], ret_V_11_reg_1402[3], ret_V_11_reg_1402[3], ret_V_11_reg_1402[3], ret_V_11_reg_1402[3], ret_V_11_reg_1402[3], ret_V_11_reg_1402[3], ret_V_11_reg_1402 } : sext_ln1118_reg_1433;
assign _012_ = ap_CS_fsm[13] ? icmp_ln1498_fu_688_p2 : icmp_ln1498_reg_1423;
assign _076_ = ap_CS_fsm[8] ? op_8[1:0] : trunc_ln731_2_reg_1321;
assign _072_ = ap_CS_fsm[8] ? { op_8[3], op_8 } : sext_ln1346_reg_1315;
assign _010_ = ap_CS_fsm[8] ? and_ln786_fu_422_p2 : and_ln786_reg_1304;
assign _036_ = ap_CS_fsm[8] ? or_ln340_1_fu_412_p2 : or_ln340_1_reg_1298;
assign _040_ = ap_CS_fsm[8] ? or_ln786_1_fu_407_p2 : or_ln786_1_reg_1292;
assign _009_ = ap_CS_fsm[4] ? and_ln785_1_fu_331_p2 : and_ln785_1_reg_1234;
assign _008_ = ap_CS_fsm[4] ? and_ln340_fu_304_p2 : and_ln340_reg_1229;
assign _055_ = ap_CS_fsm[18] ? ret_V_16_fu_891_p3 : ret_V_16_reg_1578;
assign _029_ = ap_CS_fsm[18] ? grp_fu_864_p2 : op_15_V_reg_1573;
assign _047_ = ap_CS_fsm[18] ? grp_fu_842_p2[32:11] : p_Result_4_reg_1568;
assign _007_ = ap_CS_fsm[18] ? grp_fu_855_p2 : add_ln731_reg_1562;
assign _052_ = ap_CS_fsm[18] ? grp_fu_830_p2 : ret_V_12_reg_1557;
assign _077_ = ap_CS_fsm[10] ? grp_fu_536_p2[0] : trunc_ln790_reg_1379;
assign _018_ = ap_CS_fsm[10] ? icmp_ln786_2_fu_585_p2 : icmp_ln786_2_reg_1374;
assign _015_ = ap_CS_fsm[10] ? icmp_ln768_3_fu_580_p2 : icmp_ln768_3_reg_1369;
assign _046_ = ap_CS_fsm[10] ? grp_fu_536_p2[1] : p_Result_20_reg_1363;
assign _006_ = ap_CS_fsm[10] ? grp_fu_536_p2 : add_ln731_1_reg_1358;
assign _004_ = ap_CS_fsm[20] ? grp_fu_914_p2 : add_ln69_1_reg_1614;
assign _005_ = ap_CS_fsm[20] ? grp_fu_910_p2 : add_ln69_reg_1609;
assign _021_ = ap_CS_fsm[20] ? icmp_ln850_fu_919_p2 : icmp_ln850_reg_1604;
assign _061_ = ap_CS_fsm[15] ? grp_fu_778_p2[61:30] : ret_V_7_cast_reg_1505;
assign _054_ = ap_CS_fsm[15] ? grp_fu_778_p2 : ret_V_15_reg_1500;
assign _003_ = ap_CS_fsm[15] ? grp_fu_757_p2 : add_ln691_reg_1495;
assign _002_ = _085_ ? grp_fu_1120_p2 : add_ln691_3_reg_1728;
assign _001_ = _084_ ? grp_fu_1055_p2 : add_ln691_2_reg_1691;
assign _000_ = _083_ ? grp_fu_825_p2 : add_ln691_1_reg_1552;
assign _011_ = ap_rst ? 37'h0000000001 : ap_NS_fsm;
assign icmp_ln1498_fu_688_p2 = _093_ ? 1'h1 : 1'h0;
assign icmp_ln768_1_fu_225_p2 = _222_ ? 1'h1 : 1'h0;
assign icmp_ln768_2_fu_902_p2 = _223_ ? 1'h1 : 1'h0;
assign icmp_ln768_3_fu_580_p2 = _224_ ? 1'h1 : 1'h0;
assign icmp_ln768_fu_259_p2 = _225_ ? 1'h1 : 1'h0;
assign icmp_ln786_1_fu_231_p2 = _226_ ? 1'h1 : 1'h0;
assign icmp_ln786_2_fu_585_p2 = _227_ ? 1'h1 : 1'h0;
assign icmp_ln786_fu_264_p2 = _228_ ? 1'h1 : 1'h0;
assign icmp_ln790_fu_621_p2 = _094_ ? 1'h1 : 1'h0;
assign icmp_ln850_fu_919_p2 = _229_ ? 1'h1 : 1'h0;
assign icmp_ln851_1_fu_784_p2 = _230_ ? 1'h1 : 1'h0;
assign icmp_ln851_2_fu_1040_p2 = _231_ ? 1'h1 : 1'h0;
assign icmp_ln851_3_fu_1104_p2 = _232_ ? 1'h1 : 1'h0;
assign icmp_ln851_fu_752_p2 = _233_ ? 1'h1 : 1'h0;
assign op_12_V_fu_738_p3 = or_ln384_reg_1418 ? select_ln384_fu_731_p3 : { add_ln731_1_reg_1358, 30'h00000000 };
assign op_16_V_fu_957_p2 = _234_ ? 1'h1 : 1'h0;
assign op_18_V_fu_1008_p3 = overflow_2_fu_1003_p2 ? 32'd0 : { add_ln731_reg_1562, 21'h000000 };
assign op_27 = ret_V_19_reg_1716[46] ? select_ln850_3_fu_1132_p3 : ret_V_20_cast_reg_1721;
assign op_2_V_fu_368_p3 = and_ln785_1_reg_1234 ? newsignbit_reg_1195 : select_ln340_reg_1239;
assign op_4_V_fu_594_p3 = sel_tmp18_reg_1331 ? p_Val2_2_reg_1251 : select_ln785_reg_1353;
assign p_Result_16_fu_378_p2 = op_1[0] ? 1'h1 : 1'h0;
assign ret_V_11_fu_627_p3 = op_2_V_reg_1244 ? 4'hf : op_1;
assign ret_V_16_fu_891_p3 = ret_V_15_reg_1500[62] ? select_ln850_1_fu_886_p3 : ret_V_7_cast_reg_1505;
assign ret_V_fu_818_p3 = ret_V_14_reg_1443[4] ? select_ln850_fu_813_p3 : sext_ln850_reg_1468;
assign select_ln1192_1_fu_970_p3 = op_16_V_reg_1619 ? 32'd4294967295 : 32'd0;
assign select_ln1192_fu_799_p3 = op_2_V_reg_1244 ? 32'd4294967295 : 32'd0;
assign select_ln340_1_fu_498_p3 = and_ln340_1_fu_493_p2 ? p_Val2_2_reg_1251 : { op_1[1], p_Val2_3_fu_473_p2 };
assign select_ln340_fu_362_p3 = and_ln340_reg_1229 ? newsignbit_reg_1195 : select_ln365_fu_355_p3;
assign select_ln353_fu_1072_p3 = ret_V_18_reg_1679[53] ? select_ln850_2_fu_1067_p3 : ret_V_18_cast_reg_1684;
assign select_ln365_fu_355_p3 = xor_ln365_fu_350_p2 ? ret_reg_1182[1] : newsignbit_reg_1195;
assign select_ln384_fu_731_p3 = overflow_3_reg_1391 ? 32'd2147483647 : 32'd2147483649;
assign select_ln785_fu_566_p3 = and_ln785_3_fu_561_p2 ? p_Val2_2_reg_1251 : select_ln340_1_reg_1326;
assign select_ln850_1_fu_886_p3 = icmp_ln851_1_reg_1490 ? add_ln691_1_reg_1552 : ret_V_7_cast_reg_1505;
assign select_ln850_2_fu_1067_p3 = icmp_ln851_2_reg_1674 ? add_ln691_2_reg_1691 : ret_V_18_cast_reg_1684;
assign select_ln850_3_fu_1132_p3 = icmp_ln851_3_reg_1711 ? add_ln691_3_reg_1728 : ret_V_20_cast_reg_1721;
assign select_ln850_fu_813_p3 = icmp_ln851_reg_1475 ? add_ln691_reg_1495 : sext_ln850_reg_1468;
assign select_ln874_fu_949_p3 = ret_V_13_fu_943_p2 ? 4'hf : 4'h0;
assign ret_V_13_fu_943_p2 = r_V_reg_1583[2] ^ and_ln353_fu_938_p2;
assign xor_ln365_1_fu_461_p2 = op_1[0] ^ op_1[1];
assign xor_ln365_fu_350_p2 = ret_reg_1182[1] ^ newsignbit_reg_1195;
assign ap_CS_fsm_state1 = ap_CS_fsm[0];
assign ap_CS_fsm_state10 = ap_CS_fsm[9];
assign ap_CS_fsm_state11 = ap_CS_fsm[10];
assign ap_CS_fsm_state12 = ap_CS_fsm[11];
assign ap_CS_fsm_state13 = ap_CS_fsm[12];
assign ap_CS_fsm_state14 = ap_CS_fsm[13];
assign ap_CS_fsm_state15 = ap_CS_fsm[14];
assign ap_CS_fsm_state16 = ap_CS_fsm[15];
assign ap_CS_fsm_state17 = ap_CS_fsm[16];
assign ap_CS_fsm_state18 = ap_CS_fsm[17];
assign ap_CS_fsm_state19 = ap_CS_fsm[18];
assign ap_CS_fsm_state2 = ap_CS_fsm[1];
assign ap_CS_fsm_state20 = ap_CS_fsm[19];
assign ap_CS_fsm_state21 = ap_CS_fsm[20];
assign ap_CS_fsm_state22 = ap_CS_fsm[21];
assign ap_CS_fsm_state23 = ap_CS_fsm[22];
assign ap_CS_fsm_state24 = ap_CS_fsm[23];
assign ap_CS_fsm_state25 = ap_CS_fsm[24];
assign ap_CS_fsm_state26 = ap_CS_fsm[25];
assign ap_CS_fsm_state27 = ap_CS_fsm[26];
assign ap_CS_fsm_state28 = ap_CS_fsm[27];
assign ap_CS_fsm_state29 = ap_CS_fsm[28];
assign ap_CS_fsm_state3 = ap_CS_fsm[2];
assign ap_CS_fsm_state30 = ap_CS_fsm[29];
assign ap_CS_fsm_state31 = ap_CS_fsm[30];
assign ap_CS_fsm_state32 = ap_CS_fsm[31];
assign ap_CS_fsm_state33 = ap_CS_fsm[32];
assign ap_CS_fsm_state34 = ap_CS_fsm[33];
assign ap_CS_fsm_state35 = ap_CS_fsm[34];
assign ap_CS_fsm_state36 = ap_CS_fsm[35];
assign ap_CS_fsm_state37 = ap_CS_fsm[36];
assign ap_CS_fsm_state4 = ap_CS_fsm[3];
assign ap_CS_fsm_state5 = ap_CS_fsm[4];
assign ap_CS_fsm_state6 = ap_CS_fsm[5];
assign ap_CS_fsm_state7 = ap_CS_fsm[6];
assign ap_CS_fsm_state8 = ap_CS_fsm[7];
assign ap_CS_fsm_state9 = ap_CS_fsm[8];
assign ap_done = op_27_ap_vld;
assign ap_ready = op_27_ap_vld;
assign grp_fu_1034_p0 = { op_25_V_reg_1654[31], op_25_V_reg_1654, 21'h000000 };
assign grp_fu_1034_p1 = { 22'h000000, op_18_V_reg_1649 };
assign grp_fu_1094_p0 = { select_ln353_reg_1696[31], select_ln353_reg_1696, 14'h0000 };
assign grp_fu_1094_p1 = { op_19[15], op_19[15], op_19[15], op_19[15], op_19[15], op_19[15], op_19[15], op_19[15], op_19[15], op_19[15], op_19[15], op_19[15], op_19[15], op_19[15], op_19[15], op_19[15], op_19[15], op_19[15], op_19[15], op_19[15], op_19[15], op_19[15], op_19[15], op_19[15], op_19[15], op_19[15], op_19[15], op_19[15], op_19[15], op_19[15], op_19[15], op_19 };
assign grp_fu_201_p0 = { op_0[3], op_0 };
assign grp_fu_201_p1 = { op_1[3], op_1 };
assign grp_fu_434_p0 = { op_8[3], op_8 };
assign grp_fu_434_p1 = { 4'h0, lhs_V_3_reg_1278 };
assign grp_fu_536_p1 = { 1'h0, lhs_V_3_reg_1278 };
assign grp_fu_647_p0 = { op_4_V_reg_1384[3], op_4_V_reg_1384 };
assign grp_fu_647_p1 = { 2'h0, lhs_V_3_reg_1278, 2'h0 };
assign grp_fu_704_p0 = { ret_V_11_reg_1402[3], ret_V_11_reg_1402[3], ret_V_11_reg_1402[3], ret_V_11_reg_1402[3], ret_V_11_reg_1402[3], ret_V_11_reg_1402[3], ret_V_11_reg_1402[3], ret_V_11_reg_1402[3], ret_V_11_reg_1402[3], ret_V_11_reg_1402[3], ret_V_11_reg_1402[3], ret_V_11_reg_1402[3], ret_V_11_reg_1402 };
assign grp_fu_704_p00 = { 4'h0, ret_V_11_reg_1402[3], ret_V_11_reg_1402[3], ret_V_11_reg_1402[3], ret_V_11_reg_1402[3], ret_V_11_reg_1402[3], ret_V_11_reg_1402[3], ret_V_11_reg_1402[3], ret_V_11_reg_1402[3], ret_V_11_reg_1402[3], ret_V_11_reg_1402[3], ret_V_11_reg_1402[3], ret_V_11_reg_1402[3], ret_V_11_reg_1402 };
assign grp_fu_757_p0 = { tmp_2_reg_1448[2], tmp_2_reg_1448 };
assign grp_fu_778_p0 = { op_7[31], op_7, 30'h00000000 };
assign grp_fu_778_p1 = { op_12_V_reg_1458[31], op_12_V_reg_1458[31], op_12_V_reg_1458[31], op_12_V_reg_1458[31], op_12_V_reg_1458[31], op_12_V_reg_1458[31], op_12_V_reg_1458[31], op_12_V_reg_1458[31], op_12_V_reg_1458[31], op_12_V_reg_1458[31], op_12_V_reg_1458[31], op_12_V_reg_1458[31], op_12_V_reg_1458[31], op_12_V_reg_1458[31], op_12_V_reg_1458[31], op_12_V_reg_1458[31], op_12_V_reg_1458[31], op_12_V_reg_1458[31], op_12_V_reg_1458[31], op_12_V_reg_1458[31], op_12_V_reg_1458[31], op_12_V_reg_1458[31], op_12_V_reg_1458[31], op_12_V_reg_1458[31], op_12_V_reg_1458[31], op_12_V_reg_1458[31], op_12_V_reg_1458[31], op_12_V_reg_1458[31], op_12_V_reg_1458[31], op_12_V_reg_1458[31], op_12_V_reg_1458[31], op_12_V_reg_1458 };
assign grp_fu_842_p0 = { 1'h0, op_9 };
assign grp_fu_842_p1 = { 17'h00000, sext_ln1118_reg_1433 };
assign grp_fu_855_p0 = op_9[10:0];
assign grp_fu_855_p1 = { ret_V_11_reg_1402[3], ret_V_11_reg_1402[3], ret_V_11_reg_1402[3], ret_V_11_reg_1402[3], ret_V_11_reg_1402[3], ret_V_11_reg_1402[3], ret_V_11_reg_1402[3], ret_V_11_reg_1402 };
assign grp_fu_864_p1 = { ret_V_reg_1517[3], ret_V_reg_1517 };
assign grp_fu_914_p1 = { 4'h0, icmp_ln1498_reg_1423 };
assign grp_fu_965_p0 = { add_ln69_1_reg_1614[4], add_ln69_1_reg_1614[4], add_ln69_1_reg_1614[4], add_ln69_1_reg_1614[4], add_ln69_1_reg_1614[4], add_ln69_1_reg_1614[4], add_ln69_1_reg_1614[4], add_ln69_1_reg_1614[4], add_ln69_1_reg_1614[4], add_ln69_1_reg_1614[4], add_ln69_1_reg_1614[4], add_ln69_1_reg_1614[4], add_ln69_1_reg_1614[4], add_ln69_1_reg_1614[4], add_ln69_1_reg_1614[4], add_ln69_1_reg_1614[4], add_ln69_1_reg_1614[4], add_ln69_1_reg_1614[4], add_ln69_1_reg_1614[4], add_ln69_1_reg_1614[4], add_ln69_1_reg_1614[4], add_ln69_1_reg_1614[4], add_ln69_1_reg_1614[4], add_ln69_1_reg_1614[4], add_ln69_1_reg_1614[4], add_ln69_1_reg_1614[4], add_ln69_1_reg_1614[4], add_ln69_1_reg_1614 };
assign grp_fu_984_p1 = { 31'h00000000, lhs_V_3_reg_1278 };
assign lhs_V_4_fu_763_p3 = { op_7, 30'h00000000 };
assign newsignbit_fu_245_p1 = grp_fu_201_p2[0];
assign op_16_V_fu_957_p1 = op_8;
assign p_Result_10_fu_879_p3 = ret_V_15_reg_1500[62];
assign p_Result_11_fu_1060_p3 = ret_V_18_reg_1679[53];
assign p_Result_12_fu_1125_p3 = ret_V_19_reg_1716[46];
assign p_Result_14_fu_336_p3 = ret_reg_1182[1];
assign p_Result_15_fu_207_p1 = op_1;
assign p_Result_17_fu_447_p1 = op_1;
assign p_Result_17_fu_447_p3 = op_1[1];
assign p_Result_18_fu_996_p3 = add_ln731_reg_1562[10];
assign p_Result_1_fu_215_p1 = op_1;
assign p_Result_1_fu_215_p4 = op_1[3:1];
assign p_Result_3_fu_931_p3 = r_V_reg_1583[19];
assign p_Result_6_fu_806_p3 = ret_V_14_reg_1443[4];
assign p_Result_8_fu_614_p3 = { trunc_ln790_reg_1379, 30'h00000000 };
assign p_Result_s_16_fu_478_p4 = { op_1[1], p_Val2_3_fu_473_p2 };
assign p_Val2_11_fu_724_p3 = { add_ln731_1_reg_1358, 30'h00000000 };
assign p_Val2_2_fu_373_p0 = op_1;
assign p_Val2_2_fu_373_p2 = { op_1[0], 3'h0 };
assign p_Val2_7_fu_989_p3 = { add_ln731_reg_1562, 21'h000000 };
assign ret_V_11_fu_627_p2 = op_1;
assign rhs_1_fu_636_p3 = { lhs_V_3_reg_1278, 2'h0 };
assign rhs_4_fu_1023_p3 = { op_25_V_reg_1654, 21'h000000 };
assign rhs_5_fu_1083_p3 = { select_ln353_reg_1696, 14'h0000 };
assign sext_ln1118_fu_697_p1 = { ret_V_11_reg_1402[3], ret_V_11_reg_1402[3], ret_V_11_reg_1402[3], ret_V_11_reg_1402[3], ret_V_11_reg_1402[3], ret_V_11_reg_1402[3], ret_V_11_reg_1402[3], ret_V_11_reg_1402[3], ret_V_11_reg_1402[3], ret_V_11_reg_1402[3], ret_V_11_reg_1402[3], ret_V_11_reg_1402[3], ret_V_11_reg_1402 };
assign sext_ln1346_fu_430_p0 = op_8;
assign sext_ln1346_fu_430_p1 = { op_8[3], op_8 };
assign sext_ln1347_fu_197_p0 = op_1;
assign sext_ln703_1_fu_1079_p0 = op_19;
assign sext_ln727_fu_678_p1 = { op_4_V_reg_1384[3], op_4_V_reg_1384[3], op_4_V_reg_1384 };
assign sext_ln850_fu_749_p1 = { tmp_2_reg_1448[2], tmp_2_reg_1448 };
assign shl_ln_fu_681_p1 = op_8;
assign shl_ln_fu_681_p3 = { op_8, 2'h0 };
assign tmp_5_fu_454_p1 = op_1;
assign tmp_5_fu_454_p3 = op_1[1];
assign tmp_7_fu_924_p3 = r_V_reg_1583[2];
assign tmp_fu_343_p3 = ret_reg_1182[1];
assign trunc_ln731_2_fu_440_p0 = op_8;
assign trunc_ln731_2_fu_440_p1 = op_8[1:0];
assign trunc_ln731_fu_444_p0 = op_1;
assign trunc_ln731_fu_444_p1 = op_1[0];
assign trunc_ln790_fu_590_p1 = grp_fu_536_p2[0];
assign trunc_ln851_1_fu_720_p1 = grp_fu_647_p2[1:0];
assign trunc_ln851_2_fu_745_p1 = op_12_V_fu_738_p3[29:0];
assign trunc_ln851_3_fu_1016_p1 = op_18_V_fu_1008_p3[20:0];
assign trunc_ln851_4_fu_1100_p0 = op_19;
assign trunc_ln851_4_fu_1100_p1 = op_19[13:0];
assign trunc_ln851_fu_898_p1 = grp_fu_704_p2[1:0];
assign \sub_5s_5s_5_2_1_U12.top_sub_5s_5s_5_2_1_Adder_0_U.ain_s0  = \sub_5s_5s_5_2_1_U12.top_sub_5s_5s_5_2_1_Adder_0_U.a ;
assign \sub_5s_5s_5_2_1_U12.top_sub_5s_5s_5_2_1_Adder_0_U.s  = { \sub_5s_5s_5_2_1_U12.top_sub_5s_5s_5_2_1_Adder_0_U.fas_s2 , \sub_5s_5s_5_2_1_U12.top_sub_5s_5s_5_2_1_Adder_0_U.sum_s1  };
assign \sub_5s_5s_5_2_1_U12.top_sub_5s_5s_5_2_1_Adder_0_U.u2.a  = \sub_5s_5s_5_2_1_U12.top_sub_5s_5s_5_2_1_Adder_0_U.ain_s1 ;
assign \sub_5s_5s_5_2_1_U12.top_sub_5s_5s_5_2_1_Adder_0_U.u2.b  = \sub_5s_5s_5_2_1_U12.top_sub_5s_5s_5_2_1_Adder_0_U.bin_s1 ;
assign \sub_5s_5s_5_2_1_U12.top_sub_5s_5s_5_2_1_Adder_0_U.u2.cin  = \sub_5s_5s_5_2_1_U12.top_sub_5s_5s_5_2_1_Adder_0_U.carry_s1 ;
assign \sub_5s_5s_5_2_1_U12.top_sub_5s_5s_5_2_1_Adder_0_U.facout_s2  = \sub_5s_5s_5_2_1_U12.top_sub_5s_5s_5_2_1_Adder_0_U.u2.cout ;
assign \sub_5s_5s_5_2_1_U12.top_sub_5s_5s_5_2_1_Adder_0_U.fas_s2  = \sub_5s_5s_5_2_1_U12.top_sub_5s_5s_5_2_1_Adder_0_U.u2.s ;
assign \sub_5s_5s_5_2_1_U12.top_sub_5s_5s_5_2_1_Adder_0_U.u1.a  = \sub_5s_5s_5_2_1_U12.top_sub_5s_5s_5_2_1_Adder_0_U.a [1:0];
assign \sub_5s_5s_5_2_1_U12.top_sub_5s_5s_5_2_1_Adder_0_U.u1.b  = \sub_5s_5s_5_2_1_U12.top_sub_5s_5s_5_2_1_Adder_0_U.bin_s0 [1:0];
assign \sub_5s_5s_5_2_1_U12.top_sub_5s_5s_5_2_1_Adder_0_U.u1.cin  = 1'h1;
assign \sub_5s_5s_5_2_1_U12.top_sub_5s_5s_5_2_1_Adder_0_U.facout_s1  = \sub_5s_5s_5_2_1_U12.top_sub_5s_5s_5_2_1_Adder_0_U.u1.cout ;
assign \sub_5s_5s_5_2_1_U12.top_sub_5s_5s_5_2_1_Adder_0_U.fas_s1  = \sub_5s_5s_5_2_1_U12.top_sub_5s_5s_5_2_1_Adder_0_U.u1.s ;
assign \sub_5s_5s_5_2_1_U12.top_sub_5s_5s_5_2_1_Adder_0_U.a  = \sub_5s_5s_5_2_1_U12.din0 ;
assign \sub_5s_5s_5_2_1_U12.top_sub_5s_5s_5_2_1_Adder_0_U.b  = \sub_5s_5s_5_2_1_U12.din1 ;
assign \sub_5s_5s_5_2_1_U12.top_sub_5s_5s_5_2_1_Adder_0_U.ce  = \sub_5s_5s_5_2_1_U12.ce ;
assign \sub_5s_5s_5_2_1_U12.top_sub_5s_5s_5_2_1_Adder_0_U.clk  = \sub_5s_5s_5_2_1_U12.clk ;
assign \sub_5s_5s_5_2_1_U12.top_sub_5s_5s_5_2_1_Adder_0_U.reset  = \sub_5s_5s_5_2_1_U12.reset ;
assign \sub_5s_5s_5_2_1_U12.dout  = \sub_5s_5s_5_2_1_U12.top_sub_5s_5s_5_2_1_Adder_0_U.s ;
assign \sub_5s_5s_5_2_1_U12.ce  = 1'h1;
assign \sub_5s_5s_5_2_1_U12.clk  = ap_clk;
assign \sub_5s_5s_5_2_1_U12.din0  = sext_ln1346_reg_1315;
assign \sub_5s_5s_5_2_1_U12.din1  = { ret_V_reg_1517[3], ret_V_reg_1517 };
assign grp_fu_864_p2 = \sub_5s_5s_5_2_1_U12.dout ;
assign \sub_5s_5s_5_2_1_U12.reset  = ap_rst;
assign \sub_5s_5s_5_2_1_U1.top_sub_5s_5s_5_2_1_Adder_0_U.ain_s0  = \sub_5s_5s_5_2_1_U1.top_sub_5s_5s_5_2_1_Adder_0_U.a ;
assign \sub_5s_5s_5_2_1_U1.top_sub_5s_5s_5_2_1_Adder_0_U.s  = { \sub_5s_5s_5_2_1_U1.top_sub_5s_5s_5_2_1_Adder_0_U.fas_s2 , \sub_5s_5s_5_2_1_U1.top_sub_5s_5s_5_2_1_Adder_0_U.sum_s1  };
assign \sub_5s_5s_5_2_1_U1.top_sub_5s_5s_5_2_1_Adder_0_U.u2.a  = \sub_5s_5s_5_2_1_U1.top_sub_5s_5s_5_2_1_Adder_0_U.ain_s1 ;
assign \sub_5s_5s_5_2_1_U1.top_sub_5s_5s_5_2_1_Adder_0_U.u2.b  = \sub_5s_5s_5_2_1_U1.top_sub_5s_5s_5_2_1_Adder_0_U.bin_s1 ;
assign \sub_5s_5s_5_2_1_U1.top_sub_5s_5s_5_2_1_Adder_0_U.u2.cin  = \sub_5s_5s_5_2_1_U1.top_sub_5s_5s_5_2_1_Adder_0_U.carry_s1 ;
assign \sub_5s_5s_5_2_1_U1.top_sub_5s_5s_5_2_1_Adder_0_U.facout_s2  = \sub_5s_5s_5_2_1_U1.top_sub_5s_5s_5_2_1_Adder_0_U.u2.cout ;
assign \sub_5s_5s_5_2_1_U1.top_sub_5s_5s_5_2_1_Adder_0_U.fas_s2  = \sub_5s_5s_5_2_1_U1.top_sub_5s_5s_5_2_1_Adder_0_U.u2.s ;
assign \sub_5s_5s_5_2_1_U1.top_sub_5s_5s_5_2_1_Adder_0_U.u1.a  = \sub_5s_5s_5_2_1_U1.top_sub_5s_5s_5_2_1_Adder_0_U.a [1:0];
assign \sub_5s_5s_5_2_1_U1.top_sub_5s_5s_5_2_1_Adder_0_U.u1.b  = \sub_5s_5s_5_2_1_U1.top_sub_5s_5s_5_2_1_Adder_0_U.bin_s0 [1:0];
assign \sub_5s_5s_5_2_1_U1.top_sub_5s_5s_5_2_1_Adder_0_U.u1.cin  = 1'h1;
assign \sub_5s_5s_5_2_1_U1.top_sub_5s_5s_5_2_1_Adder_0_U.facout_s1  = \sub_5s_5s_5_2_1_U1.top_sub_5s_5s_5_2_1_Adder_0_U.u1.cout ;
assign \sub_5s_5s_5_2_1_U1.top_sub_5s_5s_5_2_1_Adder_0_U.fas_s1  = \sub_5s_5s_5_2_1_U1.top_sub_5s_5s_5_2_1_Adder_0_U.u1.s ;
assign \sub_5s_5s_5_2_1_U1.top_sub_5s_5s_5_2_1_Adder_0_U.a  = \sub_5s_5s_5_2_1_U1.din0 ;
assign \sub_5s_5s_5_2_1_U1.top_sub_5s_5s_5_2_1_Adder_0_U.b  = \sub_5s_5s_5_2_1_U1.din1 ;
assign \sub_5s_5s_5_2_1_U1.top_sub_5s_5s_5_2_1_Adder_0_U.ce  = \sub_5s_5s_5_2_1_U1.ce ;
assign \sub_5s_5s_5_2_1_U1.top_sub_5s_5s_5_2_1_Adder_0_U.clk  = \sub_5s_5s_5_2_1_U1.clk ;
assign \sub_5s_5s_5_2_1_U1.top_sub_5s_5s_5_2_1_Adder_0_U.reset  = \sub_5s_5s_5_2_1_U1.reset ;
assign \sub_5s_5s_5_2_1_U1.dout  = \sub_5s_5s_5_2_1_U1.top_sub_5s_5s_5_2_1_Adder_0_U.s ;
assign \sub_5s_5s_5_2_1_U1.ce  = 1'h1;
assign \sub_5s_5s_5_2_1_U1.clk  = ap_clk;
assign \sub_5s_5s_5_2_1_U1.din0  = { op_0[3], op_0 };
assign \sub_5s_5s_5_2_1_U1.din1  = { op_1[3], op_1 };
assign grp_fu_201_p2 = \sub_5s_5s_5_2_1_U1.dout ;
assign \sub_5s_5s_5_2_1_U1.reset  = ap_rst;
assign \sub_5s_5ns_5_2_1_U4.top_sub_5s_5ns_5_2_1_Adder_3_U.ain_s0  = \sub_5s_5ns_5_2_1_U4.top_sub_5s_5ns_5_2_1_Adder_3_U.a ;
assign \sub_5s_5ns_5_2_1_U4.top_sub_5s_5ns_5_2_1_Adder_3_U.s  = { \sub_5s_5ns_5_2_1_U4.top_sub_5s_5ns_5_2_1_Adder_3_U.fas_s2 , \sub_5s_5ns_5_2_1_U4.top_sub_5s_5ns_5_2_1_Adder_3_U.sum_s1  };
assign \sub_5s_5ns_5_2_1_U4.top_sub_5s_5ns_5_2_1_Adder_3_U.u2.a  = \sub_5s_5ns_5_2_1_U4.top_sub_5s_5ns_5_2_1_Adder_3_U.ain_s1 ;
assign \sub_5s_5ns_5_2_1_U4.top_sub_5s_5ns_5_2_1_Adder_3_U.u2.b  = \sub_5s_5ns_5_2_1_U4.top_sub_5s_5ns_5_2_1_Adder_3_U.bin_s1 ;
assign \sub_5s_5ns_5_2_1_U4.top_sub_5s_5ns_5_2_1_Adder_3_U.u2.cin  = \sub_5s_5ns_5_2_1_U4.top_sub_5s_5ns_5_2_1_Adder_3_U.carry_s1 ;
assign \sub_5s_5ns_5_2_1_U4.top_sub_5s_5ns_5_2_1_Adder_3_U.facout_s2  = \sub_5s_5ns_5_2_1_U4.top_sub_5s_5ns_5_2_1_Adder_3_U.u2.cout ;
assign \sub_5s_5ns_5_2_1_U4.top_sub_5s_5ns_5_2_1_Adder_3_U.fas_s2  = \sub_5s_5ns_5_2_1_U4.top_sub_5s_5ns_5_2_1_Adder_3_U.u2.s ;
assign \sub_5s_5ns_5_2_1_U4.top_sub_5s_5ns_5_2_1_Adder_3_U.u1.a  = \sub_5s_5ns_5_2_1_U4.top_sub_5s_5ns_5_2_1_Adder_3_U.a [1:0];
assign \sub_5s_5ns_5_2_1_U4.top_sub_5s_5ns_5_2_1_Adder_3_U.u1.b  = \sub_5s_5ns_5_2_1_U4.top_sub_5s_5ns_5_2_1_Adder_3_U.bin_s0 [1:0];
assign \sub_5s_5ns_5_2_1_U4.top_sub_5s_5ns_5_2_1_Adder_3_U.u1.cin  = 1'h1;
assign \sub_5s_5ns_5_2_1_U4.top_sub_5s_5ns_5_2_1_Adder_3_U.facout_s1  = \sub_5s_5ns_5_2_1_U4.top_sub_5s_5ns_5_2_1_Adder_3_U.u1.cout ;
assign \sub_5s_5ns_5_2_1_U4.top_sub_5s_5ns_5_2_1_Adder_3_U.fas_s1  = \sub_5s_5ns_5_2_1_U4.top_sub_5s_5ns_5_2_1_Adder_3_U.u1.s ;
assign \sub_5s_5ns_5_2_1_U4.top_sub_5s_5ns_5_2_1_Adder_3_U.a  = \sub_5s_5ns_5_2_1_U4.din0 ;
assign \sub_5s_5ns_5_2_1_U4.top_sub_5s_5ns_5_2_1_Adder_3_U.b  = \sub_5s_5ns_5_2_1_U4.din1 ;
assign \sub_5s_5ns_5_2_1_U4.top_sub_5s_5ns_5_2_1_Adder_3_U.ce  = \sub_5s_5ns_5_2_1_U4.ce ;
assign \sub_5s_5ns_5_2_1_U4.top_sub_5s_5ns_5_2_1_Adder_3_U.clk  = \sub_5s_5ns_5_2_1_U4.clk ;
assign \sub_5s_5ns_5_2_1_U4.top_sub_5s_5ns_5_2_1_Adder_3_U.reset  = \sub_5s_5ns_5_2_1_U4.reset ;
assign \sub_5s_5ns_5_2_1_U4.dout  = \sub_5s_5ns_5_2_1_U4.top_sub_5s_5ns_5_2_1_Adder_3_U.s ;
assign \sub_5s_5ns_5_2_1_U4.ce  = 1'h1;
assign \sub_5s_5ns_5_2_1_U4.clk  = ap_clk;
assign \sub_5s_5ns_5_2_1_U4.din0  = { op_4_V_reg_1384[3], op_4_V_reg_1384 };
assign \sub_5s_5ns_5_2_1_U4.din1  = { 2'h0, lhs_V_3_reg_1278, 2'h0 };
assign grp_fu_647_p2 = \sub_5s_5ns_5_2_1_U4.dout ;
assign \sub_5s_5ns_5_2_1_U4.reset  = ap_rst;
assign \mul_16ns_4s_20_7_1_U5.top_mul_16ns_4s_20_7_1_Mul_DSP_0_U.p  = \mul_16ns_4s_20_7_1_U5.top_mul_16ns_4s_20_7_1_Mul_DSP_0_U.buff4 ;
assign \mul_16ns_4s_20_7_1_U5.top_mul_16ns_4s_20_7_1_Mul_DSP_0_U.a  = \mul_16ns_4s_20_7_1_U5.din0 ;
assign \mul_16ns_4s_20_7_1_U5.top_mul_16ns_4s_20_7_1_Mul_DSP_0_U.b  = \mul_16ns_4s_20_7_1_U5.din1 ;
assign \mul_16ns_4s_20_7_1_U5.top_mul_16ns_4s_20_7_1_Mul_DSP_0_U.ce  = \mul_16ns_4s_20_7_1_U5.ce ;
assign \mul_16ns_4s_20_7_1_U5.top_mul_16ns_4s_20_7_1_Mul_DSP_0_U.clk  = \mul_16ns_4s_20_7_1_U5.clk ;
assign \mul_16ns_4s_20_7_1_U5.dout  = \mul_16ns_4s_20_7_1_U5.top_mul_16ns_4s_20_7_1_Mul_DSP_0_U.p ;
assign \mul_16ns_4s_20_7_1_U5.ce  = 1'h1;
assign \mul_16ns_4s_20_7_1_U5.clk  = ap_clk;
assign \mul_16ns_4s_20_7_1_U5.din0  = { ret_V_11_reg_1402[3], ret_V_11_reg_1402[3], ret_V_11_reg_1402[3], ret_V_11_reg_1402[3], ret_V_11_reg_1402[3], ret_V_11_reg_1402[3], ret_V_11_reg_1402[3], ret_V_11_reg_1402[3], ret_V_11_reg_1402[3], ret_V_11_reg_1402[3], ret_V_11_reg_1402[3], ret_V_11_reg_1402[3], ret_V_11_reg_1402 };
assign \mul_16ns_4s_20_7_1_U5.din1  = op_4_V_reg_1384;
assign grp_fu_704_p2 = \mul_16ns_4s_20_7_1_U5.dout ;
assign \mul_16ns_4s_20_7_1_U5.reset  = ap_rst;
assign \add_63s_63s_63_2_1_U7.top_add_63s_63s_63_2_1_Adder_5_U.ain_s0  = \add_63s_63s_63_2_1_U7.top_add_63s_63s_63_2_1_Adder_5_U.a ;
assign \add_63s_63s_63_2_1_U7.top_add_63s_63s_63_2_1_Adder_5_U.bin_s0  = \add_63s_63s_63_2_1_U7.top_add_63s_63s_63_2_1_Adder_5_U.b ;
assign \add_63s_63s_63_2_1_U7.top_add_63s_63s_63_2_1_Adder_5_U.s  = { \add_63s_63s_63_2_1_U7.top_add_63s_63s_63_2_1_Adder_5_U.fas_s2 , \add_63s_63s_63_2_1_U7.top_add_63s_63s_63_2_1_Adder_5_U.sum_s1  };
assign \add_63s_63s_63_2_1_U7.top_add_63s_63s_63_2_1_Adder_5_U.u2.a  = \add_63s_63s_63_2_1_U7.top_add_63s_63s_63_2_1_Adder_5_U.ain_s1 ;
assign \add_63s_63s_63_2_1_U7.top_add_63s_63s_63_2_1_Adder_5_U.u2.b  = \add_63s_63s_63_2_1_U7.top_add_63s_63s_63_2_1_Adder_5_U.bin_s1 ;
assign \add_63s_63s_63_2_1_U7.top_add_63s_63s_63_2_1_Adder_5_U.u2.cin  = \add_63s_63s_63_2_1_U7.top_add_63s_63s_63_2_1_Adder_5_U.carry_s1 ;
assign \add_63s_63s_63_2_1_U7.top_add_63s_63s_63_2_1_Adder_5_U.facout_s2  = \add_63s_63s_63_2_1_U7.top_add_63s_63s_63_2_1_Adder_5_U.u2.cout ;
assign \add_63s_63s_63_2_1_U7.top_add_63s_63s_63_2_1_Adder_5_U.fas_s2  = \add_63s_63s_63_2_1_U7.top_add_63s_63s_63_2_1_Adder_5_U.u2.s ;
assign \add_63s_63s_63_2_1_U7.top_add_63s_63s_63_2_1_Adder_5_U.u1.a  = \add_63s_63s_63_2_1_U7.top_add_63s_63s_63_2_1_Adder_5_U.a [30:0];
assign \add_63s_63s_63_2_1_U7.top_add_63s_63s_63_2_1_Adder_5_U.u1.b  = \add_63s_63s_63_2_1_U7.top_add_63s_63s_63_2_1_Adder_5_U.b [30:0];
assign \add_63s_63s_63_2_1_U7.top_add_63s_63s_63_2_1_Adder_5_U.u1.cin  = 1'h0;
assign \add_63s_63s_63_2_1_U7.top_add_63s_63s_63_2_1_Adder_5_U.facout_s1  = \add_63s_63s_63_2_1_U7.top_add_63s_63s_63_2_1_Adder_5_U.u1.cout ;
assign \add_63s_63s_63_2_1_U7.top_add_63s_63s_63_2_1_Adder_5_U.fas_s1  = \add_63s_63s_63_2_1_U7.top_add_63s_63s_63_2_1_Adder_5_U.u1.s ;
assign \add_63s_63s_63_2_1_U7.top_add_63s_63s_63_2_1_Adder_5_U.a  = \add_63s_63s_63_2_1_U7.din0 ;
assign \add_63s_63s_63_2_1_U7.top_add_63s_63s_63_2_1_Adder_5_U.b  = \add_63s_63s_63_2_1_U7.din1 ;
assign \add_63s_63s_63_2_1_U7.top_add_63s_63s_63_2_1_Adder_5_U.ce  = \add_63s_63s_63_2_1_U7.ce ;
assign \add_63s_63s_63_2_1_U7.top_add_63s_63s_63_2_1_Adder_5_U.clk  = \add_63s_63s_63_2_1_U7.clk ;
assign \add_63s_63s_63_2_1_U7.top_add_63s_63s_63_2_1_Adder_5_U.reset  = \add_63s_63s_63_2_1_U7.reset ;
assign \add_63s_63s_63_2_1_U7.dout  = \add_63s_63s_63_2_1_U7.top_add_63s_63s_63_2_1_Adder_5_U.s ;
assign \add_63s_63s_63_2_1_U7.ce  = 1'h1;
assign \add_63s_63s_63_2_1_U7.clk  = ap_clk;
assign \add_63s_63s_63_2_1_U7.din0  = { op_7[31], op_7, 30'h00000000 };
assign \add_63s_63s_63_2_1_U7.din1  = { op_12_V_reg_1458[31], op_12_V_reg_1458[31], op_12_V_reg_1458[31], op_12_V_reg_1458[31], op_12_V_reg_1458[31], op_12_V_reg_1458[31], op_12_V_reg_1458[31], op_12_V_reg_1458[31], op_12_V_reg_1458[31], op_12_V_reg_1458[31], op_12_V_reg_1458[31], op_12_V_reg_1458[31], op_12_V_reg_1458[31], op_12_V_reg_1458[31], op_12_V_reg_1458[31], op_12_V_reg_1458[31], op_12_V_reg_1458[31], op_12_V_reg_1458[31], op_12_V_reg_1458[31], op_12_V_reg_1458[31], op_12_V_reg_1458[31], op_12_V_reg_1458[31], op_12_V_reg_1458[31], op_12_V_reg_1458[31], op_12_V_reg_1458[31], op_12_V_reg_1458[31], op_12_V_reg_1458[31], op_12_V_reg_1458[31], op_12_V_reg_1458[31], op_12_V_reg_1458[31], op_12_V_reg_1458[31], op_12_V_reg_1458 };
assign grp_fu_778_p2 = \add_63s_63s_63_2_1_U7.dout ;
assign \add_63s_63s_63_2_1_U7.reset  = ap_rst;
assign \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.ain_s0  = \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.a ;
assign \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.bin_s0  = \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.b ;
assign \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.s  = { \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.fas_s2 , \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.sum_s1  };
assign \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.u2.a  = \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.ain_s1 ;
assign \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.u2.b  = \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.bin_s1 ;
assign \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.u2.cin  = \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.carry_s1 ;
assign \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.facout_s2  = \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.u2.cout ;
assign \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.fas_s2  = \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.u2.s ;
assign \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.u1.a  = \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.a [1:0];
assign \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.u1.b  = \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.b [1:0];
assign \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.u1.cin  = 1'h0;
assign \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.facout_s1  = \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.u1.cout ;
assign \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.fas_s1  = \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.u1.s ;
assign \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.a  = \add_5s_5ns_5_2_1_U2.din0 ;
assign \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.b  = \add_5s_5ns_5_2_1_U2.din1 ;
assign \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.ce  = \add_5s_5ns_5_2_1_U2.ce ;
assign \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.clk  = \add_5s_5ns_5_2_1_U2.clk ;
assign \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.reset  = \add_5s_5ns_5_2_1_U2.reset ;
assign \add_5s_5ns_5_2_1_U2.dout  = \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.s ;
assign \add_5s_5ns_5_2_1_U2.ce  = 1'h1;
assign \add_5s_5ns_5_2_1_U2.clk  = ap_clk;
assign \add_5s_5ns_5_2_1_U2.din0  = { op_8[3], op_8 };
assign \add_5s_5ns_5_2_1_U2.din1  = { 4'h0, lhs_V_3_reg_1278 };
assign grp_fu_434_p2 = \add_5s_5ns_5_2_1_U2.dout ;
assign \add_5s_5ns_5_2_1_U2.reset  = ap_rst;
assign \add_5ns_5ns_5_2_1_U14.top_add_5ns_5ns_5_2_1_Adder_9_U.ain_s0  = \add_5ns_5ns_5_2_1_U14.top_add_5ns_5ns_5_2_1_Adder_9_U.a ;
assign \add_5ns_5ns_5_2_1_U14.top_add_5ns_5ns_5_2_1_Adder_9_U.bin_s0  = \add_5ns_5ns_5_2_1_U14.top_add_5ns_5ns_5_2_1_Adder_9_U.b ;
assign \add_5ns_5ns_5_2_1_U14.top_add_5ns_5ns_5_2_1_Adder_9_U.s  = { \add_5ns_5ns_5_2_1_U14.top_add_5ns_5ns_5_2_1_Adder_9_U.fas_s2 , \add_5ns_5ns_5_2_1_U14.top_add_5ns_5ns_5_2_1_Adder_9_U.sum_s1  };
assign \add_5ns_5ns_5_2_1_U14.top_add_5ns_5ns_5_2_1_Adder_9_U.u2.a  = \add_5ns_5ns_5_2_1_U14.top_add_5ns_5ns_5_2_1_Adder_9_U.ain_s1 ;
assign \add_5ns_5ns_5_2_1_U14.top_add_5ns_5ns_5_2_1_Adder_9_U.u2.b  = \add_5ns_5ns_5_2_1_U14.top_add_5ns_5ns_5_2_1_Adder_9_U.bin_s1 ;
assign \add_5ns_5ns_5_2_1_U14.top_add_5ns_5ns_5_2_1_Adder_9_U.u2.cin  = \add_5ns_5ns_5_2_1_U14.top_add_5ns_5ns_5_2_1_Adder_9_U.carry_s1 ;
assign \add_5ns_5ns_5_2_1_U14.top_add_5ns_5ns_5_2_1_Adder_9_U.facout_s2  = \add_5ns_5ns_5_2_1_U14.top_add_5ns_5ns_5_2_1_Adder_9_U.u2.cout ;
assign \add_5ns_5ns_5_2_1_U14.top_add_5ns_5ns_5_2_1_Adder_9_U.fas_s2  = \add_5ns_5ns_5_2_1_U14.top_add_5ns_5ns_5_2_1_Adder_9_U.u2.s ;
assign \add_5ns_5ns_5_2_1_U14.top_add_5ns_5ns_5_2_1_Adder_9_U.u1.a  = \add_5ns_5ns_5_2_1_U14.top_add_5ns_5ns_5_2_1_Adder_9_U.a [1:0];
assign \add_5ns_5ns_5_2_1_U14.top_add_5ns_5ns_5_2_1_Adder_9_U.u1.b  = \add_5ns_5ns_5_2_1_U14.top_add_5ns_5ns_5_2_1_Adder_9_U.b [1:0];
assign \add_5ns_5ns_5_2_1_U14.top_add_5ns_5ns_5_2_1_Adder_9_U.u1.cin  = 1'h0;
assign \add_5ns_5ns_5_2_1_U14.top_add_5ns_5ns_5_2_1_Adder_9_U.facout_s1  = \add_5ns_5ns_5_2_1_U14.top_add_5ns_5ns_5_2_1_Adder_9_U.u1.cout ;
assign \add_5ns_5ns_5_2_1_U14.top_add_5ns_5ns_5_2_1_Adder_9_U.fas_s1  = \add_5ns_5ns_5_2_1_U14.top_add_5ns_5ns_5_2_1_Adder_9_U.u1.s ;
assign \add_5ns_5ns_5_2_1_U14.top_add_5ns_5ns_5_2_1_Adder_9_U.a  = \add_5ns_5ns_5_2_1_U14.din0 ;
assign \add_5ns_5ns_5_2_1_U14.top_add_5ns_5ns_5_2_1_Adder_9_U.b  = \add_5ns_5ns_5_2_1_U14.din1 ;
assign \add_5ns_5ns_5_2_1_U14.top_add_5ns_5ns_5_2_1_Adder_9_U.ce  = \add_5ns_5ns_5_2_1_U14.ce ;
assign \add_5ns_5ns_5_2_1_U14.top_add_5ns_5ns_5_2_1_Adder_9_U.clk  = \add_5ns_5ns_5_2_1_U14.clk ;
assign \add_5ns_5ns_5_2_1_U14.top_add_5ns_5ns_5_2_1_Adder_9_U.reset  = \add_5ns_5ns_5_2_1_U14.reset ;
assign \add_5ns_5ns_5_2_1_U14.dout  = \add_5ns_5ns_5_2_1_U14.top_add_5ns_5ns_5_2_1_Adder_9_U.s ;
assign \add_5ns_5ns_5_2_1_U14.ce  = 1'h1;
assign \add_5ns_5ns_5_2_1_U14.clk  = ap_clk;
assign \add_5ns_5ns_5_2_1_U14.din0  = op_15_V_reg_1573;
assign \add_5ns_5ns_5_2_1_U14.din1  = { 4'h0, icmp_ln1498_reg_1423 };
assign grp_fu_914_p2 = \add_5ns_5ns_5_2_1_U14.dout ;
assign \add_5ns_5ns_5_2_1_U14.reset  = ap_rst;
assign \add_54s_54ns_54_2_1_U18.top_add_54s_54ns_54_2_1_Adder_11_U.ain_s0  = \add_54s_54ns_54_2_1_U18.top_add_54s_54ns_54_2_1_Adder_11_U.a ;
assign \add_54s_54ns_54_2_1_U18.top_add_54s_54ns_54_2_1_Adder_11_U.bin_s0  = \add_54s_54ns_54_2_1_U18.top_add_54s_54ns_54_2_1_Adder_11_U.b ;
assign \add_54s_54ns_54_2_1_U18.top_add_54s_54ns_54_2_1_Adder_11_U.s  = { \add_54s_54ns_54_2_1_U18.top_add_54s_54ns_54_2_1_Adder_11_U.fas_s2 , \add_54s_54ns_54_2_1_U18.top_add_54s_54ns_54_2_1_Adder_11_U.sum_s1  };
assign \add_54s_54ns_54_2_1_U18.top_add_54s_54ns_54_2_1_Adder_11_U.u2.a  = \add_54s_54ns_54_2_1_U18.top_add_54s_54ns_54_2_1_Adder_11_U.ain_s1 ;
assign \add_54s_54ns_54_2_1_U18.top_add_54s_54ns_54_2_1_Adder_11_U.u2.b  = \add_54s_54ns_54_2_1_U18.top_add_54s_54ns_54_2_1_Adder_11_U.bin_s1 ;
assign \add_54s_54ns_54_2_1_U18.top_add_54s_54ns_54_2_1_Adder_11_U.u2.cin  = \add_54s_54ns_54_2_1_U18.top_add_54s_54ns_54_2_1_Adder_11_U.carry_s1 ;
assign \add_54s_54ns_54_2_1_U18.top_add_54s_54ns_54_2_1_Adder_11_U.facout_s2  = \add_54s_54ns_54_2_1_U18.top_add_54s_54ns_54_2_1_Adder_11_U.u2.cout ;
assign \add_54s_54ns_54_2_1_U18.top_add_54s_54ns_54_2_1_Adder_11_U.fas_s2  = \add_54s_54ns_54_2_1_U18.top_add_54s_54ns_54_2_1_Adder_11_U.u2.s ;
assign \add_54s_54ns_54_2_1_U18.top_add_54s_54ns_54_2_1_Adder_11_U.u1.a  = \add_54s_54ns_54_2_1_U18.top_add_54s_54ns_54_2_1_Adder_11_U.a [26:0];
assign \add_54s_54ns_54_2_1_U18.top_add_54s_54ns_54_2_1_Adder_11_U.u1.b  = \add_54s_54ns_54_2_1_U18.top_add_54s_54ns_54_2_1_Adder_11_U.b [26:0];
assign \add_54s_54ns_54_2_1_U18.top_add_54s_54ns_54_2_1_Adder_11_U.u1.cin  = 1'h0;
assign \add_54s_54ns_54_2_1_U18.top_add_54s_54ns_54_2_1_Adder_11_U.facout_s1  = \add_54s_54ns_54_2_1_U18.top_add_54s_54ns_54_2_1_Adder_11_U.u1.cout ;
assign \add_54s_54ns_54_2_1_U18.top_add_54s_54ns_54_2_1_Adder_11_U.fas_s1  = \add_54s_54ns_54_2_1_U18.top_add_54s_54ns_54_2_1_Adder_11_U.u1.s ;
assign \add_54s_54ns_54_2_1_U18.top_add_54s_54ns_54_2_1_Adder_11_U.a  = \add_54s_54ns_54_2_1_U18.din0 ;
assign \add_54s_54ns_54_2_1_U18.top_add_54s_54ns_54_2_1_Adder_11_U.b  = \add_54s_54ns_54_2_1_U18.din1 ;
assign \add_54s_54ns_54_2_1_U18.top_add_54s_54ns_54_2_1_Adder_11_U.ce  = \add_54s_54ns_54_2_1_U18.ce ;
assign \add_54s_54ns_54_2_1_U18.top_add_54s_54ns_54_2_1_Adder_11_U.clk  = \add_54s_54ns_54_2_1_U18.clk ;
assign \add_54s_54ns_54_2_1_U18.top_add_54s_54ns_54_2_1_Adder_11_U.reset  = \add_54s_54ns_54_2_1_U18.reset ;
assign \add_54s_54ns_54_2_1_U18.dout  = \add_54s_54ns_54_2_1_U18.top_add_54s_54ns_54_2_1_Adder_11_U.s ;
assign \add_54s_54ns_54_2_1_U18.ce  = 1'h1;
assign \add_54s_54ns_54_2_1_U18.clk  = ap_clk;
assign \add_54s_54ns_54_2_1_U18.din0  = { op_25_V_reg_1654[31], op_25_V_reg_1654, 21'h000000 };
assign \add_54s_54ns_54_2_1_U18.din1  = { 22'h000000, op_18_V_reg_1649 };
assign grp_fu_1034_p2 = \add_54s_54ns_54_2_1_U18.dout ;
assign \add_54s_54ns_54_2_1_U18.reset  = ap_rst;
assign \add_4s_4ns_4_2_1_U6.top_add_4s_4ns_4_2_1_Adder_4_U.ain_s0  = \add_4s_4ns_4_2_1_U6.top_add_4s_4ns_4_2_1_Adder_4_U.a ;
assign \add_4s_4ns_4_2_1_U6.top_add_4s_4ns_4_2_1_Adder_4_U.bin_s0  = \add_4s_4ns_4_2_1_U6.top_add_4s_4ns_4_2_1_Adder_4_U.b ;
assign \add_4s_4ns_4_2_1_U6.top_add_4s_4ns_4_2_1_Adder_4_U.s  = { \add_4s_4ns_4_2_1_U6.top_add_4s_4ns_4_2_1_Adder_4_U.fas_s2 , \add_4s_4ns_4_2_1_U6.top_add_4s_4ns_4_2_1_Adder_4_U.sum_s1  };
assign \add_4s_4ns_4_2_1_U6.top_add_4s_4ns_4_2_1_Adder_4_U.u2.a  = \add_4s_4ns_4_2_1_U6.top_add_4s_4ns_4_2_1_Adder_4_U.ain_s1 ;
assign \add_4s_4ns_4_2_1_U6.top_add_4s_4ns_4_2_1_Adder_4_U.u2.b  = \add_4s_4ns_4_2_1_U6.top_add_4s_4ns_4_2_1_Adder_4_U.bin_s1 ;
assign \add_4s_4ns_4_2_1_U6.top_add_4s_4ns_4_2_1_Adder_4_U.u2.cin  = \add_4s_4ns_4_2_1_U6.top_add_4s_4ns_4_2_1_Adder_4_U.carry_s1 ;
assign \add_4s_4ns_4_2_1_U6.top_add_4s_4ns_4_2_1_Adder_4_U.facout_s2  = \add_4s_4ns_4_2_1_U6.top_add_4s_4ns_4_2_1_Adder_4_U.u2.cout ;
assign \add_4s_4ns_4_2_1_U6.top_add_4s_4ns_4_2_1_Adder_4_U.fas_s2  = \add_4s_4ns_4_2_1_U6.top_add_4s_4ns_4_2_1_Adder_4_U.u2.s ;
assign \add_4s_4ns_4_2_1_U6.top_add_4s_4ns_4_2_1_Adder_4_U.u1.a  = \add_4s_4ns_4_2_1_U6.top_add_4s_4ns_4_2_1_Adder_4_U.a [1:0];
assign \add_4s_4ns_4_2_1_U6.top_add_4s_4ns_4_2_1_Adder_4_U.u1.b  = \add_4s_4ns_4_2_1_U6.top_add_4s_4ns_4_2_1_Adder_4_U.b [1:0];
assign \add_4s_4ns_4_2_1_U6.top_add_4s_4ns_4_2_1_Adder_4_U.u1.cin  = 1'h0;
assign \add_4s_4ns_4_2_1_U6.top_add_4s_4ns_4_2_1_Adder_4_U.facout_s1  = \add_4s_4ns_4_2_1_U6.top_add_4s_4ns_4_2_1_Adder_4_U.u1.cout ;
assign \add_4s_4ns_4_2_1_U6.top_add_4s_4ns_4_2_1_Adder_4_U.fas_s1  = \add_4s_4ns_4_2_1_U6.top_add_4s_4ns_4_2_1_Adder_4_U.u1.s ;
assign \add_4s_4ns_4_2_1_U6.top_add_4s_4ns_4_2_1_Adder_4_U.a  = \add_4s_4ns_4_2_1_U6.din0 ;
assign \add_4s_4ns_4_2_1_U6.top_add_4s_4ns_4_2_1_Adder_4_U.b  = \add_4s_4ns_4_2_1_U6.din1 ;
assign \add_4s_4ns_4_2_1_U6.top_add_4s_4ns_4_2_1_Adder_4_U.ce  = \add_4s_4ns_4_2_1_U6.ce ;
assign \add_4s_4ns_4_2_1_U6.top_add_4s_4ns_4_2_1_Adder_4_U.clk  = \add_4s_4ns_4_2_1_U6.clk ;
assign \add_4s_4ns_4_2_1_U6.top_add_4s_4ns_4_2_1_Adder_4_U.reset  = \add_4s_4ns_4_2_1_U6.reset ;
assign \add_4s_4ns_4_2_1_U6.dout  = \add_4s_4ns_4_2_1_U6.top_add_4s_4ns_4_2_1_Adder_4_U.s ;
assign \add_4s_4ns_4_2_1_U6.ce  = 1'h1;
assign \add_4s_4ns_4_2_1_U6.clk  = ap_clk;
assign \add_4s_4ns_4_2_1_U6.din0  = { tmp_2_reg_1448[2], tmp_2_reg_1448 };
assign \add_4s_4ns_4_2_1_U6.din1  = 4'h1;
assign grp_fu_757_p2 = \add_4s_4ns_4_2_1_U6.dout ;
assign \add_4s_4ns_4_2_1_U6.reset  = ap_rst;
assign \add_47s_47s_47_2_1_U20.top_add_47s_47s_47_2_1_Adder_12_U.ain_s0  = \add_47s_47s_47_2_1_U20.top_add_47s_47s_47_2_1_Adder_12_U.a ;
assign \add_47s_47s_47_2_1_U20.top_add_47s_47s_47_2_1_Adder_12_U.bin_s0  = \add_47s_47s_47_2_1_U20.top_add_47s_47s_47_2_1_Adder_12_U.b ;
assign \add_47s_47s_47_2_1_U20.top_add_47s_47s_47_2_1_Adder_12_U.s  = { \add_47s_47s_47_2_1_U20.top_add_47s_47s_47_2_1_Adder_12_U.fas_s2 , \add_47s_47s_47_2_1_U20.top_add_47s_47s_47_2_1_Adder_12_U.sum_s1  };
assign \add_47s_47s_47_2_1_U20.top_add_47s_47s_47_2_1_Adder_12_U.u2.a  = \add_47s_47s_47_2_1_U20.top_add_47s_47s_47_2_1_Adder_12_U.ain_s1 ;
assign \add_47s_47s_47_2_1_U20.top_add_47s_47s_47_2_1_Adder_12_U.u2.b  = \add_47s_47s_47_2_1_U20.top_add_47s_47s_47_2_1_Adder_12_U.bin_s1 ;
assign \add_47s_47s_47_2_1_U20.top_add_47s_47s_47_2_1_Adder_12_U.u2.cin  = \add_47s_47s_47_2_1_U20.top_add_47s_47s_47_2_1_Adder_12_U.carry_s1 ;
assign \add_47s_47s_47_2_1_U20.top_add_47s_47s_47_2_1_Adder_12_U.facout_s2  = \add_47s_47s_47_2_1_U20.top_add_47s_47s_47_2_1_Adder_12_U.u2.cout ;
assign \add_47s_47s_47_2_1_U20.top_add_47s_47s_47_2_1_Adder_12_U.fas_s2  = \add_47s_47s_47_2_1_U20.top_add_47s_47s_47_2_1_Adder_12_U.u2.s ;
assign \add_47s_47s_47_2_1_U20.top_add_47s_47s_47_2_1_Adder_12_U.u1.a  = \add_47s_47s_47_2_1_U20.top_add_47s_47s_47_2_1_Adder_12_U.a [22:0];
assign \add_47s_47s_47_2_1_U20.top_add_47s_47s_47_2_1_Adder_12_U.u1.b  = \add_47s_47s_47_2_1_U20.top_add_47s_47s_47_2_1_Adder_12_U.b [22:0];
assign \add_47s_47s_47_2_1_U20.top_add_47s_47s_47_2_1_Adder_12_U.u1.cin  = 1'h0;
assign \add_47s_47s_47_2_1_U20.top_add_47s_47s_47_2_1_Adder_12_U.facout_s1  = \add_47s_47s_47_2_1_U20.top_add_47s_47s_47_2_1_Adder_12_U.u1.cout ;
assign \add_47s_47s_47_2_1_U20.top_add_47s_47s_47_2_1_Adder_12_U.fas_s1  = \add_47s_47s_47_2_1_U20.top_add_47s_47s_47_2_1_Adder_12_U.u1.s ;
assign \add_47s_47s_47_2_1_U20.top_add_47s_47s_47_2_1_Adder_12_U.a  = \add_47s_47s_47_2_1_U20.din0 ;
assign \add_47s_47s_47_2_1_U20.top_add_47s_47s_47_2_1_Adder_12_U.b  = \add_47s_47s_47_2_1_U20.din1 ;
assign \add_47s_47s_47_2_1_U20.top_add_47s_47s_47_2_1_Adder_12_U.ce  = \add_47s_47s_47_2_1_U20.ce ;
assign \add_47s_47s_47_2_1_U20.top_add_47s_47s_47_2_1_Adder_12_U.clk  = \add_47s_47s_47_2_1_U20.clk ;
assign \add_47s_47s_47_2_1_U20.top_add_47s_47s_47_2_1_Adder_12_U.reset  = \add_47s_47s_47_2_1_U20.reset ;
assign \add_47s_47s_47_2_1_U20.dout  = \add_47s_47s_47_2_1_U20.top_add_47s_47s_47_2_1_Adder_12_U.s ;
assign \add_47s_47s_47_2_1_U20.ce  = 1'h1;
assign \add_47s_47s_47_2_1_U20.clk  = ap_clk;
assign \add_47s_47s_47_2_1_U20.din0  = { select_ln353_reg_1696[31], select_ln353_reg_1696, 14'h0000 };
assign \add_47s_47s_47_2_1_U20.din1  = { op_19[15], op_19[15], op_19[15], op_19[15], op_19[15], op_19[15], op_19[15], op_19[15], op_19[15], op_19[15], op_19[15], op_19[15], op_19[15], op_19[15], op_19[15], op_19[15], op_19[15], op_19[15], op_19[15], op_19[15], op_19[15], op_19[15], op_19[15], op_19[15], op_19[15], op_19[15], op_19[15], op_19[15], op_19[15], op_19[15], op_19[15], op_19 };
assign grp_fu_1094_p2 = \add_47s_47s_47_2_1_U20.dout ;
assign \add_47s_47s_47_2_1_U20.reset  = ap_rst;
assign \add_33ns_33ns_33_2_1_U10.top_add_33ns_33ns_33_2_1_Adder_7_U.ain_s0  = \add_33ns_33ns_33_2_1_U10.top_add_33ns_33ns_33_2_1_Adder_7_U.a ;
assign \add_33ns_33ns_33_2_1_U10.top_add_33ns_33ns_33_2_1_Adder_7_U.bin_s0  = \add_33ns_33ns_33_2_1_U10.top_add_33ns_33ns_33_2_1_Adder_7_U.b ;
assign \add_33ns_33ns_33_2_1_U10.top_add_33ns_33ns_33_2_1_Adder_7_U.s  = { \add_33ns_33ns_33_2_1_U10.top_add_33ns_33ns_33_2_1_Adder_7_U.fas_s2 , \add_33ns_33ns_33_2_1_U10.top_add_33ns_33ns_33_2_1_Adder_7_U.sum_s1  };
assign \add_33ns_33ns_33_2_1_U10.top_add_33ns_33ns_33_2_1_Adder_7_U.u2.a  = \add_33ns_33ns_33_2_1_U10.top_add_33ns_33ns_33_2_1_Adder_7_U.ain_s1 ;
assign \add_33ns_33ns_33_2_1_U10.top_add_33ns_33ns_33_2_1_Adder_7_U.u2.b  = \add_33ns_33ns_33_2_1_U10.top_add_33ns_33ns_33_2_1_Adder_7_U.bin_s1 ;
assign \add_33ns_33ns_33_2_1_U10.top_add_33ns_33ns_33_2_1_Adder_7_U.u2.cin  = \add_33ns_33ns_33_2_1_U10.top_add_33ns_33ns_33_2_1_Adder_7_U.carry_s1 ;
assign \add_33ns_33ns_33_2_1_U10.top_add_33ns_33ns_33_2_1_Adder_7_U.facout_s2  = \add_33ns_33ns_33_2_1_U10.top_add_33ns_33ns_33_2_1_Adder_7_U.u2.cout ;
assign \add_33ns_33ns_33_2_1_U10.top_add_33ns_33ns_33_2_1_Adder_7_U.fas_s2  = \add_33ns_33ns_33_2_1_U10.top_add_33ns_33ns_33_2_1_Adder_7_U.u2.s ;
assign \add_33ns_33ns_33_2_1_U10.top_add_33ns_33ns_33_2_1_Adder_7_U.u1.a  = \add_33ns_33ns_33_2_1_U10.top_add_33ns_33ns_33_2_1_Adder_7_U.a [15:0];
assign \add_33ns_33ns_33_2_1_U10.top_add_33ns_33ns_33_2_1_Adder_7_U.u1.b  = \add_33ns_33ns_33_2_1_U10.top_add_33ns_33ns_33_2_1_Adder_7_U.b [15:0];
assign \add_33ns_33ns_33_2_1_U10.top_add_33ns_33ns_33_2_1_Adder_7_U.u1.cin  = 1'h0;
assign \add_33ns_33ns_33_2_1_U10.top_add_33ns_33ns_33_2_1_Adder_7_U.facout_s1  = \add_33ns_33ns_33_2_1_U10.top_add_33ns_33ns_33_2_1_Adder_7_U.u1.cout ;
assign \add_33ns_33ns_33_2_1_U10.top_add_33ns_33ns_33_2_1_Adder_7_U.fas_s1  = \add_33ns_33ns_33_2_1_U10.top_add_33ns_33ns_33_2_1_Adder_7_U.u1.s ;
assign \add_33ns_33ns_33_2_1_U10.top_add_33ns_33ns_33_2_1_Adder_7_U.a  = \add_33ns_33ns_33_2_1_U10.din0 ;
assign \add_33ns_33ns_33_2_1_U10.top_add_33ns_33ns_33_2_1_Adder_7_U.b  = \add_33ns_33ns_33_2_1_U10.din1 ;
assign \add_33ns_33ns_33_2_1_U10.top_add_33ns_33ns_33_2_1_Adder_7_U.ce  = \add_33ns_33ns_33_2_1_U10.ce ;
assign \add_33ns_33ns_33_2_1_U10.top_add_33ns_33ns_33_2_1_Adder_7_U.clk  = \add_33ns_33ns_33_2_1_U10.clk ;
assign \add_33ns_33ns_33_2_1_U10.top_add_33ns_33ns_33_2_1_Adder_7_U.reset  = \add_33ns_33ns_33_2_1_U10.reset ;
assign \add_33ns_33ns_33_2_1_U10.dout  = \add_33ns_33ns_33_2_1_U10.top_add_33ns_33ns_33_2_1_Adder_7_U.s ;
assign \add_33ns_33ns_33_2_1_U10.ce  = 1'h1;
assign \add_33ns_33ns_33_2_1_U10.clk  = ap_clk;
assign \add_33ns_33ns_33_2_1_U10.din0  = { 1'h0, op_9 };
assign \add_33ns_33ns_33_2_1_U10.din1  = { 17'h00000, sext_ln1118_reg_1433 };
assign grp_fu_842_p2 = \add_33ns_33ns_33_2_1_U10.dout ;
assign \add_33ns_33ns_33_2_1_U10.reset  = ap_rst;
assign \add_32s_32ns_32_2_1_U15.top_add_32s_32ns_32_2_1_Adder_10_U.ain_s0  = \add_32s_32ns_32_2_1_U15.top_add_32s_32ns_32_2_1_Adder_10_U.a ;
assign \add_32s_32ns_32_2_1_U15.top_add_32s_32ns_32_2_1_Adder_10_U.bin_s0  = \add_32s_32ns_32_2_1_U15.top_add_32s_32ns_32_2_1_Adder_10_U.b ;
assign \add_32s_32ns_32_2_1_U15.top_add_32s_32ns_32_2_1_Adder_10_U.s  = { \add_32s_32ns_32_2_1_U15.top_add_32s_32ns_32_2_1_Adder_10_U.fas_s2 , \add_32s_32ns_32_2_1_U15.top_add_32s_32ns_32_2_1_Adder_10_U.sum_s1  };
assign \add_32s_32ns_32_2_1_U15.top_add_32s_32ns_32_2_1_Adder_10_U.u2.a  = \add_32s_32ns_32_2_1_U15.top_add_32s_32ns_32_2_1_Adder_10_U.ain_s1 ;
assign \add_32s_32ns_32_2_1_U15.top_add_32s_32ns_32_2_1_Adder_10_U.u2.b  = \add_32s_32ns_32_2_1_U15.top_add_32s_32ns_32_2_1_Adder_10_U.bin_s1 ;
assign \add_32s_32ns_32_2_1_U15.top_add_32s_32ns_32_2_1_Adder_10_U.u2.cin  = \add_32s_32ns_32_2_1_U15.top_add_32s_32ns_32_2_1_Adder_10_U.carry_s1 ;
assign \add_32s_32ns_32_2_1_U15.top_add_32s_32ns_32_2_1_Adder_10_U.facout_s2  = \add_32s_32ns_32_2_1_U15.top_add_32s_32ns_32_2_1_Adder_10_U.u2.cout ;
assign \add_32s_32ns_32_2_1_U15.top_add_32s_32ns_32_2_1_Adder_10_U.fas_s2  = \add_32s_32ns_32_2_1_U15.top_add_32s_32ns_32_2_1_Adder_10_U.u2.s ;
assign \add_32s_32ns_32_2_1_U15.top_add_32s_32ns_32_2_1_Adder_10_U.u1.a  = \add_32s_32ns_32_2_1_U15.top_add_32s_32ns_32_2_1_Adder_10_U.a [15:0];
assign \add_32s_32ns_32_2_1_U15.top_add_32s_32ns_32_2_1_Adder_10_U.u1.b  = \add_32s_32ns_32_2_1_U15.top_add_32s_32ns_32_2_1_Adder_10_U.b [15:0];
assign \add_32s_32ns_32_2_1_U15.top_add_32s_32ns_32_2_1_Adder_10_U.u1.cin  = 1'h0;
assign \add_32s_32ns_32_2_1_U15.top_add_32s_32ns_32_2_1_Adder_10_U.facout_s1  = \add_32s_32ns_32_2_1_U15.top_add_32s_32ns_32_2_1_Adder_10_U.u1.cout ;
assign \add_32s_32ns_32_2_1_U15.top_add_32s_32ns_32_2_1_Adder_10_U.fas_s1  = \add_32s_32ns_32_2_1_U15.top_add_32s_32ns_32_2_1_Adder_10_U.u1.s ;
assign \add_32s_32ns_32_2_1_U15.top_add_32s_32ns_32_2_1_Adder_10_U.a  = \add_32s_32ns_32_2_1_U15.din0 ;
assign \add_32s_32ns_32_2_1_U15.top_add_32s_32ns_32_2_1_Adder_10_U.b  = \add_32s_32ns_32_2_1_U15.din1 ;
assign \add_32s_32ns_32_2_1_U15.top_add_32s_32ns_32_2_1_Adder_10_U.ce  = \add_32s_32ns_32_2_1_U15.ce ;
assign \add_32s_32ns_32_2_1_U15.top_add_32s_32ns_32_2_1_Adder_10_U.clk  = \add_32s_32ns_32_2_1_U15.clk ;
assign \add_32s_32ns_32_2_1_U15.top_add_32s_32ns_32_2_1_Adder_10_U.reset  = \add_32s_32ns_32_2_1_U15.reset ;
assign \add_32s_32ns_32_2_1_U15.dout  = \add_32s_32ns_32_2_1_U15.top_add_32s_32ns_32_2_1_Adder_10_U.s ;
assign \add_32s_32ns_32_2_1_U15.ce  = 1'h1;
assign \add_32s_32ns_32_2_1_U15.clk  = ap_clk;
assign \add_32s_32ns_32_2_1_U15.din0  = { add_ln69_1_reg_1614[4], add_ln69_1_reg_1614[4], add_ln69_1_reg_1614[4], add_ln69_1_reg_1614[4], add_ln69_1_reg_1614[4], add_ln69_1_reg_1614[4], add_ln69_1_reg_1614[4], add_ln69_1_reg_1614[4], add_ln69_1_reg_1614[4], add_ln69_1_reg_1614[4], add_ln69_1_reg_1614[4], add_ln69_1_reg_1614[4], add_ln69_1_reg_1614[4], add_ln69_1_reg_1614[4], add_ln69_1_reg_1614[4], add_ln69_1_reg_1614[4], add_ln69_1_reg_1614[4], add_ln69_1_reg_1614[4], add_ln69_1_reg_1614[4], add_ln69_1_reg_1614[4], add_ln69_1_reg_1614[4], add_ln69_1_reg_1614[4], add_ln69_1_reg_1614[4], add_ln69_1_reg_1614[4], add_ln69_1_reg_1614[4], add_ln69_1_reg_1614[4], add_ln69_1_reg_1614[4], add_ln69_1_reg_1614 };
assign \add_32s_32ns_32_2_1_U15.din1  = add_ln69_reg_1609;
assign grp_fu_965_p2 = \add_32s_32ns_32_2_1_U15.dout ;
assign \add_32s_32ns_32_2_1_U15.reset  = ap_rst;
assign \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s0  = \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.a ;
assign \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s0  = \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.b ;
assign \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.s  = { \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s2 , \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.sum_s1  };
assign \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.a  = \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s1 ;
assign \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.b  = \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s1 ;
assign \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cin  = \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.carry_s1 ;
assign \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s2  = \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cout ;
assign \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s2  = \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.s ;
assign \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.a  = \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.a [15:0];
assign \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.b  = \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.b [15:0];
assign \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cin  = 1'h0;
assign \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s1  = \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cout ;
assign \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s1  = \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.s ;
assign \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.a  = \add_32ns_32ns_32_2_1_U9.din0 ;
assign \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.b  = \add_32ns_32ns_32_2_1_U9.din1 ;
assign \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  = \add_32ns_32ns_32_2_1_U9.ce ;
assign \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.clk  = \add_32ns_32ns_32_2_1_U9.clk ;
assign \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.reset  = \add_32ns_32ns_32_2_1_U9.reset ;
assign \add_32ns_32ns_32_2_1_U9.dout  = \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_6_U.s ;
assign \add_32ns_32ns_32_2_1_U9.ce  = 1'h1;
assign \add_32ns_32ns_32_2_1_U9.clk  = ap_clk;
assign \add_32ns_32ns_32_2_1_U9.din0  = select_ln1192_reg_1512;
assign \add_32ns_32ns_32_2_1_U9.din1  = op_9;
assign grp_fu_830_p2 = \add_32ns_32ns_32_2_1_U9.dout ;
assign \add_32ns_32ns_32_2_1_U9.reset  = ap_rst;
assign \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s0  = \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.a ;
assign \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s0  = \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.b ;
assign \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.s  = { \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s2 , \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.sum_s1  };
assign \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.a  = \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s1 ;
assign \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.b  = \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s1 ;
assign \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cin  = \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.carry_s1 ;
assign \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s2  = \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cout ;
assign \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s2  = \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.s ;
assign \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.a  = \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.a [15:0];
assign \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.b  = \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.b [15:0];
assign \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cin  = 1'h0;
assign \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s1  = \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cout ;
assign \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s1  = \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.s ;
assign \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.a  = \add_32ns_32ns_32_2_1_U8.din0 ;
assign \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.b  = \add_32ns_32ns_32_2_1_U8.din1 ;
assign \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  = \add_32ns_32ns_32_2_1_U8.ce ;
assign \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.clk  = \add_32ns_32ns_32_2_1_U8.clk ;
assign \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.reset  = \add_32ns_32ns_32_2_1_U8.reset ;
assign \add_32ns_32ns_32_2_1_U8.dout  = \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_6_U.s ;
assign \add_32ns_32ns_32_2_1_U8.ce  = 1'h1;
assign \add_32ns_32ns_32_2_1_U8.clk  = ap_clk;
assign \add_32ns_32ns_32_2_1_U8.din0  = ret_V_7_cast_reg_1505;
assign \add_32ns_32ns_32_2_1_U8.din1  = 32'd1;
assign grp_fu_825_p2 = \add_32ns_32ns_32_2_1_U8.dout ;
assign \add_32ns_32ns_32_2_1_U8.reset  = ap_rst;
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s0  = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_6_U.a ;
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s0  = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_6_U.b ;
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_6_U.s  = { \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s2 , \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_6_U.sum_s1  };
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.a  = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s1 ;
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.b  = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s1 ;
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cin  = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_6_U.carry_s1 ;
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s2  = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cout ;
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s2  = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.s ;
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.a  = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_6_U.a [15:0];
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.b  = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_6_U.b [15:0];
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cin  = 1'h0;
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s1  = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cout ;
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s1  = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.s ;
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_6_U.a  = \add_32ns_32ns_32_2_1_U21.din0 ;
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_6_U.b  = \add_32ns_32ns_32_2_1_U21.din1 ;
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  = \add_32ns_32ns_32_2_1_U21.ce ;
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_6_U.clk  = \add_32ns_32ns_32_2_1_U21.clk ;
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_6_U.reset  = \add_32ns_32ns_32_2_1_U21.reset ;
assign \add_32ns_32ns_32_2_1_U21.dout  = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_6_U.s ;
assign \add_32ns_32ns_32_2_1_U21.ce  = 1'h1;
assign \add_32ns_32ns_32_2_1_U21.clk  = ap_clk;
assign \add_32ns_32ns_32_2_1_U21.din0  = ret_V_20_cast_reg_1721;
assign \add_32ns_32ns_32_2_1_U21.din1  = 32'd1;
assign grp_fu_1120_p2 = \add_32ns_32ns_32_2_1_U21.dout ;
assign \add_32ns_32ns_32_2_1_U21.reset  = ap_rst;
assign \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s0  = \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_6_U.a ;
assign \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s0  = \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_6_U.b ;
assign \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_6_U.s  = { \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s2 , \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_6_U.sum_s1  };
assign \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.a  = \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s1 ;
assign \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.b  = \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s1 ;
assign \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cin  = \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_6_U.carry_s1 ;
assign \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s2  = \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cout ;
assign \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s2  = \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.s ;
assign \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.a  = \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_6_U.a [15:0];
assign \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.b  = \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_6_U.b [15:0];
assign \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cin  = 1'h0;
assign \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s1  = \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cout ;
assign \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s1  = \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.s ;
assign \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_6_U.a  = \add_32ns_32ns_32_2_1_U19.din0 ;
assign \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_6_U.b  = \add_32ns_32ns_32_2_1_U19.din1 ;
assign \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  = \add_32ns_32ns_32_2_1_U19.ce ;
assign \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_6_U.clk  = \add_32ns_32ns_32_2_1_U19.clk ;
assign \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_6_U.reset  = \add_32ns_32ns_32_2_1_U19.reset ;
assign \add_32ns_32ns_32_2_1_U19.dout  = \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_6_U.s ;
assign \add_32ns_32ns_32_2_1_U19.ce  = 1'h1;
assign \add_32ns_32ns_32_2_1_U19.clk  = ap_clk;
assign \add_32ns_32ns_32_2_1_U19.din0  = ret_V_18_cast_reg_1684;
assign \add_32ns_32ns_32_2_1_U19.din1  = 32'd1;
assign grp_fu_1055_p2 = \add_32ns_32ns_32_2_1_U19.dout ;
assign \add_32ns_32ns_32_2_1_U19.reset  = ap_rst;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s0  = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.a ;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s0  = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.b ;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.s  = { \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s2 , \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.sum_s1  };
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.a  = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s1 ;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.b  = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s1 ;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cin  = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.carry_s1 ;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s2  = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cout ;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s2  = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.s ;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.a  = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.a [15:0];
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.b  = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.b [15:0];
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cin  = 1'h0;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s1  = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cout ;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s1  = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.s ;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.a  = \add_32ns_32ns_32_2_1_U17.din0 ;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.b  = \add_32ns_32ns_32_2_1_U17.din1 ;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  = \add_32ns_32ns_32_2_1_U17.ce ;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.clk  = \add_32ns_32ns_32_2_1_U17.clk ;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.reset  = \add_32ns_32ns_32_2_1_U17.reset ;
assign \add_32ns_32ns_32_2_1_U17.dout  = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.s ;
assign \add_32ns_32ns_32_2_1_U17.ce  = 1'h1;
assign \add_32ns_32ns_32_2_1_U17.clk  = ap_clk;
assign \add_32ns_32ns_32_2_1_U17.din0  = ret_V_17_reg_1639;
assign \add_32ns_32ns_32_2_1_U17.din1  = { 31'h00000000, lhs_V_3_reg_1278 };
assign grp_fu_984_p2 = \add_32ns_32ns_32_2_1_U17.dout ;
assign \add_32ns_32ns_32_2_1_U17.reset  = ap_rst;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s0  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.a ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s0  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.b ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.s  = { \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s2 , \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.sum_s1  };
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.a  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s1 ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.b  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s1 ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cin  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.carry_s1 ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s2  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cout ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s2  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.s ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.a  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.a [15:0];
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.b  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.b [15:0];
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cin  = 1'h0;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s1  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cout ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s1  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.s ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.a  = \add_32ns_32ns_32_2_1_U16.din0 ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.b  = \add_32ns_32ns_32_2_1_U16.din1 ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  = \add_32ns_32ns_32_2_1_U16.ce ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.clk  = \add_32ns_32ns_32_2_1_U16.clk ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.reset  = \add_32ns_32ns_32_2_1_U16.reset ;
assign \add_32ns_32ns_32_2_1_U16.dout  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_6_U.s ;
assign \add_32ns_32ns_32_2_1_U16.ce  = 1'h1;
assign \add_32ns_32ns_32_2_1_U16.clk  = ap_clk;
assign \add_32ns_32ns_32_2_1_U16.din0  = op_23_V_reg_1629;
assign \add_32ns_32ns_32_2_1_U16.din1  = select_ln1192_1_reg_1634;
assign grp_fu_977_p2 = \add_32ns_32ns_32_2_1_U16.dout ;
assign \add_32ns_32ns_32_2_1_U16.reset  = ap_rst;
assign \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s0  = \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.a ;
assign \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s0  = \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.b ;
assign \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.s  = { \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s2 , \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.sum_s1  };
assign \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.a  = \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s1 ;
assign \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.b  = \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s1 ;
assign \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cin  = \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.carry_s1 ;
assign \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s2  = \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cout ;
assign \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s2  = \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.s ;
assign \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.a  = \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.a [15:0];
assign \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.b  = \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.b [15:0];
assign \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cin  = 1'h0;
assign \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s1  = \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cout ;
assign \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s1  = \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.s ;
assign \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.a  = \add_32ns_32ns_32_2_1_U13.din0 ;
assign \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.b  = \add_32ns_32ns_32_2_1_U13.din1 ;
assign \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  = \add_32ns_32ns_32_2_1_U13.ce ;
assign \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.clk  = \add_32ns_32ns_32_2_1_U13.clk ;
assign \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.reset  = \add_32ns_32ns_32_2_1_U13.reset ;
assign \add_32ns_32ns_32_2_1_U13.dout  = \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_6_U.s ;
assign \add_32ns_32ns_32_2_1_U13.ce  = 1'h1;
assign \add_32ns_32ns_32_2_1_U13.clk  = ap_clk;
assign \add_32ns_32ns_32_2_1_U13.din0  = ret_V_12_reg_1557;
assign \add_32ns_32ns_32_2_1_U13.din1  = ret_V_16_reg_1578;
assign grp_fu_910_p2 = \add_32ns_32ns_32_2_1_U13.dout ;
assign \add_32ns_32ns_32_2_1_U13.reset  = ap_rst;
assign \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_2_U.ain_s0  = \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_2_U.a ;
assign \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_2_U.bin_s0  = \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_2_U.b ;
assign \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_2_U.s  = { \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_2_U.fas_s2 , \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_2_U.sum_s1  };
assign \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_2_U.u2.a  = \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_2_U.ain_s1 ;
assign \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_2_U.u2.b  = \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_2_U.bin_s1 ;
assign \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_2_U.u2.cin  = \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_2_U.carry_s1 ;
assign \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_2_U.facout_s2  = \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_2_U.u2.cout ;
assign \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_2_U.fas_s2  = \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_2_U.u2.s ;
assign \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_2_U.u1.a  = \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_2_U.a [0];
assign \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_2_U.u1.b  = \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_2_U.b [0];
assign \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_2_U.u1.cin  = 1'h0;
assign \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_2_U.facout_s1  = \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_2_U.u1.cout ;
assign \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_2_U.fas_s1  = \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_2_U.u1.s ;
assign \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_2_U.a  = \add_2ns_2ns_2_2_1_U3.din0 ;
assign \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_2_U.b  = \add_2ns_2ns_2_2_1_U3.din1 ;
assign \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_2_U.ce  = \add_2ns_2ns_2_2_1_U3.ce ;
assign \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_2_U.clk  = \add_2ns_2ns_2_2_1_U3.clk ;
assign \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_2_U.reset  = \add_2ns_2ns_2_2_1_U3.reset ;
assign \add_2ns_2ns_2_2_1_U3.dout  = \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_2_U.s ;
assign \add_2ns_2ns_2_2_1_U3.ce  = 1'h1;
assign \add_2ns_2ns_2_2_1_U3.clk  = ap_clk;
assign \add_2ns_2ns_2_2_1_U3.din0  = trunc_ln731_2_reg_1321;
assign \add_2ns_2ns_2_2_1_U3.din1  = { 1'h0, lhs_V_3_reg_1278 };
assign grp_fu_536_p2 = \add_2ns_2ns_2_2_1_U3.dout ;
assign \add_2ns_2ns_2_2_1_U3.reset  = ap_rst;
assign \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_8_U.ain_s0  = \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_8_U.a ;
assign \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_8_U.bin_s0  = \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_8_U.b ;
assign \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_8_U.s  = { \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_8_U.fas_s2 , \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_8_U.sum_s1  };
assign \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_8_U.u2.a  = \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_8_U.ain_s1 ;
assign \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_8_U.u2.b  = \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_8_U.bin_s1 ;
assign \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_8_U.u2.cin  = \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_8_U.carry_s1 ;
assign \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_8_U.facout_s2  = \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_8_U.u2.cout ;
assign \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_8_U.fas_s2  = \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_8_U.u2.s ;
assign \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_8_U.u1.a  = \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_8_U.a [4:0];
assign \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_8_U.u1.b  = \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_8_U.b [4:0];
assign \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_8_U.u1.cin  = 1'h0;
assign \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_8_U.facout_s1  = \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_8_U.u1.cout ;
assign \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_8_U.fas_s1  = \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_8_U.u1.s ;
assign \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_8_U.a  = \add_11ns_11s_11_2_1_U11.din0 ;
assign \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_8_U.b  = \add_11ns_11s_11_2_1_U11.din1 ;
assign \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_8_U.ce  = \add_11ns_11s_11_2_1_U11.ce ;
assign \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_8_U.clk  = \add_11ns_11s_11_2_1_U11.clk ;
assign \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_8_U.reset  = \add_11ns_11s_11_2_1_U11.reset ;
assign \add_11ns_11s_11_2_1_U11.dout  = \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_8_U.s ;
assign \add_11ns_11s_11_2_1_U11.ce  = 1'h1;
assign \add_11ns_11s_11_2_1_U11.clk  = ap_clk;
assign \add_11ns_11s_11_2_1_U11.din0  = op_9[10:0];
assign \add_11ns_11s_11_2_1_U11.din1  = { ret_V_11_reg_1402[3], ret_V_11_reg_1402[3], ret_V_11_reg_1402[3], ret_V_11_reg_1402[3], ret_V_11_reg_1402[3], ret_V_11_reg_1402[3], ret_V_11_reg_1402[3], ret_V_11_reg_1402 };
assign grp_fu_855_p2 = \add_11ns_11s_11_2_1_U11.dout ;
assign \add_11ns_11s_11_2_1_U11.reset  = ap_rst;
endmodule


// Product machine:
module top_A_times_top_B (ap_start, op_0, op_1, op_19, op_7, op_8, op_9, ap_clk, unsafe_signal);
input ap_start;
input [3:0] op_0;
input [3:0] op_1;
input [15:0] op_19;
input [31:0] op_7;
input [3:0] op_8;
input [31:0] op_9;
input ap_clk;
output unsafe_signal;
reg _setup;
initial _setup = 1'b0;
always @ (posedge ap_clk) _setup <= 1'b1;
reg ap_start_internal;
always @ (posedge ap_clk) if (!_setup) ap_start_internal <= ap_start;
reg [3:0] op_0_internal;
always @ (posedge ap_clk) if (!_setup) op_0_internal <= op_0;
reg [3:0] op_1_internal;
always @ (posedge ap_clk) if (!_setup) op_1_internal <= op_1;
reg [15:0] op_19_internal;
always @ (posedge ap_clk) if (!_setup) op_19_internal <= op_19;
reg [31:0] op_7_internal;
always @ (posedge ap_clk) if (!_setup) op_7_internal <= op_7;
reg [3:0] op_8_internal;
always @ (posedge ap_clk) if (!_setup) op_8_internal <= op_8;
reg [31:0] op_9_internal;
always @ (posedge ap_clk) if (!_setup) op_9_internal <= op_9;
wire ap_done_A;
wire ap_done_B;
wire ap_done_eq;
assign ap_done_eq = ap_done_A == ap_done_B;
wire ap_idle_A;
wire ap_idle_B;
wire ap_idle_eq;
assign ap_idle_eq = ap_idle_A == ap_idle_B;
wire ap_ready_A;
wire ap_ready_B;
wire ap_ready_eq;
assign ap_ready_eq = ap_ready_A == ap_ready_B;
wire [31:0] op_27_A;
wire [31:0] op_27_B;
wire op_27_eq;
assign op_27_eq = op_27_A == op_27_B;
wire op_27_ap_vld_A;
wire op_27_ap_vld_B;
wire clk_enable_A;
wire clk_enable_B;
assign clk_enable_A = _setup & (~op_27_ap_vld_A | op_27_ap_vld_B);
assign clk_enable_B = _setup;
wire divergent;
assign divergent = ~(ap_done_eq & ap_idle_eq & ap_ready_eq & op_27_eq);
assign unsafe_signal = op_27_ap_vld_A & op_27_ap_vld_B & divergent;
top_A instance_A (
    .ap_clk(ap_clk),
    .clk_enable(clk_enable_A),
    .ap_start(ap_start_internal),
    .op_0(op_0_internal),
    .op_1(op_1_internal),
    .op_19(op_19_internal),
    .op_7(op_7_internal),
    .op_8(op_8_internal),
    .op_9(op_9_internal),
    .ap_done(ap_done_A),
    .ap_idle(ap_idle_A),
    .ap_ready(ap_ready_A),
    .op_27(op_27_A),
    .op_27_ap_vld(op_27_ap_vld_A)
);
top_B instance_B (
    .ap_clk(ap_clk),
    .clk_enable(clk_enable_B),
    .ap_start(ap_start_internal),
    .op_0(op_0_internal),
    .op_1(op_1_internal),
    .op_19(op_19_internal),
    .op_7(op_7_internal),
    .op_8(op_8_internal),
    .op_9(op_9_internal),
    .ap_done(ap_done_B),
    .ap_idle(ap_idle_B),
    .ap_ready(ap_ready_B),
    .op_27(op_27_B),
    .op_27_ap_vld(op_27_ap_vld_B)
);
endmodule
