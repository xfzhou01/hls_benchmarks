// Processed by function `construct_kairos` in `verilog_tricks.py`.
// Machine A:
// Processed by function `add_clk_enable_signal` in `verilog_tricks.py`.
// Processed by function `remove_reset_signal` in `verilog_tricks.py`.
module top_A (
  ap_clk,
  ap_start,
  ap_done,
  ap_idle,
  ap_ready,
  op_0,
  op_2,
  op_3,
  op_4,
  op_5,
  op_7,
  op_8,
  op_9,
  op_10,
  op_11,
  op_17,
  op_18,
  op_19,
  op_31,
  op_31_ap_vld,
clk_enable
);
input clk_enable;


input ap_clk;
wire ap_rst;
assign ap_rst = op_31_ap_vld;
input ap_start;
input [1:0] op_0;
input [31:0] op_10;
input [1:0] op_11;
input [3:0] op_17;
input [7:0] op_18;
input [7:0] op_19;
input [1:0] op_2;
input [3:0] op_3;
input [7:0] op_4;
input [3:0] op_5;
input op_7;
input [15:0] op_8;
input [3:0] op_9;
output ap_done;
output ap_idle;
output ap_ready;
output [31:0] op_31;
output op_31_ap_vld;


reg [11:0] \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.ain_s1 ;
reg [11:0] \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.bin_s1 ;
reg \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.carry_s1 ;
reg [10:0] \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.sum_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.ain_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.bin_s1 ;
reg \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.carry_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.sum_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.ain_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.bin_s1 ;
reg \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.carry_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.sum_s1 ;
reg [15:0] \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.ain_s1 ;
reg [15:0] \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.bin_s1 ;
reg \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.carry_s1 ;
reg [15:0] \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.sum_s1 ;
reg [15:0] \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.ain_s1 ;
reg [15:0] \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.bin_s1 ;
reg \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.carry_s1 ;
reg [15:0] \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.sum_s1 ;
reg [15:0] \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.ain_s1 ;
reg [15:0] \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.bin_s1 ;
reg \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.carry_s1 ;
reg [15:0] \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.sum_s1 ;
reg [16:0] \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.ain_s1 ;
reg [16:0] \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.bin_s1 ;
reg \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.carry_s1 ;
reg [15:0] \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.sum_s1 ;
reg [16:0] \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.ain_s1 ;
reg [16:0] \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.bin_s1 ;
reg \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.carry_s1 ;
reg [15:0] \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.sum_s1 ;
reg [16:0] \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.ain_s1 ;
reg [16:0] \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.bin_s1 ;
reg \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.carry_s1 ;
reg [16:0] \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.sum_s1 ;
reg [17:0] \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.ain_s1 ;
reg [17:0] \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.bin_s1 ;
reg \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.carry_s1 ;
reg [17:0] \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.sum_s1 ;
reg [31:0] add_ln691_1_reg_1147;
reg [31:0] add_ln691_4_reg_1259;
reg [22:0] add_ln691_reg_1034;
reg [1:0] add_ln69_1_reg_1182;
reg [9:0] add_ln69_3_reg_1217;
reg [31:0] add_ln69_reg_1177;
reg and_ln785_reg_1078;
reg [24:0] ap_CS_fsm = 25'h0000001;
reg icmp_ln1496_reg_1162;
reg icmp_ln768_reg_1023;
reg icmp_ln786_reg_1028;
reg icmp_ln851_1_reg_1137;
reg icmp_ln851_2_reg_965;
reg icmp_ln851_3_reg_1242;
reg icmp_ln851_reg_940;
reg [3:0] newSel22_reg_1088;
reg op_15_V_reg_1167;
reg [6:0] op_21_V_reg_950;
reg [31:0] op_27_V_reg_1197;
reg [31:0] op_28_V_reg_1212;
reg [31:0] op_30_V_reg_1227;
reg or_ln785_reg_1051;
reg p_Result_6_reg_1003;
reg p_Result_7_reg_1045;
reg [5:0] p_Result_s_reg_1010;
reg [3:0] p_Val2_1_reg_1073;
reg [4:0] r_V_reg_1125;
reg [31:0] ret_V_12_cast_reg_1113;
reg [31:0] ret_V_16_cast_reg_1252;
reg [32:0] ret_V_16_reg_970;
reg [33:0] ret_V_17_reg_1108;
reg [31:0] ret_V_18_reg_1157;
reg [35:0] ret_V_19_reg_1247;
reg [6:0] ret_V_3_reg_945;
reg [2:0] ret_V_5_reg_1130;
reg [2:0] ret_V_6_reg_1142;
reg [2:0] ret_V_7_reg_1152;
reg [8:0] ret_V_reg_1192;
reg sel_tmp11_reg_1083;
reg [22:0] select_ln353_reg_1063;
reg [6:0] sext_ln831_reg_934;
reg [22:0] sext_ln850_reg_1016;
reg [4:0] sub_ln1118_reg_1103;
reg [21:0] tmp_reg_975;
reg [2:0] trunc_ln1196_1_reg_998;
reg [1:0] trunc_ln1196_reg_993;
reg [1:0] xor_ln731_reg_1039;
reg xor_ln785_reg_1057;
wire [31:0] _000_;
wire [31:0] _001_;
wire [22:0] _002_;
wire [1:0] _003_;
wire [9:0] _004_;
wire [31:0] _005_;
wire _006_;
wire [24:0] _007_;
wire _008_;
wire _009_;
wire _010_;
wire _011_;
wire _012_;
wire _013_;
wire _014_;
wire [3:0] _015_;
wire _016_;
wire [6:0] _017_;
wire [31:0] _018_;
wire [31:0] _019_;
wire [31:0] _020_;
wire _021_;
wire _022_;
wire _023_;
wire [5:0] _024_;
wire [1:0] _025_;
wire [4:0] _026_;
wire [31:0] _027_;
wire [31:0] _028_;
wire [32:0] _029_;
wire [33:0] _030_;
wire [31:0] _031_;
wire [35:0] _032_;
wire [6:0] _033_;
wire [2:0] _034_;
wire [2:0] _035_;
wire [2:0] _036_;
wire [8:0] _037_;
wire _038_;
wire [22:0] _039_;
wire [6:0] _040_;
wire [22:0] _041_;
wire [4:0] _042_;
wire [21:0] _043_;
wire [2:0] _044_;
wire [1:0] _045_;
wire [1:0] _046_;
wire _047_;
wire [1:0] _048_;
wire _049_;
wire _050_;
wire _051_;
wire _052_;
wire _053_;
wire _054_;
wire _055_;
wire _056_;
wire _057_;
wire _058_;
wire [11:0] _059_;
wire [11:0] _060_;
wire _061_;
wire [10:0] _062_;
wire [11:0] _063_;
wire [12:0] _064_;
wire [15:0] _065_;
wire [15:0] _066_;
wire _067_;
wire [15:0] _068_;
wire [16:0] _069_;
wire [16:0] _070_;
wire [15:0] _071_;
wire [15:0] _072_;
wire _073_;
wire [15:0] _074_;
wire [16:0] _075_;
wire [16:0] _076_;
wire [15:0] _077_;
wire [15:0] _078_;
wire _079_;
wire [15:0] _080_;
wire [16:0] _081_;
wire [16:0] _082_;
wire [15:0] _083_;
wire [15:0] _084_;
wire _085_;
wire [15:0] _086_;
wire [16:0] _087_;
wire [16:0] _088_;
wire [15:0] _089_;
wire [15:0] _090_;
wire _091_;
wire [15:0] _092_;
wire [16:0] _093_;
wire [16:0] _094_;
wire [16:0] _095_;
wire [16:0] _096_;
wire _097_;
wire [15:0] _098_;
wire [16:0] _099_;
wire [17:0] _100_;
wire [16:0] _101_;
wire [16:0] _102_;
wire _103_;
wire [15:0] _104_;
wire [16:0] _105_;
wire [17:0] _106_;
wire [16:0] _107_;
wire [16:0] _108_;
wire _109_;
wire [16:0] _110_;
wire [17:0] _111_;
wire [17:0] _112_;
wire [17:0] _113_;
wire [17:0] _114_;
wire _115_;
wire [17:0] _116_;
wire [18:0] _117_;
wire [18:0] _118_;
wire _119_;
wire _120_;
wire _121_;
wire _122_;
wire _123_;
wire _124_;
wire _125_;
wire _126_;
wire _127_;
wire _128_;
wire _129_;
wire _130_;
wire _131_;
wire _132_;
wire _133_;
wire _134_;
wire _135_;
wire _136_;
wire _137_;
wire _138_;
wire _139_;
wire _140_;
wire _141_;
wire _142_;
wire _143_;
wire _144_;
wire _145_;
wire _146_;
wire _147_;
wire _148_;
wire \add_23s_23ns_23_2_1_U2.ce ;
wire \add_23s_23ns_23_2_1_U2.clk ;
wire [22:0] \add_23s_23ns_23_2_1_U2.din0 ;
wire [22:0] \add_23s_23ns_23_2_1_U2.din1 ;
wire [22:0] \add_23s_23ns_23_2_1_U2.dout ;
wire \add_23s_23ns_23_2_1_U2.reset ;
wire [22:0] \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.a ;
wire [22:0] \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.ain_s0 ;
wire [22:0] \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.b ;
wire [22:0] \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.bin_s0 ;
wire \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.ce ;
wire \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.clk ;
wire \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.facout_s1 ;
wire \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.facout_s2 ;
wire [10:0] \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.fas_s1 ;
wire [11:0] \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.fas_s2 ;
wire \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.reset ;
wire [22:0] \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.s ;
wire [10:0] \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.u1.a ;
wire [10:0] \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.u1.b ;
wire \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.u1.cin ;
wire \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.u1.cout ;
wire [10:0] \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.u1.s ;
wire [11:0] \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.u2.a ;
wire [11:0] \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.u2.b ;
wire \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.u2.cin ;
wire \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.u2.cout ;
wire [11:0] \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.u2.s ;
wire \add_32ns_32ns_32_2_1_U10.ce ;
wire \add_32ns_32ns_32_2_1_U10.clk ;
wire [31:0] \add_32ns_32ns_32_2_1_U10.din0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U10.din1 ;
wire [31:0] \add_32ns_32ns_32_2_1_U10.dout ;
wire \add_32ns_32ns_32_2_1_U10.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.a ;
wire [31:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.ain_s0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.b ;
wire [31:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.bin_s0 ;
wire \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.ce ;
wire \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.clk ;
wire \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.facout_s1 ;
wire \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.facout_s2 ;
wire [15:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.fas_s1 ;
wire [15:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.fas_s2 ;
wire \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.u1.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.u1.b ;
wire \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.u1.cin ;
wire \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.u1.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.u1.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.u2.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.u2.b ;
wire \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.u2.cin ;
wire \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.u2.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.u2.s ;
wire \add_32ns_32ns_32_2_1_U4.ce ;
wire \add_32ns_32ns_32_2_1_U4.clk ;
wire [31:0] \add_32ns_32ns_32_2_1_U4.din0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U4.din1 ;
wire [31:0] \add_32ns_32ns_32_2_1_U4.dout ;
wire \add_32ns_32ns_32_2_1_U4.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.a ;
wire [31:0] \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.ain_s0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.b ;
wire [31:0] \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.bin_s0 ;
wire \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.ce ;
wire \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.clk ;
wire \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.facout_s1 ;
wire \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.facout_s2 ;
wire [15:0] \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.fas_s1 ;
wire [15:0] \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.fas_s2 ;
wire \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.u1.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.u1.b ;
wire \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.u1.cin ;
wire \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.u1.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.u1.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.u2.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.u2.b ;
wire \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.u2.cin ;
wire \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.u2.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.u2.s ;
wire \add_32ns_32s_32_2_1_U5.ce ;
wire \add_32ns_32s_32_2_1_U5.clk ;
wire [31:0] \add_32ns_32s_32_2_1_U5.din0 ;
wire [31:0] \add_32ns_32s_32_2_1_U5.din1 ;
wire [31:0] \add_32ns_32s_32_2_1_U5.dout ;
wire \add_32ns_32s_32_2_1_U5.reset ;
wire [31:0] \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.a ;
wire [31:0] \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.ain_s0 ;
wire [31:0] \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.b ;
wire [31:0] \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.bin_s0 ;
wire \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.ce ;
wire \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.clk ;
wire \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.facout_s1 ;
wire \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.facout_s2 ;
wire [15:0] \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.fas_s1 ;
wire [15:0] \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.fas_s2 ;
wire \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.reset ;
wire [31:0] \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.s ;
wire [15:0] \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.u1.a ;
wire [15:0] \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.u1.b ;
wire \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.u1.cin ;
wire \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.u1.cout ;
wire [15:0] \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.u1.s ;
wire [15:0] \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.u2.a ;
wire [15:0] \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.u2.b ;
wire \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.u2.cin ;
wire \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.u2.cout ;
wire [15:0] \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.u2.s ;
wire \add_32s_32ns_32_2_1_U6.ce ;
wire \add_32s_32ns_32_2_1_U6.clk ;
wire [31:0] \add_32s_32ns_32_2_1_U6.din0 ;
wire [31:0] \add_32s_32ns_32_2_1_U6.din1 ;
wire [31:0] \add_32s_32ns_32_2_1_U6.dout ;
wire \add_32s_32ns_32_2_1_U6.reset ;
wire [31:0] \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.a ;
wire [31:0] \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.ain_s0 ;
wire [31:0] \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.b ;
wire [31:0] \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.bin_s0 ;
wire \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.ce ;
wire \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.clk ;
wire \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.facout_s1 ;
wire \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.facout_s2 ;
wire [15:0] \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.fas_s1 ;
wire [15:0] \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.fas_s2 ;
wire \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.reset ;
wire [31:0] \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.s ;
wire [15:0] \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.u1.a ;
wire [15:0] \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.u1.b ;
wire \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.u1.cin ;
wire \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.u1.cout ;
wire [15:0] \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.u1.s ;
wire [15:0] \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.u2.a ;
wire [15:0] \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.u2.b ;
wire \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.u2.cin ;
wire \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.u2.cout ;
wire [15:0] \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.u2.s ;
wire \add_32s_32ns_32_2_1_U8.ce ;
wire \add_32s_32ns_32_2_1_U8.clk ;
wire [31:0] \add_32s_32ns_32_2_1_U8.din0 ;
wire [31:0] \add_32s_32ns_32_2_1_U8.din1 ;
wire [31:0] \add_32s_32ns_32_2_1_U8.dout ;
wire \add_32s_32ns_32_2_1_U8.reset ;
wire [31:0] \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.a ;
wire [31:0] \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.ain_s0 ;
wire [31:0] \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.b ;
wire [31:0] \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.bin_s0 ;
wire \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.ce ;
wire \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.clk ;
wire \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.facout_s1 ;
wire \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.facout_s2 ;
wire [15:0] \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.fas_s1 ;
wire [15:0] \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.fas_s2 ;
wire \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.reset ;
wire [31:0] \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.s ;
wire [15:0] \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.u1.a ;
wire [15:0] \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.u1.b ;
wire \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.u1.cin ;
wire \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.u1.cout ;
wire [15:0] \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.u1.s ;
wire [15:0] \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.u2.a ;
wire [15:0] \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.u2.b ;
wire \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.u2.cin ;
wire \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.u2.cout ;
wire [15:0] \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.u2.s ;
wire \add_33ns_33s_33_2_1_U7.ce ;
wire \add_33ns_33s_33_2_1_U7.clk ;
wire [32:0] \add_33ns_33s_33_2_1_U7.din0 ;
wire [32:0] \add_33ns_33s_33_2_1_U7.din1 ;
wire [32:0] \add_33ns_33s_33_2_1_U7.dout ;
wire \add_33ns_33s_33_2_1_U7.reset ;
wire [32:0] \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.a ;
wire [32:0] \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.ain_s0 ;
wire [32:0] \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.b ;
wire [32:0] \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.bin_s0 ;
wire \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.ce ;
wire \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.clk ;
wire \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.facout_s1 ;
wire \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.facout_s2 ;
wire [15:0] \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.fas_s1 ;
wire [16:0] \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.fas_s2 ;
wire \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.reset ;
wire [32:0] \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.s ;
wire [15:0] \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.u1.a ;
wire [15:0] \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.u1.b ;
wire \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.u1.cin ;
wire \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.u1.cout ;
wire [15:0] \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.u1.s ;
wire [16:0] \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.u2.a ;
wire [16:0] \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.u2.b ;
wire \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.u2.cin ;
wire \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.u2.cout ;
wire [16:0] \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.u2.s ;
wire \add_33s_33s_33_2_1_U1.ce ;
wire \add_33s_33s_33_2_1_U1.clk ;
wire [32:0] \add_33s_33s_33_2_1_U1.din0 ;
wire [32:0] \add_33s_33s_33_2_1_U1.din1 ;
wire [32:0] \add_33s_33s_33_2_1_U1.dout ;
wire \add_33s_33s_33_2_1_U1.reset ;
wire [32:0] \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.a ;
wire [32:0] \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.ain_s0 ;
wire [32:0] \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.b ;
wire [32:0] \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.bin_s0 ;
wire \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.ce ;
wire \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.clk ;
wire \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.facout_s1 ;
wire \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.facout_s2 ;
wire [15:0] \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.fas_s1 ;
wire [16:0] \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.fas_s2 ;
wire \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.reset ;
wire [32:0] \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.s ;
wire [15:0] \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.u1.a ;
wire [15:0] \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.u1.b ;
wire \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.u1.cin ;
wire \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.u1.cout ;
wire [15:0] \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.u1.s ;
wire [16:0] \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.u2.a ;
wire [16:0] \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.u2.b ;
wire \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.u2.cin ;
wire \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.u2.cout ;
wire [16:0] \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.u2.s ;
wire \add_34s_34s_34_2_1_U3.ce ;
wire \add_34s_34s_34_2_1_U3.clk ;
wire [33:0] \add_34s_34s_34_2_1_U3.din0 ;
wire [33:0] \add_34s_34s_34_2_1_U3.din1 ;
wire [33:0] \add_34s_34s_34_2_1_U3.dout ;
wire \add_34s_34s_34_2_1_U3.reset ;
wire [33:0] \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.a ;
wire [33:0] \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.ain_s0 ;
wire [33:0] \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.b ;
wire [33:0] \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.bin_s0 ;
wire \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.ce ;
wire \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.clk ;
wire \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.facout_s1 ;
wire \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.facout_s2 ;
wire [16:0] \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.fas_s1 ;
wire [16:0] \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.fas_s2 ;
wire \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.reset ;
wire [33:0] \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.s ;
wire [16:0] \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.u1.a ;
wire [16:0] \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.u1.b ;
wire \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.u1.cin ;
wire \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.u1.cout ;
wire [16:0] \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.u1.s ;
wire [16:0] \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.u2.a ;
wire [16:0] \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.u2.b ;
wire \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.u2.cin ;
wire \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.u2.cout ;
wire [16:0] \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.u2.s ;
wire \add_36s_36s_36_2_1_U9.ce ;
wire \add_36s_36s_36_2_1_U9.clk ;
wire [35:0] \add_36s_36s_36_2_1_U9.din0 ;
wire [35:0] \add_36s_36s_36_2_1_U9.din1 ;
wire [35:0] \add_36s_36s_36_2_1_U9.dout ;
wire \add_36s_36s_36_2_1_U9.reset ;
wire [35:0] \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.a ;
wire [35:0] \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.ain_s0 ;
wire [35:0] \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.b ;
wire [35:0] \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.bin_s0 ;
wire \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.ce ;
wire \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.clk ;
wire \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.facout_s1 ;
wire \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.facout_s2 ;
wire [17:0] \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.fas_s1 ;
wire [17:0] \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.fas_s2 ;
wire \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.reset ;
wire [35:0] \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.s ;
wire [17:0] \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.u1.a ;
wire [17:0] \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.u1.b ;
wire \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.u1.cin ;
wire \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.u1.cout ;
wire [17:0] \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.u1.s ;
wire [17:0] \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.u2.a ;
wire [17:0] \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.u2.b ;
wire \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.u2.cin ;
wire \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.u2.cout ;
wire [17:0] \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.u2.s ;
wire [1:0] add_ln69_1_fu_777_p2;
wire [9:0] add_ln69_3_fu_849_p2;
wire and_ln340_1_fu_558_p2;
wire and_ln340_fu_526_p2;
wire and_ln785_1_fu_564_p2;
wire and_ln785_fu_552_p2;
wire and_ln786_fu_537_p2;
wire ap_CS_fsm_state1;
wire ap_CS_fsm_state10;
wire ap_CS_fsm_state11;
wire ap_CS_fsm_state12;
wire ap_CS_fsm_state13;
wire ap_CS_fsm_state14;
wire ap_CS_fsm_state15;
wire ap_CS_fsm_state16;
wire ap_CS_fsm_state17;
wire ap_CS_fsm_state18;
wire ap_CS_fsm_state19;
wire ap_CS_fsm_state2;
wire ap_CS_fsm_state20;
wire ap_CS_fsm_state21;
wire ap_CS_fsm_state22;
wire ap_CS_fsm_state23;
wire ap_CS_fsm_state24;
wire ap_CS_fsm_state25;
wire ap_CS_fsm_state3;
wire ap_CS_fsm_state4;
wire ap_CS_fsm_state5;
wire ap_CS_fsm_state6;
wire ap_CS_fsm_state7;
wire ap_CS_fsm_state8;
wire ap_CS_fsm_state9;
wire [24:0] ap_NS_fsm;
wire ap_clk;
wire ap_done;
wire ap_idle;
wire ap_ready;
wire ap_rst;
wire ap_start;
wire [32:0] grp_fu_313_p0;
wire [32:0] grp_fu_313_p1;
wire [32:0] grp_fu_313_p2;
wire [22:0] grp_fu_378_p0;
wire [22:0] grp_fu_378_p2;
wire [33:0] grp_fu_604_p0;
wire [33:0] grp_fu_604_p1;
wire [33:0] grp_fu_604_p2;
wire [31:0] grp_fu_667_p2;
wire [31:0] grp_fu_756_p1;
wire [31:0] grp_fu_756_p2;
wire [31:0] grp_fu_786_p0;
wire [31:0] grp_fu_786_p2;
wire [32:0] grp_fu_825_p0;
wire [32:0] grp_fu_825_p1;
wire [32:0] grp_fu_825_p2;
wire [31:0] grp_fu_858_p0;
wire [31:0] grp_fu_858_p2;
wire [35:0] grp_fu_878_p0;
wire [35:0] grp_fu_878_p1;
wire [35:0] grp_fu_878_p2;
wire [31:0] grp_fu_904_p2;
wire icmp_ln1496_fu_730_p2;
wire icmp_ln768_fu_384_p2;
wire icmp_ln786_fu_389_p2;
wire icmp_ln851_1_fu_661_p2;
wire icmp_ln851_2_fu_323_p2;
wire icmp_ln851_3_fu_888_p2;
wire icmp_ln851_fu_257_p2;
wire [3:0] newSel22_fu_581_p3;
wire [1:0] op_0;
wire [31:0] op_10;
wire [1:0] op_11;
wire op_15_V_fu_747_p2;
wire [9:0] op_16_V_fu_807_p3;
wire [3:0] op_17;
wire [7:0] op_18;
wire [7:0] op_19;
wire [1:0] op_2;
wire [6:0] op_21_V_fu_292_p2;
wire [3:0] op_3;
wire [31:0] op_31;
wire op_31_ap_vld;
wire [7:0] op_4;
wire [3:0] op_5;
wire [3:0] op_6_V_fu_614_p3;
wire op_7;
wire [15:0] op_8;
wire [3:0] op_9;
wire or_cond_fu_610_p2;
wire or_ln340_fu_472_p2;
wire or_ln785_1_fu_547_p2;
wire or_ln785_2_fu_569_p2;
wire or_ln785_fu_406_p2;
wire or_ln786_fu_467_p2;
wire overflow_fu_458_p2;
wire p_Result_1_fu_269_p3;
wire p_Result_2_fu_677_p3;
wire p_Result_3_fu_416_p3;
wire p_Result_4_fu_696_p3;
wire p_Result_5_fu_909_p3;
wire p_Result_7_fu_398_p3;
wire p_Result_8_fu_450_p3;
wire [3:0] p_Result_s_16_fu_510_p4;
wire [3:0] p_Val2_1_fu_443_p3;
wire [2:0] p_Val2_2_fu_504_p2;
wire [4:0] r_V_fu_640_p3;
wire [7:0] ret_V_14_fu_351_p1;
wire [7:0] ret_V_14_fu_351_p2;
wire [6:0] ret_V_15_fu_281_p3;
wire [31:0] ret_V_18_fu_712_p3;
wire [5:0] ret_V_2_fu_239_p4;
wire [6:0] ret_V_3_fu_263_p2;
wire [2:0] ret_V_6_fu_672_p2;
wire [2:0] ret_V_7_fu_689_p3;
wire [8:0] ret_V_fu_801_p2;
wire [17:0] rhs_1_fu_302_p3;
wire [34:0] rhs_5_fu_867_p3;
wire sel_tmp11_fu_575_p2;
wire [22:0] select_ln353_fu_428_p3;
wire [1:0] select_ln69_fu_770_p3;
wire [8:0] select_ln703_fu_794_p3;
wire [2:0] select_ln850_1_fu_684_p3;
wire [31:0] select_ln850_3_fu_706_p3;
wire [31:0] select_ln850_4_fu_916_p3;
wire [22:0] select_ln850_6_fu_423_p3;
wire [6:0] select_ln850_fu_276_p3;
wire [4:0] sext_ln1116_fu_620_p1;
wire [31:0] sext_ln1192_fu_298_p0;
wire [1:0] sext_ln1196_fu_435_p0;
wire [2:0] sext_ln1196_fu_435_p1;
wire [3:0] sext_ln1496_fu_726_p1;
wire [4:0] sext_ln1498_fu_743_p1;
wire [9:0] sext_ln69_3_fu_841_p1;
wire [6:0] sext_ln69_fu_288_p1;
wire [7:0] sext_ln703_1_fu_791_p0;
wire [8:0] sext_ln703_1_fu_791_p1;
wire [1:0] sext_ln703_2_fu_589_p0;
wire [7:0] sext_ln703_3_fu_863_p0;
wire [1:0] sext_ln703_fu_339_p0;
wire [7:0] sext_ln703_fu_339_p1;
wire [6:0] sext_ln831_fu_249_p1;
wire [22:0] sext_ln850_fu_375_p1;
wire [1:0] shl_ln728_1_fu_736_p1;
wire [4:0] shl_ln728_1_fu_736_p3;
wire [1:0] shl_ln_fu_719_p1;
wire [2:0] shl_ln_fu_719_p3;
wire [4:0] sub_ln1118_fu_624_p2;
wire [23:0] tmp_10_fu_593_p3;
wire tmp_4_fu_477_p3;
wire tmp_5_fu_485_p3;
wire [7:0] trunc_ln1196_1_fu_347_p0;
wire [2:0] trunc_ln1196_1_fu_347_p1;
wire [7:0] trunc_ln1196_fu_343_p0;
wire [1:0] trunc_ln1196_fu_343_p1;
wire [1:0] trunc_ln851_1_fu_657_p1;
wire [31:0] trunc_ln851_2_fu_319_p0;
wire [10:0] trunc_ln851_2_fu_319_p1;
wire [1:0] trunc_ln851_3_fu_703_p0;
wire trunc_ln851_3_fu_703_p1;
wire [7:0] trunc_ln851_4_fu_884_p0;
wire [2:0] trunc_ln851_4_fu_884_p1;
wire [9:0] trunc_ln851_fu_253_p1;
wire [2:0] xor_ln1196_1_fu_438_p2;
wire xor_ln1496_fu_761_p2;
wire xor_ln340_fu_520_p2;
wire xor_ln365_1_fu_498_p2;
wire xor_ln365_fu_492_p2;
wire [1:0] xor_ln731_fu_394_p1;
wire [1:0] xor_ln731_fu_394_p2;
wire xor_ln785_1_fu_542_p2;
wire xor_ln785_fu_411_p2;
wire xor_ln786_1_fu_532_p2;
wire xor_ln786_fu_462_p2;
wire [9:0] zext_ln69_1_fu_845_p1;
wire [1:0] zext_ln69_fu_766_p1;


assign add_ln69_1_fu_777_p2 = select_ln69_fu_770_p3 + xor_ln1496_fu_761_p2;
assign add_ln69_3_fu_849_p2 = $signed({ 1'h0, op_18 }) + $signed(op_17);
assign op_21_V_fu_292_p2 = $signed(ret_V_15_fu_281_p3) + $signed(op_9);
assign ret_V_3_fu_263_p2 = $signed(op_8[15:10]) + $signed(2'h1);
assign ret_V_6_fu_672_p2 = ret_V_5_reg_1130 + 1'h1;
assign ret_V_fu_801_p2 = $signed(op_4) + $signed(select_ln703_fu_794_p3);
assign _049_ = icmp_ln851_3_reg_1242 & ap_CS_fsm[23];
assign _050_ = icmp_ln851_2_reg_965 & ap_CS_fsm[5];
assign _051_ = ap_CS_fsm[10] & _054_;
assign _052_ = _055_ & ap_CS_fsm[0];
assign _053_ = ap_start & ap_CS_fsm[0];
assign and_ln340_1_fu_558_p2 = or_ln786_fu_467_p2 & or_ln340_fu_472_p2;
assign and_ln340_fu_526_p2 = xor_ln340_fu_520_p2 & or_ln786_fu_467_p2;
assign and_ln785_1_fu_564_p2 = xor_ln785_reg_1057 & and_ln786_fu_537_p2;
assign and_ln785_fu_552_p2 = or_ln785_1_fu_547_p2 & and_ln786_fu_537_p2;
assign and_ln786_fu_537_p2 = xor_ln786_1_fu_532_p2 & p_Result_7_reg_1045;
assign overflow_fu_458_p2 = xor_ln785_reg_1057 & or_ln785_reg_1051;
assign sel_tmp11_fu_575_p2 = xor_ln365_1_fu_498_p2 & or_ln785_2_fu_569_p2;
assign xor_ln1496_fu_761_p2 = ~ icmp_ln1496_reg_1162;
assign xor_ln786_fu_462_p2 = ~ p_Result_7_reg_1045;
assign xor_ln340_fu_520_p2 = ~ or_ln340_fu_472_p2;
assign xor_ln786_1_fu_532_p2 = ~ icmp_ln786_reg_1028;
assign xor_ln785_1_fu_542_p2 = ~ or_ln785_reg_1051;
assign xor_ln365_1_fu_498_p2 = ~ xor_ln365_fu_492_p2;
assign xor_ln785_fu_411_p2 = ~ p_Result_6_reg_1003;
assign p_Val2_2_fu_504_p2 = ~ { xor_ln731_reg_1039[0], 2'h0 };
assign _054_ = ~ icmp_ln851_1_reg_1137;
assign _055_ = ~ ap_start;
assign _056_ = ! r_V_fu_640_p3[1:0];
assign _057_ = ! op_8[9:0];
assign _058_ = { op_2, 3'h0 } == { op_5[3], op_5 };
always @(posedge \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.clk )
\add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.bin_s1  <= _060_;
always @(posedge \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.clk )
\add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.ain_s1  <= _059_;
always @(posedge \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.clk )
\add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.sum_s1  <= _062_;
always @(posedge \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.clk )
\add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.carry_s1  <= _061_;
assign _060_ = \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.ce  ? \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.b [22:11] : \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.bin_s1 ;
assign _059_ = \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.ce  ? \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.a [22:11] : \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.ain_s1 ;
assign _061_ = \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.ce  ? \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.facout_s1  : \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.carry_s1 ;
assign _062_ = \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.ce  ? \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.fas_s1  : \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.sum_s1 ;
assign _063_ = \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.u1.a  + \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.u1.b ;
assign { \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.u1.cout , \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.u1.s  } = _063_ + \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.u1.cin ;
assign _064_ = \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.u2.a  + \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.u2.b ;
assign { \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.u2.cout , \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.u2.s  } = _064_ + \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.u2.cin ;
always @(posedge \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.clk )
\add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.bin_s1  <= _066_;
always @(posedge \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.clk )
\add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.ain_s1  <= _065_;
always @(posedge \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.clk )
\add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.sum_s1  <= _068_;
always @(posedge \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.clk )
\add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.carry_s1  <= _067_;
assign _066_ = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.ce  ? \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.b [31:16] : \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.bin_s1 ;
assign _065_ = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.ce  ? \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.a [31:16] : \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.ain_s1 ;
assign _067_ = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.ce  ? \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.facout_s1  : \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.carry_s1 ;
assign _068_ = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.ce  ? \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.fas_s1  : \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.sum_s1 ;
assign _069_ = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.u1.a  + \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.u1.b ;
assign { \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.u1.cout , \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.u1.s  } = _069_ + \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.u1.cin ;
assign _070_ = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.u2.a  + \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.u2.b ;
assign { \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.u2.cout , \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.u2.s  } = _070_ + \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.u2.cin ;
always @(posedge \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.clk )
\add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.bin_s1  <= _072_;
always @(posedge \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.clk )
\add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.ain_s1  <= _071_;
always @(posedge \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.clk )
\add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.sum_s1  <= _074_;
always @(posedge \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.clk )
\add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.carry_s1  <= _073_;
assign _072_ = \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.ce  ? \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.b [31:16] : \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.bin_s1 ;
assign _071_ = \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.ce  ? \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.a [31:16] : \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.ain_s1 ;
assign _073_ = \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.ce  ? \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.facout_s1  : \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.carry_s1 ;
assign _074_ = \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.ce  ? \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.fas_s1  : \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.sum_s1 ;
assign _075_ = \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.u1.a  + \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.u1.b ;
assign { \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.u1.cout , \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.u1.s  } = _075_ + \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.u1.cin ;
assign _076_ = \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.u2.a  + \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.u2.b ;
assign { \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.u2.cout , \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.u2.s  } = _076_ + \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.u2.cin ;
always @(posedge \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.clk )
\add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.bin_s1  <= _078_;
always @(posedge \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.clk )
\add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.ain_s1  <= _077_;
always @(posedge \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.clk )
\add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.sum_s1  <= _080_;
always @(posedge \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.clk )
\add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.carry_s1  <= _079_;
assign _078_ = \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.ce  ? \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.b [31:16] : \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.bin_s1 ;
assign _077_ = \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.ce  ? \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.a [31:16] : \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.ain_s1 ;
assign _079_ = \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.ce  ? \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.facout_s1  : \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.carry_s1 ;
assign _080_ = \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.ce  ? \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.fas_s1  : \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.sum_s1 ;
assign _081_ = \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.u1.a  + \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.u1.b ;
assign { \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.u1.cout , \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.u1.s  } = _081_ + \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.u1.cin ;
assign _082_ = \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.u2.a  + \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.u2.b ;
assign { \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.u2.cout , \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.u2.s  } = _082_ + \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.u2.cin ;
always @(posedge \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.clk )
\add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.bin_s1  <= _084_;
always @(posedge \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.clk )
\add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.ain_s1  <= _083_;
always @(posedge \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.clk )
\add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.sum_s1  <= _086_;
always @(posedge \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.clk )
\add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.carry_s1  <= _085_;
assign _084_ = \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.ce  ? \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.b [31:16] : \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.bin_s1 ;
assign _083_ = \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.ce  ? \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.a [31:16] : \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.ain_s1 ;
assign _085_ = \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.ce  ? \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.facout_s1  : \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.carry_s1 ;
assign _086_ = \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.ce  ? \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.fas_s1  : \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.sum_s1 ;
assign _087_ = \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.u1.a  + \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.u1.b ;
assign { \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.u1.cout , \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.u1.s  } = _087_ + \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.u1.cin ;
assign _088_ = \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.u2.a  + \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.u2.b ;
assign { \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.u2.cout , \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.u2.s  } = _088_ + \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.u2.cin ;
always @(posedge \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.clk )
\add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.bin_s1  <= _090_;
always @(posedge \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.clk )
\add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.ain_s1  <= _089_;
always @(posedge \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.clk )
\add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.sum_s1  <= _092_;
always @(posedge \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.clk )
\add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.carry_s1  <= _091_;
assign _090_ = \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.ce  ? \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.b [31:16] : \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.bin_s1 ;
assign _089_ = \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.ce  ? \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.a [31:16] : \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.ain_s1 ;
assign _091_ = \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.ce  ? \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.facout_s1  : \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.carry_s1 ;
assign _092_ = \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.ce  ? \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.fas_s1  : \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.sum_s1 ;
assign _093_ = \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.u1.a  + \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.u1.b ;
assign { \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.u1.cout , \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.u1.s  } = _093_ + \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.u1.cin ;
assign _094_ = \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.u2.a  + \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.u2.b ;
assign { \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.u2.cout , \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.u2.s  } = _094_ + \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.u2.cin ;
always @(posedge \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.clk )
\add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.bin_s1  <= _096_;
always @(posedge \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.clk )
\add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.ain_s1  <= _095_;
always @(posedge \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.clk )
\add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.sum_s1  <= _098_;
always @(posedge \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.clk )
\add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.carry_s1  <= _097_;
assign _096_ = \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.ce  ? \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.b [32:16] : \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.bin_s1 ;
assign _095_ = \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.ce  ? \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.a [32:16] : \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.ain_s1 ;
assign _097_ = \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.ce  ? \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.facout_s1  : \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.carry_s1 ;
assign _098_ = \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.ce  ? \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.fas_s1  : \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.sum_s1 ;
assign _099_ = \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.u1.a  + \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.u1.b ;
assign { \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.u1.cout , \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.u1.s  } = _099_ + \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.u1.cin ;
assign _100_ = \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.u2.a  + \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.u2.b ;
assign { \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.u2.cout , \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.u2.s  } = _100_ + \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.u2.cin ;
always @(posedge \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.clk )
\add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.bin_s1  <= _102_;
always @(posedge \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.clk )
\add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.ain_s1  <= _101_;
always @(posedge \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.clk )
\add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.sum_s1  <= _104_;
always @(posedge \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.clk )
\add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.carry_s1  <= _103_;
assign _102_ = \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.ce  ? \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.b [32:16] : \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.bin_s1 ;
assign _101_ = \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.ce  ? \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.a [32:16] : \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.ain_s1 ;
assign _103_ = \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.ce  ? \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.facout_s1  : \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.carry_s1 ;
assign _104_ = \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.ce  ? \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.fas_s1  : \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.sum_s1 ;
assign _105_ = \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.u1.a  + \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.u1.b ;
assign { \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.u1.cout , \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.u1.s  } = _105_ + \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.u1.cin ;
assign _106_ = \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.u2.a  + \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.u2.b ;
assign { \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.u2.cout , \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.u2.s  } = _106_ + \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.u2.cin ;
always @(posedge \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.clk )
\add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.bin_s1  <= _108_;
always @(posedge \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.clk )
\add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.ain_s1  <= _107_;
always @(posedge \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.clk )
\add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.sum_s1  <= _110_;
always @(posedge \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.clk )
\add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.carry_s1  <= _109_;
assign _108_ = \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.ce  ? \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.b [33:17] : \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.bin_s1 ;
assign _107_ = \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.ce  ? \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.a [33:17] : \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.ain_s1 ;
assign _109_ = \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.ce  ? \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.facout_s1  : \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.carry_s1 ;
assign _110_ = \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.ce  ? \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.fas_s1  : \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.sum_s1 ;
assign _111_ = \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.u1.a  + \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.u1.b ;
assign { \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.u1.cout , \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.u1.s  } = _111_ + \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.u1.cin ;
assign _112_ = \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.u2.a  + \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.u2.b ;
assign { \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.u2.cout , \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.u2.s  } = _112_ + \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.u2.cin ;
always @(posedge \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.clk )
\add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.bin_s1  <= _114_;
always @(posedge \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.clk )
\add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.ain_s1  <= _113_;
always @(posedge \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.clk )
\add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.sum_s1  <= _116_;
always @(posedge \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.clk )
\add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.carry_s1  <= _115_;
assign _114_ = \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.ce  ? \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.b [35:18] : \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.bin_s1 ;
assign _113_ = \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.ce  ? \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.a [35:18] : \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.ain_s1 ;
assign _115_ = \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.ce  ? \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.facout_s1  : \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.carry_s1 ;
assign _116_ = \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.ce  ? \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.fas_s1  : \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.sum_s1 ;
assign _117_ = \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.u1.a  + \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.u1.b ;
assign { \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.u1.cout , \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.u1.s  } = _117_ + \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.u1.cin ;
assign _118_ = \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.u2.a  + \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.u2.b ;
assign { \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.u2.cout , \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.u2.s  } = _118_ + \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.u2.cin ;
assign _119_ = $signed({ op_2, 1'h0 }) < $signed(op_3);
assign _120_ = | p_Result_s_reg_1010;
assign _121_ = p_Result_s_reg_1010 != 6'h3f;
assign _122_ = | op_10[10:0];
assign _123_ = | op_19[2:0];
assign or_cond_fu_610_p2 = sel_tmp11_reg_1083 | and_ln785_reg_1078;
assign or_ln340_fu_472_p2 = p_Result_6_reg_1003 | overflow_fu_458_p2;
assign or_ln785_1_fu_547_p2 = xor_ln785_1_fu_542_p2 | p_Result_6_reg_1003;
assign or_ln785_2_fu_569_p2 = and_ln785_1_fu_564_p2 | and_ln340_1_fu_558_p2;
assign or_ln785_fu_406_p2 = xor_ln731_fu_394_p2[1] | icmp_ln768_reg_1023;
assign or_ln786_fu_467_p2 = xor_ln786_fu_462_p2 | icmp_ln786_reg_1028;
always @(posedge ap_clk)
p_Val2_1_reg_1073[1:0] <= 2'h0;
always @(posedge ap_clk)
ret_V_6_reg_1142 <= _035_;
always @(posedge ap_clk)
ret_V_7_reg_1152 <= _036_;
always @(posedge ap_clk)
ret_V_18_reg_1157 <= _031_;
always @(posedge ap_clk)
ret_V_16_reg_970 <= _029_;
always @(posedge ap_clk)
tmp_reg_975 <= _043_;
always @(posedge ap_clk)
ret_V_19_reg_1247 <= _032_;
always @(posedge ap_clk)
ret_V_16_cast_reg_1252 <= _028_;
always @(posedge ap_clk)
sub_ln1118_reg_1103 <= _042_;
always @(posedge ap_clk)
ret_V_17_reg_1108 <= _030_;
always @(posedge ap_clk)
ret_V_12_cast_reg_1113 <= _027_;
always @(posedge ap_clk)
trunc_ln1196_reg_993 <= _045_;
always @(posedge ap_clk)
trunc_ln1196_1_reg_998 <= _044_;
always @(posedge ap_clk)
p_Result_6_reg_1003 <= _022_;
always @(posedge ap_clk)
p_Result_s_reg_1010 <= _024_;
always @(posedge ap_clk)
sext_ln850_reg_1016 <= _041_;
always @(posedge ap_clk)
xor_ln731_reg_1039 <= _046_;
always @(posedge ap_clk)
p_Result_7_reg_1045 <= _023_;
always @(posedge ap_clk)
or_ln785_reg_1051 <= _021_;
always @(posedge ap_clk)
xor_ln785_reg_1057 <= _047_;
always @(posedge ap_clk)
select_ln353_reg_1063 <= _039_;
always @(posedge ap_clk)
op_30_V_reg_1227 <= _020_;
always @(posedge ap_clk)
ret_V_reg_1192 <= _037_;
always @(posedge ap_clk)
op_27_V_reg_1197 <= _018_;
always @(posedge ap_clk)
op_21_V_reg_950 <= _017_;
always @(posedge ap_clk)
sext_ln831_reg_934 <= _040_;
always @(posedge ap_clk)
icmp_ln851_reg_940 <= _014_;
always @(posedge ap_clk)
ret_V_3_reg_945 <= _033_;
always @(posedge ap_clk)
icmp_ln851_3_reg_1242 <= _013_;
always @(posedge ap_clk)
icmp_ln851_2_reg_965 <= _012_;
always @(posedge ap_clk)
r_V_reg_1125 <= _026_;
always @(posedge ap_clk)
ret_V_5_reg_1130 <= _034_;
always @(posedge ap_clk)
icmp_ln851_1_reg_1137 <= _011_;
always @(posedge ap_clk)
icmp_ln768_reg_1023 <= _009_;
always @(posedge ap_clk)
icmp_ln786_reg_1028 <= _010_;
always @(posedge ap_clk)
icmp_ln1496_reg_1162 <= _008_;
always @(posedge ap_clk)
op_15_V_reg_1167 <= _016_;
always @(posedge ap_clk)
p_Val2_1_reg_1073[3:2] <= _025_;
always @(posedge ap_clk)
and_ln785_reg_1078 <= _006_;
always @(posedge ap_clk)
sel_tmp11_reg_1083 <= _038_;
always @(posedge ap_clk)
newSel22_reg_1088 <= _015_;
always @(posedge ap_clk)
op_28_V_reg_1212 <= _019_;
always @(posedge ap_clk)
add_ln69_3_reg_1217 <= _004_;
always @(posedge ap_clk)
add_ln69_reg_1177 <= _005_;
always @(posedge ap_clk)
add_ln69_1_reg_1182 <= _003_;
always @(posedge ap_clk)
add_ln691_reg_1034 <= _002_;
always @(posedge ap_clk)
add_ln691_4_reg_1259 <= _001_;
always @(posedge ap_clk)
add_ln691_1_reg_1147 <= _000_;
always @(posedge ap_clk)
ap_CS_fsm <= _007_;
assign _048_ = _053_ ? 2'h2 : 2'h1;
assign _124_ = ap_CS_fsm == 1'h1;
function [24:0] _362_;
input [24:0] a;
input [624:0] b;
input [24:0] s;
case (s)
25'b0000000000000000000000001:
_362_ = b[24:0];
25'b0000000000000000000000010:
_362_ = b[49:25];
25'b0000000000000000000000100:
_362_ = b[74:50];
25'b0000000000000000000001000:
_362_ = b[99:75];
25'b0000000000000000000010000:
_362_ = b[124:100];
25'b0000000000000000000100000:
_362_ = b[149:125];
25'b0000000000000000001000000:
_362_ = b[174:150];
25'b0000000000000000010000000:
_362_ = b[199:175];
25'b0000000000000000100000000:
_362_ = b[224:200];
25'b0000000000000001000000000:
_362_ = b[249:225];
25'b0000000000000010000000000:
_362_ = b[274:250];
25'b0000000000000100000000000:
_362_ = b[299:275];
25'b0000000000001000000000000:
_362_ = b[324:300];
25'b0000000000010000000000000:
_362_ = b[349:325];
25'b0000000000100000000000000:
_362_ = b[374:350];
25'b0000000001000000000000000:
_362_ = b[399:375];
25'b0000000010000000000000000:
_362_ = b[424:400];
25'b0000000100000000000000000:
_362_ = b[449:425];
25'b0000001000000000000000000:
_362_ = b[474:450];
25'b0000010000000000000000000:
_362_ = b[499:475];
25'b0000100000000000000000000:
_362_ = b[524:500];
25'b0001000000000000000000000:
_362_ = b[549:525];
25'b0010000000000000000000000:
_362_ = b[574:550];
25'b0100000000000000000000000:
_362_ = b[599:575];
25'b1000000000000000000000000:
_362_ = b[624:600];
25'b0000000000000000000000000:
_362_ = a;
default:
_362_ = 25'bx;
endcase
endfunction
assign ap_NS_fsm = _362_(25'hxxxxxxx, { 23'h000000, _048_, 600'h000002000002000002000002000002000002000002000002000002000002000002000002000002000002000002000002000002000002000002000002000002000002000002000000000001 }, { _124_, _148_, _147_, _146_, _145_, _144_, _143_, _142_, _141_, _140_, _139_, _138_, _137_, _136_, _135_, _134_, _133_, _132_, _131_, _130_, _129_, _128_, _127_, _126_, _125_ });
assign _125_ = ap_CS_fsm == 25'h1000000;
assign _126_ = ap_CS_fsm == 24'h800000;
assign _127_ = ap_CS_fsm == 23'h400000;
assign _128_ = ap_CS_fsm == 22'h200000;
assign _129_ = ap_CS_fsm == 21'h100000;
assign _130_ = ap_CS_fsm == 20'h80000;
assign _131_ = ap_CS_fsm == 19'h40000;
assign _132_ = ap_CS_fsm == 18'h20000;
assign _133_ = ap_CS_fsm == 17'h10000;
assign _134_ = ap_CS_fsm == 16'h8000;
assign _135_ = ap_CS_fsm == 15'h4000;
assign _136_ = ap_CS_fsm == 14'h2000;
assign _137_ = ap_CS_fsm == 13'h1000;
assign _138_ = ap_CS_fsm == 12'h800;
assign _139_ = ap_CS_fsm == 11'h400;
assign _140_ = ap_CS_fsm == 10'h200;
assign _141_ = ap_CS_fsm == 9'h100;
assign _142_ = ap_CS_fsm == 8'h80;
assign _143_ = ap_CS_fsm == 7'h40;
assign _144_ = ap_CS_fsm == 6'h20;
assign _145_ = ap_CS_fsm == 5'h10;
assign _146_ = ap_CS_fsm == 4'h8;
assign _147_ = ap_CS_fsm == 3'h4;
assign _148_ = ap_CS_fsm == 2'h2;
assign op_31_ap_vld = ap_CS_fsm[24] ? 1'h1 : 1'h0;
assign ap_idle = _052_ ? 1'h1 : 1'h0;
assign _035_ = _051_ ? ret_V_6_fu_672_p2 : ret_V_6_reg_1142;
assign _031_ = ap_CS_fsm[11] ? ret_V_18_fu_712_p3 : ret_V_18_reg_1157;
assign _036_ = ap_CS_fsm[11] ? ret_V_7_fu_689_p3 : ret_V_7_reg_1152;
assign _043_ = ap_CS_fsm[3] ? grp_fu_313_p2[32:11] : tmp_reg_975;
assign _029_ = ap_CS_fsm[3] ? grp_fu_313_p2 : ret_V_16_reg_970;
assign _028_ = ap_CS_fsm[21] ? grp_fu_878_p2[34:3] : ret_V_16_cast_reg_1252;
assign _032_ = ap_CS_fsm[21] ? grp_fu_878_p2 : ret_V_19_reg_1247;
assign _027_ = ap_CS_fsm[8] ? grp_fu_604_p2[32:1] : ret_V_12_cast_reg_1113;
assign _030_ = ap_CS_fsm[8] ? grp_fu_604_p2 : ret_V_17_reg_1108;
assign _042_ = ap_CS_fsm[8] ? sub_ln1118_fu_624_p2 : sub_ln1118_reg_1103;
assign _041_ = ap_CS_fsm[4] ? { tmp_reg_975[21], tmp_reg_975 } : sext_ln850_reg_1016;
assign _024_ = ap_CS_fsm[4] ? ret_V_14_fu_351_p2[7:2] : p_Result_s_reg_1010;
assign _022_ = ap_CS_fsm[4] ? ret_V_14_fu_351_p2[7] : p_Result_6_reg_1003;
assign _044_ = ap_CS_fsm[4] ? op_4[2:0] : trunc_ln1196_1_reg_998;
assign _045_ = ap_CS_fsm[4] ? op_4[1:0] : trunc_ln1196_reg_993;
assign _039_ = ap_CS_fsm[6] ? select_ln353_fu_428_p3 : select_ln353_reg_1063;
assign _047_ = ap_CS_fsm[6] ? xor_ln785_fu_411_p2 : xor_ln785_reg_1057;
assign _021_ = ap_CS_fsm[6] ? or_ln785_fu_406_p2 : or_ln785_reg_1051;
assign _023_ = ap_CS_fsm[6] ? xor_ln731_fu_394_p2[1] : p_Result_7_reg_1045;
assign _046_ = ap_CS_fsm[6] ? xor_ln731_fu_394_p2 : xor_ln731_reg_1039;
assign _020_ = ap_CS_fsm[19] ? grp_fu_858_p2 : op_30_V_reg_1227;
assign _018_ = ap_CS_fsm[15] ? grp_fu_786_p2 : op_27_V_reg_1197;
assign _037_ = ap_CS_fsm[15] ? ret_V_fu_801_p2 : ret_V_reg_1192;
assign _017_ = ap_CS_fsm[1] ? op_21_V_fu_292_p2 : op_21_V_reg_950;
assign _033_ = ap_CS_fsm[0] ? ret_V_3_fu_263_p2 : ret_V_3_reg_945;
assign _014_ = ap_CS_fsm[0] ? icmp_ln851_fu_257_p2 : icmp_ln851_reg_940;
assign _040_ = ap_CS_fsm[0] ? { op_8[15], op_8[15:10] } : sext_ln831_reg_934;
assign _013_ = ap_CS_fsm[20] ? icmp_ln851_3_fu_888_p2 : icmp_ln851_3_reg_1242;
assign _012_ = ap_CS_fsm[2] ? icmp_ln851_2_fu_323_p2 : icmp_ln851_2_reg_965;
assign _011_ = ap_CS_fsm[9] ? icmp_ln851_1_fu_661_p2 : icmp_ln851_1_reg_1137;
assign _034_ = ap_CS_fsm[9] ? r_V_fu_640_p3[4:2] : ret_V_5_reg_1130;
assign _026_ = ap_CS_fsm[9] ? r_V_fu_640_p3 : r_V_reg_1125;
assign _010_ = ap_CS_fsm[5] ? icmp_ln786_fu_389_p2 : icmp_ln786_reg_1028;
assign _009_ = ap_CS_fsm[5] ? icmp_ln768_fu_384_p2 : icmp_ln768_reg_1023;
assign _016_ = ap_CS_fsm[12] ? op_15_V_fu_747_p2 : op_15_V_reg_1167;
assign _008_ = ap_CS_fsm[12] ? icmp_ln1496_fu_730_p2 : icmp_ln1496_reg_1162;
assign _015_ = ap_CS_fsm[7] ? newSel22_fu_581_p3 : newSel22_reg_1088;
assign _038_ = ap_CS_fsm[7] ? sel_tmp11_fu_575_p2 : sel_tmp11_reg_1083;
assign _006_ = ap_CS_fsm[7] ? and_ln785_fu_552_p2 : and_ln785_reg_1078;
assign _025_ = ap_CS_fsm[7] ? xor_ln731_reg_1039 : p_Val2_1_reg_1073[3:2];
assign _004_ = ap_CS_fsm[17] ? add_ln69_3_fu_849_p2 : add_ln69_3_reg_1217;
assign _019_ = ap_CS_fsm[17] ? grp_fu_825_p2[32:1] : op_28_V_reg_1212;
assign _003_ = ap_CS_fsm[13] ? add_ln69_1_fu_777_p2 : add_ln69_1_reg_1182;
assign _005_ = ap_CS_fsm[13] ? grp_fu_756_p2 : add_ln69_reg_1177;
assign _002_ = _050_ ? grp_fu_378_p2 : add_ln691_reg_1034;
assign _001_ = _049_ ? grp_fu_904_p2 : add_ln691_4_reg_1259;
assign _000_ = ap_CS_fsm[10] ? grp_fu_667_p2 : add_ln691_1_reg_1147;
assign _007_ = ap_rst ? 25'h0000001 : ap_NS_fsm;
assign sub_ln1118_fu_624_p2 = $signed(1'h0) - $signed(op_6_V_fu_614_p3);
assign icmp_ln1496_fu_730_p2 = _119_ ? 1'h1 : 1'h0;
assign icmp_ln768_fu_384_p2 = _120_ ? 1'h1 : 1'h0;
assign icmp_ln786_fu_389_p2 = _121_ ? 1'h1 : 1'h0;
assign icmp_ln851_1_fu_661_p2 = _056_ ? 1'h1 : 1'h0;
assign icmp_ln851_2_fu_323_p2 = _122_ ? 1'h1 : 1'h0;
assign icmp_ln851_3_fu_888_p2 = _123_ ? 1'h1 : 1'h0;
assign icmp_ln851_fu_257_p2 = _057_ ? 1'h1 : 1'h0;
assign newSel22_fu_581_p3 = and_ln340_fu_526_p2 ? { xor_ln731_reg_1039, 2'h0 } : { xor_ln1196_1_fu_438_p2[2], p_Val2_2_fu_504_p2 };
assign op_15_V_fu_747_p2 = _058_ ? 1'h1 : 1'h0;
assign op_31 = ret_V_19_reg_1247[35] ? select_ln850_4_fu_916_p3 : ret_V_16_cast_reg_1252;
assign op_6_V_fu_614_p3 = or_cond_fu_610_p2 ? p_Val2_1_reg_1073 : newSel22_reg_1088;
assign r_V_fu_640_p3 = op_7 ? sub_ln1118_reg_1103 : 5'h00;
assign ret_V_15_fu_281_p3 = op_8[15] ? select_ln850_fu_276_p3 : sext_ln831_reg_934;
assign ret_V_18_fu_712_p3 = ret_V_17_reg_1108[33] ? select_ln850_3_fu_706_p3 : ret_V_12_cast_reg_1113;
assign ret_V_7_fu_689_p3 = r_V_reg_1125[4] ? select_ln850_1_fu_684_p3 : ret_V_5_reg_1130;
assign select_ln353_fu_428_p3 = ret_V_16_reg_970[32] ? select_ln850_6_fu_423_p3 : sext_ln850_reg_1016;
assign select_ln69_fu_770_p3 = op_15_V_reg_1167 ? 2'h3 : 2'h0;
assign select_ln703_fu_794_p3 = op_7 ? 9'h1ff : 9'h000;
assign select_ln850_1_fu_684_p3 = icmp_ln851_1_reg_1137 ? ret_V_5_reg_1130 : ret_V_6_reg_1142;
assign select_ln850_3_fu_706_p3 = op_11[0] ? add_ln691_1_reg_1147 : ret_V_12_cast_reg_1113;
assign select_ln850_4_fu_916_p3 = icmp_ln851_3_reg_1242 ? add_ln691_4_reg_1259 : ret_V_16_cast_reg_1252;
assign select_ln850_6_fu_423_p3 = icmp_ln851_2_reg_965 ? add_ln691_reg_1034 : sext_ln850_reg_1016;
assign select_ln850_fu_276_p3 = icmp_ln851_reg_940 ? sext_ln831_reg_934 : ret_V_3_reg_945;
assign ret_V_14_fu_351_p2 = $signed(op_2) ^ $signed(op_4);
assign xor_ln1196_1_fu_438_p2 = trunc_ln1196_1_reg_998 ^ { op_2[1], op_2 };
assign xor_ln365_fu_492_p2 = xor_ln731_reg_1039[1] ^ xor_ln1196_1_fu_438_p2[2];
assign xor_ln731_fu_394_p2 = op_2 ^ trunc_ln1196_reg_993;
assign ap_CS_fsm_state1 = ap_CS_fsm[0];
assign ap_CS_fsm_state10 = ap_CS_fsm[9];
assign ap_CS_fsm_state11 = ap_CS_fsm[10];
assign ap_CS_fsm_state12 = ap_CS_fsm[11];
assign ap_CS_fsm_state13 = ap_CS_fsm[12];
assign ap_CS_fsm_state14 = ap_CS_fsm[13];
assign ap_CS_fsm_state15 = ap_CS_fsm[14];
assign ap_CS_fsm_state16 = ap_CS_fsm[15];
assign ap_CS_fsm_state17 = ap_CS_fsm[16];
assign ap_CS_fsm_state18 = ap_CS_fsm[17];
assign ap_CS_fsm_state19 = ap_CS_fsm[18];
assign ap_CS_fsm_state2 = ap_CS_fsm[1];
assign ap_CS_fsm_state20 = ap_CS_fsm[19];
assign ap_CS_fsm_state21 = ap_CS_fsm[20];
assign ap_CS_fsm_state22 = ap_CS_fsm[21];
assign ap_CS_fsm_state23 = ap_CS_fsm[22];
assign ap_CS_fsm_state24 = ap_CS_fsm[23];
assign ap_CS_fsm_state25 = ap_CS_fsm[24];
assign ap_CS_fsm_state3 = ap_CS_fsm[2];
assign ap_CS_fsm_state4 = ap_CS_fsm[3];
assign ap_CS_fsm_state5 = ap_CS_fsm[4];
assign ap_CS_fsm_state6 = ap_CS_fsm[5];
assign ap_CS_fsm_state7 = ap_CS_fsm[6];
assign ap_CS_fsm_state8 = ap_CS_fsm[7];
assign ap_CS_fsm_state9 = ap_CS_fsm[8];
assign ap_done = op_31_ap_vld;
assign ap_ready = op_31_ap_vld;
assign grp_fu_313_p0 = { op_21_V_reg_950[6], op_21_V_reg_950[6], op_21_V_reg_950[6], op_21_V_reg_950[6], op_21_V_reg_950[6], op_21_V_reg_950[6], op_21_V_reg_950[6], op_21_V_reg_950[6], op_21_V_reg_950[6], op_21_V_reg_950[6], op_21_V_reg_950[6], op_21_V_reg_950[6], op_21_V_reg_950[6], op_21_V_reg_950[6], op_21_V_reg_950[6], op_21_V_reg_950, 11'h000 };
assign grp_fu_313_p1 = { op_10[31], op_10 };
assign grp_fu_378_p0 = { tmp_reg_975[21], tmp_reg_975 };
assign grp_fu_604_p0 = { select_ln353_reg_1063[22], select_ln353_reg_1063[22], select_ln353_reg_1063[22], select_ln353_reg_1063[22], select_ln353_reg_1063[22], select_ln353_reg_1063[22], select_ln353_reg_1063[22], select_ln353_reg_1063[22], select_ln353_reg_1063[22], select_ln353_reg_1063[22], select_ln353_reg_1063, 1'h0 };
assign grp_fu_604_p1 = { op_11[1], op_11[1], op_11[1], op_11[1], op_11[1], op_11[1], op_11[1], op_11[1], op_11[1], op_11[1], op_11[1], op_11[1], op_11[1], op_11[1], op_11[1], op_11[1], op_11[1], op_11[1], op_11[1], op_11[1], op_11[1], op_11[1], op_11[1], op_11[1], op_11[1], op_11[1], op_11[1], op_11[1], op_11[1], op_11[1], op_11[1], op_11[1], op_11 };
assign grp_fu_756_p1 = { ret_V_7_reg_1152[2], ret_V_7_reg_1152[2], ret_V_7_reg_1152[2], ret_V_7_reg_1152[2], ret_V_7_reg_1152[2], ret_V_7_reg_1152[2], ret_V_7_reg_1152[2], ret_V_7_reg_1152[2], ret_V_7_reg_1152[2], ret_V_7_reg_1152[2], ret_V_7_reg_1152[2], ret_V_7_reg_1152[2], ret_V_7_reg_1152[2], ret_V_7_reg_1152[2], ret_V_7_reg_1152[2], ret_V_7_reg_1152[2], ret_V_7_reg_1152[2], ret_V_7_reg_1152[2], ret_V_7_reg_1152[2], ret_V_7_reg_1152[2], ret_V_7_reg_1152[2], ret_V_7_reg_1152[2], ret_V_7_reg_1152[2], ret_V_7_reg_1152[2], ret_V_7_reg_1152[2], ret_V_7_reg_1152[2], ret_V_7_reg_1152[2], ret_V_7_reg_1152[2], ret_V_7_reg_1152[2], ret_V_7_reg_1152 };
assign grp_fu_786_p0 = { add_ln69_1_reg_1182[1], add_ln69_1_reg_1182[1], add_ln69_1_reg_1182[1], add_ln69_1_reg_1182[1], add_ln69_1_reg_1182[1], add_ln69_1_reg_1182[1], add_ln69_1_reg_1182[1], add_ln69_1_reg_1182[1], add_ln69_1_reg_1182[1], add_ln69_1_reg_1182[1], add_ln69_1_reg_1182[1], add_ln69_1_reg_1182[1], add_ln69_1_reg_1182[1], add_ln69_1_reg_1182[1], add_ln69_1_reg_1182[1], add_ln69_1_reg_1182[1], add_ln69_1_reg_1182[1], add_ln69_1_reg_1182[1], add_ln69_1_reg_1182[1], add_ln69_1_reg_1182[1], add_ln69_1_reg_1182[1], add_ln69_1_reg_1182[1], add_ln69_1_reg_1182[1], add_ln69_1_reg_1182[1], add_ln69_1_reg_1182[1], add_ln69_1_reg_1182[1], add_ln69_1_reg_1182[1], add_ln69_1_reg_1182[1], add_ln69_1_reg_1182[1], add_ln69_1_reg_1182[1], add_ln69_1_reg_1182 };
assign grp_fu_825_p0 = { op_27_V_reg_1197, 1'h0 };
assign grp_fu_825_p1 = { ret_V_reg_1192[8], ret_V_reg_1192[8], ret_V_reg_1192[8], ret_V_reg_1192[8], ret_V_reg_1192[8], ret_V_reg_1192[8], ret_V_reg_1192[8], ret_V_reg_1192[8], ret_V_reg_1192[8], ret_V_reg_1192[8], ret_V_reg_1192[8], ret_V_reg_1192[8], ret_V_reg_1192[8], ret_V_reg_1192[8], ret_V_reg_1192[8], ret_V_reg_1192[8], ret_V_reg_1192[8], ret_V_reg_1192[8], ret_V_reg_1192[8], ret_V_reg_1192[8], ret_V_reg_1192[8], ret_V_reg_1192[8], ret_V_reg_1192[8], ret_V_reg_1192, 1'h0 };
assign grp_fu_858_p0 = { add_ln69_3_reg_1217[9], add_ln69_3_reg_1217[9], add_ln69_3_reg_1217[9], add_ln69_3_reg_1217[9], add_ln69_3_reg_1217[9], add_ln69_3_reg_1217[9], add_ln69_3_reg_1217[9], add_ln69_3_reg_1217[9], add_ln69_3_reg_1217[9], add_ln69_3_reg_1217[9], add_ln69_3_reg_1217[9], add_ln69_3_reg_1217[9], add_ln69_3_reg_1217[9], add_ln69_3_reg_1217[9], add_ln69_3_reg_1217[9], add_ln69_3_reg_1217[9], add_ln69_3_reg_1217[9], add_ln69_3_reg_1217[9], add_ln69_3_reg_1217[9], add_ln69_3_reg_1217[9], add_ln69_3_reg_1217[9], add_ln69_3_reg_1217[9], add_ln69_3_reg_1217 };
assign grp_fu_878_p0 = { op_30_V_reg_1227[31], op_30_V_reg_1227, 3'h0 };
assign grp_fu_878_p1 = { op_19[7], op_19[7], op_19[7], op_19[7], op_19[7], op_19[7], op_19[7], op_19[7], op_19[7], op_19[7], op_19[7], op_19[7], op_19[7], op_19[7], op_19[7], op_19[7], op_19[7], op_19[7], op_19[7], op_19[7], op_19[7], op_19[7], op_19[7], op_19[7], op_19[7], op_19[7], op_19[7], op_19[7], op_19 };
assign op_16_V_fu_807_p3 = { ret_V_reg_1192, 1'h0 };
assign p_Result_1_fu_269_p3 = op_8[15];
assign p_Result_2_fu_677_p3 = r_V_reg_1125[4];
assign p_Result_3_fu_416_p3 = ret_V_16_reg_970[32];
assign p_Result_4_fu_696_p3 = ret_V_17_reg_1108[33];
assign p_Result_5_fu_909_p3 = ret_V_19_reg_1247[35];
assign p_Result_7_fu_398_p3 = xor_ln731_fu_394_p2[1];
assign p_Result_8_fu_450_p3 = xor_ln1196_1_fu_438_p2[2];
assign p_Result_s_16_fu_510_p4 = { xor_ln1196_1_fu_438_p2[2], p_Val2_2_fu_504_p2 };
assign p_Val2_1_fu_443_p3 = { xor_ln731_reg_1039, 2'h0 };
assign ret_V_14_fu_351_p1 = op_4;
assign ret_V_2_fu_239_p4 = op_8[15:10];
assign rhs_1_fu_302_p3 = { op_21_V_reg_950, 11'h000 };
assign rhs_5_fu_867_p3 = { op_30_V_reg_1227, 3'h0 };
assign sext_ln1116_fu_620_p1 = { op_6_V_fu_614_p3[3], op_6_V_fu_614_p3 };
assign sext_ln1192_fu_298_p0 = op_10;
assign sext_ln1196_fu_435_p0 = op_2;
assign sext_ln1196_fu_435_p1 = { op_2[1], op_2 };
assign sext_ln1496_fu_726_p1 = { op_2[1], op_2, 1'h0 };
assign sext_ln1498_fu_743_p1 = { op_5[3], op_5 };
assign sext_ln69_3_fu_841_p1 = { op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17 };
assign sext_ln69_fu_288_p1 = { op_9[3], op_9[3], op_9[3], op_9 };
assign sext_ln703_1_fu_791_p0 = op_4;
assign sext_ln703_1_fu_791_p1 = { op_4[7], op_4 };
assign sext_ln703_2_fu_589_p0 = op_11;
assign sext_ln703_3_fu_863_p0 = op_19;
assign sext_ln703_fu_339_p0 = op_2;
assign sext_ln703_fu_339_p1 = { op_2[1], op_2[1], op_2[1], op_2[1], op_2[1], op_2[1], op_2 };
assign sext_ln831_fu_249_p1 = { op_8[15], op_8[15:10] };
assign sext_ln850_fu_375_p1 = { tmp_reg_975[21], tmp_reg_975 };
assign shl_ln728_1_fu_736_p1 = op_2;
assign shl_ln728_1_fu_736_p3 = { op_2, 3'h0 };
assign shl_ln_fu_719_p1 = op_2;
assign shl_ln_fu_719_p3 = { op_2, 1'h0 };
assign tmp_10_fu_593_p3 = { select_ln353_reg_1063, 1'h0 };
assign tmp_4_fu_477_p3 = xor_ln1196_1_fu_438_p2[2];
assign tmp_5_fu_485_p3 = xor_ln731_reg_1039[1];
assign trunc_ln1196_1_fu_347_p0 = op_4;
assign trunc_ln1196_1_fu_347_p1 = op_4[2:0];
assign trunc_ln1196_fu_343_p0 = op_4;
assign trunc_ln1196_fu_343_p1 = op_4[1:0];
assign trunc_ln851_1_fu_657_p1 = r_V_fu_640_p3[1:0];
assign trunc_ln851_2_fu_319_p0 = op_10;
assign trunc_ln851_2_fu_319_p1 = op_10[10:0];
assign trunc_ln851_3_fu_703_p0 = op_11;
assign trunc_ln851_3_fu_703_p1 = op_11[0];
assign trunc_ln851_4_fu_884_p0 = op_19;
assign trunc_ln851_4_fu_884_p1 = op_19[2:0];
assign trunc_ln851_fu_253_p1 = op_8[9:0];
assign xor_ln731_fu_394_p1 = op_2;
assign zext_ln69_1_fu_845_p1 = { 2'h0, op_18 };
assign zext_ln69_fu_766_p1 = { 1'h0, xor_ln1496_fu_761_p2 };
assign \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.ain_s0  = \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.a ;
assign \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.bin_s0  = \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.b ;
assign \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.s  = { \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.fas_s2 , \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.sum_s1  };
assign \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.u2.a  = \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.ain_s1 ;
assign \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.u2.b  = \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.bin_s1 ;
assign \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.u2.cin  = \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.carry_s1 ;
assign \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.facout_s2  = \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.u2.cout ;
assign \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.fas_s2  = \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.u2.s ;
assign \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.u1.a  = \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.a [17:0];
assign \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.u1.b  = \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.b [17:0];
assign \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.u1.cin  = 1'h0;
assign \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.facout_s1  = \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.u1.cout ;
assign \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.fas_s1  = \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.u1.s ;
assign \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.a  = \add_36s_36s_36_2_1_U9.din0 ;
assign \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.b  = \add_36s_36s_36_2_1_U9.din1 ;
assign \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.ce  = \add_36s_36s_36_2_1_U9.ce ;
assign \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.clk  = \add_36s_36s_36_2_1_U9.clk ;
assign \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.reset  = \add_36s_36s_36_2_1_U9.reset ;
assign \add_36s_36s_36_2_1_U9.dout  = \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.s ;
assign \add_36s_36s_36_2_1_U9.ce  = 1'h1;
assign \add_36s_36s_36_2_1_U9.clk  = ap_clk;
assign \add_36s_36s_36_2_1_U9.din0  = { op_30_V_reg_1227[31], op_30_V_reg_1227, 3'h0 };
assign \add_36s_36s_36_2_1_U9.din1  = { op_19[7], op_19[7], op_19[7], op_19[7], op_19[7], op_19[7], op_19[7], op_19[7], op_19[7], op_19[7], op_19[7], op_19[7], op_19[7], op_19[7], op_19[7], op_19[7], op_19[7], op_19[7], op_19[7], op_19[7], op_19[7], op_19[7], op_19[7], op_19[7], op_19[7], op_19[7], op_19[7], op_19[7], op_19 };
assign grp_fu_878_p2 = \add_36s_36s_36_2_1_U9.dout ;
assign \add_36s_36s_36_2_1_U9.reset  = ap_rst;
assign \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.ain_s0  = \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.a ;
assign \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.bin_s0  = \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.b ;
assign \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.s  = { \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.fas_s2 , \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.sum_s1  };
assign \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.u2.a  = \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.ain_s1 ;
assign \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.u2.b  = \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.bin_s1 ;
assign \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.u2.cin  = \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.carry_s1 ;
assign \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.facout_s2  = \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.u2.cout ;
assign \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.fas_s2  = \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.u2.s ;
assign \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.u1.a  = \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.a [16:0];
assign \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.u1.b  = \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.b [16:0];
assign \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.u1.cin  = 1'h0;
assign \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.facout_s1  = \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.u1.cout ;
assign \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.fas_s1  = \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.u1.s ;
assign \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.a  = \add_34s_34s_34_2_1_U3.din0 ;
assign \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.b  = \add_34s_34s_34_2_1_U3.din1 ;
assign \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.ce  = \add_34s_34s_34_2_1_U3.ce ;
assign \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.clk  = \add_34s_34s_34_2_1_U3.clk ;
assign \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.reset  = \add_34s_34s_34_2_1_U3.reset ;
assign \add_34s_34s_34_2_1_U3.dout  = \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.s ;
assign \add_34s_34s_34_2_1_U3.ce  = 1'h1;
assign \add_34s_34s_34_2_1_U3.clk  = ap_clk;
assign \add_34s_34s_34_2_1_U3.din0  = { select_ln353_reg_1063[22], select_ln353_reg_1063[22], select_ln353_reg_1063[22], select_ln353_reg_1063[22], select_ln353_reg_1063[22], select_ln353_reg_1063[22], select_ln353_reg_1063[22], select_ln353_reg_1063[22], select_ln353_reg_1063[22], select_ln353_reg_1063[22], select_ln353_reg_1063, 1'h0 };
assign \add_34s_34s_34_2_1_U3.din1  = { op_11[1], op_11[1], op_11[1], op_11[1], op_11[1], op_11[1], op_11[1], op_11[1], op_11[1], op_11[1], op_11[1], op_11[1], op_11[1], op_11[1], op_11[1], op_11[1], op_11[1], op_11[1], op_11[1], op_11[1], op_11[1], op_11[1], op_11[1], op_11[1], op_11[1], op_11[1], op_11[1], op_11[1], op_11[1], op_11[1], op_11[1], op_11[1], op_11 };
assign grp_fu_604_p2 = \add_34s_34s_34_2_1_U3.dout ;
assign \add_34s_34s_34_2_1_U3.reset  = ap_rst;
assign \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.ain_s0  = \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.a ;
assign \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.bin_s0  = \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.b ;
assign \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.s  = { \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.fas_s2 , \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.sum_s1  };
assign \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.u2.a  = \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.ain_s1 ;
assign \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.u2.b  = \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.bin_s1 ;
assign \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.u2.cin  = \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.carry_s1 ;
assign \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.facout_s2  = \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.u2.cout ;
assign \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.fas_s2  = \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.u2.s ;
assign \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.u1.a  = \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.a [15:0];
assign \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.u1.b  = \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.b [15:0];
assign \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.u1.cin  = 1'h0;
assign \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.facout_s1  = \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.u1.cout ;
assign \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.fas_s1  = \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.u1.s ;
assign \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.a  = \add_33s_33s_33_2_1_U1.din0 ;
assign \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.b  = \add_33s_33s_33_2_1_U1.din1 ;
assign \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.ce  = \add_33s_33s_33_2_1_U1.ce ;
assign \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.clk  = \add_33s_33s_33_2_1_U1.clk ;
assign \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.reset  = \add_33s_33s_33_2_1_U1.reset ;
assign \add_33s_33s_33_2_1_U1.dout  = \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.s ;
assign \add_33s_33s_33_2_1_U1.ce  = 1'h1;
assign \add_33s_33s_33_2_1_U1.clk  = ap_clk;
assign \add_33s_33s_33_2_1_U1.din0  = { op_21_V_reg_950[6], op_21_V_reg_950[6], op_21_V_reg_950[6], op_21_V_reg_950[6], op_21_V_reg_950[6], op_21_V_reg_950[6], op_21_V_reg_950[6], op_21_V_reg_950[6], op_21_V_reg_950[6], op_21_V_reg_950[6], op_21_V_reg_950[6], op_21_V_reg_950[6], op_21_V_reg_950[6], op_21_V_reg_950[6], op_21_V_reg_950[6], op_21_V_reg_950, 11'h000 };
assign \add_33s_33s_33_2_1_U1.din1  = { op_10[31], op_10 };
assign grp_fu_313_p2 = \add_33s_33s_33_2_1_U1.dout ;
assign \add_33s_33s_33_2_1_U1.reset  = ap_rst;
assign \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.ain_s0  = \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.a ;
assign \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.bin_s0  = \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.b ;
assign \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.s  = { \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.fas_s2 , \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.sum_s1  };
assign \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.u2.a  = \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.ain_s1 ;
assign \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.u2.b  = \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.bin_s1 ;
assign \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.u2.cin  = \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.carry_s1 ;
assign \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.facout_s2  = \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.u2.cout ;
assign \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.fas_s2  = \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.u2.s ;
assign \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.u1.a  = \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.a [15:0];
assign \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.u1.b  = \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.b [15:0];
assign \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.u1.cin  = 1'h0;
assign \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.facout_s1  = \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.u1.cout ;
assign \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.fas_s1  = \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.u1.s ;
assign \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.a  = \add_33ns_33s_33_2_1_U7.din0 ;
assign \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.b  = \add_33ns_33s_33_2_1_U7.din1 ;
assign \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.ce  = \add_33ns_33s_33_2_1_U7.ce ;
assign \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.clk  = \add_33ns_33s_33_2_1_U7.clk ;
assign \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.reset  = \add_33ns_33s_33_2_1_U7.reset ;
assign \add_33ns_33s_33_2_1_U7.dout  = \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.s ;
assign \add_33ns_33s_33_2_1_U7.ce  = 1'h1;
assign \add_33ns_33s_33_2_1_U7.clk  = ap_clk;
assign \add_33ns_33s_33_2_1_U7.din0  = { op_27_V_reg_1197, 1'h0 };
assign \add_33ns_33s_33_2_1_U7.din1  = { ret_V_reg_1192[8], ret_V_reg_1192[8], ret_V_reg_1192[8], ret_V_reg_1192[8], ret_V_reg_1192[8], ret_V_reg_1192[8], ret_V_reg_1192[8], ret_V_reg_1192[8], ret_V_reg_1192[8], ret_V_reg_1192[8], ret_V_reg_1192[8], ret_V_reg_1192[8], ret_V_reg_1192[8], ret_V_reg_1192[8], ret_V_reg_1192[8], ret_V_reg_1192[8], ret_V_reg_1192[8], ret_V_reg_1192[8], ret_V_reg_1192[8], ret_V_reg_1192[8], ret_V_reg_1192[8], ret_V_reg_1192[8], ret_V_reg_1192[8], ret_V_reg_1192, 1'h0 };
assign grp_fu_825_p2 = \add_33ns_33s_33_2_1_U7.dout ;
assign \add_33ns_33s_33_2_1_U7.reset  = ap_rst;
assign \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.ain_s0  = \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.a ;
assign \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.bin_s0  = \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.b ;
assign \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.s  = { \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.fas_s2 , \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.sum_s1  };
assign \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.u2.a  = \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.ain_s1 ;
assign \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.u2.b  = \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.bin_s1 ;
assign \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.u2.cin  = \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.carry_s1 ;
assign \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.facout_s2  = \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.u2.cout ;
assign \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.fas_s2  = \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.u2.s ;
assign \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.u1.a  = \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.a [15:0];
assign \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.u1.b  = \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.b [15:0];
assign \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.u1.cin  = 1'h0;
assign \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.facout_s1  = \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.u1.cout ;
assign \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.fas_s1  = \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.u1.s ;
assign \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.a  = \add_32s_32ns_32_2_1_U8.din0 ;
assign \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.b  = \add_32s_32ns_32_2_1_U8.din1 ;
assign \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.ce  = \add_32s_32ns_32_2_1_U8.ce ;
assign \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.clk  = \add_32s_32ns_32_2_1_U8.clk ;
assign \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.reset  = \add_32s_32ns_32_2_1_U8.reset ;
assign \add_32s_32ns_32_2_1_U8.dout  = \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.s ;
assign \add_32s_32ns_32_2_1_U8.ce  = 1'h1;
assign \add_32s_32ns_32_2_1_U8.clk  = ap_clk;
assign \add_32s_32ns_32_2_1_U8.din0  = { add_ln69_3_reg_1217[9], add_ln69_3_reg_1217[9], add_ln69_3_reg_1217[9], add_ln69_3_reg_1217[9], add_ln69_3_reg_1217[9], add_ln69_3_reg_1217[9], add_ln69_3_reg_1217[9], add_ln69_3_reg_1217[9], add_ln69_3_reg_1217[9], add_ln69_3_reg_1217[9], add_ln69_3_reg_1217[9], add_ln69_3_reg_1217[9], add_ln69_3_reg_1217[9], add_ln69_3_reg_1217[9], add_ln69_3_reg_1217[9], add_ln69_3_reg_1217[9], add_ln69_3_reg_1217[9], add_ln69_3_reg_1217[9], add_ln69_3_reg_1217[9], add_ln69_3_reg_1217[9], add_ln69_3_reg_1217[9], add_ln69_3_reg_1217[9], add_ln69_3_reg_1217 };
assign \add_32s_32ns_32_2_1_U8.din1  = op_28_V_reg_1212;
assign grp_fu_858_p2 = \add_32s_32ns_32_2_1_U8.dout ;
assign \add_32s_32ns_32_2_1_U8.reset  = ap_rst;
assign \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.ain_s0  = \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.a ;
assign \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.bin_s0  = \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.b ;
assign \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.s  = { \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.fas_s2 , \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.sum_s1  };
assign \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.u2.a  = \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.ain_s1 ;
assign \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.u2.b  = \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.bin_s1 ;
assign \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.u2.cin  = \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.carry_s1 ;
assign \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.facout_s2  = \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.u2.cout ;
assign \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.fas_s2  = \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.u2.s ;
assign \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.u1.a  = \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.a [15:0];
assign \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.u1.b  = \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.b [15:0];
assign \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.u1.cin  = 1'h0;
assign \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.facout_s1  = \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.u1.cout ;
assign \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.fas_s1  = \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.u1.s ;
assign \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.a  = \add_32s_32ns_32_2_1_U6.din0 ;
assign \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.b  = \add_32s_32ns_32_2_1_U6.din1 ;
assign \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.ce  = \add_32s_32ns_32_2_1_U6.ce ;
assign \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.clk  = \add_32s_32ns_32_2_1_U6.clk ;
assign \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.reset  = \add_32s_32ns_32_2_1_U6.reset ;
assign \add_32s_32ns_32_2_1_U6.dout  = \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.s ;
assign \add_32s_32ns_32_2_1_U6.ce  = 1'h1;
assign \add_32s_32ns_32_2_1_U6.clk  = ap_clk;
assign \add_32s_32ns_32_2_1_U6.din0  = { add_ln69_1_reg_1182[1], add_ln69_1_reg_1182[1], add_ln69_1_reg_1182[1], add_ln69_1_reg_1182[1], add_ln69_1_reg_1182[1], add_ln69_1_reg_1182[1], add_ln69_1_reg_1182[1], add_ln69_1_reg_1182[1], add_ln69_1_reg_1182[1], add_ln69_1_reg_1182[1], add_ln69_1_reg_1182[1], add_ln69_1_reg_1182[1], add_ln69_1_reg_1182[1], add_ln69_1_reg_1182[1], add_ln69_1_reg_1182[1], add_ln69_1_reg_1182[1], add_ln69_1_reg_1182[1], add_ln69_1_reg_1182[1], add_ln69_1_reg_1182[1], add_ln69_1_reg_1182[1], add_ln69_1_reg_1182[1], add_ln69_1_reg_1182[1], add_ln69_1_reg_1182[1], add_ln69_1_reg_1182[1], add_ln69_1_reg_1182[1], add_ln69_1_reg_1182[1], add_ln69_1_reg_1182[1], add_ln69_1_reg_1182[1], add_ln69_1_reg_1182[1], add_ln69_1_reg_1182[1], add_ln69_1_reg_1182 };
assign \add_32s_32ns_32_2_1_U6.din1  = add_ln69_reg_1177;
assign grp_fu_786_p2 = \add_32s_32ns_32_2_1_U6.dout ;
assign \add_32s_32ns_32_2_1_U6.reset  = ap_rst;
assign \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.ain_s0  = \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.a ;
assign \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.bin_s0  = \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.b ;
assign \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.s  = { \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.fas_s2 , \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.sum_s1  };
assign \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.u2.a  = \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.ain_s1 ;
assign \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.u2.b  = \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.bin_s1 ;
assign \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.u2.cin  = \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.carry_s1 ;
assign \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.facout_s2  = \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.u2.cout ;
assign \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.fas_s2  = \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.u2.s ;
assign \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.u1.a  = \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.a [15:0];
assign \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.u1.b  = \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.b [15:0];
assign \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.u1.cin  = 1'h0;
assign \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.facout_s1  = \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.u1.cout ;
assign \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.fas_s1  = \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.u1.s ;
assign \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.a  = \add_32ns_32s_32_2_1_U5.din0 ;
assign \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.b  = \add_32ns_32s_32_2_1_U5.din1 ;
assign \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.ce  = \add_32ns_32s_32_2_1_U5.ce ;
assign \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.clk  = \add_32ns_32s_32_2_1_U5.clk ;
assign \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.reset  = \add_32ns_32s_32_2_1_U5.reset ;
assign \add_32ns_32s_32_2_1_U5.dout  = \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.s ;
assign \add_32ns_32s_32_2_1_U5.ce  = 1'h1;
assign \add_32ns_32s_32_2_1_U5.clk  = ap_clk;
assign \add_32ns_32s_32_2_1_U5.din0  = ret_V_18_reg_1157;
assign \add_32ns_32s_32_2_1_U5.din1  = { ret_V_7_reg_1152[2], ret_V_7_reg_1152[2], ret_V_7_reg_1152[2], ret_V_7_reg_1152[2], ret_V_7_reg_1152[2], ret_V_7_reg_1152[2], ret_V_7_reg_1152[2], ret_V_7_reg_1152[2], ret_V_7_reg_1152[2], ret_V_7_reg_1152[2], ret_V_7_reg_1152[2], ret_V_7_reg_1152[2], ret_V_7_reg_1152[2], ret_V_7_reg_1152[2], ret_V_7_reg_1152[2], ret_V_7_reg_1152[2], ret_V_7_reg_1152[2], ret_V_7_reg_1152[2], ret_V_7_reg_1152[2], ret_V_7_reg_1152[2], ret_V_7_reg_1152[2], ret_V_7_reg_1152[2], ret_V_7_reg_1152[2], ret_V_7_reg_1152[2], ret_V_7_reg_1152[2], ret_V_7_reg_1152[2], ret_V_7_reg_1152[2], ret_V_7_reg_1152[2], ret_V_7_reg_1152[2], ret_V_7_reg_1152 };
assign grp_fu_756_p2 = \add_32ns_32s_32_2_1_U5.dout ;
assign \add_32ns_32s_32_2_1_U5.reset  = ap_rst;
assign \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.ain_s0  = \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.a ;
assign \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.bin_s0  = \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.b ;
assign \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.s  = { \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.fas_s2 , \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.sum_s1  };
assign \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.u2.a  = \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.ain_s1 ;
assign \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.u2.b  = \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.bin_s1 ;
assign \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.u2.cin  = \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.carry_s1 ;
assign \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.facout_s2  = \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.u2.cout ;
assign \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.fas_s2  = \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.u2.s ;
assign \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.u1.a  = \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.a [15:0];
assign \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.u1.b  = \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.b [15:0];
assign \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.u1.cin  = 1'h0;
assign \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.facout_s1  = \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.u1.cout ;
assign \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.fas_s1  = \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.u1.s ;
assign \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.a  = \add_32ns_32ns_32_2_1_U4.din0 ;
assign \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.b  = \add_32ns_32ns_32_2_1_U4.din1 ;
assign \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.ce  = \add_32ns_32ns_32_2_1_U4.ce ;
assign \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.clk  = \add_32ns_32ns_32_2_1_U4.clk ;
assign \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.reset  = \add_32ns_32ns_32_2_1_U4.reset ;
assign \add_32ns_32ns_32_2_1_U4.dout  = \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.s ;
assign \add_32ns_32ns_32_2_1_U4.ce  = 1'h1;
assign \add_32ns_32ns_32_2_1_U4.clk  = ap_clk;
assign \add_32ns_32ns_32_2_1_U4.din0  = ret_V_12_cast_reg_1113;
assign \add_32ns_32ns_32_2_1_U4.din1  = 32'd1;
assign grp_fu_667_p2 = \add_32ns_32ns_32_2_1_U4.dout ;
assign \add_32ns_32ns_32_2_1_U4.reset  = ap_rst;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.ain_s0  = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.a ;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.bin_s0  = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.b ;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.s  = { \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.fas_s2 , \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.sum_s1  };
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.u2.a  = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.ain_s1 ;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.u2.b  = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.bin_s1 ;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.u2.cin  = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.carry_s1 ;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.facout_s2  = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.u2.cout ;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.fas_s2  = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.u2.s ;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.u1.a  = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.a [15:0];
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.u1.b  = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.b [15:0];
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.u1.cin  = 1'h0;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.facout_s1  = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.u1.cout ;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.fas_s1  = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.u1.s ;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.a  = \add_32ns_32ns_32_2_1_U10.din0 ;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.b  = \add_32ns_32ns_32_2_1_U10.din1 ;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.ce  = \add_32ns_32ns_32_2_1_U10.ce ;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.clk  = \add_32ns_32ns_32_2_1_U10.clk ;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.reset  = \add_32ns_32ns_32_2_1_U10.reset ;
assign \add_32ns_32ns_32_2_1_U10.dout  = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.s ;
assign \add_32ns_32ns_32_2_1_U10.ce  = 1'h1;
assign \add_32ns_32ns_32_2_1_U10.clk  = ap_clk;
assign \add_32ns_32ns_32_2_1_U10.din0  = ret_V_16_cast_reg_1252;
assign \add_32ns_32ns_32_2_1_U10.din1  = 32'd1;
assign grp_fu_904_p2 = \add_32ns_32ns_32_2_1_U10.dout ;
assign \add_32ns_32ns_32_2_1_U10.reset  = ap_rst;
assign \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.ain_s0  = \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.a ;
assign \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.bin_s0  = \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.b ;
assign \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.s  = { \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.fas_s2 , \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.sum_s1  };
assign \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.u2.a  = \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.ain_s1 ;
assign \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.u2.b  = \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.bin_s1 ;
assign \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.u2.cin  = \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.carry_s1 ;
assign \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.facout_s2  = \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.u2.cout ;
assign \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.fas_s2  = \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.u2.s ;
assign \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.u1.a  = \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.a [10:0];
assign \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.u1.b  = \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.b [10:0];
assign \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.u1.cin  = 1'h0;
assign \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.facout_s1  = \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.u1.cout ;
assign \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.fas_s1  = \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.u1.s ;
assign \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.a  = \add_23s_23ns_23_2_1_U2.din0 ;
assign \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.b  = \add_23s_23ns_23_2_1_U2.din1 ;
assign \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.ce  = \add_23s_23ns_23_2_1_U2.ce ;
assign \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.clk  = \add_23s_23ns_23_2_1_U2.clk ;
assign \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.reset  = \add_23s_23ns_23_2_1_U2.reset ;
assign \add_23s_23ns_23_2_1_U2.dout  = \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.s ;
assign \add_23s_23ns_23_2_1_U2.ce  = 1'h1;
assign \add_23s_23ns_23_2_1_U2.clk  = ap_clk;
assign \add_23s_23ns_23_2_1_U2.din0  = { tmp_reg_975[21], tmp_reg_975 };
assign \add_23s_23ns_23_2_1_U2.din1  = 23'h000001;
assign grp_fu_378_p2 = \add_23s_23ns_23_2_1_U2.dout ;
assign \add_23s_23ns_23_2_1_U2.reset  = ap_rst;
endmodule


// Machine B:
// Processed by function `add_clk_enable_signal` in `verilog_tricks.py`.
// Processed by function `remove_reset_signal` in `verilog_tricks.py`.
module top_B (
  ap_clk,
  ap_start,
  ap_done,
  ap_idle,
  ap_ready,
  op_0,
  op_2,
  op_3,
  op_4,
  op_5,
  op_7,
  op_8,
  op_9,
  op_10,
  op_11,
  op_17,
  op_18,
  op_19,
  op_31,
  op_31_ap_vld,
clk_enable
);
input clk_enable;


input ap_clk;
wire ap_rst;
assign ap_rst = op_31_ap_vld;
input ap_start;
input [1:0] op_0;
input [31:0] op_10;
input [1:0] op_11;
input [3:0] op_17;
input [7:0] op_18;
input [7:0] op_19;
input [1:0] op_2;
input [3:0] op_3;
input [7:0] op_4;
input [3:0] op_5;
input op_7;
input [15:0] op_8;
input [3:0] op_9;
output ap_done;
output ap_idle;
output ap_ready;
output [31:0] op_31;
output op_31_ap_vld;


reg [11:0] \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.ain_s1 ;
reg [11:0] \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.bin_s1 ;
reg \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.carry_s1 ;
reg [10:0] \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.sum_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.ain_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.bin_s1 ;
reg \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.carry_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.sum_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.ain_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.bin_s1 ;
reg \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.carry_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.sum_s1 ;
reg [15:0] \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.ain_s1 ;
reg [15:0] \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.bin_s1 ;
reg \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.carry_s1 ;
reg [15:0] \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.sum_s1 ;
reg [15:0] \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.ain_s1 ;
reg [15:0] \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.bin_s1 ;
reg \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.carry_s1 ;
reg [15:0] \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.sum_s1 ;
reg [15:0] \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.ain_s1 ;
reg [15:0] \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.bin_s1 ;
reg \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.carry_s1 ;
reg [15:0] \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.sum_s1 ;
reg [16:0] \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.ain_s1 ;
reg [16:0] \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.bin_s1 ;
reg \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.carry_s1 ;
reg [15:0] \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.sum_s1 ;
reg [16:0] \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.ain_s1 ;
reg [16:0] \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.bin_s1 ;
reg \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.carry_s1 ;
reg [15:0] \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.sum_s1 ;
reg [16:0] \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.ain_s1 ;
reg [16:0] \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.bin_s1 ;
reg \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.carry_s1 ;
reg [16:0] \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.sum_s1 ;
reg [17:0] \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.ain_s1 ;
reg [17:0] \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.bin_s1 ;
reg \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.carry_s1 ;
reg [17:0] \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.sum_s1 ;
reg [31:0] add_ln691_1_reg_1147;
reg [31:0] add_ln691_4_reg_1259;
reg [22:0] add_ln691_reg_1034;
reg [1:0] add_ln69_1_reg_1182;
reg [9:0] add_ln69_3_reg_1217;
reg [31:0] add_ln69_reg_1177;
reg and_ln785_reg_1078;
reg [24:0] ap_CS_fsm = 25'h0000001;
reg icmp_ln1496_reg_1162;
reg icmp_ln768_reg_1023;
reg icmp_ln786_reg_1028;
reg icmp_ln851_1_reg_1137;
reg icmp_ln851_2_reg_965;
reg icmp_ln851_3_reg_1242;
reg icmp_ln851_reg_940;
reg [3:0] newSel22_reg_1088;
reg op_15_V_reg_1167;
reg [6:0] op_21_V_reg_950;
reg [31:0] op_27_V_reg_1197;
reg [31:0] op_28_V_reg_1212;
reg [31:0] op_30_V_reg_1227;
reg or_ln785_reg_1051;
reg p_Result_6_reg_1003;
reg p_Result_7_reg_1045;
reg [5:0] p_Result_s_reg_1010;
reg [3:0] p_Val2_1_reg_1073;
reg [4:0] r_V_reg_1125;
reg [31:0] ret_V_12_cast_reg_1113;
reg [31:0] ret_V_16_cast_reg_1252;
reg [32:0] ret_V_16_reg_970;
reg [33:0] ret_V_17_reg_1108;
reg [31:0] ret_V_18_reg_1157;
reg [35:0] ret_V_19_reg_1247;
reg [6:0] ret_V_3_reg_945;
reg [2:0] ret_V_5_reg_1130;
reg [2:0] ret_V_6_reg_1142;
reg [2:0] ret_V_7_reg_1152;
reg [8:0] ret_V_reg_1192;
reg sel_tmp11_reg_1083;
reg [22:0] select_ln353_reg_1063;
reg [6:0] sext_ln831_reg_934;
reg [22:0] sext_ln850_reg_1016;
reg [4:0] sub_ln1118_reg_1103;
reg [21:0] tmp_reg_975;
reg [2:0] trunc_ln1196_1_reg_998;
reg [1:0] trunc_ln1196_reg_993;
reg [1:0] xor_ln731_reg_1039;
reg xor_ln785_reg_1057;
wire [31:0] _000_;
wire [31:0] _001_;
wire [22:0] _002_;
wire [1:0] _003_;
wire [9:0] _004_;
wire [31:0] _005_;
wire _006_;
wire [24:0] _007_;
wire _008_;
wire _009_;
wire _010_;
wire _011_;
wire _012_;
wire _013_;
wire _014_;
wire [3:0] _015_;
wire _016_;
wire [6:0] _017_;
wire [31:0] _018_;
wire [31:0] _019_;
wire [31:0] _020_;
wire _021_;
wire _022_;
wire _023_;
wire [5:0] _024_;
wire [1:0] _025_;
wire [4:0] _026_;
wire [31:0] _027_;
wire [31:0] _028_;
wire [32:0] _029_;
wire [33:0] _030_;
wire [31:0] _031_;
wire [35:0] _032_;
wire [6:0] _033_;
wire [2:0] _034_;
wire [2:0] _035_;
wire [2:0] _036_;
wire [8:0] _037_;
wire _038_;
wire [22:0] _039_;
wire [6:0] _040_;
wire [22:0] _041_;
wire [4:0] _042_;
wire [21:0] _043_;
wire [2:0] _044_;
wire [1:0] _045_;
wire [1:0] _046_;
wire _047_;
wire [1:0] _048_;
wire _049_;
wire _050_;
wire _051_;
wire _052_;
wire _053_;
wire _054_;
wire _055_;
wire _056_;
wire _057_;
wire _058_;
wire [11:0] _059_;
wire [11:0] _060_;
wire _061_;
wire [10:0] _062_;
wire [11:0] _063_;
wire [12:0] _064_;
wire [15:0] _065_;
wire [15:0] _066_;
wire _067_;
wire [15:0] _068_;
wire [16:0] _069_;
wire [16:0] _070_;
wire [15:0] _071_;
wire [15:0] _072_;
wire _073_;
wire [15:0] _074_;
wire [16:0] _075_;
wire [16:0] _076_;
wire [15:0] _077_;
wire [15:0] _078_;
wire _079_;
wire [15:0] _080_;
wire [16:0] _081_;
wire [16:0] _082_;
wire [15:0] _083_;
wire [15:0] _084_;
wire _085_;
wire [15:0] _086_;
wire [16:0] _087_;
wire [16:0] _088_;
wire [15:0] _089_;
wire [15:0] _090_;
wire _091_;
wire [15:0] _092_;
wire [16:0] _093_;
wire [16:0] _094_;
wire [16:0] _095_;
wire [16:0] _096_;
wire _097_;
wire [15:0] _098_;
wire [16:0] _099_;
wire [17:0] _100_;
wire [16:0] _101_;
wire [16:0] _102_;
wire _103_;
wire [15:0] _104_;
wire [16:0] _105_;
wire [17:0] _106_;
wire [16:0] _107_;
wire [16:0] _108_;
wire _109_;
wire [16:0] _110_;
wire [17:0] _111_;
wire [17:0] _112_;
wire [17:0] _113_;
wire [17:0] _114_;
wire _115_;
wire [17:0] _116_;
wire [18:0] _117_;
wire [18:0] _118_;
wire _119_;
wire _120_;
wire _121_;
wire _122_;
wire _123_;
wire _124_;
wire _125_;
wire _126_;
wire _127_;
wire _128_;
wire _129_;
wire _130_;
wire _131_;
wire _132_;
wire _133_;
wire _134_;
wire _135_;
wire _136_;
wire _137_;
wire _138_;
wire _139_;
wire _140_;
wire _141_;
wire _142_;
wire _143_;
wire _144_;
wire _145_;
wire _146_;
wire _147_;
wire _148_;
wire \add_23s_23ns_23_2_1_U2.ce ;
wire \add_23s_23ns_23_2_1_U2.clk ;
wire [22:0] \add_23s_23ns_23_2_1_U2.din0 ;
wire [22:0] \add_23s_23ns_23_2_1_U2.din1 ;
wire [22:0] \add_23s_23ns_23_2_1_U2.dout ;
wire \add_23s_23ns_23_2_1_U2.reset ;
wire [22:0] \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.a ;
wire [22:0] \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.ain_s0 ;
wire [22:0] \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.b ;
wire [22:0] \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.bin_s0 ;
wire \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.ce ;
wire \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.clk ;
wire \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.facout_s1 ;
wire \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.facout_s2 ;
wire [10:0] \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.fas_s1 ;
wire [11:0] \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.fas_s2 ;
wire \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.reset ;
wire [22:0] \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.s ;
wire [10:0] \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.u1.a ;
wire [10:0] \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.u1.b ;
wire \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.u1.cin ;
wire \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.u1.cout ;
wire [10:0] \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.u1.s ;
wire [11:0] \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.u2.a ;
wire [11:0] \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.u2.b ;
wire \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.u2.cin ;
wire \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.u2.cout ;
wire [11:0] \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.u2.s ;
wire \add_32ns_32ns_32_2_1_U10.ce ;
wire \add_32ns_32ns_32_2_1_U10.clk ;
wire [31:0] \add_32ns_32ns_32_2_1_U10.din0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U10.din1 ;
wire [31:0] \add_32ns_32ns_32_2_1_U10.dout ;
wire \add_32ns_32ns_32_2_1_U10.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.a ;
wire [31:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.ain_s0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.b ;
wire [31:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.bin_s0 ;
wire \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.ce ;
wire \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.clk ;
wire \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.facout_s1 ;
wire \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.facout_s2 ;
wire [15:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.fas_s1 ;
wire [15:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.fas_s2 ;
wire \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.u1.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.u1.b ;
wire \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.u1.cin ;
wire \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.u1.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.u1.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.u2.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.u2.b ;
wire \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.u2.cin ;
wire \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.u2.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.u2.s ;
wire \add_32ns_32ns_32_2_1_U4.ce ;
wire \add_32ns_32ns_32_2_1_U4.clk ;
wire [31:0] \add_32ns_32ns_32_2_1_U4.din0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U4.din1 ;
wire [31:0] \add_32ns_32ns_32_2_1_U4.dout ;
wire \add_32ns_32ns_32_2_1_U4.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.a ;
wire [31:0] \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.ain_s0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.b ;
wire [31:0] \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.bin_s0 ;
wire \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.ce ;
wire \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.clk ;
wire \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.facout_s1 ;
wire \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.facout_s2 ;
wire [15:0] \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.fas_s1 ;
wire [15:0] \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.fas_s2 ;
wire \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.u1.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.u1.b ;
wire \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.u1.cin ;
wire \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.u1.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.u1.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.u2.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.u2.b ;
wire \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.u2.cin ;
wire \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.u2.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.u2.s ;
wire \add_32ns_32s_32_2_1_U5.ce ;
wire \add_32ns_32s_32_2_1_U5.clk ;
wire [31:0] \add_32ns_32s_32_2_1_U5.din0 ;
wire [31:0] \add_32ns_32s_32_2_1_U5.din1 ;
wire [31:0] \add_32ns_32s_32_2_1_U5.dout ;
wire \add_32ns_32s_32_2_1_U5.reset ;
wire [31:0] \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.a ;
wire [31:0] \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.ain_s0 ;
wire [31:0] \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.b ;
wire [31:0] \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.bin_s0 ;
wire \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.ce ;
wire \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.clk ;
wire \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.facout_s1 ;
wire \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.facout_s2 ;
wire [15:0] \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.fas_s1 ;
wire [15:0] \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.fas_s2 ;
wire \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.reset ;
wire [31:0] \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.s ;
wire [15:0] \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.u1.a ;
wire [15:0] \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.u1.b ;
wire \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.u1.cin ;
wire \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.u1.cout ;
wire [15:0] \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.u1.s ;
wire [15:0] \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.u2.a ;
wire [15:0] \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.u2.b ;
wire \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.u2.cin ;
wire \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.u2.cout ;
wire [15:0] \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.u2.s ;
wire \add_32s_32ns_32_2_1_U6.ce ;
wire \add_32s_32ns_32_2_1_U6.clk ;
wire [31:0] \add_32s_32ns_32_2_1_U6.din0 ;
wire [31:0] \add_32s_32ns_32_2_1_U6.din1 ;
wire [31:0] \add_32s_32ns_32_2_1_U6.dout ;
wire \add_32s_32ns_32_2_1_U6.reset ;
wire [31:0] \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.a ;
wire [31:0] \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.ain_s0 ;
wire [31:0] \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.b ;
wire [31:0] \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.bin_s0 ;
wire \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.ce ;
wire \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.clk ;
wire \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.facout_s1 ;
wire \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.facout_s2 ;
wire [15:0] \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.fas_s1 ;
wire [15:0] \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.fas_s2 ;
wire \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.reset ;
wire [31:0] \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.s ;
wire [15:0] \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.u1.a ;
wire [15:0] \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.u1.b ;
wire \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.u1.cin ;
wire \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.u1.cout ;
wire [15:0] \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.u1.s ;
wire [15:0] \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.u2.a ;
wire [15:0] \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.u2.b ;
wire \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.u2.cin ;
wire \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.u2.cout ;
wire [15:0] \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.u2.s ;
wire \add_32s_32ns_32_2_1_U8.ce ;
wire \add_32s_32ns_32_2_1_U8.clk ;
wire [31:0] \add_32s_32ns_32_2_1_U8.din0 ;
wire [31:0] \add_32s_32ns_32_2_1_U8.din1 ;
wire [31:0] \add_32s_32ns_32_2_1_U8.dout ;
wire \add_32s_32ns_32_2_1_U8.reset ;
wire [31:0] \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.a ;
wire [31:0] \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.ain_s0 ;
wire [31:0] \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.b ;
wire [31:0] \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.bin_s0 ;
wire \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.ce ;
wire \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.clk ;
wire \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.facout_s1 ;
wire \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.facout_s2 ;
wire [15:0] \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.fas_s1 ;
wire [15:0] \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.fas_s2 ;
wire \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.reset ;
wire [31:0] \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.s ;
wire [15:0] \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.u1.a ;
wire [15:0] \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.u1.b ;
wire \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.u1.cin ;
wire \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.u1.cout ;
wire [15:0] \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.u1.s ;
wire [15:0] \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.u2.a ;
wire [15:0] \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.u2.b ;
wire \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.u2.cin ;
wire \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.u2.cout ;
wire [15:0] \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.u2.s ;
wire \add_33ns_33s_33_2_1_U7.ce ;
wire \add_33ns_33s_33_2_1_U7.clk ;
wire [32:0] \add_33ns_33s_33_2_1_U7.din0 ;
wire [32:0] \add_33ns_33s_33_2_1_U7.din1 ;
wire [32:0] \add_33ns_33s_33_2_1_U7.dout ;
wire \add_33ns_33s_33_2_1_U7.reset ;
wire [32:0] \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.a ;
wire [32:0] \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.ain_s0 ;
wire [32:0] \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.b ;
wire [32:0] \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.bin_s0 ;
wire \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.ce ;
wire \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.clk ;
wire \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.facout_s1 ;
wire \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.facout_s2 ;
wire [15:0] \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.fas_s1 ;
wire [16:0] \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.fas_s2 ;
wire \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.reset ;
wire [32:0] \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.s ;
wire [15:0] \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.u1.a ;
wire [15:0] \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.u1.b ;
wire \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.u1.cin ;
wire \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.u1.cout ;
wire [15:0] \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.u1.s ;
wire [16:0] \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.u2.a ;
wire [16:0] \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.u2.b ;
wire \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.u2.cin ;
wire \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.u2.cout ;
wire [16:0] \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.u2.s ;
wire \add_33s_33s_33_2_1_U1.ce ;
wire \add_33s_33s_33_2_1_U1.clk ;
wire [32:0] \add_33s_33s_33_2_1_U1.din0 ;
wire [32:0] \add_33s_33s_33_2_1_U1.din1 ;
wire [32:0] \add_33s_33s_33_2_1_U1.dout ;
wire \add_33s_33s_33_2_1_U1.reset ;
wire [32:0] \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.a ;
wire [32:0] \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.ain_s0 ;
wire [32:0] \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.b ;
wire [32:0] \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.bin_s0 ;
wire \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.ce ;
wire \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.clk ;
wire \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.facout_s1 ;
wire \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.facout_s2 ;
wire [15:0] \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.fas_s1 ;
wire [16:0] \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.fas_s2 ;
wire \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.reset ;
wire [32:0] \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.s ;
wire [15:0] \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.u1.a ;
wire [15:0] \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.u1.b ;
wire \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.u1.cin ;
wire \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.u1.cout ;
wire [15:0] \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.u1.s ;
wire [16:0] \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.u2.a ;
wire [16:0] \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.u2.b ;
wire \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.u2.cin ;
wire \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.u2.cout ;
wire [16:0] \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.u2.s ;
wire \add_34s_34s_34_2_1_U3.ce ;
wire \add_34s_34s_34_2_1_U3.clk ;
wire [33:0] \add_34s_34s_34_2_1_U3.din0 ;
wire [33:0] \add_34s_34s_34_2_1_U3.din1 ;
wire [33:0] \add_34s_34s_34_2_1_U3.dout ;
wire \add_34s_34s_34_2_1_U3.reset ;
wire [33:0] \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.a ;
wire [33:0] \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.ain_s0 ;
wire [33:0] \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.b ;
wire [33:0] \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.bin_s0 ;
wire \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.ce ;
wire \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.clk ;
wire \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.facout_s1 ;
wire \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.facout_s2 ;
wire [16:0] \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.fas_s1 ;
wire [16:0] \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.fas_s2 ;
wire \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.reset ;
wire [33:0] \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.s ;
wire [16:0] \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.u1.a ;
wire [16:0] \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.u1.b ;
wire \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.u1.cin ;
wire \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.u1.cout ;
wire [16:0] \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.u1.s ;
wire [16:0] \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.u2.a ;
wire [16:0] \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.u2.b ;
wire \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.u2.cin ;
wire \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.u2.cout ;
wire [16:0] \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.u2.s ;
wire \add_36s_36s_36_2_1_U9.ce ;
wire \add_36s_36s_36_2_1_U9.clk ;
wire [35:0] \add_36s_36s_36_2_1_U9.din0 ;
wire [35:0] \add_36s_36s_36_2_1_U9.din1 ;
wire [35:0] \add_36s_36s_36_2_1_U9.dout ;
wire \add_36s_36s_36_2_1_U9.reset ;
wire [35:0] \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.a ;
wire [35:0] \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.ain_s0 ;
wire [35:0] \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.b ;
wire [35:0] \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.bin_s0 ;
wire \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.ce ;
wire \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.clk ;
wire \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.facout_s1 ;
wire \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.facout_s2 ;
wire [17:0] \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.fas_s1 ;
wire [17:0] \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.fas_s2 ;
wire \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.reset ;
wire [35:0] \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.s ;
wire [17:0] \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.u1.a ;
wire [17:0] \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.u1.b ;
wire \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.u1.cin ;
wire \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.u1.cout ;
wire [17:0] \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.u1.s ;
wire [17:0] \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.u2.a ;
wire [17:0] \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.u2.b ;
wire \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.u2.cin ;
wire \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.u2.cout ;
wire [17:0] \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.u2.s ;
wire [1:0] add_ln69_1_fu_777_p2;
wire [9:0] add_ln69_3_fu_849_p2;
wire and_ln340_1_fu_558_p2;
wire and_ln340_fu_526_p2;
wire and_ln785_1_fu_564_p2;
wire and_ln785_fu_552_p2;
wire and_ln786_fu_537_p2;
wire ap_CS_fsm_state1;
wire ap_CS_fsm_state10;
wire ap_CS_fsm_state11;
wire ap_CS_fsm_state12;
wire ap_CS_fsm_state13;
wire ap_CS_fsm_state14;
wire ap_CS_fsm_state15;
wire ap_CS_fsm_state16;
wire ap_CS_fsm_state17;
wire ap_CS_fsm_state18;
wire ap_CS_fsm_state19;
wire ap_CS_fsm_state2;
wire ap_CS_fsm_state20;
wire ap_CS_fsm_state21;
wire ap_CS_fsm_state22;
wire ap_CS_fsm_state23;
wire ap_CS_fsm_state24;
wire ap_CS_fsm_state25;
wire ap_CS_fsm_state3;
wire ap_CS_fsm_state4;
wire ap_CS_fsm_state5;
wire ap_CS_fsm_state6;
wire ap_CS_fsm_state7;
wire ap_CS_fsm_state8;
wire ap_CS_fsm_state9;
wire [24:0] ap_NS_fsm;
wire ap_clk;
wire ap_done;
wire ap_idle;
wire ap_ready;
wire ap_rst;
wire ap_start;
wire [32:0] grp_fu_313_p0;
wire [32:0] grp_fu_313_p1;
wire [32:0] grp_fu_313_p2;
wire [22:0] grp_fu_378_p0;
wire [22:0] grp_fu_378_p2;
wire [33:0] grp_fu_604_p0;
wire [33:0] grp_fu_604_p1;
wire [33:0] grp_fu_604_p2;
wire [31:0] grp_fu_667_p2;
wire [31:0] grp_fu_756_p1;
wire [31:0] grp_fu_756_p2;
wire [31:0] grp_fu_786_p0;
wire [31:0] grp_fu_786_p2;
wire [32:0] grp_fu_825_p0;
wire [32:0] grp_fu_825_p1;
wire [32:0] grp_fu_825_p2;
wire [31:0] grp_fu_858_p0;
wire [31:0] grp_fu_858_p2;
wire [35:0] grp_fu_878_p0;
wire [35:0] grp_fu_878_p1;
wire [35:0] grp_fu_878_p2;
wire [31:0] grp_fu_904_p2;
wire icmp_ln1496_fu_730_p2;
wire icmp_ln768_fu_384_p2;
wire icmp_ln786_fu_389_p2;
wire icmp_ln851_1_fu_661_p2;
wire icmp_ln851_2_fu_323_p2;
wire icmp_ln851_3_fu_888_p2;
wire icmp_ln851_fu_257_p2;
wire [3:0] newSel22_fu_581_p3;
wire [1:0] op_0;
wire [31:0] op_10;
wire [1:0] op_11;
wire op_15_V_fu_747_p2;
wire [9:0] op_16_V_fu_807_p3;
wire [3:0] op_17;
wire [7:0] op_18;
wire [7:0] op_19;
wire [1:0] op_2;
wire [6:0] op_21_V_fu_292_p2;
wire [3:0] op_3;
wire [31:0] op_31;
wire op_31_ap_vld;
wire [7:0] op_4;
wire [3:0] op_5;
wire [3:0] op_6_V_fu_614_p3;
wire op_7;
wire [15:0] op_8;
wire [3:0] op_9;
wire or_cond_fu_610_p2;
wire or_ln340_fu_472_p2;
wire or_ln785_1_fu_547_p2;
wire or_ln785_2_fu_569_p2;
wire or_ln785_fu_406_p2;
wire or_ln786_fu_467_p2;
wire overflow_fu_458_p2;
wire p_Result_1_fu_269_p3;
wire p_Result_2_fu_677_p3;
wire p_Result_3_fu_416_p3;
wire p_Result_4_fu_696_p3;
wire p_Result_5_fu_909_p3;
wire p_Result_7_fu_398_p3;
wire p_Result_8_fu_450_p3;
wire [3:0] p_Result_s_16_fu_510_p4;
wire [3:0] p_Val2_1_fu_443_p3;
wire [2:0] p_Val2_2_fu_504_p2;
wire [4:0] r_V_fu_640_p3;
wire [7:0] ret_V_14_fu_351_p1;
wire [7:0] ret_V_14_fu_351_p2;
wire [6:0] ret_V_15_fu_281_p3;
wire [31:0] ret_V_18_fu_712_p3;
wire [5:0] ret_V_2_fu_239_p4;
wire [6:0] ret_V_3_fu_263_p2;
wire [2:0] ret_V_6_fu_672_p2;
wire [2:0] ret_V_7_fu_689_p3;
wire [8:0] ret_V_fu_801_p2;
wire [17:0] rhs_1_fu_302_p3;
wire [34:0] rhs_5_fu_867_p3;
wire sel_tmp11_fu_575_p2;
wire [22:0] select_ln353_fu_428_p3;
wire [1:0] select_ln69_fu_770_p3;
wire [8:0] select_ln703_fu_794_p3;
wire [2:0] select_ln850_1_fu_684_p3;
wire [31:0] select_ln850_3_fu_706_p3;
wire [31:0] select_ln850_4_fu_916_p3;
wire [22:0] select_ln850_6_fu_423_p3;
wire [6:0] select_ln850_fu_276_p3;
wire [4:0] sext_ln1116_fu_620_p1;
wire [31:0] sext_ln1192_fu_298_p0;
wire [1:0] sext_ln1196_fu_435_p0;
wire [2:0] sext_ln1196_fu_435_p1;
wire [3:0] sext_ln1496_fu_726_p1;
wire [4:0] sext_ln1498_fu_743_p1;
wire [9:0] sext_ln69_3_fu_841_p1;
wire [6:0] sext_ln69_fu_288_p1;
wire [7:0] sext_ln703_1_fu_791_p0;
wire [8:0] sext_ln703_1_fu_791_p1;
wire [1:0] sext_ln703_2_fu_589_p0;
wire [7:0] sext_ln703_3_fu_863_p0;
wire [1:0] sext_ln703_fu_339_p0;
wire [7:0] sext_ln703_fu_339_p1;
wire [6:0] sext_ln831_fu_249_p1;
wire [22:0] sext_ln850_fu_375_p1;
wire [1:0] shl_ln728_1_fu_736_p1;
wire [4:0] shl_ln728_1_fu_736_p3;
wire [1:0] shl_ln_fu_719_p1;
wire [2:0] shl_ln_fu_719_p3;
wire [4:0] sub_ln1118_fu_624_p2;
wire [23:0] tmp_10_fu_593_p3;
wire tmp_4_fu_477_p3;
wire tmp_5_fu_485_p3;
wire [7:0] trunc_ln1196_1_fu_347_p0;
wire [2:0] trunc_ln1196_1_fu_347_p1;
wire [7:0] trunc_ln1196_fu_343_p0;
wire [1:0] trunc_ln1196_fu_343_p1;
wire [1:0] trunc_ln851_1_fu_657_p1;
wire [31:0] trunc_ln851_2_fu_319_p0;
wire [10:0] trunc_ln851_2_fu_319_p1;
wire [1:0] trunc_ln851_3_fu_703_p0;
wire trunc_ln851_3_fu_703_p1;
wire [7:0] trunc_ln851_4_fu_884_p0;
wire [2:0] trunc_ln851_4_fu_884_p1;
wire [9:0] trunc_ln851_fu_253_p1;
wire [2:0] xor_ln1196_1_fu_438_p2;
wire xor_ln1496_fu_761_p2;
wire xor_ln340_fu_520_p2;
wire xor_ln365_1_fu_498_p2;
wire xor_ln365_fu_492_p2;
wire [1:0] xor_ln731_fu_394_p1;
wire [1:0] xor_ln731_fu_394_p2;
wire xor_ln785_1_fu_542_p2;
wire xor_ln785_fu_411_p2;
wire xor_ln786_1_fu_532_p2;
wire xor_ln786_fu_462_p2;
wire [9:0] zext_ln69_1_fu_845_p1;
wire [1:0] zext_ln69_fu_766_p1;


assign add_ln69_1_fu_777_p2 = select_ln69_fu_770_p3 + xor_ln1496_fu_761_p2;
assign add_ln69_3_fu_849_p2 = $signed({ 1'h0, op_18 }) + $signed(op_17);
assign op_21_V_fu_292_p2 = $signed(ret_V_15_fu_281_p3) + $signed(op_9);
assign ret_V_3_fu_263_p2 = $signed(op_8[15:10]) + $signed(2'h1);
assign ret_V_6_fu_672_p2 = ret_V_5_reg_1130 + 1'h1;
assign ret_V_fu_801_p2 = $signed(op_4) + $signed(select_ln703_fu_794_p3);
assign _049_ = icmp_ln851_3_reg_1242 & ap_CS_fsm[23];
assign _050_ = icmp_ln851_2_reg_965 & ap_CS_fsm[5];
assign _051_ = ap_CS_fsm[10] & _054_;
assign _052_ = _055_ & ap_CS_fsm[0];
assign _053_ = ap_start & ap_CS_fsm[0];
assign and_ln340_1_fu_558_p2 = or_ln786_fu_467_p2 & or_ln340_fu_472_p2;
assign and_ln340_fu_526_p2 = xor_ln340_fu_520_p2 & or_ln786_fu_467_p2;
assign and_ln785_1_fu_564_p2 = xor_ln785_reg_1057 & and_ln786_fu_537_p2;
assign and_ln785_fu_552_p2 = or_ln785_1_fu_547_p2 & and_ln786_fu_537_p2;
assign and_ln786_fu_537_p2 = xor_ln786_1_fu_532_p2 & p_Result_7_reg_1045;
assign overflow_fu_458_p2 = xor_ln785_reg_1057 & or_ln785_reg_1051;
assign sel_tmp11_fu_575_p2 = xor_ln365_1_fu_498_p2 & or_ln785_2_fu_569_p2;
assign xor_ln1496_fu_761_p2 = ~ icmp_ln1496_reg_1162;
assign xor_ln786_fu_462_p2 = ~ p_Result_7_reg_1045;
assign xor_ln340_fu_520_p2 = ~ or_ln340_fu_472_p2;
assign xor_ln786_1_fu_532_p2 = ~ icmp_ln786_reg_1028;
assign xor_ln785_1_fu_542_p2 = ~ or_ln785_reg_1051;
assign xor_ln365_1_fu_498_p2 = ~ xor_ln365_fu_492_p2;
assign xor_ln785_fu_411_p2 = ~ p_Result_6_reg_1003;
assign p_Val2_2_fu_504_p2 = ~ { xor_ln731_reg_1039[0], 2'h0 };
assign _054_ = ~ icmp_ln851_1_reg_1137;
assign _055_ = ~ ap_start;
assign _056_ = ! r_V_fu_640_p3[1:0];
assign _057_ = ! op_8[9:0];
assign _058_ = { op_2, 3'h0 } == { op_5[3], op_5 };
always @(posedge \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.clk )
\add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.bin_s1  <= _060_;
always @(posedge \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.clk )
\add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.ain_s1  <= _059_;
always @(posedge \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.clk )
\add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.sum_s1  <= _062_;
always @(posedge \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.clk )
\add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.carry_s1  <= _061_;
assign _060_ = \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.ce  ? \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.b [22:11] : \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.bin_s1 ;
assign _059_ = \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.ce  ? \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.a [22:11] : \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.ain_s1 ;
assign _061_ = \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.ce  ? \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.facout_s1  : \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.carry_s1 ;
assign _062_ = \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.ce  ? \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.fas_s1  : \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.sum_s1 ;
assign _063_ = \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.u1.a  + \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.u1.b ;
assign { \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.u1.cout , \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.u1.s  } = _063_ + \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.u1.cin ;
assign _064_ = \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.u2.a  + \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.u2.b ;
assign { \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.u2.cout , \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.u2.s  } = _064_ + \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.u2.cin ;
always @(posedge \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.clk )
\add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.bin_s1  <= _066_;
always @(posedge \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.clk )
\add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.ain_s1  <= _065_;
always @(posedge \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.clk )
\add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.sum_s1  <= _068_;
always @(posedge \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.clk )
\add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.carry_s1  <= _067_;
assign _066_ = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.ce  ? \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.b [31:16] : \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.bin_s1 ;
assign _065_ = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.ce  ? \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.a [31:16] : \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.ain_s1 ;
assign _067_ = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.ce  ? \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.facout_s1  : \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.carry_s1 ;
assign _068_ = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.ce  ? \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.fas_s1  : \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.sum_s1 ;
assign _069_ = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.u1.a  + \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.u1.b ;
assign { \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.u1.cout , \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.u1.s  } = _069_ + \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.u1.cin ;
assign _070_ = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.u2.a  + \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.u2.b ;
assign { \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.u2.cout , \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.u2.s  } = _070_ + \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.u2.cin ;
always @(posedge \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.clk )
\add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.bin_s1  <= _072_;
always @(posedge \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.clk )
\add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.ain_s1  <= _071_;
always @(posedge \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.clk )
\add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.sum_s1  <= _074_;
always @(posedge \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.clk )
\add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.carry_s1  <= _073_;
assign _072_ = \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.ce  ? \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.b [31:16] : \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.bin_s1 ;
assign _071_ = \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.ce  ? \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.a [31:16] : \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.ain_s1 ;
assign _073_ = \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.ce  ? \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.facout_s1  : \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.carry_s1 ;
assign _074_ = \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.ce  ? \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.fas_s1  : \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.sum_s1 ;
assign _075_ = \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.u1.a  + \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.u1.b ;
assign { \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.u1.cout , \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.u1.s  } = _075_ + \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.u1.cin ;
assign _076_ = \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.u2.a  + \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.u2.b ;
assign { \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.u2.cout , \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.u2.s  } = _076_ + \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.u2.cin ;
always @(posedge \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.clk )
\add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.bin_s1  <= _078_;
always @(posedge \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.clk )
\add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.ain_s1  <= _077_;
always @(posedge \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.clk )
\add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.sum_s1  <= _080_;
always @(posedge \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.clk )
\add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.carry_s1  <= _079_;
assign _078_ = \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.ce  ? \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.b [31:16] : \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.bin_s1 ;
assign _077_ = \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.ce  ? \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.a [31:16] : \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.ain_s1 ;
assign _079_ = \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.ce  ? \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.facout_s1  : \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.carry_s1 ;
assign _080_ = \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.ce  ? \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.fas_s1  : \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.sum_s1 ;
assign _081_ = \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.u1.a  + \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.u1.b ;
assign { \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.u1.cout , \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.u1.s  } = _081_ + \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.u1.cin ;
assign _082_ = \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.u2.a  + \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.u2.b ;
assign { \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.u2.cout , \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.u2.s  } = _082_ + \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.u2.cin ;
always @(posedge \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.clk )
\add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.bin_s1  <= _084_;
always @(posedge \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.clk )
\add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.ain_s1  <= _083_;
always @(posedge \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.clk )
\add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.sum_s1  <= _086_;
always @(posedge \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.clk )
\add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.carry_s1  <= _085_;
assign _084_ = \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.ce  ? \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.b [31:16] : \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.bin_s1 ;
assign _083_ = \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.ce  ? \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.a [31:16] : \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.ain_s1 ;
assign _085_ = \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.ce  ? \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.facout_s1  : \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.carry_s1 ;
assign _086_ = \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.ce  ? \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.fas_s1  : \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.sum_s1 ;
assign _087_ = \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.u1.a  + \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.u1.b ;
assign { \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.u1.cout , \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.u1.s  } = _087_ + \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.u1.cin ;
assign _088_ = \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.u2.a  + \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.u2.b ;
assign { \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.u2.cout , \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.u2.s  } = _088_ + \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.u2.cin ;
always @(posedge \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.clk )
\add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.bin_s1  <= _090_;
always @(posedge \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.clk )
\add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.ain_s1  <= _089_;
always @(posedge \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.clk )
\add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.sum_s1  <= _092_;
always @(posedge \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.clk )
\add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.carry_s1  <= _091_;
assign _090_ = \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.ce  ? \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.b [31:16] : \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.bin_s1 ;
assign _089_ = \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.ce  ? \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.a [31:16] : \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.ain_s1 ;
assign _091_ = \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.ce  ? \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.facout_s1  : \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.carry_s1 ;
assign _092_ = \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.ce  ? \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.fas_s1  : \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.sum_s1 ;
assign _093_ = \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.u1.a  + \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.u1.b ;
assign { \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.u1.cout , \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.u1.s  } = _093_ + \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.u1.cin ;
assign _094_ = \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.u2.a  + \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.u2.b ;
assign { \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.u2.cout , \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.u2.s  } = _094_ + \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.u2.cin ;
always @(posedge \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.clk )
\add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.bin_s1  <= _096_;
always @(posedge \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.clk )
\add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.ain_s1  <= _095_;
always @(posedge \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.clk )
\add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.sum_s1  <= _098_;
always @(posedge \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.clk )
\add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.carry_s1  <= _097_;
assign _096_ = \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.ce  ? \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.b [32:16] : \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.bin_s1 ;
assign _095_ = \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.ce  ? \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.a [32:16] : \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.ain_s1 ;
assign _097_ = \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.ce  ? \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.facout_s1  : \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.carry_s1 ;
assign _098_ = \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.ce  ? \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.fas_s1  : \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.sum_s1 ;
assign _099_ = \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.u1.a  + \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.u1.b ;
assign { \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.u1.cout , \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.u1.s  } = _099_ + \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.u1.cin ;
assign _100_ = \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.u2.a  + \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.u2.b ;
assign { \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.u2.cout , \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.u2.s  } = _100_ + \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.u2.cin ;
always @(posedge \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.clk )
\add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.bin_s1  <= _102_;
always @(posedge \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.clk )
\add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.ain_s1  <= _101_;
always @(posedge \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.clk )
\add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.sum_s1  <= _104_;
always @(posedge \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.clk )
\add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.carry_s1  <= _103_;
assign _102_ = \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.ce  ? \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.b [32:16] : \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.bin_s1 ;
assign _101_ = \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.ce  ? \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.a [32:16] : \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.ain_s1 ;
assign _103_ = \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.ce  ? \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.facout_s1  : \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.carry_s1 ;
assign _104_ = \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.ce  ? \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.fas_s1  : \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.sum_s1 ;
assign _105_ = \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.u1.a  + \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.u1.b ;
assign { \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.u1.cout , \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.u1.s  } = _105_ + \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.u1.cin ;
assign _106_ = \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.u2.a  + \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.u2.b ;
assign { \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.u2.cout , \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.u2.s  } = _106_ + \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.u2.cin ;
always @(posedge \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.clk )
\add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.bin_s1  <= _108_;
always @(posedge \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.clk )
\add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.ain_s1  <= _107_;
always @(posedge \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.clk )
\add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.sum_s1  <= _110_;
always @(posedge \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.clk )
\add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.carry_s1  <= _109_;
assign _108_ = \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.ce  ? \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.b [33:17] : \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.bin_s1 ;
assign _107_ = \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.ce  ? \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.a [33:17] : \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.ain_s1 ;
assign _109_ = \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.ce  ? \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.facout_s1  : \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.carry_s1 ;
assign _110_ = \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.ce  ? \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.fas_s1  : \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.sum_s1 ;
assign _111_ = \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.u1.a  + \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.u1.b ;
assign { \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.u1.cout , \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.u1.s  } = _111_ + \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.u1.cin ;
assign _112_ = \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.u2.a  + \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.u2.b ;
assign { \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.u2.cout , \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.u2.s  } = _112_ + \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.u2.cin ;
always @(posedge \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.clk )
\add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.bin_s1  <= _114_;
always @(posedge \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.clk )
\add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.ain_s1  <= _113_;
always @(posedge \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.clk )
\add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.sum_s1  <= _116_;
always @(posedge \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.clk )
\add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.carry_s1  <= _115_;
assign _114_ = \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.ce  ? \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.b [35:18] : \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.bin_s1 ;
assign _113_ = \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.ce  ? \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.a [35:18] : \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.ain_s1 ;
assign _115_ = \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.ce  ? \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.facout_s1  : \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.carry_s1 ;
assign _116_ = \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.ce  ? \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.fas_s1  : \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.sum_s1 ;
assign _117_ = \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.u1.a  + \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.u1.b ;
assign { \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.u1.cout , \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.u1.s  } = _117_ + \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.u1.cin ;
assign _118_ = \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.u2.a  + \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.u2.b ;
assign { \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.u2.cout , \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.u2.s  } = _118_ + \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.u2.cin ;
assign _119_ = $signed({ op_2, 1'h0 }) < $signed(op_3);
assign _120_ = | p_Result_s_reg_1010;
assign _121_ = p_Result_s_reg_1010 != 6'h3f;
assign _122_ = | op_10[10:0];
assign _123_ = | op_19[2:0];
assign or_cond_fu_610_p2 = sel_tmp11_reg_1083 | and_ln785_reg_1078;
assign or_ln340_fu_472_p2 = p_Result_6_reg_1003 | overflow_fu_458_p2;
assign or_ln785_1_fu_547_p2 = xor_ln785_1_fu_542_p2 | p_Result_6_reg_1003;
assign or_ln785_2_fu_569_p2 = and_ln785_1_fu_564_p2 | and_ln340_1_fu_558_p2;
assign or_ln785_fu_406_p2 = xor_ln731_fu_394_p2[1] | icmp_ln768_reg_1023;
assign or_ln786_fu_467_p2 = xor_ln786_fu_462_p2 | icmp_ln786_reg_1028;
always @(posedge ap_clk)
p_Val2_1_reg_1073[1:0] <= 2'h0;
always @(posedge ap_clk)
ret_V_6_reg_1142 <= _035_;
always @(posedge ap_clk)
ret_V_7_reg_1152 <= _036_;
always @(posedge ap_clk)
ret_V_18_reg_1157 <= _031_;
always @(posedge ap_clk)
ret_V_16_reg_970 <= _029_;
always @(posedge ap_clk)
tmp_reg_975 <= _043_;
always @(posedge ap_clk)
ret_V_19_reg_1247 <= _032_;
always @(posedge ap_clk)
ret_V_16_cast_reg_1252 <= _028_;
always @(posedge ap_clk)
sub_ln1118_reg_1103 <= _042_;
always @(posedge ap_clk)
ret_V_17_reg_1108 <= _030_;
always @(posedge ap_clk)
ret_V_12_cast_reg_1113 <= _027_;
always @(posedge ap_clk)
trunc_ln1196_reg_993 <= _045_;
always @(posedge ap_clk)
trunc_ln1196_1_reg_998 <= _044_;
always @(posedge ap_clk)
p_Result_6_reg_1003 <= _022_;
always @(posedge ap_clk)
p_Result_s_reg_1010 <= _024_;
always @(posedge ap_clk)
sext_ln850_reg_1016 <= _041_;
always @(posedge ap_clk)
xor_ln731_reg_1039 <= _046_;
always @(posedge ap_clk)
p_Result_7_reg_1045 <= _023_;
always @(posedge ap_clk)
or_ln785_reg_1051 <= _021_;
always @(posedge ap_clk)
xor_ln785_reg_1057 <= _047_;
always @(posedge ap_clk)
select_ln353_reg_1063 <= _039_;
always @(posedge ap_clk)
op_30_V_reg_1227 <= _020_;
always @(posedge ap_clk)
ret_V_reg_1192 <= _037_;
always @(posedge ap_clk)
op_27_V_reg_1197 <= _018_;
always @(posedge ap_clk)
op_21_V_reg_950 <= _017_;
always @(posedge ap_clk)
sext_ln831_reg_934 <= _040_;
always @(posedge ap_clk)
icmp_ln851_reg_940 <= _014_;
always @(posedge ap_clk)
ret_V_3_reg_945 <= _033_;
always @(posedge ap_clk)
icmp_ln851_3_reg_1242 <= _013_;
always @(posedge ap_clk)
icmp_ln851_2_reg_965 <= _012_;
always @(posedge ap_clk)
r_V_reg_1125 <= _026_;
always @(posedge ap_clk)
ret_V_5_reg_1130 <= _034_;
always @(posedge ap_clk)
icmp_ln851_1_reg_1137 <= _011_;
always @(posedge ap_clk)
icmp_ln768_reg_1023 <= _009_;
always @(posedge ap_clk)
icmp_ln786_reg_1028 <= _010_;
always @(posedge ap_clk)
icmp_ln1496_reg_1162 <= _008_;
always @(posedge ap_clk)
op_15_V_reg_1167 <= _016_;
always @(posedge ap_clk)
p_Val2_1_reg_1073[3:2] <= _025_;
always @(posedge ap_clk)
and_ln785_reg_1078 <= _006_;
always @(posedge ap_clk)
sel_tmp11_reg_1083 <= _038_;
always @(posedge ap_clk)
newSel22_reg_1088 <= _015_;
always @(posedge ap_clk)
op_28_V_reg_1212 <= _019_;
always @(posedge ap_clk)
add_ln69_3_reg_1217 <= _004_;
always @(posedge ap_clk)
add_ln69_reg_1177 <= _005_;
always @(posedge ap_clk)
add_ln69_1_reg_1182 <= _003_;
always @(posedge ap_clk)
add_ln691_reg_1034 <= _002_;
always @(posedge ap_clk)
add_ln691_4_reg_1259 <= _001_;
always @(posedge ap_clk)
add_ln691_1_reg_1147 <= _000_;
always @(posedge ap_clk)
ap_CS_fsm <= _007_;
assign _048_ = _053_ ? 2'h2 : 2'h1;
assign _124_ = ap_CS_fsm == 1'h1;
function [24:0] _362_;
input [24:0] a;
input [624:0] b;
input [24:0] s;
case (s)
25'b0000000000000000000000001:
_362_ = b[24:0];
25'b0000000000000000000000010:
_362_ = b[49:25];
25'b0000000000000000000000100:
_362_ = b[74:50];
25'b0000000000000000000001000:
_362_ = b[99:75];
25'b0000000000000000000010000:
_362_ = b[124:100];
25'b0000000000000000000100000:
_362_ = b[149:125];
25'b0000000000000000001000000:
_362_ = b[174:150];
25'b0000000000000000010000000:
_362_ = b[199:175];
25'b0000000000000000100000000:
_362_ = b[224:200];
25'b0000000000000001000000000:
_362_ = b[249:225];
25'b0000000000000010000000000:
_362_ = b[274:250];
25'b0000000000000100000000000:
_362_ = b[299:275];
25'b0000000000001000000000000:
_362_ = b[324:300];
25'b0000000000010000000000000:
_362_ = b[349:325];
25'b0000000000100000000000000:
_362_ = b[374:350];
25'b0000000001000000000000000:
_362_ = b[399:375];
25'b0000000010000000000000000:
_362_ = b[424:400];
25'b0000000100000000000000000:
_362_ = b[449:425];
25'b0000001000000000000000000:
_362_ = b[474:450];
25'b0000010000000000000000000:
_362_ = b[499:475];
25'b0000100000000000000000000:
_362_ = b[524:500];
25'b0001000000000000000000000:
_362_ = b[549:525];
25'b0010000000000000000000000:
_362_ = b[574:550];
25'b0100000000000000000000000:
_362_ = b[599:575];
25'b1000000000000000000000000:
_362_ = b[624:600];
25'b0000000000000000000000000:
_362_ = a;
default:
_362_ = 25'bx;
endcase
endfunction
assign ap_NS_fsm = _362_(25'hxxxxxxx, { 23'h000000, _048_, 600'h000002000002000002000002000002000002000002000002000002000002000002000002000002000002000002000002000002000002000002000002000002000002000002000000000001 }, { _124_, _148_, _147_, _146_, _145_, _144_, _143_, _142_, _141_, _140_, _139_, _138_, _137_, _136_, _135_, _134_, _133_, _132_, _131_, _130_, _129_, _128_, _127_, _126_, _125_ });
assign _125_ = ap_CS_fsm == 25'h1000000;
assign _126_ = ap_CS_fsm == 24'h800000;
assign _127_ = ap_CS_fsm == 23'h400000;
assign _128_ = ap_CS_fsm == 22'h200000;
assign _129_ = ap_CS_fsm == 21'h100000;
assign _130_ = ap_CS_fsm == 20'h80000;
assign _131_ = ap_CS_fsm == 19'h40000;
assign _132_ = ap_CS_fsm == 18'h20000;
assign _133_ = ap_CS_fsm == 17'h10000;
assign _134_ = ap_CS_fsm == 16'h8000;
assign _135_ = ap_CS_fsm == 15'h4000;
assign _136_ = ap_CS_fsm == 14'h2000;
assign _137_ = ap_CS_fsm == 13'h1000;
assign _138_ = ap_CS_fsm == 12'h800;
assign _139_ = ap_CS_fsm == 11'h400;
assign _140_ = ap_CS_fsm == 10'h200;
assign _141_ = ap_CS_fsm == 9'h100;
assign _142_ = ap_CS_fsm == 8'h80;
assign _143_ = ap_CS_fsm == 7'h40;
assign _144_ = ap_CS_fsm == 6'h20;
assign _145_ = ap_CS_fsm == 5'h10;
assign _146_ = ap_CS_fsm == 4'h8;
assign _147_ = ap_CS_fsm == 3'h4;
assign _148_ = ap_CS_fsm == 2'h2;
assign op_31_ap_vld = ap_CS_fsm[24] ? 1'h1 : 1'h0;
assign ap_idle = _052_ ? 1'h1 : 1'h0;
assign _035_ = _051_ ? ret_V_6_fu_672_p2 : ret_V_6_reg_1142;
assign _031_ = ap_CS_fsm[11] ? ret_V_18_fu_712_p3 : ret_V_18_reg_1157;
assign _036_ = ap_CS_fsm[11] ? ret_V_7_fu_689_p3 : ret_V_7_reg_1152;
assign _043_ = ap_CS_fsm[3] ? grp_fu_313_p2[32:11] : tmp_reg_975;
assign _029_ = ap_CS_fsm[3] ? grp_fu_313_p2 : ret_V_16_reg_970;
assign _028_ = ap_CS_fsm[21] ? grp_fu_878_p2[34:3] : ret_V_16_cast_reg_1252;
assign _032_ = ap_CS_fsm[21] ? grp_fu_878_p2 : ret_V_19_reg_1247;
assign _027_ = ap_CS_fsm[8] ? grp_fu_604_p2[32:1] : ret_V_12_cast_reg_1113;
assign _030_ = ap_CS_fsm[8] ? grp_fu_604_p2 : ret_V_17_reg_1108;
assign _042_ = ap_CS_fsm[8] ? sub_ln1118_fu_624_p2 : sub_ln1118_reg_1103;
assign _041_ = ap_CS_fsm[4] ? { tmp_reg_975[21], tmp_reg_975 } : sext_ln850_reg_1016;
assign _024_ = ap_CS_fsm[4] ? ret_V_14_fu_351_p2[7:2] : p_Result_s_reg_1010;
assign _022_ = ap_CS_fsm[4] ? ret_V_14_fu_351_p2[7] : p_Result_6_reg_1003;
assign _044_ = ap_CS_fsm[4] ? op_4[2:0] : trunc_ln1196_1_reg_998;
assign _045_ = ap_CS_fsm[4] ? op_4[1:0] : trunc_ln1196_reg_993;
assign _039_ = ap_CS_fsm[6] ? select_ln353_fu_428_p3 : select_ln353_reg_1063;
assign _047_ = ap_CS_fsm[6] ? xor_ln785_fu_411_p2 : xor_ln785_reg_1057;
assign _021_ = ap_CS_fsm[6] ? or_ln785_fu_406_p2 : or_ln785_reg_1051;
assign _023_ = ap_CS_fsm[6] ? xor_ln731_fu_394_p2[1] : p_Result_7_reg_1045;
assign _046_ = ap_CS_fsm[6] ? xor_ln731_fu_394_p2 : xor_ln731_reg_1039;
assign _020_ = ap_CS_fsm[19] ? grp_fu_858_p2 : op_30_V_reg_1227;
assign _018_ = ap_CS_fsm[15] ? grp_fu_786_p2 : op_27_V_reg_1197;
assign _037_ = ap_CS_fsm[15] ? ret_V_fu_801_p2 : ret_V_reg_1192;
assign _017_ = ap_CS_fsm[1] ? op_21_V_fu_292_p2 : op_21_V_reg_950;
assign _033_ = ap_CS_fsm[0] ? ret_V_3_fu_263_p2 : ret_V_3_reg_945;
assign _014_ = ap_CS_fsm[0] ? icmp_ln851_fu_257_p2 : icmp_ln851_reg_940;
assign _040_ = ap_CS_fsm[0] ? { op_8[15], op_8[15:10] } : sext_ln831_reg_934;
assign _013_ = ap_CS_fsm[20] ? icmp_ln851_3_fu_888_p2 : icmp_ln851_3_reg_1242;
assign _012_ = ap_CS_fsm[2] ? icmp_ln851_2_fu_323_p2 : icmp_ln851_2_reg_965;
assign _011_ = ap_CS_fsm[9] ? icmp_ln851_1_fu_661_p2 : icmp_ln851_1_reg_1137;
assign _034_ = ap_CS_fsm[9] ? r_V_fu_640_p3[4:2] : ret_V_5_reg_1130;
assign _026_ = ap_CS_fsm[9] ? r_V_fu_640_p3 : r_V_reg_1125;
assign _010_ = ap_CS_fsm[5] ? icmp_ln786_fu_389_p2 : icmp_ln786_reg_1028;
assign _009_ = ap_CS_fsm[5] ? icmp_ln768_fu_384_p2 : icmp_ln768_reg_1023;
assign _016_ = ap_CS_fsm[12] ? op_15_V_fu_747_p2 : op_15_V_reg_1167;
assign _008_ = ap_CS_fsm[12] ? icmp_ln1496_fu_730_p2 : icmp_ln1496_reg_1162;
assign _015_ = ap_CS_fsm[7] ? newSel22_fu_581_p3 : newSel22_reg_1088;
assign _038_ = ap_CS_fsm[7] ? sel_tmp11_fu_575_p2 : sel_tmp11_reg_1083;
assign _006_ = ap_CS_fsm[7] ? and_ln785_fu_552_p2 : and_ln785_reg_1078;
assign _025_ = ap_CS_fsm[7] ? xor_ln731_reg_1039 : p_Val2_1_reg_1073[3:2];
assign _004_ = ap_CS_fsm[17] ? add_ln69_3_fu_849_p2 : add_ln69_3_reg_1217;
assign _019_ = ap_CS_fsm[17] ? grp_fu_825_p2[32:1] : op_28_V_reg_1212;
assign _003_ = ap_CS_fsm[13] ? add_ln69_1_fu_777_p2 : add_ln69_1_reg_1182;
assign _005_ = ap_CS_fsm[13] ? grp_fu_756_p2 : add_ln69_reg_1177;
assign _002_ = _050_ ? grp_fu_378_p2 : add_ln691_reg_1034;
assign _001_ = _049_ ? grp_fu_904_p2 : add_ln691_4_reg_1259;
assign _000_ = ap_CS_fsm[10] ? grp_fu_667_p2 : add_ln691_1_reg_1147;
assign _007_ = ap_rst ? 25'h0000001 : ap_NS_fsm;
assign sub_ln1118_fu_624_p2 = $signed(1'h0) - $signed(op_6_V_fu_614_p3);
assign icmp_ln1496_fu_730_p2 = _119_ ? 1'h1 : 1'h0;
assign icmp_ln768_fu_384_p2 = _120_ ? 1'h1 : 1'h0;
assign icmp_ln786_fu_389_p2 = _121_ ? 1'h1 : 1'h0;
assign icmp_ln851_1_fu_661_p2 = _056_ ? 1'h1 : 1'h0;
assign icmp_ln851_2_fu_323_p2 = _122_ ? 1'h1 : 1'h0;
assign icmp_ln851_3_fu_888_p2 = _123_ ? 1'h1 : 1'h0;
assign icmp_ln851_fu_257_p2 = _057_ ? 1'h1 : 1'h0;
assign newSel22_fu_581_p3 = and_ln340_fu_526_p2 ? { xor_ln731_reg_1039, 2'h0 } : { xor_ln1196_1_fu_438_p2[2], p_Val2_2_fu_504_p2 };
assign op_15_V_fu_747_p2 = _058_ ? 1'h1 : 1'h0;
assign op_31 = ret_V_19_reg_1247[35] ? select_ln850_4_fu_916_p3 : ret_V_16_cast_reg_1252;
assign op_6_V_fu_614_p3 = or_cond_fu_610_p2 ? p_Val2_1_reg_1073 : newSel22_reg_1088;
assign r_V_fu_640_p3 = op_7 ? sub_ln1118_reg_1103 : 5'h00;
assign ret_V_15_fu_281_p3 = op_8[15] ? select_ln850_fu_276_p3 : sext_ln831_reg_934;
assign ret_V_18_fu_712_p3 = ret_V_17_reg_1108[33] ? select_ln850_3_fu_706_p3 : ret_V_12_cast_reg_1113;
assign ret_V_7_fu_689_p3 = r_V_reg_1125[4] ? select_ln850_1_fu_684_p3 : ret_V_5_reg_1130;
assign select_ln353_fu_428_p3 = ret_V_16_reg_970[32] ? select_ln850_6_fu_423_p3 : sext_ln850_reg_1016;
assign select_ln69_fu_770_p3 = op_15_V_reg_1167 ? 2'h3 : 2'h0;
assign select_ln703_fu_794_p3 = op_7 ? 9'h1ff : 9'h000;
assign select_ln850_1_fu_684_p3 = icmp_ln851_1_reg_1137 ? ret_V_5_reg_1130 : ret_V_6_reg_1142;
assign select_ln850_3_fu_706_p3 = op_11[0] ? add_ln691_1_reg_1147 : ret_V_12_cast_reg_1113;
assign select_ln850_4_fu_916_p3 = icmp_ln851_3_reg_1242 ? add_ln691_4_reg_1259 : ret_V_16_cast_reg_1252;
assign select_ln850_6_fu_423_p3 = icmp_ln851_2_reg_965 ? add_ln691_reg_1034 : sext_ln850_reg_1016;
assign select_ln850_fu_276_p3 = icmp_ln851_reg_940 ? sext_ln831_reg_934 : ret_V_3_reg_945;
assign ret_V_14_fu_351_p2 = $signed(op_2) ^ $signed(op_4);
assign xor_ln1196_1_fu_438_p2 = trunc_ln1196_1_reg_998 ^ { op_2[1], op_2 };
assign xor_ln365_fu_492_p2 = xor_ln731_reg_1039[1] ^ xor_ln1196_1_fu_438_p2[2];
assign xor_ln731_fu_394_p2 = op_2 ^ trunc_ln1196_reg_993;
assign ap_CS_fsm_state1 = ap_CS_fsm[0];
assign ap_CS_fsm_state10 = ap_CS_fsm[9];
assign ap_CS_fsm_state11 = ap_CS_fsm[10];
assign ap_CS_fsm_state12 = ap_CS_fsm[11];
assign ap_CS_fsm_state13 = ap_CS_fsm[12];
assign ap_CS_fsm_state14 = ap_CS_fsm[13];
assign ap_CS_fsm_state15 = ap_CS_fsm[14];
assign ap_CS_fsm_state16 = ap_CS_fsm[15];
assign ap_CS_fsm_state17 = ap_CS_fsm[16];
assign ap_CS_fsm_state18 = ap_CS_fsm[17];
assign ap_CS_fsm_state19 = ap_CS_fsm[18];
assign ap_CS_fsm_state2 = ap_CS_fsm[1];
assign ap_CS_fsm_state20 = ap_CS_fsm[19];
assign ap_CS_fsm_state21 = ap_CS_fsm[20];
assign ap_CS_fsm_state22 = ap_CS_fsm[21];
assign ap_CS_fsm_state23 = ap_CS_fsm[22];
assign ap_CS_fsm_state24 = ap_CS_fsm[23];
assign ap_CS_fsm_state25 = ap_CS_fsm[24];
assign ap_CS_fsm_state3 = ap_CS_fsm[2];
assign ap_CS_fsm_state4 = ap_CS_fsm[3];
assign ap_CS_fsm_state5 = ap_CS_fsm[4];
assign ap_CS_fsm_state6 = ap_CS_fsm[5];
assign ap_CS_fsm_state7 = ap_CS_fsm[6];
assign ap_CS_fsm_state8 = ap_CS_fsm[7];
assign ap_CS_fsm_state9 = ap_CS_fsm[8];
assign ap_done = op_31_ap_vld;
assign ap_ready = op_31_ap_vld;
assign grp_fu_313_p0 = { op_21_V_reg_950[6], op_21_V_reg_950[6], op_21_V_reg_950[6], op_21_V_reg_950[6], op_21_V_reg_950[6], op_21_V_reg_950[6], op_21_V_reg_950[6], op_21_V_reg_950[6], op_21_V_reg_950[6], op_21_V_reg_950[6], op_21_V_reg_950[6], op_21_V_reg_950[6], op_21_V_reg_950[6], op_21_V_reg_950[6], op_21_V_reg_950[6], op_21_V_reg_950, 11'h000 };
assign grp_fu_313_p1 = { op_10[31], op_10 };
assign grp_fu_378_p0 = { tmp_reg_975[21], tmp_reg_975 };
assign grp_fu_604_p0 = { select_ln353_reg_1063[22], select_ln353_reg_1063[22], select_ln353_reg_1063[22], select_ln353_reg_1063[22], select_ln353_reg_1063[22], select_ln353_reg_1063[22], select_ln353_reg_1063[22], select_ln353_reg_1063[22], select_ln353_reg_1063[22], select_ln353_reg_1063[22], select_ln353_reg_1063, 1'h0 };
assign grp_fu_604_p1 = { op_11[1], op_11[1], op_11[1], op_11[1], op_11[1], op_11[1], op_11[1], op_11[1], op_11[1], op_11[1], op_11[1], op_11[1], op_11[1], op_11[1], op_11[1], op_11[1], op_11[1], op_11[1], op_11[1], op_11[1], op_11[1], op_11[1], op_11[1], op_11[1], op_11[1], op_11[1], op_11[1], op_11[1], op_11[1], op_11[1], op_11[1], op_11[1], op_11 };
assign grp_fu_756_p1 = { ret_V_7_reg_1152[2], ret_V_7_reg_1152[2], ret_V_7_reg_1152[2], ret_V_7_reg_1152[2], ret_V_7_reg_1152[2], ret_V_7_reg_1152[2], ret_V_7_reg_1152[2], ret_V_7_reg_1152[2], ret_V_7_reg_1152[2], ret_V_7_reg_1152[2], ret_V_7_reg_1152[2], ret_V_7_reg_1152[2], ret_V_7_reg_1152[2], ret_V_7_reg_1152[2], ret_V_7_reg_1152[2], ret_V_7_reg_1152[2], ret_V_7_reg_1152[2], ret_V_7_reg_1152[2], ret_V_7_reg_1152[2], ret_V_7_reg_1152[2], ret_V_7_reg_1152[2], ret_V_7_reg_1152[2], ret_V_7_reg_1152[2], ret_V_7_reg_1152[2], ret_V_7_reg_1152[2], ret_V_7_reg_1152[2], ret_V_7_reg_1152[2], ret_V_7_reg_1152[2], ret_V_7_reg_1152[2], ret_V_7_reg_1152 };
assign grp_fu_786_p0 = { add_ln69_1_reg_1182[1], add_ln69_1_reg_1182[1], add_ln69_1_reg_1182[1], add_ln69_1_reg_1182[1], add_ln69_1_reg_1182[1], add_ln69_1_reg_1182[1], add_ln69_1_reg_1182[1], add_ln69_1_reg_1182[1], add_ln69_1_reg_1182[1], add_ln69_1_reg_1182[1], add_ln69_1_reg_1182[1], add_ln69_1_reg_1182[1], add_ln69_1_reg_1182[1], add_ln69_1_reg_1182[1], add_ln69_1_reg_1182[1], add_ln69_1_reg_1182[1], add_ln69_1_reg_1182[1], add_ln69_1_reg_1182[1], add_ln69_1_reg_1182[1], add_ln69_1_reg_1182[1], add_ln69_1_reg_1182[1], add_ln69_1_reg_1182[1], add_ln69_1_reg_1182[1], add_ln69_1_reg_1182[1], add_ln69_1_reg_1182[1], add_ln69_1_reg_1182[1], add_ln69_1_reg_1182[1], add_ln69_1_reg_1182[1], add_ln69_1_reg_1182[1], add_ln69_1_reg_1182[1], add_ln69_1_reg_1182 };
assign grp_fu_825_p0 = { op_27_V_reg_1197, 1'h0 };
assign grp_fu_825_p1 = { ret_V_reg_1192[8], ret_V_reg_1192[8], ret_V_reg_1192[8], ret_V_reg_1192[8], ret_V_reg_1192[8], ret_V_reg_1192[8], ret_V_reg_1192[8], ret_V_reg_1192[8], ret_V_reg_1192[8], ret_V_reg_1192[8], ret_V_reg_1192[8], ret_V_reg_1192[8], ret_V_reg_1192[8], ret_V_reg_1192[8], ret_V_reg_1192[8], ret_V_reg_1192[8], ret_V_reg_1192[8], ret_V_reg_1192[8], ret_V_reg_1192[8], ret_V_reg_1192[8], ret_V_reg_1192[8], ret_V_reg_1192[8], ret_V_reg_1192[8], ret_V_reg_1192, 1'h0 };
assign grp_fu_858_p0 = { add_ln69_3_reg_1217[9], add_ln69_3_reg_1217[9], add_ln69_3_reg_1217[9], add_ln69_3_reg_1217[9], add_ln69_3_reg_1217[9], add_ln69_3_reg_1217[9], add_ln69_3_reg_1217[9], add_ln69_3_reg_1217[9], add_ln69_3_reg_1217[9], add_ln69_3_reg_1217[9], add_ln69_3_reg_1217[9], add_ln69_3_reg_1217[9], add_ln69_3_reg_1217[9], add_ln69_3_reg_1217[9], add_ln69_3_reg_1217[9], add_ln69_3_reg_1217[9], add_ln69_3_reg_1217[9], add_ln69_3_reg_1217[9], add_ln69_3_reg_1217[9], add_ln69_3_reg_1217[9], add_ln69_3_reg_1217[9], add_ln69_3_reg_1217[9], add_ln69_3_reg_1217 };
assign grp_fu_878_p0 = { op_30_V_reg_1227[31], op_30_V_reg_1227, 3'h0 };
assign grp_fu_878_p1 = { op_19[7], op_19[7], op_19[7], op_19[7], op_19[7], op_19[7], op_19[7], op_19[7], op_19[7], op_19[7], op_19[7], op_19[7], op_19[7], op_19[7], op_19[7], op_19[7], op_19[7], op_19[7], op_19[7], op_19[7], op_19[7], op_19[7], op_19[7], op_19[7], op_19[7], op_19[7], op_19[7], op_19[7], op_19 };
assign op_16_V_fu_807_p3 = { ret_V_reg_1192, 1'h0 };
assign p_Result_1_fu_269_p3 = op_8[15];
assign p_Result_2_fu_677_p3 = r_V_reg_1125[4];
assign p_Result_3_fu_416_p3 = ret_V_16_reg_970[32];
assign p_Result_4_fu_696_p3 = ret_V_17_reg_1108[33];
assign p_Result_5_fu_909_p3 = ret_V_19_reg_1247[35];
assign p_Result_7_fu_398_p3 = xor_ln731_fu_394_p2[1];
assign p_Result_8_fu_450_p3 = xor_ln1196_1_fu_438_p2[2];
assign p_Result_s_16_fu_510_p4 = { xor_ln1196_1_fu_438_p2[2], p_Val2_2_fu_504_p2 };
assign p_Val2_1_fu_443_p3 = { xor_ln731_reg_1039, 2'h0 };
assign ret_V_14_fu_351_p1 = op_4;
assign ret_V_2_fu_239_p4 = op_8[15:10];
assign rhs_1_fu_302_p3 = { op_21_V_reg_950, 11'h000 };
assign rhs_5_fu_867_p3 = { op_30_V_reg_1227, 3'h0 };
assign sext_ln1116_fu_620_p1 = { op_6_V_fu_614_p3[3], op_6_V_fu_614_p3 };
assign sext_ln1192_fu_298_p0 = op_10;
assign sext_ln1196_fu_435_p0 = op_2;
assign sext_ln1196_fu_435_p1 = { op_2[1], op_2 };
assign sext_ln1496_fu_726_p1 = { op_2[1], op_2, 1'h0 };
assign sext_ln1498_fu_743_p1 = { op_5[3], op_5 };
assign sext_ln69_3_fu_841_p1 = { op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17 };
assign sext_ln69_fu_288_p1 = { op_9[3], op_9[3], op_9[3], op_9 };
assign sext_ln703_1_fu_791_p0 = op_4;
assign sext_ln703_1_fu_791_p1 = { op_4[7], op_4 };
assign sext_ln703_2_fu_589_p0 = op_11;
assign sext_ln703_3_fu_863_p0 = op_19;
assign sext_ln703_fu_339_p0 = op_2;
assign sext_ln703_fu_339_p1 = { op_2[1], op_2[1], op_2[1], op_2[1], op_2[1], op_2[1], op_2 };
assign sext_ln831_fu_249_p1 = { op_8[15], op_8[15:10] };
assign sext_ln850_fu_375_p1 = { tmp_reg_975[21], tmp_reg_975 };
assign shl_ln728_1_fu_736_p1 = op_2;
assign shl_ln728_1_fu_736_p3 = { op_2, 3'h0 };
assign shl_ln_fu_719_p1 = op_2;
assign shl_ln_fu_719_p3 = { op_2, 1'h0 };
assign tmp_10_fu_593_p3 = { select_ln353_reg_1063, 1'h0 };
assign tmp_4_fu_477_p3 = xor_ln1196_1_fu_438_p2[2];
assign tmp_5_fu_485_p3 = xor_ln731_reg_1039[1];
assign trunc_ln1196_1_fu_347_p0 = op_4;
assign trunc_ln1196_1_fu_347_p1 = op_4[2:0];
assign trunc_ln1196_fu_343_p0 = op_4;
assign trunc_ln1196_fu_343_p1 = op_4[1:0];
assign trunc_ln851_1_fu_657_p1 = r_V_fu_640_p3[1:0];
assign trunc_ln851_2_fu_319_p0 = op_10;
assign trunc_ln851_2_fu_319_p1 = op_10[10:0];
assign trunc_ln851_3_fu_703_p0 = op_11;
assign trunc_ln851_3_fu_703_p1 = op_11[0];
assign trunc_ln851_4_fu_884_p0 = op_19;
assign trunc_ln851_4_fu_884_p1 = op_19[2:0];
assign trunc_ln851_fu_253_p1 = op_8[9:0];
assign xor_ln731_fu_394_p1 = op_2;
assign zext_ln69_1_fu_845_p1 = { 2'h0, op_18 };
assign zext_ln69_fu_766_p1 = { 1'h0, xor_ln1496_fu_761_p2 };
assign \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.ain_s0  = \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.a ;
assign \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.bin_s0  = \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.b ;
assign \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.s  = { \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.fas_s2 , \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.sum_s1  };
assign \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.u2.a  = \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.ain_s1 ;
assign \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.u2.b  = \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.bin_s1 ;
assign \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.u2.cin  = \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.carry_s1 ;
assign \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.facout_s2  = \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.u2.cout ;
assign \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.fas_s2  = \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.u2.s ;
assign \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.u1.a  = \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.a [17:0];
assign \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.u1.b  = \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.b [17:0];
assign \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.u1.cin  = 1'h0;
assign \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.facout_s1  = \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.u1.cout ;
assign \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.fas_s1  = \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.u1.s ;
assign \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.a  = \add_36s_36s_36_2_1_U9.din0 ;
assign \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.b  = \add_36s_36s_36_2_1_U9.din1 ;
assign \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.ce  = \add_36s_36s_36_2_1_U9.ce ;
assign \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.clk  = \add_36s_36s_36_2_1_U9.clk ;
assign \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.reset  = \add_36s_36s_36_2_1_U9.reset ;
assign \add_36s_36s_36_2_1_U9.dout  = \add_36s_36s_36_2_1_U9.top_add_36s_36s_36_2_1_Adder_7_U.s ;
assign \add_36s_36s_36_2_1_U9.ce  = 1'h1;
assign \add_36s_36s_36_2_1_U9.clk  = ap_clk;
assign \add_36s_36s_36_2_1_U9.din0  = { op_30_V_reg_1227[31], op_30_V_reg_1227, 3'h0 };
assign \add_36s_36s_36_2_1_U9.din1  = { op_19[7], op_19[7], op_19[7], op_19[7], op_19[7], op_19[7], op_19[7], op_19[7], op_19[7], op_19[7], op_19[7], op_19[7], op_19[7], op_19[7], op_19[7], op_19[7], op_19[7], op_19[7], op_19[7], op_19[7], op_19[7], op_19[7], op_19[7], op_19[7], op_19[7], op_19[7], op_19[7], op_19[7], op_19 };
assign grp_fu_878_p2 = \add_36s_36s_36_2_1_U9.dout ;
assign \add_36s_36s_36_2_1_U9.reset  = ap_rst;
assign \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.ain_s0  = \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.a ;
assign \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.bin_s0  = \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.b ;
assign \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.s  = { \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.fas_s2 , \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.sum_s1  };
assign \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.u2.a  = \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.ain_s1 ;
assign \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.u2.b  = \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.bin_s1 ;
assign \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.u2.cin  = \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.carry_s1 ;
assign \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.facout_s2  = \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.u2.cout ;
assign \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.fas_s2  = \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.u2.s ;
assign \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.u1.a  = \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.a [16:0];
assign \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.u1.b  = \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.b [16:0];
assign \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.u1.cin  = 1'h0;
assign \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.facout_s1  = \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.u1.cout ;
assign \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.fas_s1  = \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.u1.s ;
assign \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.a  = \add_34s_34s_34_2_1_U3.din0 ;
assign \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.b  = \add_34s_34s_34_2_1_U3.din1 ;
assign \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.ce  = \add_34s_34s_34_2_1_U3.ce ;
assign \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.clk  = \add_34s_34s_34_2_1_U3.clk ;
assign \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.reset  = \add_34s_34s_34_2_1_U3.reset ;
assign \add_34s_34s_34_2_1_U3.dout  = \add_34s_34s_34_2_1_U3.top_add_34s_34s_34_2_1_Adder_2_U.s ;
assign \add_34s_34s_34_2_1_U3.ce  = 1'h1;
assign \add_34s_34s_34_2_1_U3.clk  = ap_clk;
assign \add_34s_34s_34_2_1_U3.din0  = { select_ln353_reg_1063[22], select_ln353_reg_1063[22], select_ln353_reg_1063[22], select_ln353_reg_1063[22], select_ln353_reg_1063[22], select_ln353_reg_1063[22], select_ln353_reg_1063[22], select_ln353_reg_1063[22], select_ln353_reg_1063[22], select_ln353_reg_1063[22], select_ln353_reg_1063, 1'h0 };
assign \add_34s_34s_34_2_1_U3.din1  = { op_11[1], op_11[1], op_11[1], op_11[1], op_11[1], op_11[1], op_11[1], op_11[1], op_11[1], op_11[1], op_11[1], op_11[1], op_11[1], op_11[1], op_11[1], op_11[1], op_11[1], op_11[1], op_11[1], op_11[1], op_11[1], op_11[1], op_11[1], op_11[1], op_11[1], op_11[1], op_11[1], op_11[1], op_11[1], op_11[1], op_11[1], op_11[1], op_11 };
assign grp_fu_604_p2 = \add_34s_34s_34_2_1_U3.dout ;
assign \add_34s_34s_34_2_1_U3.reset  = ap_rst;
assign \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.ain_s0  = \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.a ;
assign \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.bin_s0  = \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.b ;
assign \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.s  = { \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.fas_s2 , \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.sum_s1  };
assign \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.u2.a  = \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.ain_s1 ;
assign \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.u2.b  = \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.bin_s1 ;
assign \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.u2.cin  = \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.carry_s1 ;
assign \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.facout_s2  = \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.u2.cout ;
assign \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.fas_s2  = \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.u2.s ;
assign \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.u1.a  = \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.a [15:0];
assign \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.u1.b  = \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.b [15:0];
assign \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.u1.cin  = 1'h0;
assign \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.facout_s1  = \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.u1.cout ;
assign \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.fas_s1  = \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.u1.s ;
assign \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.a  = \add_33s_33s_33_2_1_U1.din0 ;
assign \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.b  = \add_33s_33s_33_2_1_U1.din1 ;
assign \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.ce  = \add_33s_33s_33_2_1_U1.ce ;
assign \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.clk  = \add_33s_33s_33_2_1_U1.clk ;
assign \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.reset  = \add_33s_33s_33_2_1_U1.reset ;
assign \add_33s_33s_33_2_1_U1.dout  = \add_33s_33s_33_2_1_U1.top_add_33s_33s_33_2_1_Adder_0_U.s ;
assign \add_33s_33s_33_2_1_U1.ce  = 1'h1;
assign \add_33s_33s_33_2_1_U1.clk  = ap_clk;
assign \add_33s_33s_33_2_1_U1.din0  = { op_21_V_reg_950[6], op_21_V_reg_950[6], op_21_V_reg_950[6], op_21_V_reg_950[6], op_21_V_reg_950[6], op_21_V_reg_950[6], op_21_V_reg_950[6], op_21_V_reg_950[6], op_21_V_reg_950[6], op_21_V_reg_950[6], op_21_V_reg_950[6], op_21_V_reg_950[6], op_21_V_reg_950[6], op_21_V_reg_950[6], op_21_V_reg_950[6], op_21_V_reg_950, 11'h000 };
assign \add_33s_33s_33_2_1_U1.din1  = { op_10[31], op_10 };
assign grp_fu_313_p2 = \add_33s_33s_33_2_1_U1.dout ;
assign \add_33s_33s_33_2_1_U1.reset  = ap_rst;
assign \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.ain_s0  = \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.a ;
assign \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.bin_s0  = \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.b ;
assign \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.s  = { \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.fas_s2 , \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.sum_s1  };
assign \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.u2.a  = \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.ain_s1 ;
assign \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.u2.b  = \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.bin_s1 ;
assign \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.u2.cin  = \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.carry_s1 ;
assign \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.facout_s2  = \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.u2.cout ;
assign \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.fas_s2  = \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.u2.s ;
assign \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.u1.a  = \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.a [15:0];
assign \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.u1.b  = \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.b [15:0];
assign \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.u1.cin  = 1'h0;
assign \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.facout_s1  = \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.u1.cout ;
assign \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.fas_s1  = \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.u1.s ;
assign \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.a  = \add_33ns_33s_33_2_1_U7.din0 ;
assign \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.b  = \add_33ns_33s_33_2_1_U7.din1 ;
assign \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.ce  = \add_33ns_33s_33_2_1_U7.ce ;
assign \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.clk  = \add_33ns_33s_33_2_1_U7.clk ;
assign \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.reset  = \add_33ns_33s_33_2_1_U7.reset ;
assign \add_33ns_33s_33_2_1_U7.dout  = \add_33ns_33s_33_2_1_U7.top_add_33ns_33s_33_2_1_Adder_6_U.s ;
assign \add_33ns_33s_33_2_1_U7.ce  = 1'h1;
assign \add_33ns_33s_33_2_1_U7.clk  = ap_clk;
assign \add_33ns_33s_33_2_1_U7.din0  = { op_27_V_reg_1197, 1'h0 };
assign \add_33ns_33s_33_2_1_U7.din1  = { ret_V_reg_1192[8], ret_V_reg_1192[8], ret_V_reg_1192[8], ret_V_reg_1192[8], ret_V_reg_1192[8], ret_V_reg_1192[8], ret_V_reg_1192[8], ret_V_reg_1192[8], ret_V_reg_1192[8], ret_V_reg_1192[8], ret_V_reg_1192[8], ret_V_reg_1192[8], ret_V_reg_1192[8], ret_V_reg_1192[8], ret_V_reg_1192[8], ret_V_reg_1192[8], ret_V_reg_1192[8], ret_V_reg_1192[8], ret_V_reg_1192[8], ret_V_reg_1192[8], ret_V_reg_1192[8], ret_V_reg_1192[8], ret_V_reg_1192[8], ret_V_reg_1192, 1'h0 };
assign grp_fu_825_p2 = \add_33ns_33s_33_2_1_U7.dout ;
assign \add_33ns_33s_33_2_1_U7.reset  = ap_rst;
assign \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.ain_s0  = \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.a ;
assign \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.bin_s0  = \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.b ;
assign \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.s  = { \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.fas_s2 , \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.sum_s1  };
assign \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.u2.a  = \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.ain_s1 ;
assign \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.u2.b  = \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.bin_s1 ;
assign \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.u2.cin  = \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.carry_s1 ;
assign \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.facout_s2  = \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.u2.cout ;
assign \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.fas_s2  = \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.u2.s ;
assign \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.u1.a  = \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.a [15:0];
assign \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.u1.b  = \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.b [15:0];
assign \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.u1.cin  = 1'h0;
assign \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.facout_s1  = \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.u1.cout ;
assign \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.fas_s1  = \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.u1.s ;
assign \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.a  = \add_32s_32ns_32_2_1_U8.din0 ;
assign \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.b  = \add_32s_32ns_32_2_1_U8.din1 ;
assign \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.ce  = \add_32s_32ns_32_2_1_U8.ce ;
assign \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.clk  = \add_32s_32ns_32_2_1_U8.clk ;
assign \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.reset  = \add_32s_32ns_32_2_1_U8.reset ;
assign \add_32s_32ns_32_2_1_U8.dout  = \add_32s_32ns_32_2_1_U8.top_add_32s_32ns_32_2_1_Adder_5_U.s ;
assign \add_32s_32ns_32_2_1_U8.ce  = 1'h1;
assign \add_32s_32ns_32_2_1_U8.clk  = ap_clk;
assign \add_32s_32ns_32_2_1_U8.din0  = { add_ln69_3_reg_1217[9], add_ln69_3_reg_1217[9], add_ln69_3_reg_1217[9], add_ln69_3_reg_1217[9], add_ln69_3_reg_1217[9], add_ln69_3_reg_1217[9], add_ln69_3_reg_1217[9], add_ln69_3_reg_1217[9], add_ln69_3_reg_1217[9], add_ln69_3_reg_1217[9], add_ln69_3_reg_1217[9], add_ln69_3_reg_1217[9], add_ln69_3_reg_1217[9], add_ln69_3_reg_1217[9], add_ln69_3_reg_1217[9], add_ln69_3_reg_1217[9], add_ln69_3_reg_1217[9], add_ln69_3_reg_1217[9], add_ln69_3_reg_1217[9], add_ln69_3_reg_1217[9], add_ln69_3_reg_1217[9], add_ln69_3_reg_1217[9], add_ln69_3_reg_1217 };
assign \add_32s_32ns_32_2_1_U8.din1  = op_28_V_reg_1212;
assign grp_fu_858_p2 = \add_32s_32ns_32_2_1_U8.dout ;
assign \add_32s_32ns_32_2_1_U8.reset  = ap_rst;
assign \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.ain_s0  = \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.a ;
assign \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.bin_s0  = \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.b ;
assign \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.s  = { \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.fas_s2 , \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.sum_s1  };
assign \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.u2.a  = \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.ain_s1 ;
assign \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.u2.b  = \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.bin_s1 ;
assign \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.u2.cin  = \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.carry_s1 ;
assign \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.facout_s2  = \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.u2.cout ;
assign \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.fas_s2  = \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.u2.s ;
assign \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.u1.a  = \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.a [15:0];
assign \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.u1.b  = \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.b [15:0];
assign \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.u1.cin  = 1'h0;
assign \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.facout_s1  = \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.u1.cout ;
assign \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.fas_s1  = \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.u1.s ;
assign \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.a  = \add_32s_32ns_32_2_1_U6.din0 ;
assign \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.b  = \add_32s_32ns_32_2_1_U6.din1 ;
assign \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.ce  = \add_32s_32ns_32_2_1_U6.ce ;
assign \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.clk  = \add_32s_32ns_32_2_1_U6.clk ;
assign \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.reset  = \add_32s_32ns_32_2_1_U6.reset ;
assign \add_32s_32ns_32_2_1_U6.dout  = \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.s ;
assign \add_32s_32ns_32_2_1_U6.ce  = 1'h1;
assign \add_32s_32ns_32_2_1_U6.clk  = ap_clk;
assign \add_32s_32ns_32_2_1_U6.din0  = { add_ln69_1_reg_1182[1], add_ln69_1_reg_1182[1], add_ln69_1_reg_1182[1], add_ln69_1_reg_1182[1], add_ln69_1_reg_1182[1], add_ln69_1_reg_1182[1], add_ln69_1_reg_1182[1], add_ln69_1_reg_1182[1], add_ln69_1_reg_1182[1], add_ln69_1_reg_1182[1], add_ln69_1_reg_1182[1], add_ln69_1_reg_1182[1], add_ln69_1_reg_1182[1], add_ln69_1_reg_1182[1], add_ln69_1_reg_1182[1], add_ln69_1_reg_1182[1], add_ln69_1_reg_1182[1], add_ln69_1_reg_1182[1], add_ln69_1_reg_1182[1], add_ln69_1_reg_1182[1], add_ln69_1_reg_1182[1], add_ln69_1_reg_1182[1], add_ln69_1_reg_1182[1], add_ln69_1_reg_1182[1], add_ln69_1_reg_1182[1], add_ln69_1_reg_1182[1], add_ln69_1_reg_1182[1], add_ln69_1_reg_1182[1], add_ln69_1_reg_1182[1], add_ln69_1_reg_1182[1], add_ln69_1_reg_1182 };
assign \add_32s_32ns_32_2_1_U6.din1  = add_ln69_reg_1177;
assign grp_fu_786_p2 = \add_32s_32ns_32_2_1_U6.dout ;
assign \add_32s_32ns_32_2_1_U6.reset  = ap_rst;
assign \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.ain_s0  = \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.a ;
assign \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.bin_s0  = \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.b ;
assign \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.s  = { \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.fas_s2 , \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.sum_s1  };
assign \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.u2.a  = \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.ain_s1 ;
assign \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.u2.b  = \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.bin_s1 ;
assign \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.u2.cin  = \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.carry_s1 ;
assign \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.facout_s2  = \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.u2.cout ;
assign \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.fas_s2  = \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.u2.s ;
assign \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.u1.a  = \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.a [15:0];
assign \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.u1.b  = \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.b [15:0];
assign \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.u1.cin  = 1'h0;
assign \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.facout_s1  = \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.u1.cout ;
assign \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.fas_s1  = \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.u1.s ;
assign \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.a  = \add_32ns_32s_32_2_1_U5.din0 ;
assign \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.b  = \add_32ns_32s_32_2_1_U5.din1 ;
assign \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.ce  = \add_32ns_32s_32_2_1_U5.ce ;
assign \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.clk  = \add_32ns_32s_32_2_1_U5.clk ;
assign \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.reset  = \add_32ns_32s_32_2_1_U5.reset ;
assign \add_32ns_32s_32_2_1_U5.dout  = \add_32ns_32s_32_2_1_U5.top_add_32ns_32s_32_2_1_Adder_4_U.s ;
assign \add_32ns_32s_32_2_1_U5.ce  = 1'h1;
assign \add_32ns_32s_32_2_1_U5.clk  = ap_clk;
assign \add_32ns_32s_32_2_1_U5.din0  = ret_V_18_reg_1157;
assign \add_32ns_32s_32_2_1_U5.din1  = { ret_V_7_reg_1152[2], ret_V_7_reg_1152[2], ret_V_7_reg_1152[2], ret_V_7_reg_1152[2], ret_V_7_reg_1152[2], ret_V_7_reg_1152[2], ret_V_7_reg_1152[2], ret_V_7_reg_1152[2], ret_V_7_reg_1152[2], ret_V_7_reg_1152[2], ret_V_7_reg_1152[2], ret_V_7_reg_1152[2], ret_V_7_reg_1152[2], ret_V_7_reg_1152[2], ret_V_7_reg_1152[2], ret_V_7_reg_1152[2], ret_V_7_reg_1152[2], ret_V_7_reg_1152[2], ret_V_7_reg_1152[2], ret_V_7_reg_1152[2], ret_V_7_reg_1152[2], ret_V_7_reg_1152[2], ret_V_7_reg_1152[2], ret_V_7_reg_1152[2], ret_V_7_reg_1152[2], ret_V_7_reg_1152[2], ret_V_7_reg_1152[2], ret_V_7_reg_1152[2], ret_V_7_reg_1152[2], ret_V_7_reg_1152 };
assign grp_fu_756_p2 = \add_32ns_32s_32_2_1_U5.dout ;
assign \add_32ns_32s_32_2_1_U5.reset  = ap_rst;
assign \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.ain_s0  = \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.a ;
assign \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.bin_s0  = \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.b ;
assign \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.s  = { \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.fas_s2 , \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.sum_s1  };
assign \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.u2.a  = \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.ain_s1 ;
assign \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.u2.b  = \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.bin_s1 ;
assign \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.u2.cin  = \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.carry_s1 ;
assign \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.facout_s2  = \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.u2.cout ;
assign \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.fas_s2  = \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.u2.s ;
assign \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.u1.a  = \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.a [15:0];
assign \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.u1.b  = \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.b [15:0];
assign \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.u1.cin  = 1'h0;
assign \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.facout_s1  = \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.u1.cout ;
assign \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.fas_s1  = \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.u1.s ;
assign \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.a  = \add_32ns_32ns_32_2_1_U4.din0 ;
assign \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.b  = \add_32ns_32ns_32_2_1_U4.din1 ;
assign \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.ce  = \add_32ns_32ns_32_2_1_U4.ce ;
assign \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.clk  = \add_32ns_32ns_32_2_1_U4.clk ;
assign \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.reset  = \add_32ns_32ns_32_2_1_U4.reset ;
assign \add_32ns_32ns_32_2_1_U4.dout  = \add_32ns_32ns_32_2_1_U4.top_add_32ns_32ns_32_2_1_Adder_3_U.s ;
assign \add_32ns_32ns_32_2_1_U4.ce  = 1'h1;
assign \add_32ns_32ns_32_2_1_U4.clk  = ap_clk;
assign \add_32ns_32ns_32_2_1_U4.din0  = ret_V_12_cast_reg_1113;
assign \add_32ns_32ns_32_2_1_U4.din1  = 32'd1;
assign grp_fu_667_p2 = \add_32ns_32ns_32_2_1_U4.dout ;
assign \add_32ns_32ns_32_2_1_U4.reset  = ap_rst;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.ain_s0  = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.a ;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.bin_s0  = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.b ;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.s  = { \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.fas_s2 , \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.sum_s1  };
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.u2.a  = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.ain_s1 ;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.u2.b  = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.bin_s1 ;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.u2.cin  = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.carry_s1 ;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.facout_s2  = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.u2.cout ;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.fas_s2  = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.u2.s ;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.u1.a  = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.a [15:0];
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.u1.b  = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.b [15:0];
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.u1.cin  = 1'h0;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.facout_s1  = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.u1.cout ;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.fas_s1  = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.u1.s ;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.a  = \add_32ns_32ns_32_2_1_U10.din0 ;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.b  = \add_32ns_32ns_32_2_1_U10.din1 ;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.ce  = \add_32ns_32ns_32_2_1_U10.ce ;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.clk  = \add_32ns_32ns_32_2_1_U10.clk ;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.reset  = \add_32ns_32ns_32_2_1_U10.reset ;
assign \add_32ns_32ns_32_2_1_U10.dout  = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_3_U.s ;
assign \add_32ns_32ns_32_2_1_U10.ce  = 1'h1;
assign \add_32ns_32ns_32_2_1_U10.clk  = ap_clk;
assign \add_32ns_32ns_32_2_1_U10.din0  = ret_V_16_cast_reg_1252;
assign \add_32ns_32ns_32_2_1_U10.din1  = 32'd1;
assign grp_fu_904_p2 = \add_32ns_32ns_32_2_1_U10.dout ;
assign \add_32ns_32ns_32_2_1_U10.reset  = ap_rst;
assign \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.ain_s0  = \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.a ;
assign \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.bin_s0  = \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.b ;
assign \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.s  = { \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.fas_s2 , \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.sum_s1  };
assign \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.u2.a  = \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.ain_s1 ;
assign \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.u2.b  = \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.bin_s1 ;
assign \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.u2.cin  = \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.carry_s1 ;
assign \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.facout_s2  = \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.u2.cout ;
assign \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.fas_s2  = \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.u2.s ;
assign \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.u1.a  = \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.a [10:0];
assign \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.u1.b  = \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.b [10:0];
assign \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.u1.cin  = 1'h0;
assign \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.facout_s1  = \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.u1.cout ;
assign \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.fas_s1  = \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.u1.s ;
assign \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.a  = \add_23s_23ns_23_2_1_U2.din0 ;
assign \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.b  = \add_23s_23ns_23_2_1_U2.din1 ;
assign \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.ce  = \add_23s_23ns_23_2_1_U2.ce ;
assign \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.clk  = \add_23s_23ns_23_2_1_U2.clk ;
assign \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.reset  = \add_23s_23ns_23_2_1_U2.reset ;
assign \add_23s_23ns_23_2_1_U2.dout  = \add_23s_23ns_23_2_1_U2.top_add_23s_23ns_23_2_1_Adder_1_U.s ;
assign \add_23s_23ns_23_2_1_U2.ce  = 1'h1;
assign \add_23s_23ns_23_2_1_U2.clk  = ap_clk;
assign \add_23s_23ns_23_2_1_U2.din0  = { tmp_reg_975[21], tmp_reg_975 };
assign \add_23s_23ns_23_2_1_U2.din1  = 23'h000001;
assign grp_fu_378_p2 = \add_23s_23ns_23_2_1_U2.dout ;
assign \add_23s_23ns_23_2_1_U2.reset  = ap_rst;
endmodule


// Product machine:
module top_A_times_top_B (ap_start, op_0, op_10, op_11, op_17, op_18, op_19, op_2, op_3, op_4, op_5, op_7, op_8, op_9, ap_clk, unsafe_signal);
input ap_start;
input [1:0] op_0;
input [31:0] op_10;
input [1:0] op_11;
input [3:0] op_17;
input [7:0] op_18;
input [7:0] op_19;
input [1:0] op_2;
input [3:0] op_3;
input [7:0] op_4;
input [3:0] op_5;
input op_7;
input [15:0] op_8;
input [3:0] op_9;
input ap_clk;
output unsafe_signal;
reg _setup;
initial _setup = 1'b0;
always @ (posedge ap_clk) _setup <= 1'b1;
reg ap_start_internal;
always @ (posedge ap_clk) if (!_setup) ap_start_internal <= ap_start;
reg [1:0] op_0_internal;
always @ (posedge ap_clk) if (!_setup) op_0_internal <= op_0;
reg [31:0] op_10_internal;
always @ (posedge ap_clk) if (!_setup) op_10_internal <= op_10;
reg [1:0] op_11_internal;
always @ (posedge ap_clk) if (!_setup) op_11_internal <= op_11;
reg [3:0] op_17_internal;
always @ (posedge ap_clk) if (!_setup) op_17_internal <= op_17;
reg [7:0] op_18_internal;
always @ (posedge ap_clk) if (!_setup) op_18_internal <= op_18;
reg [7:0] op_19_internal;
always @ (posedge ap_clk) if (!_setup) op_19_internal <= op_19;
reg [1:0] op_2_internal;
always @ (posedge ap_clk) if (!_setup) op_2_internal <= op_2;
reg [3:0] op_3_internal;
always @ (posedge ap_clk) if (!_setup) op_3_internal <= op_3;
reg [7:0] op_4_internal;
always @ (posedge ap_clk) if (!_setup) op_4_internal <= op_4;
reg [3:0] op_5_internal;
always @ (posedge ap_clk) if (!_setup) op_5_internal <= op_5;
reg op_7_internal;
always @ (posedge ap_clk) if (!_setup) op_7_internal <= op_7;
reg [15:0] op_8_internal;
always @ (posedge ap_clk) if (!_setup) op_8_internal <= op_8;
reg [3:0] op_9_internal;
always @ (posedge ap_clk) if (!_setup) op_9_internal <= op_9;
wire ap_done_A;
wire ap_done_B;
wire ap_done_eq;
assign ap_done_eq = ap_done_A == ap_done_B;
wire ap_idle_A;
wire ap_idle_B;
wire ap_idle_eq;
assign ap_idle_eq = ap_idle_A == ap_idle_B;
wire ap_ready_A;
wire ap_ready_B;
wire ap_ready_eq;
assign ap_ready_eq = ap_ready_A == ap_ready_B;
wire [31:0] op_31_A;
wire [31:0] op_31_B;
wire op_31_eq;
assign op_31_eq = op_31_A == op_31_B;
wire op_31_ap_vld_A;
wire op_31_ap_vld_B;
wire clk_enable_A;
wire clk_enable_B;
assign clk_enable_A = _setup & (~op_31_ap_vld_A | op_31_ap_vld_B);
assign clk_enable_B = _setup;
wire divergent;
assign divergent = ~(ap_done_eq & ap_idle_eq & ap_ready_eq & op_31_eq);
assign unsafe_signal = op_31_ap_vld_A & op_31_ap_vld_B & divergent;
top_A instance_A (
    .ap_clk(ap_clk),
    .clk_enable(clk_enable_A),
    .ap_start(ap_start_internal),
    .op_0(op_0_internal),
    .op_10(op_10_internal),
    .op_11(op_11_internal),
    .op_17(op_17_internal),
    .op_18(op_18_internal),
    .op_19(op_19_internal),
    .op_2(op_2_internal),
    .op_3(op_3_internal),
    .op_4(op_4_internal),
    .op_5(op_5_internal),
    .op_7(op_7_internal),
    .op_8(op_8_internal),
    .op_9(op_9_internal),
    .ap_done(ap_done_A),
    .ap_idle(ap_idle_A),
    .ap_ready(ap_ready_A),
    .op_31(op_31_A),
    .op_31_ap_vld(op_31_ap_vld_A)
);
top_B instance_B (
    .ap_clk(ap_clk),
    .clk_enable(clk_enable_B),
    .ap_start(ap_start_internal),
    .op_0(op_0_internal),
    .op_10(op_10_internal),
    .op_11(op_11_internal),
    .op_17(op_17_internal),
    .op_18(op_18_internal),
    .op_19(op_19_internal),
    .op_2(op_2_internal),
    .op_3(op_3_internal),
    .op_4(op_4_internal),
    .op_5(op_5_internal),
    .op_7(op_7_internal),
    .op_8(op_8_internal),
    .op_9(op_9_internal),
    .ap_done(ap_done_B),
    .ap_idle(ap_idle_B),
    .ap_ready(ap_ready_B),
    .op_31(op_31_B),
    .op_31_ap_vld(op_31_ap_vld_B)
);
endmodule
