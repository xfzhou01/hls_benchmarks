// Processed by function `construct_kairos` in `verilog_tricks.py`.
// Machine A:
// Processed by function `add_clk_enable_signal` in `verilog_tricks.py`.
// Processed by function `remove_reset_signal` in `verilog_tricks.py`.
module top_A (
  ap_clk,
  ap_start,
  ap_done,
  ap_idle,
  ap_ready,
  op_0,
  op_1,
  op_2,
  op_3,
  op_4,
  op_5,
  op_7,
  op_8,
  op_13,
  op_15,
  op_16,
  op_17,
  op_30,
  op_30_ap_vld,
clk_enable
);
input clk_enable;


input ap_clk;
wire ap_rst;
assign ap_rst = op_30_ap_vld;
input ap_start;
input [1:0] op_0;
input [7:0] op_1;
input [7:0] op_13;
input [7:0] op_15;
input [3:0] op_16;
input [3:0] op_17;
input [1:0] op_2;
input [7:0] op_3;
input [15:0] op_4;
input [3:0] op_5;
input [1:0] op_7;
input [1:0] op_8;
output ap_done;
output ap_idle;
output ap_ready;
output [31:0] op_30;
output op_30_ap_vld;


reg [4:0] \add_10ns_10s_10_2_1_U18.top_add_10ns_10s_10_2_1_Adder_12_U.ain_s1 ;
reg [4:0] \add_10ns_10s_10_2_1_U18.top_add_10ns_10s_10_2_1_Adder_12_U.bin_s1 ;
reg \add_10ns_10s_10_2_1_U18.top_add_10ns_10s_10_2_1_Adder_12_U.carry_s1 ;
reg [4:0] \add_10ns_10s_10_2_1_U18.top_add_10ns_10s_10_2_1_Adder_12_U.sum_s1 ;
reg [5:0] \add_11s_11s_11_2_1_U17.top_add_11s_11s_11_2_1_Adder_11_U.ain_s1 ;
reg [5:0] \add_11s_11s_11_2_1_U17.top_add_11s_11s_11_2_1_Adder_11_U.bin_s1 ;
reg \add_11s_11s_11_2_1_U17.top_add_11s_11s_11_2_1_Adder_11_U.carry_s1 ;
reg [4:0] \add_11s_11s_11_2_1_U17.top_add_11s_11s_11_2_1_Adder_11_U.sum_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.ain_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.bin_s1 ;
reg \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.carry_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.sum_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.ain_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.bin_s1 ;
reg \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.carry_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.sum_s1 ;
reg [15:0] \add_32ns_32s_32_2_1_U24.top_add_32ns_32s_32_2_1_Adder_17_U.ain_s1 ;
reg [15:0] \add_32ns_32s_32_2_1_U24.top_add_32ns_32s_32_2_1_Adder_17_U.bin_s1 ;
reg \add_32ns_32s_32_2_1_U24.top_add_32ns_32s_32_2_1_Adder_17_U.carry_s1 ;
reg [15:0] \add_32ns_32s_32_2_1_U24.top_add_32ns_32s_32_2_1_Adder_17_U.sum_s1 ;
reg [15:0] \add_32ns_32s_32_2_1_U25.top_add_32ns_32s_32_2_1_Adder_17_U.ain_s1 ;
reg [15:0] \add_32ns_32s_32_2_1_U25.top_add_32ns_32s_32_2_1_Adder_17_U.bin_s1 ;
reg \add_32ns_32s_32_2_1_U25.top_add_32ns_32s_32_2_1_Adder_17_U.carry_s1 ;
reg [15:0] \add_32ns_32s_32_2_1_U25.top_add_32ns_32s_32_2_1_Adder_17_U.sum_s1 ;
reg [15:0] \add_32s_32ns_32_2_1_U26.top_add_32s_32ns_32_2_1_Adder_18_U.ain_s1 ;
reg [15:0] \add_32s_32ns_32_2_1_U26.top_add_32s_32ns_32_2_1_Adder_18_U.bin_s1 ;
reg \add_32s_32ns_32_2_1_U26.top_add_32s_32ns_32_2_1_Adder_18_U.carry_s1 ;
reg [15:0] \add_32s_32ns_32_2_1_U26.top_add_32s_32ns_32_2_1_Adder_18_U.sum_s1 ;
reg [18:0] \add_38s_38s_38_2_1_U22.top_add_38s_38s_38_2_1_Adder_16_U.ain_s1 ;
reg [18:0] \add_38s_38s_38_2_1_U22.top_add_38s_38s_38_2_1_Adder_16_U.bin_s1 ;
reg \add_38s_38s_38_2_1_U22.top_add_38s_38s_38_2_1_Adder_16_U.carry_s1 ;
reg [18:0] \add_38s_38s_38_2_1_U22.top_add_38s_38s_38_2_1_Adder_16_U.sum_s1 ;
reg [1:0] \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_9_U.ain_s1 ;
reg [1:0] \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_9_U.bin_s1 ;
reg \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_9_U.carry_s1 ;
reg \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_9_U.sum_s1 ;
reg [1:0] \add_3s_3s_3_2_1_U6.top_add_3s_3s_3_2_1_Adder_2_U.ain_s1 ;
reg [1:0] \add_3s_3s_3_2_1_U6.top_add_3s_3s_3_2_1_Adder_2_U.bin_s1 ;
reg \add_3s_3s_3_2_1_U6.top_add_3s_3s_3_2_1_Adder_2_U.carry_s1 ;
reg \add_3s_3s_3_2_1_U6.top_add_3s_3s_3_2_1_Adder_2_U.sum_s1 ;
reg [19:0] \add_40s_40s_40_2_1_U20.top_add_40s_40s_40_2_1_Adder_14_U.ain_s1 ;
reg [19:0] \add_40s_40s_40_2_1_U20.top_add_40s_40s_40_2_1_Adder_14_U.bin_s1 ;
reg \add_40s_40s_40_2_1_U20.top_add_40s_40s_40_2_1_Adder_14_U.carry_s1 ;
reg [19:0] \add_40s_40s_40_2_1_U20.top_add_40s_40s_40_2_1_Adder_14_U.sum_s1 ;
reg [1:0] \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_7_U.ain_s1 ;
reg [1:0] \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_7_U.bin_s1 ;
reg \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_7_U.carry_s1 ;
reg [1:0] \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_7_U.sum_s1 ;
reg [2:0] \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_3_U.ain_s1 ;
reg [2:0] \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_3_U.bin_s1 ;
reg \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_3_U.carry_s1 ;
reg [1:0] \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_3_U.sum_s1 ;
reg [2:0] \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_6_U.ain_s1 ;
reg [2:0] \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_6_U.bin_s1 ;
reg \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_6_U.carry_s1 ;
reg [2:0] \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_6_U.sum_s1 ;
reg [3:0] \add_7ns_7ns_7_2_1_U16.top_add_7ns_7ns_7_2_1_Adder_10_U.ain_s1 ;
reg [3:0] \add_7ns_7ns_7_2_1_U16.top_add_7ns_7ns_7_2_1_Adder_10_U.bin_s1 ;
reg \add_7ns_7ns_7_2_1_U16.top_add_7ns_7ns_7_2_1_Adder_10_U.carry_s1 ;
reg [2:0] \add_7ns_7ns_7_2_1_U16.top_add_7ns_7ns_7_2_1_Adder_10_U.sum_s1 ;
reg [3:0] \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_8_U.ain_s1 ;
reg [3:0] \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_8_U.bin_s1 ;
reg \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_8_U.carry_s1 ;
reg [2:0] \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_8_U.sum_s1 ;
reg [4:0] \add_9ns_9s_9_2_1_U9.top_add_9ns_9s_9_2_1_Adder_5_U.ain_s1 ;
reg [4:0] \add_9ns_9s_9_2_1_U9.top_add_9ns_9s_9_2_1_Adder_5_U.bin_s1 ;
reg \add_9ns_9s_9_2_1_U9.top_add_9ns_9s_9_2_1_Adder_5_U.carry_s1 ;
reg [3:0] \add_9ns_9s_9_2_1_U9.top_add_9ns_9s_9_2_1_Adder_5_U.sum_s1 ;
reg [4:0] \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_13_U.ain_s1 ;
reg [4:0] \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_13_U.bin_s1 ;
reg \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_13_U.carry_s1 ;
reg [3:0] \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_13_U.sum_s1 ;
reg [31:0] add_ln691_1_reg_1491;
reg [31:0] add_ln691_2_reg_1528;
reg [8:0] add_ln691_reg_1454;
reg [2:0] add_ln69_1_reg_1362;
reg [9:0] add_ln69_3_reg_1442;
reg [6:0] add_ln69_reg_1357;
reg and_ln786_reg_1326;
reg [37:0] ap_CS_fsm = 38'h0000000001;
reg [3:0] \ashr_16s_4ns_16_7_1_U4.din1_cast_array[0] ;
reg [3:0] \ashr_16s_4ns_16_7_1_U4.din1_cast_array[1] ;
reg [3:0] \ashr_16s_4ns_16_7_1_U4.din1_cast_array[2] ;
reg [3:0] \ashr_16s_4ns_16_7_1_U4.din1_cast_array[3] ;
reg [3:0] \ashr_16s_4ns_16_7_1_U4.din1_cast_array[4] ;
reg [3:0] \ashr_16s_4ns_16_7_1_U4.din1_cast_array[5] ;
reg [15:0] \ashr_16s_4ns_16_7_1_U4.dout_array[0] ;
reg [15:0] \ashr_16s_4ns_16_7_1_U4.dout_array[1] ;
reg [15:0] \ashr_16s_4ns_16_7_1_U4.dout_array[2] ;
reg [15:0] \ashr_16s_4ns_16_7_1_U4.dout_array[3] ;
reg [15:0] \ashr_16s_4ns_16_7_1_U4.dout_array[4] ;
reg [15:0] \ashr_16s_4ns_16_7_1_U4.dout_array[5] ;
reg [7:0] \ashr_8ns_8s_8_7_1_U11.din1_cast_array[0] ;
reg [7:0] \ashr_8ns_8s_8_7_1_U11.din1_cast_array[1] ;
reg [7:0] \ashr_8ns_8s_8_7_1_U11.din1_cast_array[2] ;
reg [7:0] \ashr_8ns_8s_8_7_1_U11.din1_cast_array[3] ;
reg [7:0] \ashr_8ns_8s_8_7_1_U11.din1_cast_array[4] ;
reg [7:0] \ashr_8ns_8s_8_7_1_U11.din1_cast_array[5] ;
reg [7:0] \ashr_8ns_8s_8_7_1_U11.dout_array[0] ;
reg [7:0] \ashr_8ns_8s_8_7_1_U11.dout_array[1] ;
reg [7:0] \ashr_8ns_8s_8_7_1_U11.dout_array[2] ;
reg [7:0] \ashr_8ns_8s_8_7_1_U11.dout_array[3] ;
reg [7:0] \ashr_8ns_8s_8_7_1_U11.dout_array[4] ;
reg [7:0] \ashr_8ns_8s_8_7_1_U11.dout_array[5] ;
reg [15:0] ashr_ln1333_reg_1194;
reg [7:0] ashr_ln799_reg_1377;
reg icmp_ln1494_reg_1131;
reg icmp_ln1499_reg_1082;
reg icmp_ln768_reg_1271;
reg icmp_ln786_reg_1276;
reg icmp_ln851_1_reg_1261;
reg icmp_ln851_2_reg_1422;
reg icmp_ln851_3_reg_1474;
reg icmp_ln851_4_reg_1511;
reg icmp_ln851_reg_1167;
reg isNeg_reg_1033;
reg [15:0] \mul_16s_2s_18_7_1_U5.top_mul_16s_2s_18_7_1_Mul_DSP_0_U.a_reg0 ;
reg [1:0] \mul_16s_2s_18_7_1_U5.top_mul_16s_2s_18_7_1_Mul_DSP_0_U.b_reg0 ;
reg [17:0] \mul_16s_2s_18_7_1_U5.top_mul_16s_2s_18_7_1_Mul_DSP_0_U.buff0 ;
reg [17:0] \mul_16s_2s_18_7_1_U5.top_mul_16s_2s_18_7_1_Mul_DSP_0_U.buff1 ;
reg [17:0] \mul_16s_2s_18_7_1_U5.top_mul_16s_2s_18_7_1_Mul_DSP_0_U.buff2 ;
reg [17:0] \mul_16s_2s_18_7_1_U5.top_mul_16s_2s_18_7_1_Mul_DSP_0_U.buff3 ;
reg [17:0] \mul_16s_2s_18_7_1_U5.top_mul_16s_2s_18_7_1_Mul_DSP_0_U.buff4 ;
reg [7:0] op_12_V_reg_1387;
reg [6:0] op_23_V_reg_1397;
reg or_ln340_reg_1320;
reg or_ln785_reg_1292;
reg or_ln786_reg_1314;
reg p_Result_11_reg_1233;
reg p_Result_12_reg_1248;
reg p_Result_14_reg_1147;
reg [4:0] p_Result_s_18_reg_1255;
reg [7:0] p_Val2_2_reg_1240;
reg [17:0] r_V_1_reg_1199;
reg [15:0] r_V_reg_1226;
reg [7:0] r_reg_1392;
reg [8:0] ret_V_16_reg_1177;
reg [5:0] ret_V_17_reg_1287;
reg [3:0] ret_V_18_reg_1304;
reg [5:0] ret_V_19_reg_1113;
reg [4:0] ret_V_20_reg_1141;
reg [10:0] ret_V_21_reg_1432;
reg [39:0] ret_V_22_reg_1479;
reg [31:0] ret_V_23_cast_reg_1484;
reg [37:0] ret_V_23_reg_1516;
reg [31:0] ret_V_24_reg_1533;
reg [31:0] ret_V_25_cast_reg_1521;
reg [31:0] ret_V_25_reg_1543;
reg [31:0] ret_V_26_reg_1553;
reg [5:0] ret_V_2_reg_1266;
reg [3:0] ret_V_3_cast_reg_1204;
reg [3:0] ret_V_4_reg_1282;
reg [4:0] ret_V_7_reg_1119;
reg [4:0] ret_V_8_reg_1136;
reg [5:0] ret_V_reg_1182;
reg [2:0] ret_reg_1126;
reg sel_tmp11_reg_1352;
reg [7:0] select_ln340_reg_1347;
reg [31:0] select_ln353_1_reg_1496;
reg [8:0] select_ln353_reg_1459;
reg [7:0] select_ln785_reg_1367;
reg [8:0] sext_ln850_reg_1447;
reg [5:0] sh_V_1_reg_1172;
reg [3:0] \shl_16s_4ns_16_7_1_U3.din1_cast_array[0] ;
reg [3:0] \shl_16s_4ns_16_7_1_U3.din1_cast_array[1] ;
reg [3:0] \shl_16s_4ns_16_7_1_U3.din1_cast_array[2] ;
reg [3:0] \shl_16s_4ns_16_7_1_U3.din1_cast_array[3] ;
reg [3:0] \shl_16s_4ns_16_7_1_U3.din1_cast_array[4] ;
reg [3:0] \shl_16s_4ns_16_7_1_U3.din1_cast_array[5] ;
reg [15:0] \shl_16s_4ns_16_7_1_U3.dout_array[0] ;
reg [15:0] \shl_16s_4ns_16_7_1_U3.dout_array[1] ;
reg [15:0] \shl_16s_4ns_16_7_1_U3.dout_array[2] ;
reg [15:0] \shl_16s_4ns_16_7_1_U3.dout_array[3] ;
reg [15:0] \shl_16s_4ns_16_7_1_U3.dout_array[4] ;
reg [15:0] \shl_16s_4ns_16_7_1_U3.dout_array[5] ;
reg [7:0] \shl_8ns_8s_8_7_1_U10.din1_cast_array[0] ;
reg [7:0] \shl_8ns_8s_8_7_1_U10.din1_cast_array[1] ;
reg [7:0] \shl_8ns_8s_8_7_1_U10.din1_cast_array[2] ;
reg [7:0] \shl_8ns_8s_8_7_1_U10.din1_cast_array[3] ;
reg [7:0] \shl_8ns_8s_8_7_1_U10.din1_cast_array[4] ;
reg [7:0] \shl_8ns_8s_8_7_1_U10.din1_cast_array[5] ;
reg [7:0] \shl_8ns_8s_8_7_1_U10.dout_array[0] ;
reg [7:0] \shl_8ns_8s_8_7_1_U10.dout_array[1] ;
reg [7:0] \shl_8ns_8s_8_7_1_U10.dout_array[2] ;
reg [7:0] \shl_8ns_8s_8_7_1_U10.dout_array[3] ;
reg [7:0] \shl_8ns_8s_8_7_1_U10.dout_array[4] ;
reg [7:0] \shl_8ns_8s_8_7_1_U10.dout_array[5] ;
reg [15:0] shl_ln1299_reg_1189;
reg [7:0] shl_ln781_reg_1372;
reg signbit_reg_1049;
reg [1:0] \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.ain_s1 ;
reg [1:0] \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.bin_s1 ;
reg \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.carry_s1 ;
reg [1:0] \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.sum_s1 ;
reg [2:0] \sub_6ns_6s_6_2_1_U8.top_sub_6ns_6s_6_2_1_Adder_4_U.ain_s1 ;
reg [2:0] \sub_6ns_6s_6_2_1_U8.top_sub_6ns_6s_6_2_1_Adder_4_U.bin_s1 ;
reg \sub_6ns_6s_6_2_1_U8.top_sub_6ns_6s_6_2_1_Adder_4_U.carry_s1 ;
reg [2:0] \sub_6ns_6s_6_2_1_U8.top_sub_6ns_6s_6_2_1_Adder_4_U.sum_s1 ;
reg [2:0] \sub_6s_6ns_6_2_1_U2.top_sub_6s_6ns_6_2_1_Adder_1_U.ain_s1 ;
reg [2:0] \sub_6s_6ns_6_2_1_U2.top_sub_6s_6ns_6_2_1_Adder_1_U.bin_s1 ;
reg \sub_6s_6ns_6_2_1_U2.top_sub_6s_6ns_6_2_1_Adder_1_U.carry_s1 ;
reg [2:0] \sub_6s_6ns_6_2_1_U2.top_sub_6s_6ns_6_2_1_Adder_1_U.sum_s1 ;
reg [3:0] sub_ln1367_reg_1044;
reg [7:0] tmp_reg_1437;
reg [5:0] trunc_ln851_1_reg_1211;
reg [2:0] trunc_ln851_3_reg_1402;
reg [3:0] ush_reg_1054;
reg xor_ln785_reg_1298;
wire [31:0] _0000_;
wire [31:0] _0001_;
wire [8:0] _0002_;
wire [2:0] _0003_;
wire [9:0] _0004_;
wire [6:0] _0005_;
wire _0006_;
wire [37:0] _0007_;
wire [15:0] _0008_;
wire [7:0] _0009_;
wire _0010_;
wire _0011_;
wire _0012_;
wire _0013_;
wire _0014_;
wire _0015_;
wire _0016_;
wire _0017_;
wire _0018_;
wire _0019_;
wire [7:0] _0020_;
wire [6:0] _0021_;
wire _0022_;
wire _0023_;
wire _0024_;
wire _0025_;
wire _0026_;
wire _0027_;
wire [4:0] _0028_;
wire [7:0] _0029_;
wire [17:0] _0030_;
wire [15:0] _0031_;
wire [7:0] _0032_;
wire [8:0] _0033_;
wire [5:0] _0034_;
wire [3:0] _0035_;
wire [5:0] _0036_;
wire [4:0] _0037_;
wire [10:0] _0038_;
wire [39:0] _0039_;
wire [31:0] _0040_;
wire [37:0] _0041_;
wire [31:0] _0042_;
wire [31:0] _0043_;
wire [31:0] _0044_;
wire [31:0] _0045_;
wire [5:0] _0046_;
wire [3:0] _0047_;
wire [3:0] _0048_;
wire [4:0] _0049_;
wire [4:0] _0050_;
wire [5:0] _0051_;
wire [2:0] _0052_;
wire _0053_;
wire [7:0] _0054_;
wire [31:0] _0055_;
wire [8:0] _0056_;
wire [7:0] _0057_;
wire [8:0] _0058_;
wire [5:0] _0059_;
wire [15:0] _0060_;
wire [7:0] _0061_;
wire _0062_;
wire [3:0] _0063_;
wire [7:0] _0064_;
wire [5:0] _0065_;
wire [2:0] _0066_;
wire [3:0] _0067_;
wire _0068_;
wire [1:0] _0069_;
wire _0070_;
wire _0071_;
wire _0072_;
wire _0073_;
wire _0074_;
wire _0075_;
wire _0076_;
wire _0077_;
wire _0078_;
wire _0079_;
wire _0080_;
wire _0081_;
wire _0082_;
wire _0083_;
wire _0084_;
wire _0085_;
wire _0086_;
wire _0087_;
wire _0088_;
wire [4:0] _0089_;
wire [4:0] _0090_;
wire _0091_;
wire [4:0] _0092_;
wire [5:0] _0093_;
wire [5:0] _0094_;
wire [5:0] _0095_;
wire [5:0] _0096_;
wire _0097_;
wire [4:0] _0098_;
wire [5:0] _0099_;
wire [6:0] _0100_;
wire [15:0] _0101_;
wire [15:0] _0102_;
wire _0103_;
wire [15:0] _0104_;
wire [16:0] _0105_;
wire [16:0] _0106_;
wire [15:0] _0107_;
wire [15:0] _0108_;
wire _0109_;
wire [15:0] _0110_;
wire [16:0] _0111_;
wire [16:0] _0112_;
wire [15:0] _0113_;
wire [15:0] _0114_;
wire _0115_;
wire [15:0] _0116_;
wire [16:0] _0117_;
wire [16:0] _0118_;
wire [15:0] _0119_;
wire [15:0] _0120_;
wire _0121_;
wire [15:0] _0122_;
wire [16:0] _0123_;
wire [16:0] _0124_;
wire [15:0] _0125_;
wire [15:0] _0126_;
wire _0127_;
wire [15:0] _0128_;
wire [16:0] _0129_;
wire [16:0] _0130_;
wire [18:0] _0131_;
wire [18:0] _0132_;
wire _0133_;
wire [18:0] _0134_;
wire [19:0] _0135_;
wire [19:0] _0136_;
wire [1:0] _0137_;
wire [1:0] _0138_;
wire _0139_;
wire _0140_;
wire [1:0] _0141_;
wire [2:0] _0142_;
wire [1:0] _0143_;
wire [1:0] _0144_;
wire _0145_;
wire _0146_;
wire [1:0] _0147_;
wire [2:0] _0148_;
wire [19:0] _0149_;
wire [19:0] _0150_;
wire _0151_;
wire [19:0] _0152_;
wire [20:0] _0153_;
wire [20:0] _0154_;
wire [1:0] _0155_;
wire [1:0] _0156_;
wire _0157_;
wire [1:0] _0158_;
wire [2:0] _0159_;
wire [2:0] _0160_;
wire [2:0] _0161_;
wire [2:0] _0162_;
wire _0163_;
wire [1:0] _0164_;
wire [2:0] _0165_;
wire [3:0] _0166_;
wire [2:0] _0167_;
wire [2:0] _0168_;
wire _0169_;
wire [2:0] _0170_;
wire [3:0] _0171_;
wire [3:0] _0172_;
wire [3:0] _0173_;
wire [3:0] _0174_;
wire _0175_;
wire [2:0] _0176_;
wire [3:0] _0177_;
wire [4:0] _0178_;
wire [3:0] _0179_;
wire [3:0] _0180_;
wire _0181_;
wire [2:0] _0182_;
wire [3:0] _0183_;
wire [4:0] _0184_;
wire [4:0] _0185_;
wire [4:0] _0186_;
wire _0187_;
wire [3:0] _0188_;
wire [4:0] _0189_;
wire [5:0] _0190_;
wire [4:0] _0191_;
wire [4:0] _0192_;
wire _0193_;
wire [3:0] _0194_;
wire [4:0] _0195_;
wire [5:0] _0196_;
wire [3:0] _0197_;
wire [3:0] _0198_;
wire [3:0] _0199_;
wire [3:0] _0200_;
wire [3:0] _0201_;
wire [3:0] _0202_;
wire [15:0] _0203_;
wire [15:0] _0204_;
wire [15:0] _0205_;
wire [15:0] _0206_;
wire [15:0] _0207_;
wire [15:0] _0208_;
wire [3:0] _0209_;
wire [15:0] _0210_;
wire [3:0] _0211_;
wire [15:0] _0212_;
wire [3:0] _0213_;
wire [15:0] _0214_;
wire [3:0] _0215_;
wire [15:0] _0216_;
wire [3:0] _0217_;
wire [15:0] _0218_;
wire [3:0] _0219_;
wire [15:0] _0220_;
wire [15:0] _0221_;
wire [15:0] _0222_;
wire [15:0] _0223_;
wire [7:0] _0224_;
wire [7:0] _0225_;
wire [7:0] _0226_;
wire [7:0] _0227_;
wire [7:0] _0228_;
wire [7:0] _0229_;
wire [7:0] _0230_;
wire [7:0] _0231_;
wire [7:0] _0232_;
wire [7:0] _0233_;
wire [7:0] _0234_;
wire [7:0] _0235_;
wire [7:0] _0236_;
wire [7:0] _0237_;
wire [7:0] _0238_;
wire [7:0] _0239_;
wire [7:0] _0240_;
wire [7:0] _0241_;
wire [7:0] _0242_;
wire [7:0] _0243_;
wire [7:0] _0244_;
wire [7:0] _0245_;
wire [7:0] _0246_;
wire [7:0] _0247_;
wire [7:0] _0248_;
wire [7:0] _0249_;
wire [7:0] _0250_;
wire [15:0] _0251_;
wire [1:0] _0252_;
wire [17:0] _0253_;
wire [17:0] _0254_;
wire [17:0] _0255_;
wire [17:0] _0256_;
wire [17:0] _0257_;
wire [3:0] _0258_;
wire [3:0] _0259_;
wire [3:0] _0260_;
wire [3:0] _0261_;
wire [3:0] _0262_;
wire [3:0] _0263_;
wire [15:0] _0264_;
wire [15:0] _0265_;
wire [15:0] _0266_;
wire [15:0] _0267_;
wire [15:0] _0268_;
wire [15:0] _0269_;
wire [3:0] _0270_;
wire [15:0] _0271_;
wire [3:0] _0272_;
wire [15:0] _0273_;
wire [3:0] _0274_;
wire [15:0] _0275_;
wire [3:0] _0276_;
wire [15:0] _0277_;
wire [3:0] _0278_;
wire [15:0] _0279_;
wire [3:0] _0280_;
wire [15:0] _0281_;
wire [15:0] _0282_;
wire [15:0] _0283_;
wire [15:0] _0284_;
wire [7:0] _0285_;
wire [7:0] _0286_;
wire [7:0] _0287_;
wire [7:0] _0288_;
wire [7:0] _0289_;
wire [7:0] _0290_;
wire [7:0] _0291_;
wire [7:0] _0292_;
wire [7:0] _0293_;
wire [7:0] _0294_;
wire [7:0] _0295_;
wire [7:0] _0296_;
wire [7:0] _0297_;
wire [7:0] _0298_;
wire [7:0] _0299_;
wire [7:0] _0300_;
wire [7:0] _0301_;
wire [7:0] _0302_;
wire [7:0] _0303_;
wire [7:0] _0304_;
wire [7:0] _0305_;
wire [7:0] _0306_;
wire [7:0] _0307_;
wire [7:0] _0308_;
wire [7:0] _0309_;
wire [7:0] _0310_;
wire [7:0] _0311_;
wire [1:0] _0312_;
wire [1:0] _0313_;
wire _0314_;
wire [1:0] _0315_;
wire [2:0] _0316_;
wire [2:0] _0317_;
wire [2:0] _0318_;
wire [2:0] _0319_;
wire _0320_;
wire [2:0] _0321_;
wire [3:0] _0322_;
wire [3:0] _0323_;
wire [2:0] _0324_;
wire [2:0] _0325_;
wire _0326_;
wire [2:0] _0327_;
wire [3:0] _0328_;
wire [3:0] _0329_;
wire _0330_;
wire _0331_;
wire _0332_;
wire _0333_;
wire _0334_;
wire _0335_;
wire _0336_;
wire _0337_;
wire _0338_;
wire _0339_;
wire _0340_;
wire _0341_;
wire _0342_;
wire _0343_;
wire _0344_;
wire _0345_;
wire _0346_;
wire _0347_;
wire _0348_;
wire _0349_;
wire _0350_;
wire _0351_;
wire _0352_;
wire _0353_;
wire _0354_;
wire _0355_;
wire _0356_;
wire _0357_;
wire _0358_;
wire _0359_;
wire _0360_;
wire _0361_;
wire _0362_;
wire _0363_;
wire _0364_;
wire _0365_;
wire _0366_;
wire _0367_;
wire _0368_;
wire _0369_;
wire _0370_;
wire _0371_;
wire _0372_;
wire _0373_;
wire _0374_;
wire _0375_;
wire \add_10ns_10s_10_2_1_U18.ce ;
wire \add_10ns_10s_10_2_1_U18.clk ;
wire [9:0] \add_10ns_10s_10_2_1_U18.din0 ;
wire [9:0] \add_10ns_10s_10_2_1_U18.din1 ;
wire [9:0] \add_10ns_10s_10_2_1_U18.dout ;
wire \add_10ns_10s_10_2_1_U18.reset ;
wire [9:0] \add_10ns_10s_10_2_1_U18.top_add_10ns_10s_10_2_1_Adder_12_U.a ;
wire [9:0] \add_10ns_10s_10_2_1_U18.top_add_10ns_10s_10_2_1_Adder_12_U.ain_s0 ;
wire [9:0] \add_10ns_10s_10_2_1_U18.top_add_10ns_10s_10_2_1_Adder_12_U.b ;
wire [9:0] \add_10ns_10s_10_2_1_U18.top_add_10ns_10s_10_2_1_Adder_12_U.bin_s0 ;
wire \add_10ns_10s_10_2_1_U18.top_add_10ns_10s_10_2_1_Adder_12_U.ce ;
wire \add_10ns_10s_10_2_1_U18.top_add_10ns_10s_10_2_1_Adder_12_U.clk ;
wire \add_10ns_10s_10_2_1_U18.top_add_10ns_10s_10_2_1_Adder_12_U.facout_s1 ;
wire \add_10ns_10s_10_2_1_U18.top_add_10ns_10s_10_2_1_Adder_12_U.facout_s2 ;
wire [4:0] \add_10ns_10s_10_2_1_U18.top_add_10ns_10s_10_2_1_Adder_12_U.fas_s1 ;
wire [4:0] \add_10ns_10s_10_2_1_U18.top_add_10ns_10s_10_2_1_Adder_12_U.fas_s2 ;
wire \add_10ns_10s_10_2_1_U18.top_add_10ns_10s_10_2_1_Adder_12_U.reset ;
wire [9:0] \add_10ns_10s_10_2_1_U18.top_add_10ns_10s_10_2_1_Adder_12_U.s ;
wire [4:0] \add_10ns_10s_10_2_1_U18.top_add_10ns_10s_10_2_1_Adder_12_U.u1.a ;
wire [4:0] \add_10ns_10s_10_2_1_U18.top_add_10ns_10s_10_2_1_Adder_12_U.u1.b ;
wire \add_10ns_10s_10_2_1_U18.top_add_10ns_10s_10_2_1_Adder_12_U.u1.cin ;
wire \add_10ns_10s_10_2_1_U18.top_add_10ns_10s_10_2_1_Adder_12_U.u1.cout ;
wire [4:0] \add_10ns_10s_10_2_1_U18.top_add_10ns_10s_10_2_1_Adder_12_U.u1.s ;
wire [4:0] \add_10ns_10s_10_2_1_U18.top_add_10ns_10s_10_2_1_Adder_12_U.u2.a ;
wire [4:0] \add_10ns_10s_10_2_1_U18.top_add_10ns_10s_10_2_1_Adder_12_U.u2.b ;
wire \add_10ns_10s_10_2_1_U18.top_add_10ns_10s_10_2_1_Adder_12_U.u2.cin ;
wire \add_10ns_10s_10_2_1_U18.top_add_10ns_10s_10_2_1_Adder_12_U.u2.cout ;
wire [4:0] \add_10ns_10s_10_2_1_U18.top_add_10ns_10s_10_2_1_Adder_12_U.u2.s ;
wire \add_11s_11s_11_2_1_U17.ce ;
wire \add_11s_11s_11_2_1_U17.clk ;
wire [10:0] \add_11s_11s_11_2_1_U17.din0 ;
wire [10:0] \add_11s_11s_11_2_1_U17.din1 ;
wire [10:0] \add_11s_11s_11_2_1_U17.dout ;
wire \add_11s_11s_11_2_1_U17.reset ;
wire [10:0] \add_11s_11s_11_2_1_U17.top_add_11s_11s_11_2_1_Adder_11_U.a ;
wire [10:0] \add_11s_11s_11_2_1_U17.top_add_11s_11s_11_2_1_Adder_11_U.ain_s0 ;
wire [10:0] \add_11s_11s_11_2_1_U17.top_add_11s_11s_11_2_1_Adder_11_U.b ;
wire [10:0] \add_11s_11s_11_2_1_U17.top_add_11s_11s_11_2_1_Adder_11_U.bin_s0 ;
wire \add_11s_11s_11_2_1_U17.top_add_11s_11s_11_2_1_Adder_11_U.ce ;
wire \add_11s_11s_11_2_1_U17.top_add_11s_11s_11_2_1_Adder_11_U.clk ;
wire \add_11s_11s_11_2_1_U17.top_add_11s_11s_11_2_1_Adder_11_U.facout_s1 ;
wire \add_11s_11s_11_2_1_U17.top_add_11s_11s_11_2_1_Adder_11_U.facout_s2 ;
wire [4:0] \add_11s_11s_11_2_1_U17.top_add_11s_11s_11_2_1_Adder_11_U.fas_s1 ;
wire [5:0] \add_11s_11s_11_2_1_U17.top_add_11s_11s_11_2_1_Adder_11_U.fas_s2 ;
wire \add_11s_11s_11_2_1_U17.top_add_11s_11s_11_2_1_Adder_11_U.reset ;
wire [10:0] \add_11s_11s_11_2_1_U17.top_add_11s_11s_11_2_1_Adder_11_U.s ;
wire [4:0] \add_11s_11s_11_2_1_U17.top_add_11s_11s_11_2_1_Adder_11_U.u1.a ;
wire [4:0] \add_11s_11s_11_2_1_U17.top_add_11s_11s_11_2_1_Adder_11_U.u1.b ;
wire \add_11s_11s_11_2_1_U17.top_add_11s_11s_11_2_1_Adder_11_U.u1.cin ;
wire \add_11s_11s_11_2_1_U17.top_add_11s_11s_11_2_1_Adder_11_U.u1.cout ;
wire [4:0] \add_11s_11s_11_2_1_U17.top_add_11s_11s_11_2_1_Adder_11_U.u1.s ;
wire [5:0] \add_11s_11s_11_2_1_U17.top_add_11s_11s_11_2_1_Adder_11_U.u2.a ;
wire [5:0] \add_11s_11s_11_2_1_U17.top_add_11s_11s_11_2_1_Adder_11_U.u2.b ;
wire \add_11s_11s_11_2_1_U17.top_add_11s_11s_11_2_1_Adder_11_U.u2.cin ;
wire \add_11s_11s_11_2_1_U17.top_add_11s_11s_11_2_1_Adder_11_U.u2.cout ;
wire [5:0] \add_11s_11s_11_2_1_U17.top_add_11s_11s_11_2_1_Adder_11_U.u2.s ;
wire \add_32ns_32ns_32_2_1_U21.ce ;
wire \add_32ns_32ns_32_2_1_U21.clk ;
wire [31:0] \add_32ns_32ns_32_2_1_U21.din0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U21.din1 ;
wire [31:0] \add_32ns_32ns_32_2_1_U21.dout ;
wire \add_32ns_32ns_32_2_1_U21.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.a ;
wire [31:0] \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.ain_s0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.b ;
wire [31:0] \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.bin_s0 ;
wire \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.ce ;
wire \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.clk ;
wire \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.facout_s1 ;
wire \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.facout_s2 ;
wire [15:0] \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.fas_s1 ;
wire [15:0] \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.fas_s2 ;
wire \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.b ;
wire \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.cin ;
wire \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.b ;
wire \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.cin ;
wire \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.s ;
wire \add_32ns_32ns_32_2_1_U23.ce ;
wire \add_32ns_32ns_32_2_1_U23.clk ;
wire [31:0] \add_32ns_32ns_32_2_1_U23.din0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U23.din1 ;
wire [31:0] \add_32ns_32ns_32_2_1_U23.dout ;
wire \add_32ns_32ns_32_2_1_U23.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.a ;
wire [31:0] \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.ain_s0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.b ;
wire [31:0] \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.bin_s0 ;
wire \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.ce ;
wire \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.clk ;
wire \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.facout_s1 ;
wire \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.facout_s2 ;
wire [15:0] \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.fas_s1 ;
wire [15:0] \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.fas_s2 ;
wire \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.b ;
wire \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.cin ;
wire \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.b ;
wire \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.cin ;
wire \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.s ;
wire \add_32ns_32s_32_2_1_U24.ce ;
wire \add_32ns_32s_32_2_1_U24.clk ;
wire [31:0] \add_32ns_32s_32_2_1_U24.din0 ;
wire [31:0] \add_32ns_32s_32_2_1_U24.din1 ;
wire [31:0] \add_32ns_32s_32_2_1_U24.dout ;
wire \add_32ns_32s_32_2_1_U24.reset ;
wire [31:0] \add_32ns_32s_32_2_1_U24.top_add_32ns_32s_32_2_1_Adder_17_U.a ;
wire [31:0] \add_32ns_32s_32_2_1_U24.top_add_32ns_32s_32_2_1_Adder_17_U.ain_s0 ;
wire [31:0] \add_32ns_32s_32_2_1_U24.top_add_32ns_32s_32_2_1_Adder_17_U.b ;
wire [31:0] \add_32ns_32s_32_2_1_U24.top_add_32ns_32s_32_2_1_Adder_17_U.bin_s0 ;
wire \add_32ns_32s_32_2_1_U24.top_add_32ns_32s_32_2_1_Adder_17_U.ce ;
wire \add_32ns_32s_32_2_1_U24.top_add_32ns_32s_32_2_1_Adder_17_U.clk ;
wire \add_32ns_32s_32_2_1_U24.top_add_32ns_32s_32_2_1_Adder_17_U.facout_s1 ;
wire \add_32ns_32s_32_2_1_U24.top_add_32ns_32s_32_2_1_Adder_17_U.facout_s2 ;
wire [15:0] \add_32ns_32s_32_2_1_U24.top_add_32ns_32s_32_2_1_Adder_17_U.fas_s1 ;
wire [15:0] \add_32ns_32s_32_2_1_U24.top_add_32ns_32s_32_2_1_Adder_17_U.fas_s2 ;
wire \add_32ns_32s_32_2_1_U24.top_add_32ns_32s_32_2_1_Adder_17_U.reset ;
wire [31:0] \add_32ns_32s_32_2_1_U24.top_add_32ns_32s_32_2_1_Adder_17_U.s ;
wire [15:0] \add_32ns_32s_32_2_1_U24.top_add_32ns_32s_32_2_1_Adder_17_U.u1.a ;
wire [15:0] \add_32ns_32s_32_2_1_U24.top_add_32ns_32s_32_2_1_Adder_17_U.u1.b ;
wire \add_32ns_32s_32_2_1_U24.top_add_32ns_32s_32_2_1_Adder_17_U.u1.cin ;
wire \add_32ns_32s_32_2_1_U24.top_add_32ns_32s_32_2_1_Adder_17_U.u1.cout ;
wire [15:0] \add_32ns_32s_32_2_1_U24.top_add_32ns_32s_32_2_1_Adder_17_U.u1.s ;
wire [15:0] \add_32ns_32s_32_2_1_U24.top_add_32ns_32s_32_2_1_Adder_17_U.u2.a ;
wire [15:0] \add_32ns_32s_32_2_1_U24.top_add_32ns_32s_32_2_1_Adder_17_U.u2.b ;
wire \add_32ns_32s_32_2_1_U24.top_add_32ns_32s_32_2_1_Adder_17_U.u2.cin ;
wire \add_32ns_32s_32_2_1_U24.top_add_32ns_32s_32_2_1_Adder_17_U.u2.cout ;
wire [15:0] \add_32ns_32s_32_2_1_U24.top_add_32ns_32s_32_2_1_Adder_17_U.u2.s ;
wire \add_32ns_32s_32_2_1_U25.ce ;
wire \add_32ns_32s_32_2_1_U25.clk ;
wire [31:0] \add_32ns_32s_32_2_1_U25.din0 ;
wire [31:0] \add_32ns_32s_32_2_1_U25.din1 ;
wire [31:0] \add_32ns_32s_32_2_1_U25.dout ;
wire \add_32ns_32s_32_2_1_U25.reset ;
wire [31:0] \add_32ns_32s_32_2_1_U25.top_add_32ns_32s_32_2_1_Adder_17_U.a ;
wire [31:0] \add_32ns_32s_32_2_1_U25.top_add_32ns_32s_32_2_1_Adder_17_U.ain_s0 ;
wire [31:0] \add_32ns_32s_32_2_1_U25.top_add_32ns_32s_32_2_1_Adder_17_U.b ;
wire [31:0] \add_32ns_32s_32_2_1_U25.top_add_32ns_32s_32_2_1_Adder_17_U.bin_s0 ;
wire \add_32ns_32s_32_2_1_U25.top_add_32ns_32s_32_2_1_Adder_17_U.ce ;
wire \add_32ns_32s_32_2_1_U25.top_add_32ns_32s_32_2_1_Adder_17_U.clk ;
wire \add_32ns_32s_32_2_1_U25.top_add_32ns_32s_32_2_1_Adder_17_U.facout_s1 ;
wire \add_32ns_32s_32_2_1_U25.top_add_32ns_32s_32_2_1_Adder_17_U.facout_s2 ;
wire [15:0] \add_32ns_32s_32_2_1_U25.top_add_32ns_32s_32_2_1_Adder_17_U.fas_s1 ;
wire [15:0] \add_32ns_32s_32_2_1_U25.top_add_32ns_32s_32_2_1_Adder_17_U.fas_s2 ;
wire \add_32ns_32s_32_2_1_U25.top_add_32ns_32s_32_2_1_Adder_17_U.reset ;
wire [31:0] \add_32ns_32s_32_2_1_U25.top_add_32ns_32s_32_2_1_Adder_17_U.s ;
wire [15:0] \add_32ns_32s_32_2_1_U25.top_add_32ns_32s_32_2_1_Adder_17_U.u1.a ;
wire [15:0] \add_32ns_32s_32_2_1_U25.top_add_32ns_32s_32_2_1_Adder_17_U.u1.b ;
wire \add_32ns_32s_32_2_1_U25.top_add_32ns_32s_32_2_1_Adder_17_U.u1.cin ;
wire \add_32ns_32s_32_2_1_U25.top_add_32ns_32s_32_2_1_Adder_17_U.u1.cout ;
wire [15:0] \add_32ns_32s_32_2_1_U25.top_add_32ns_32s_32_2_1_Adder_17_U.u1.s ;
wire [15:0] \add_32ns_32s_32_2_1_U25.top_add_32ns_32s_32_2_1_Adder_17_U.u2.a ;
wire [15:0] \add_32ns_32s_32_2_1_U25.top_add_32ns_32s_32_2_1_Adder_17_U.u2.b ;
wire \add_32ns_32s_32_2_1_U25.top_add_32ns_32s_32_2_1_Adder_17_U.u2.cin ;
wire \add_32ns_32s_32_2_1_U25.top_add_32ns_32s_32_2_1_Adder_17_U.u2.cout ;
wire [15:0] \add_32ns_32s_32_2_1_U25.top_add_32ns_32s_32_2_1_Adder_17_U.u2.s ;
wire \add_32s_32ns_32_2_1_U26.ce ;
wire \add_32s_32ns_32_2_1_U26.clk ;
wire [31:0] \add_32s_32ns_32_2_1_U26.din0 ;
wire [31:0] \add_32s_32ns_32_2_1_U26.din1 ;
wire [31:0] \add_32s_32ns_32_2_1_U26.dout ;
wire \add_32s_32ns_32_2_1_U26.reset ;
wire [31:0] \add_32s_32ns_32_2_1_U26.top_add_32s_32ns_32_2_1_Adder_18_U.a ;
wire [31:0] \add_32s_32ns_32_2_1_U26.top_add_32s_32ns_32_2_1_Adder_18_U.ain_s0 ;
wire [31:0] \add_32s_32ns_32_2_1_U26.top_add_32s_32ns_32_2_1_Adder_18_U.b ;
wire [31:0] \add_32s_32ns_32_2_1_U26.top_add_32s_32ns_32_2_1_Adder_18_U.bin_s0 ;
wire \add_32s_32ns_32_2_1_U26.top_add_32s_32ns_32_2_1_Adder_18_U.ce ;
wire \add_32s_32ns_32_2_1_U26.top_add_32s_32ns_32_2_1_Adder_18_U.clk ;
wire \add_32s_32ns_32_2_1_U26.top_add_32s_32ns_32_2_1_Adder_18_U.facout_s1 ;
wire \add_32s_32ns_32_2_1_U26.top_add_32s_32ns_32_2_1_Adder_18_U.facout_s2 ;
wire [15:0] \add_32s_32ns_32_2_1_U26.top_add_32s_32ns_32_2_1_Adder_18_U.fas_s1 ;
wire [15:0] \add_32s_32ns_32_2_1_U26.top_add_32s_32ns_32_2_1_Adder_18_U.fas_s2 ;
wire \add_32s_32ns_32_2_1_U26.top_add_32s_32ns_32_2_1_Adder_18_U.reset ;
wire [31:0] \add_32s_32ns_32_2_1_U26.top_add_32s_32ns_32_2_1_Adder_18_U.s ;
wire [15:0] \add_32s_32ns_32_2_1_U26.top_add_32s_32ns_32_2_1_Adder_18_U.u1.a ;
wire [15:0] \add_32s_32ns_32_2_1_U26.top_add_32s_32ns_32_2_1_Adder_18_U.u1.b ;
wire \add_32s_32ns_32_2_1_U26.top_add_32s_32ns_32_2_1_Adder_18_U.u1.cin ;
wire \add_32s_32ns_32_2_1_U26.top_add_32s_32ns_32_2_1_Adder_18_U.u1.cout ;
wire [15:0] \add_32s_32ns_32_2_1_U26.top_add_32s_32ns_32_2_1_Adder_18_U.u1.s ;
wire [15:0] \add_32s_32ns_32_2_1_U26.top_add_32s_32ns_32_2_1_Adder_18_U.u2.a ;
wire [15:0] \add_32s_32ns_32_2_1_U26.top_add_32s_32ns_32_2_1_Adder_18_U.u2.b ;
wire \add_32s_32ns_32_2_1_U26.top_add_32s_32ns_32_2_1_Adder_18_U.u2.cin ;
wire \add_32s_32ns_32_2_1_U26.top_add_32s_32ns_32_2_1_Adder_18_U.u2.cout ;
wire [15:0] \add_32s_32ns_32_2_1_U26.top_add_32s_32ns_32_2_1_Adder_18_U.u2.s ;
wire \add_38s_38s_38_2_1_U22.ce ;
wire \add_38s_38s_38_2_1_U22.clk ;
wire [37:0] \add_38s_38s_38_2_1_U22.din0 ;
wire [37:0] \add_38s_38s_38_2_1_U22.din1 ;
wire [37:0] \add_38s_38s_38_2_1_U22.dout ;
wire \add_38s_38s_38_2_1_U22.reset ;
wire [37:0] \add_38s_38s_38_2_1_U22.top_add_38s_38s_38_2_1_Adder_16_U.a ;
wire [37:0] \add_38s_38s_38_2_1_U22.top_add_38s_38s_38_2_1_Adder_16_U.ain_s0 ;
wire [37:0] \add_38s_38s_38_2_1_U22.top_add_38s_38s_38_2_1_Adder_16_U.b ;
wire [37:0] \add_38s_38s_38_2_1_U22.top_add_38s_38s_38_2_1_Adder_16_U.bin_s0 ;
wire \add_38s_38s_38_2_1_U22.top_add_38s_38s_38_2_1_Adder_16_U.ce ;
wire \add_38s_38s_38_2_1_U22.top_add_38s_38s_38_2_1_Adder_16_U.clk ;
wire \add_38s_38s_38_2_1_U22.top_add_38s_38s_38_2_1_Adder_16_U.facout_s1 ;
wire \add_38s_38s_38_2_1_U22.top_add_38s_38s_38_2_1_Adder_16_U.facout_s2 ;
wire [18:0] \add_38s_38s_38_2_1_U22.top_add_38s_38s_38_2_1_Adder_16_U.fas_s1 ;
wire [18:0] \add_38s_38s_38_2_1_U22.top_add_38s_38s_38_2_1_Adder_16_U.fas_s2 ;
wire \add_38s_38s_38_2_1_U22.top_add_38s_38s_38_2_1_Adder_16_U.reset ;
wire [37:0] \add_38s_38s_38_2_1_U22.top_add_38s_38s_38_2_1_Adder_16_U.s ;
wire [18:0] \add_38s_38s_38_2_1_U22.top_add_38s_38s_38_2_1_Adder_16_U.u1.a ;
wire [18:0] \add_38s_38s_38_2_1_U22.top_add_38s_38s_38_2_1_Adder_16_U.u1.b ;
wire \add_38s_38s_38_2_1_U22.top_add_38s_38s_38_2_1_Adder_16_U.u1.cin ;
wire \add_38s_38s_38_2_1_U22.top_add_38s_38s_38_2_1_Adder_16_U.u1.cout ;
wire [18:0] \add_38s_38s_38_2_1_U22.top_add_38s_38s_38_2_1_Adder_16_U.u1.s ;
wire [18:0] \add_38s_38s_38_2_1_U22.top_add_38s_38s_38_2_1_Adder_16_U.u2.a ;
wire [18:0] \add_38s_38s_38_2_1_U22.top_add_38s_38s_38_2_1_Adder_16_U.u2.b ;
wire \add_38s_38s_38_2_1_U22.top_add_38s_38s_38_2_1_Adder_16_U.u2.cin ;
wire \add_38s_38s_38_2_1_U22.top_add_38s_38s_38_2_1_Adder_16_U.u2.cout ;
wire [18:0] \add_38s_38s_38_2_1_U22.top_add_38s_38s_38_2_1_Adder_16_U.u2.s ;
wire \add_3ns_3ns_3_2_1_U15.ce ;
wire \add_3ns_3ns_3_2_1_U15.clk ;
wire [2:0] \add_3ns_3ns_3_2_1_U15.din0 ;
wire [2:0] \add_3ns_3ns_3_2_1_U15.din1 ;
wire [2:0] \add_3ns_3ns_3_2_1_U15.dout ;
wire \add_3ns_3ns_3_2_1_U15.reset ;
wire [2:0] \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_9_U.a ;
wire [2:0] \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_9_U.ain_s0 ;
wire [2:0] \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_9_U.b ;
wire [2:0] \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_9_U.bin_s0 ;
wire \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_9_U.ce ;
wire \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_9_U.clk ;
wire \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_9_U.facout_s1 ;
wire \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_9_U.facout_s2 ;
wire \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_9_U.fas_s1 ;
wire [1:0] \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_9_U.fas_s2 ;
wire \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_9_U.reset ;
wire [2:0] \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_9_U.s ;
wire \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_9_U.u1.a ;
wire \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_9_U.u1.b ;
wire \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_9_U.u1.cin ;
wire \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_9_U.u1.cout ;
wire \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_9_U.u1.s ;
wire [1:0] \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_9_U.u2.a ;
wire [1:0] \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_9_U.u2.b ;
wire \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_9_U.u2.cin ;
wire \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_9_U.u2.cout ;
wire [1:0] \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_9_U.u2.s ;
wire \add_3s_3s_3_2_1_U6.ce ;
wire \add_3s_3s_3_2_1_U6.clk ;
wire [2:0] \add_3s_3s_3_2_1_U6.din0 ;
wire [2:0] \add_3s_3s_3_2_1_U6.din1 ;
wire [2:0] \add_3s_3s_3_2_1_U6.dout ;
wire \add_3s_3s_3_2_1_U6.reset ;
wire [2:0] \add_3s_3s_3_2_1_U6.top_add_3s_3s_3_2_1_Adder_2_U.a ;
wire [2:0] \add_3s_3s_3_2_1_U6.top_add_3s_3s_3_2_1_Adder_2_U.ain_s0 ;
wire [2:0] \add_3s_3s_3_2_1_U6.top_add_3s_3s_3_2_1_Adder_2_U.b ;
wire [2:0] \add_3s_3s_3_2_1_U6.top_add_3s_3s_3_2_1_Adder_2_U.bin_s0 ;
wire \add_3s_3s_3_2_1_U6.top_add_3s_3s_3_2_1_Adder_2_U.ce ;
wire \add_3s_3s_3_2_1_U6.top_add_3s_3s_3_2_1_Adder_2_U.clk ;
wire \add_3s_3s_3_2_1_U6.top_add_3s_3s_3_2_1_Adder_2_U.facout_s1 ;
wire \add_3s_3s_3_2_1_U6.top_add_3s_3s_3_2_1_Adder_2_U.facout_s2 ;
wire \add_3s_3s_3_2_1_U6.top_add_3s_3s_3_2_1_Adder_2_U.fas_s1 ;
wire [1:0] \add_3s_3s_3_2_1_U6.top_add_3s_3s_3_2_1_Adder_2_U.fas_s2 ;
wire \add_3s_3s_3_2_1_U6.top_add_3s_3s_3_2_1_Adder_2_U.reset ;
wire [2:0] \add_3s_3s_3_2_1_U6.top_add_3s_3s_3_2_1_Adder_2_U.s ;
wire \add_3s_3s_3_2_1_U6.top_add_3s_3s_3_2_1_Adder_2_U.u1.a ;
wire \add_3s_3s_3_2_1_U6.top_add_3s_3s_3_2_1_Adder_2_U.u1.b ;
wire \add_3s_3s_3_2_1_U6.top_add_3s_3s_3_2_1_Adder_2_U.u1.cin ;
wire \add_3s_3s_3_2_1_U6.top_add_3s_3s_3_2_1_Adder_2_U.u1.cout ;
wire \add_3s_3s_3_2_1_U6.top_add_3s_3s_3_2_1_Adder_2_U.u1.s ;
wire [1:0] \add_3s_3s_3_2_1_U6.top_add_3s_3s_3_2_1_Adder_2_U.u2.a ;
wire [1:0] \add_3s_3s_3_2_1_U6.top_add_3s_3s_3_2_1_Adder_2_U.u2.b ;
wire \add_3s_3s_3_2_1_U6.top_add_3s_3s_3_2_1_Adder_2_U.u2.cin ;
wire \add_3s_3s_3_2_1_U6.top_add_3s_3s_3_2_1_Adder_2_U.u2.cout ;
wire [1:0] \add_3s_3s_3_2_1_U6.top_add_3s_3s_3_2_1_Adder_2_U.u2.s ;
wire \add_40s_40s_40_2_1_U20.ce ;
wire \add_40s_40s_40_2_1_U20.clk ;
wire [39:0] \add_40s_40s_40_2_1_U20.din0 ;
wire [39:0] \add_40s_40s_40_2_1_U20.din1 ;
wire [39:0] \add_40s_40s_40_2_1_U20.dout ;
wire \add_40s_40s_40_2_1_U20.reset ;
wire [39:0] \add_40s_40s_40_2_1_U20.top_add_40s_40s_40_2_1_Adder_14_U.a ;
wire [39:0] \add_40s_40s_40_2_1_U20.top_add_40s_40s_40_2_1_Adder_14_U.ain_s0 ;
wire [39:0] \add_40s_40s_40_2_1_U20.top_add_40s_40s_40_2_1_Adder_14_U.b ;
wire [39:0] \add_40s_40s_40_2_1_U20.top_add_40s_40s_40_2_1_Adder_14_U.bin_s0 ;
wire \add_40s_40s_40_2_1_U20.top_add_40s_40s_40_2_1_Adder_14_U.ce ;
wire \add_40s_40s_40_2_1_U20.top_add_40s_40s_40_2_1_Adder_14_U.clk ;
wire \add_40s_40s_40_2_1_U20.top_add_40s_40s_40_2_1_Adder_14_U.facout_s1 ;
wire \add_40s_40s_40_2_1_U20.top_add_40s_40s_40_2_1_Adder_14_U.facout_s2 ;
wire [19:0] \add_40s_40s_40_2_1_U20.top_add_40s_40s_40_2_1_Adder_14_U.fas_s1 ;
wire [19:0] \add_40s_40s_40_2_1_U20.top_add_40s_40s_40_2_1_Adder_14_U.fas_s2 ;
wire \add_40s_40s_40_2_1_U20.top_add_40s_40s_40_2_1_Adder_14_U.reset ;
wire [39:0] \add_40s_40s_40_2_1_U20.top_add_40s_40s_40_2_1_Adder_14_U.s ;
wire [19:0] \add_40s_40s_40_2_1_U20.top_add_40s_40s_40_2_1_Adder_14_U.u1.a ;
wire [19:0] \add_40s_40s_40_2_1_U20.top_add_40s_40s_40_2_1_Adder_14_U.u1.b ;
wire \add_40s_40s_40_2_1_U20.top_add_40s_40s_40_2_1_Adder_14_U.u1.cin ;
wire \add_40s_40s_40_2_1_U20.top_add_40s_40s_40_2_1_Adder_14_U.u1.cout ;
wire [19:0] \add_40s_40s_40_2_1_U20.top_add_40s_40s_40_2_1_Adder_14_U.u1.s ;
wire [19:0] \add_40s_40s_40_2_1_U20.top_add_40s_40s_40_2_1_Adder_14_U.u2.a ;
wire [19:0] \add_40s_40s_40_2_1_U20.top_add_40s_40s_40_2_1_Adder_14_U.u2.b ;
wire \add_40s_40s_40_2_1_U20.top_add_40s_40s_40_2_1_Adder_14_U.u2.cin ;
wire \add_40s_40s_40_2_1_U20.top_add_40s_40s_40_2_1_Adder_14_U.u2.cout ;
wire [19:0] \add_40s_40s_40_2_1_U20.top_add_40s_40s_40_2_1_Adder_14_U.u2.s ;
wire \add_4ns_4ns_4_2_1_U13.ce ;
wire \add_4ns_4ns_4_2_1_U13.clk ;
wire [3:0] \add_4ns_4ns_4_2_1_U13.din0 ;
wire [3:0] \add_4ns_4ns_4_2_1_U13.din1 ;
wire [3:0] \add_4ns_4ns_4_2_1_U13.dout ;
wire \add_4ns_4ns_4_2_1_U13.reset ;
wire [3:0] \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_7_U.a ;
wire [3:0] \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_7_U.ain_s0 ;
wire [3:0] \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_7_U.b ;
wire [3:0] \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_7_U.bin_s0 ;
wire \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_7_U.ce ;
wire \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_7_U.clk ;
wire \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_7_U.facout_s1 ;
wire \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_7_U.facout_s2 ;
wire [1:0] \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_7_U.fas_s1 ;
wire [1:0] \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_7_U.fas_s2 ;
wire \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_7_U.reset ;
wire [3:0] \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_7_U.s ;
wire [1:0] \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_7_U.u1.a ;
wire [1:0] \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_7_U.u1.b ;
wire \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_7_U.u1.cin ;
wire \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_7_U.u1.cout ;
wire [1:0] \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_7_U.u1.s ;
wire [1:0] \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_7_U.u2.a ;
wire [1:0] \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_7_U.u2.b ;
wire \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_7_U.u2.cin ;
wire \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_7_U.u2.cout ;
wire [1:0] \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_7_U.u2.s ;
wire \add_5ns_5ns_5_2_1_U7.ce ;
wire \add_5ns_5ns_5_2_1_U7.clk ;
wire [4:0] \add_5ns_5ns_5_2_1_U7.din0 ;
wire [4:0] \add_5ns_5ns_5_2_1_U7.din1 ;
wire [4:0] \add_5ns_5ns_5_2_1_U7.dout ;
wire \add_5ns_5ns_5_2_1_U7.reset ;
wire [4:0] \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_3_U.a ;
wire [4:0] \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_3_U.ain_s0 ;
wire [4:0] \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_3_U.b ;
wire [4:0] \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_3_U.bin_s0 ;
wire \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_3_U.ce ;
wire \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_3_U.clk ;
wire \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_3_U.facout_s1 ;
wire \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_3_U.facout_s2 ;
wire [1:0] \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_3_U.fas_s1 ;
wire [2:0] \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_3_U.fas_s2 ;
wire \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_3_U.reset ;
wire [4:0] \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_3_U.s ;
wire [1:0] \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_3_U.u1.a ;
wire [1:0] \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_3_U.u1.b ;
wire \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_3_U.u1.cin ;
wire \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_3_U.u1.cout ;
wire [1:0] \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_3_U.u1.s ;
wire [2:0] \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_3_U.u2.a ;
wire [2:0] \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_3_U.u2.b ;
wire \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_3_U.u2.cin ;
wire \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_3_U.u2.cout ;
wire [2:0] \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_3_U.u2.s ;
wire \add_6ns_6ns_6_2_1_U12.ce ;
wire \add_6ns_6ns_6_2_1_U12.clk ;
wire [5:0] \add_6ns_6ns_6_2_1_U12.din0 ;
wire [5:0] \add_6ns_6ns_6_2_1_U12.din1 ;
wire [5:0] \add_6ns_6ns_6_2_1_U12.dout ;
wire \add_6ns_6ns_6_2_1_U12.reset ;
wire [5:0] \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_6_U.a ;
wire [5:0] \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_6_U.ain_s0 ;
wire [5:0] \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_6_U.b ;
wire [5:0] \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_6_U.bin_s0 ;
wire \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_6_U.ce ;
wire \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_6_U.clk ;
wire \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_6_U.facout_s1 ;
wire \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_6_U.facout_s2 ;
wire [2:0] \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_6_U.fas_s1 ;
wire [2:0] \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_6_U.fas_s2 ;
wire \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_6_U.reset ;
wire [5:0] \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_6_U.s ;
wire [2:0] \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_6_U.u1.a ;
wire [2:0] \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_6_U.u1.b ;
wire \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_6_U.u1.cin ;
wire \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_6_U.u1.cout ;
wire [2:0] \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_6_U.u1.s ;
wire [2:0] \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_6_U.u2.a ;
wire [2:0] \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_6_U.u2.b ;
wire \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_6_U.u2.cin ;
wire \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_6_U.u2.cout ;
wire [2:0] \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_6_U.u2.s ;
wire \add_7ns_7ns_7_2_1_U16.ce ;
wire \add_7ns_7ns_7_2_1_U16.clk ;
wire [6:0] \add_7ns_7ns_7_2_1_U16.din0 ;
wire [6:0] \add_7ns_7ns_7_2_1_U16.din1 ;
wire [6:0] \add_7ns_7ns_7_2_1_U16.dout ;
wire \add_7ns_7ns_7_2_1_U16.reset ;
wire [6:0] \add_7ns_7ns_7_2_1_U16.top_add_7ns_7ns_7_2_1_Adder_10_U.a ;
wire [6:0] \add_7ns_7ns_7_2_1_U16.top_add_7ns_7ns_7_2_1_Adder_10_U.ain_s0 ;
wire [6:0] \add_7ns_7ns_7_2_1_U16.top_add_7ns_7ns_7_2_1_Adder_10_U.b ;
wire [6:0] \add_7ns_7ns_7_2_1_U16.top_add_7ns_7ns_7_2_1_Adder_10_U.bin_s0 ;
wire \add_7ns_7ns_7_2_1_U16.top_add_7ns_7ns_7_2_1_Adder_10_U.ce ;
wire \add_7ns_7ns_7_2_1_U16.top_add_7ns_7ns_7_2_1_Adder_10_U.clk ;
wire \add_7ns_7ns_7_2_1_U16.top_add_7ns_7ns_7_2_1_Adder_10_U.facout_s1 ;
wire \add_7ns_7ns_7_2_1_U16.top_add_7ns_7ns_7_2_1_Adder_10_U.facout_s2 ;
wire [2:0] \add_7ns_7ns_7_2_1_U16.top_add_7ns_7ns_7_2_1_Adder_10_U.fas_s1 ;
wire [3:0] \add_7ns_7ns_7_2_1_U16.top_add_7ns_7ns_7_2_1_Adder_10_U.fas_s2 ;
wire \add_7ns_7ns_7_2_1_U16.top_add_7ns_7ns_7_2_1_Adder_10_U.reset ;
wire [6:0] \add_7ns_7ns_7_2_1_U16.top_add_7ns_7ns_7_2_1_Adder_10_U.s ;
wire [2:0] \add_7ns_7ns_7_2_1_U16.top_add_7ns_7ns_7_2_1_Adder_10_U.u1.a ;
wire [2:0] \add_7ns_7ns_7_2_1_U16.top_add_7ns_7ns_7_2_1_Adder_10_U.u1.b ;
wire \add_7ns_7ns_7_2_1_U16.top_add_7ns_7ns_7_2_1_Adder_10_U.u1.cin ;
wire \add_7ns_7ns_7_2_1_U16.top_add_7ns_7ns_7_2_1_Adder_10_U.u1.cout ;
wire [2:0] \add_7ns_7ns_7_2_1_U16.top_add_7ns_7ns_7_2_1_Adder_10_U.u1.s ;
wire [3:0] \add_7ns_7ns_7_2_1_U16.top_add_7ns_7ns_7_2_1_Adder_10_U.u2.a ;
wire [3:0] \add_7ns_7ns_7_2_1_U16.top_add_7ns_7ns_7_2_1_Adder_10_U.u2.b ;
wire \add_7ns_7ns_7_2_1_U16.top_add_7ns_7ns_7_2_1_Adder_10_U.u2.cin ;
wire \add_7ns_7ns_7_2_1_U16.top_add_7ns_7ns_7_2_1_Adder_10_U.u2.cout ;
wire [3:0] \add_7ns_7ns_7_2_1_U16.top_add_7ns_7ns_7_2_1_Adder_10_U.u2.s ;
wire \add_7s_7ns_7_2_1_U14.ce ;
wire \add_7s_7ns_7_2_1_U14.clk ;
wire [6:0] \add_7s_7ns_7_2_1_U14.din0 ;
wire [6:0] \add_7s_7ns_7_2_1_U14.din1 ;
wire [6:0] \add_7s_7ns_7_2_1_U14.dout ;
wire \add_7s_7ns_7_2_1_U14.reset ;
wire [6:0] \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_8_U.a ;
wire [6:0] \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_8_U.ain_s0 ;
wire [6:0] \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_8_U.b ;
wire [6:0] \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_8_U.bin_s0 ;
wire \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_8_U.ce ;
wire \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_8_U.clk ;
wire \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_8_U.facout_s1 ;
wire \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_8_U.facout_s2 ;
wire [2:0] \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_8_U.fas_s1 ;
wire [3:0] \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_8_U.fas_s2 ;
wire \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_8_U.reset ;
wire [6:0] \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_8_U.s ;
wire [2:0] \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_8_U.u1.a ;
wire [2:0] \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_8_U.u1.b ;
wire \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_8_U.u1.cin ;
wire \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_8_U.u1.cout ;
wire [2:0] \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_8_U.u1.s ;
wire [3:0] \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_8_U.u2.a ;
wire [3:0] \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_8_U.u2.b ;
wire \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_8_U.u2.cin ;
wire \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_8_U.u2.cout ;
wire [3:0] \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_8_U.u2.s ;
wire \add_9ns_9s_9_2_1_U9.ce ;
wire \add_9ns_9s_9_2_1_U9.clk ;
wire [8:0] \add_9ns_9s_9_2_1_U9.din0 ;
wire [8:0] \add_9ns_9s_9_2_1_U9.din1 ;
wire [8:0] \add_9ns_9s_9_2_1_U9.dout ;
wire \add_9ns_9s_9_2_1_U9.reset ;
wire [8:0] \add_9ns_9s_9_2_1_U9.top_add_9ns_9s_9_2_1_Adder_5_U.a ;
wire [8:0] \add_9ns_9s_9_2_1_U9.top_add_9ns_9s_9_2_1_Adder_5_U.ain_s0 ;
wire [8:0] \add_9ns_9s_9_2_1_U9.top_add_9ns_9s_9_2_1_Adder_5_U.b ;
wire [8:0] \add_9ns_9s_9_2_1_U9.top_add_9ns_9s_9_2_1_Adder_5_U.bin_s0 ;
wire \add_9ns_9s_9_2_1_U9.top_add_9ns_9s_9_2_1_Adder_5_U.ce ;
wire \add_9ns_9s_9_2_1_U9.top_add_9ns_9s_9_2_1_Adder_5_U.clk ;
wire \add_9ns_9s_9_2_1_U9.top_add_9ns_9s_9_2_1_Adder_5_U.facout_s1 ;
wire \add_9ns_9s_9_2_1_U9.top_add_9ns_9s_9_2_1_Adder_5_U.facout_s2 ;
wire [3:0] \add_9ns_9s_9_2_1_U9.top_add_9ns_9s_9_2_1_Adder_5_U.fas_s1 ;
wire [4:0] \add_9ns_9s_9_2_1_U9.top_add_9ns_9s_9_2_1_Adder_5_U.fas_s2 ;
wire \add_9ns_9s_9_2_1_U9.top_add_9ns_9s_9_2_1_Adder_5_U.reset ;
wire [8:0] \add_9ns_9s_9_2_1_U9.top_add_9ns_9s_9_2_1_Adder_5_U.s ;
wire [3:0] \add_9ns_9s_9_2_1_U9.top_add_9ns_9s_9_2_1_Adder_5_U.u1.a ;
wire [3:0] \add_9ns_9s_9_2_1_U9.top_add_9ns_9s_9_2_1_Adder_5_U.u1.b ;
wire \add_9ns_9s_9_2_1_U9.top_add_9ns_9s_9_2_1_Adder_5_U.u1.cin ;
wire \add_9ns_9s_9_2_1_U9.top_add_9ns_9s_9_2_1_Adder_5_U.u1.cout ;
wire [3:0] \add_9ns_9s_9_2_1_U9.top_add_9ns_9s_9_2_1_Adder_5_U.u1.s ;
wire [4:0] \add_9ns_9s_9_2_1_U9.top_add_9ns_9s_9_2_1_Adder_5_U.u2.a ;
wire [4:0] \add_9ns_9s_9_2_1_U9.top_add_9ns_9s_9_2_1_Adder_5_U.u2.b ;
wire \add_9ns_9s_9_2_1_U9.top_add_9ns_9s_9_2_1_Adder_5_U.u2.cin ;
wire \add_9ns_9s_9_2_1_U9.top_add_9ns_9s_9_2_1_Adder_5_U.u2.cout ;
wire [4:0] \add_9ns_9s_9_2_1_U9.top_add_9ns_9s_9_2_1_Adder_5_U.u2.s ;
wire \add_9s_9ns_9_2_1_U19.ce ;
wire \add_9s_9ns_9_2_1_U19.clk ;
wire [8:0] \add_9s_9ns_9_2_1_U19.din0 ;
wire [8:0] \add_9s_9ns_9_2_1_U19.din1 ;
wire [8:0] \add_9s_9ns_9_2_1_U19.dout ;
wire \add_9s_9ns_9_2_1_U19.reset ;
wire [8:0] \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_13_U.a ;
wire [8:0] \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_13_U.ain_s0 ;
wire [8:0] \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_13_U.b ;
wire [8:0] \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_13_U.bin_s0 ;
wire \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_13_U.ce ;
wire \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_13_U.clk ;
wire \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_13_U.facout_s1 ;
wire \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_13_U.facout_s2 ;
wire [3:0] \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_13_U.fas_s1 ;
wire [4:0] \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_13_U.fas_s2 ;
wire \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_13_U.reset ;
wire [8:0] \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_13_U.s ;
wire [3:0] \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_13_U.u1.a ;
wire [3:0] \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_13_U.u1.b ;
wire \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_13_U.u1.cin ;
wire \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_13_U.u1.cout ;
wire [3:0] \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_13_U.u1.s ;
wire [4:0] \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_13_U.u2.a ;
wire [4:0] \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_13_U.u2.b ;
wire \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_13_U.u2.cin ;
wire \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_13_U.u2.cout ;
wire [4:0] \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_13_U.u2.s ;
wire and_ln340_1_fu_730_p2;
wire and_ln340_fu_718_p2;
wire and_ln785_1_fu_734_p2;
wire and_ln785_fu_760_p2;
wire and_ln786_fu_638_p2;
wire ap_CS_fsm_state1;
wire ap_CS_fsm_state10;
wire ap_CS_fsm_state11;
wire ap_CS_fsm_state12;
wire ap_CS_fsm_state13;
wire ap_CS_fsm_state14;
wire ap_CS_fsm_state15;
wire ap_CS_fsm_state16;
wire ap_CS_fsm_state17;
wire ap_CS_fsm_state18;
wire ap_CS_fsm_state19;
wire ap_CS_fsm_state2;
wire ap_CS_fsm_state20;
wire ap_CS_fsm_state21;
wire ap_CS_fsm_state22;
wire ap_CS_fsm_state23;
wire ap_CS_fsm_state24;
wire ap_CS_fsm_state25;
wire ap_CS_fsm_state26;
wire ap_CS_fsm_state27;
wire ap_CS_fsm_state28;
wire ap_CS_fsm_state29;
wire ap_CS_fsm_state3;
wire ap_CS_fsm_state30;
wire ap_CS_fsm_state31;
wire ap_CS_fsm_state32;
wire ap_CS_fsm_state33;
wire ap_CS_fsm_state34;
wire ap_CS_fsm_state35;
wire ap_CS_fsm_state36;
wire ap_CS_fsm_state37;
wire ap_CS_fsm_state38;
wire ap_CS_fsm_state4;
wire ap_CS_fsm_state5;
wire ap_CS_fsm_state6;
wire ap_CS_fsm_state7;
wire ap_CS_fsm_state8;
wire ap_CS_fsm_state9;
wire [37:0] ap_NS_fsm;
wire ap_clk;
wire ap_done;
wire ap_idle;
wire ap_ready;
wire ap_rst;
wire ap_start;
wire \ashr_16s_4ns_16_7_1_U4.ce ;
wire \ashr_16s_4ns_16_7_1_U4.clk ;
wire [15:0] \ashr_16s_4ns_16_7_1_U4.din0 ;
wire [15:0] \ashr_16s_4ns_16_7_1_U4.din1 ;
wire [3:0] \ashr_16s_4ns_16_7_1_U4.din1_cast ;
wire [3:0] \ashr_16s_4ns_16_7_1_U4.din1_mask ;
wire [15:0] \ashr_16s_4ns_16_7_1_U4.dout ;
wire \ashr_16s_4ns_16_7_1_U4.reset ;
wire \ashr_8ns_8s_8_7_1_U11.ce ;
wire \ashr_8ns_8s_8_7_1_U11.clk ;
wire [7:0] \ashr_8ns_8s_8_7_1_U11.din0 ;
wire [7:0] \ashr_8ns_8s_8_7_1_U11.din1 ;
wire [7:0] \ashr_8ns_8s_8_7_1_U11.din1_cast ;
wire [7:0] \ashr_8ns_8s_8_7_1_U11.din1_mask ;
wire [7:0] \ashr_8ns_8s_8_7_1_U11.dout ;
wire \ashr_8ns_8s_8_7_1_U11.reset ;
wire [31:0] grp_fu_1002_p1;
wire [31:0] grp_fu_1002_p2;
wire [31:0] grp_fu_1011_p1;
wire [31:0] grp_fu_1011_p2;
wire [31:0] grp_fu_1019_p0;
wire [31:0] grp_fu_1019_p2;
wire [3:0] grp_fu_247_p2;
wire [5:0] grp_fu_289_p0;
wire [5:0] grp_fu_289_p1;
wire [5:0] grp_fu_289_p2;
wire [15:0] grp_fu_316_p2;
wire [15:0] grp_fu_322_p2;
wire [17:0] grp_fu_336_p2;
wire [2:0] grp_fu_349_p0;
wire [2:0] grp_fu_349_p1;
wire [2:0] grp_fu_349_p2;
wire [4:0] grp_fu_381_p2;
wire [5:0] grp_fu_420_p1;
wire [5:0] grp_fu_420_p2;
wire [8:0] grp_fu_442_p0;
wire [8:0] grp_fu_442_p1;
wire [8:0] grp_fu_442_p2;
wire [7:0] grp_fu_485_p1;
wire [7:0] grp_fu_485_p2;
wire [7:0] grp_fu_493_p1;
wire [7:0] grp_fu_493_p2;
wire [5:0] grp_fu_498_p2;
wire [3:0] grp_fu_549_p2;
wire [6:0] grp_fu_653_p0;
wire [6:0] grp_fu_653_p1;
wire [6:0] grp_fu_653_p2;
wire [2:0] grp_fu_659_p0;
wire [2:0] grp_fu_659_p1;
wire [2:0] grp_fu_659_p2;
wire [6:0] grp_fu_774_p0;
wire [6:0] grp_fu_774_p2;
wire [10:0] grp_fu_810_p0;
wire [10:0] grp_fu_810_p1;
wire [10:0] grp_fu_810_p2;
wire [9:0] grp_fu_824_p0;
wire [9:0] grp_fu_824_p1;
wire [9:0] grp_fu_824_p2;
wire [8:0] grp_fu_843_p0;
wire [8:0] grp_fu_843_p2;
wire [39:0] grp_fu_883_p0;
wire [39:0] grp_fu_883_p1;
wire [39:0] grp_fu_883_p2;
wire [31:0] grp_fu_909_p2;
wire [37:0] grp_fu_948_p0;
wire [37:0] grp_fu_948_p1;
wire [37:0] grp_fu_948_p2;
wire [31:0] grp_fu_974_p2;
wire [15:0] icmp_ln1494_fu_376_p1;
wire icmp_ln1494_fu_376_p2;
wire [15:0] icmp_ln1499_fu_307_p1;
wire icmp_ln1499_fu_307_p2;
wire icmp_ln768_fu_554_p2;
wire icmp_ln786_fu_559_p2;
wire icmp_ln851_1_fu_544_p2;
wire icmp_ln851_2_fu_816_p2;
wire icmp_ln851_3_fu_893_p2;
wire icmp_ln851_4_fu_958_p2;
wire icmp_ln851_fu_452_p2;
wire [4:0] lhs_V_fu_274_p3;
wire [4:0] lhs_fu_426_p3;
wire \mul_16s_2s_18_7_1_U5.ce ;
wire \mul_16s_2s_18_7_1_U5.clk ;
wire [15:0] \mul_16s_2s_18_7_1_U5.din0 ;
wire [1:0] \mul_16s_2s_18_7_1_U5.din1 ;
wire [17:0] \mul_16s_2s_18_7_1_U5.dout ;
wire \mul_16s_2s_18_7_1_U5.reset ;
wire [15:0] \mul_16s_2s_18_7_1_U5.top_mul_16s_2s_18_7_1_Mul_DSP_0_U.a ;
wire [1:0] \mul_16s_2s_18_7_1_U5.top_mul_16s_2s_18_7_1_Mul_DSP_0_U.b ;
wire \mul_16s_2s_18_7_1_U5.top_mul_16s_2s_18_7_1_Mul_DSP_0_U.ce ;
wire \mul_16s_2s_18_7_1_U5.top_mul_16s_2s_18_7_1_Mul_DSP_0_U.clk ;
wire [17:0] \mul_16s_2s_18_7_1_U5.top_mul_16s_2s_18_7_1_Mul_DSP_0_U.p ;
wire [17:0] \mul_16s_2s_18_7_1_U5.top_mul_16s_2s_18_7_1_Mul_DSP_0_U.tmp_product ;
wire [1:0] op_0;
wire [7:0] op_1;
wire [7:0] op_12_V_fu_779_p3;
wire [7:0] op_13;
wire [7:0] op_15;
wire [3:0] op_16;
wire [3:0] op_17;
wire [1:0] op_2;
wire [7:0] op_3;
wire [31:0] op_30;
wire op_30_ap_vld;
wire [15:0] op_4;
wire [3:0] op_5;
wire [1:0] op_7;
wire [1:0] op_8;
wire [1:0] op_9_V_fu_267_p3;
wire or_ln340_fu_628_p2;
wire or_ln785_1_fu_755_p2;
wire or_ln785_2_fu_738_p2;
wire or_ln785_fu_583_p2;
wire or_ln786_fu_623_p2;
wire overflow_fu_614_p2;
wire p_Result_10_fu_979_p3;
wire p_Result_13_fu_665_p3;
wire [7:0] p_Result_4_fu_703_p4;
wire p_Result_5_fu_592_p3;
wire p_Result_6_fu_386_p3;
wire p_Result_8_fu_849_p3;
wire p_Result_9_fu_914_p3;
wire p_Result_s_fu_564_p3;
wire [6:0] p_Val2_3_fu_698_p2;
wire [15:0] r_V_fu_503_p3;
wire [7:0] r_fu_784_p3;
wire [5:0] ret_V_17_fu_576_p3;
wire [3:0] ret_V_18_fu_604_p3;
wire [4:0] ret_V_20_fu_402_p3;
wire [31:0] ret_V_24_fu_991_p3;
wire [9:0] rhs_2_fu_799_p3;
wire [36:0] rhs_3_fu_937_p3;
wire sel_tmp11_fu_744_p2;
wire [7:0] select_ln340_fu_723_p3;
wire [31:0] select_ln353_1_fu_926_p3;
wire [8:0] select_ln353_fu_861_p3;
wire [7:0] select_ln785_fu_765_p3;
wire [3:0] select_ln850_1_fu_599_p3;
wire [4:0] select_ln850_2_fu_396_p3;
wire [31:0] select_ln850_5_fu_986_p3;
wire [8:0] select_ln850_6_fu_856_p3;
wire [31:0] select_ln850_7_fu_921_p3;
wire [5:0] select_ln850_fu_571_p3;
wire [15:0] sext_ln1499_fu_303_p1;
wire [1:0] sext_ln215_1_fu_346_p0;
wire [1:0] sext_ln215_fu_342_p0;
wire [7:0] sext_ln703_1_fu_868_p0;
wire [7:0] sext_ln703_2_fu_933_p0;
wire [7:0] sext_ln703_fu_438_p0;
wire [8:0] sext_ln850_fu_840_p1;
wire [1:0] sext_ln886_fu_253_p0;
wire [3:0] sext_ln886_fu_253_p1;
wire \shl_16s_4ns_16_7_1_U3.ce ;
wire \shl_16s_4ns_16_7_1_U3.clk ;
wire [15:0] \shl_16s_4ns_16_7_1_U3.din0 ;
wire [15:0] \shl_16s_4ns_16_7_1_U3.din1 ;
wire [3:0] \shl_16s_4ns_16_7_1_U3.din1_cast ;
wire [3:0] \shl_16s_4ns_16_7_1_U3.din1_mask ;
wire [15:0] \shl_16s_4ns_16_7_1_U3.dout ;
wire \shl_16s_4ns_16_7_1_U3.reset ;
wire \shl_8ns_8s_8_7_1_U10.ce ;
wire \shl_8ns_8s_8_7_1_U10.clk ;
wire [7:0] \shl_8ns_8s_8_7_1_U10.din0 ;
wire [7:0] \shl_8ns_8s_8_7_1_U10.din1 ;
wire [7:0] \shl_8ns_8s_8_7_1_U10.din1_cast ;
wire [7:0] \shl_8ns_8s_8_7_1_U10.din1_mask ;
wire [7:0] \shl_8ns_8s_8_7_1_U10.dout ;
wire \shl_8ns_8s_8_7_1_U10.reset ;
wire [6:0] shl_ln728_2_fu_365_p3;
wire [13:0] shl_ln_fu_295_p3;
wire signbit_fu_257_p2;
wire \sub_4ns_4ns_4_2_1_U1.ce ;
wire \sub_4ns_4ns_4_2_1_U1.clk ;
wire [3:0] \sub_4ns_4ns_4_2_1_U1.din0 ;
wire [3:0] \sub_4ns_4ns_4_2_1_U1.din1 ;
wire [3:0] \sub_4ns_4ns_4_2_1_U1.dout ;
wire \sub_4ns_4ns_4_2_1_U1.reset ;
wire [3:0] \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.a ;
wire [3:0] \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.ain_s0 ;
wire [3:0] \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.b ;
wire [3:0] \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.bin_s0 ;
wire \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.ce ;
wire \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.clk ;
wire \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.facout_s1 ;
wire \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.facout_s2 ;
wire [1:0] \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.fas_s1 ;
wire [1:0] \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.fas_s2 ;
wire \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.reset ;
wire [3:0] \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.s ;
wire [1:0] \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.u1.a ;
wire [1:0] \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.u1.b ;
wire \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.u1.cin ;
wire \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.u1.cout ;
wire [1:0] \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.u1.s ;
wire [1:0] \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.u2.a ;
wire [1:0] \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.u2.b ;
wire \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.u2.cin ;
wire \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.u2.cout ;
wire [1:0] \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.u2.s ;
wire \sub_6ns_6s_6_2_1_U8.ce ;
wire \sub_6ns_6s_6_2_1_U8.clk ;
wire [5:0] \sub_6ns_6s_6_2_1_U8.din0 ;
wire [5:0] \sub_6ns_6s_6_2_1_U8.din1 ;
wire [5:0] \sub_6ns_6s_6_2_1_U8.dout ;
wire \sub_6ns_6s_6_2_1_U8.reset ;
wire [5:0] \sub_6ns_6s_6_2_1_U8.top_sub_6ns_6s_6_2_1_Adder_4_U.a ;
wire [5:0] \sub_6ns_6s_6_2_1_U8.top_sub_6ns_6s_6_2_1_Adder_4_U.ain_s0 ;
wire [5:0] \sub_6ns_6s_6_2_1_U8.top_sub_6ns_6s_6_2_1_Adder_4_U.b ;
wire [5:0] \sub_6ns_6s_6_2_1_U8.top_sub_6ns_6s_6_2_1_Adder_4_U.bin_s0 ;
wire \sub_6ns_6s_6_2_1_U8.top_sub_6ns_6s_6_2_1_Adder_4_U.ce ;
wire \sub_6ns_6s_6_2_1_U8.top_sub_6ns_6s_6_2_1_Adder_4_U.clk ;
wire \sub_6ns_6s_6_2_1_U8.top_sub_6ns_6s_6_2_1_Adder_4_U.facout_s1 ;
wire \sub_6ns_6s_6_2_1_U8.top_sub_6ns_6s_6_2_1_Adder_4_U.facout_s2 ;
wire [2:0] \sub_6ns_6s_6_2_1_U8.top_sub_6ns_6s_6_2_1_Adder_4_U.fas_s1 ;
wire [2:0] \sub_6ns_6s_6_2_1_U8.top_sub_6ns_6s_6_2_1_Adder_4_U.fas_s2 ;
wire \sub_6ns_6s_6_2_1_U8.top_sub_6ns_6s_6_2_1_Adder_4_U.reset ;
wire [5:0] \sub_6ns_6s_6_2_1_U8.top_sub_6ns_6s_6_2_1_Adder_4_U.s ;
wire [2:0] \sub_6ns_6s_6_2_1_U8.top_sub_6ns_6s_6_2_1_Adder_4_U.u1.a ;
wire [2:0] \sub_6ns_6s_6_2_1_U8.top_sub_6ns_6s_6_2_1_Adder_4_U.u1.b ;
wire \sub_6ns_6s_6_2_1_U8.top_sub_6ns_6s_6_2_1_Adder_4_U.u1.cin ;
wire \sub_6ns_6s_6_2_1_U8.top_sub_6ns_6s_6_2_1_Adder_4_U.u1.cout ;
wire [2:0] \sub_6ns_6s_6_2_1_U8.top_sub_6ns_6s_6_2_1_Adder_4_U.u1.s ;
wire [2:0] \sub_6ns_6s_6_2_1_U8.top_sub_6ns_6s_6_2_1_Adder_4_U.u2.a ;
wire [2:0] \sub_6ns_6s_6_2_1_U8.top_sub_6ns_6s_6_2_1_Adder_4_U.u2.b ;
wire \sub_6ns_6s_6_2_1_U8.top_sub_6ns_6s_6_2_1_Adder_4_U.u2.cin ;
wire \sub_6ns_6s_6_2_1_U8.top_sub_6ns_6s_6_2_1_Adder_4_U.u2.cout ;
wire [2:0] \sub_6ns_6s_6_2_1_U8.top_sub_6ns_6s_6_2_1_Adder_4_U.u2.s ;
wire \sub_6s_6ns_6_2_1_U2.ce ;
wire \sub_6s_6ns_6_2_1_U2.clk ;
wire [5:0] \sub_6s_6ns_6_2_1_U2.din0 ;
wire [5:0] \sub_6s_6ns_6_2_1_U2.din1 ;
wire [5:0] \sub_6s_6ns_6_2_1_U2.dout ;
wire \sub_6s_6ns_6_2_1_U2.reset ;
wire [5:0] \sub_6s_6ns_6_2_1_U2.top_sub_6s_6ns_6_2_1_Adder_1_U.a ;
wire [5:0] \sub_6s_6ns_6_2_1_U2.top_sub_6s_6ns_6_2_1_Adder_1_U.ain_s0 ;
wire [5:0] \sub_6s_6ns_6_2_1_U2.top_sub_6s_6ns_6_2_1_Adder_1_U.b ;
wire [5:0] \sub_6s_6ns_6_2_1_U2.top_sub_6s_6ns_6_2_1_Adder_1_U.bin_s0 ;
wire \sub_6s_6ns_6_2_1_U2.top_sub_6s_6ns_6_2_1_Adder_1_U.ce ;
wire \sub_6s_6ns_6_2_1_U2.top_sub_6s_6ns_6_2_1_Adder_1_U.clk ;
wire \sub_6s_6ns_6_2_1_U2.top_sub_6s_6ns_6_2_1_Adder_1_U.facout_s1 ;
wire \sub_6s_6ns_6_2_1_U2.top_sub_6s_6ns_6_2_1_Adder_1_U.facout_s2 ;
wire [2:0] \sub_6s_6ns_6_2_1_U2.top_sub_6s_6ns_6_2_1_Adder_1_U.fas_s1 ;
wire [2:0] \sub_6s_6ns_6_2_1_U2.top_sub_6s_6ns_6_2_1_Adder_1_U.fas_s2 ;
wire \sub_6s_6ns_6_2_1_U2.top_sub_6s_6ns_6_2_1_Adder_1_U.reset ;
wire [5:0] \sub_6s_6ns_6_2_1_U2.top_sub_6s_6ns_6_2_1_Adder_1_U.s ;
wire [2:0] \sub_6s_6ns_6_2_1_U2.top_sub_6s_6ns_6_2_1_Adder_1_U.u1.a ;
wire [2:0] \sub_6s_6ns_6_2_1_U2.top_sub_6s_6ns_6_2_1_Adder_1_U.u1.b ;
wire \sub_6s_6ns_6_2_1_U2.top_sub_6s_6ns_6_2_1_Adder_1_U.u1.cin ;
wire \sub_6s_6ns_6_2_1_U2.top_sub_6s_6ns_6_2_1_Adder_1_U.u1.cout ;
wire [2:0] \sub_6s_6ns_6_2_1_U2.top_sub_6s_6ns_6_2_1_Adder_1_U.u1.s ;
wire [2:0] \sub_6s_6ns_6_2_1_U2.top_sub_6s_6ns_6_2_1_Adder_1_U.u2.a ;
wire [2:0] \sub_6s_6ns_6_2_1_U2.top_sub_6s_6ns_6_2_1_Adder_1_U.u2.b ;
wire \sub_6s_6ns_6_2_1_U2.top_sub_6s_6ns_6_2_1_Adder_1_U.u2.cin ;
wire \sub_6s_6ns_6_2_1_U2.top_sub_6s_6ns_6_2_1_Adder_1_U.u2.cout ;
wire [2:0] \sub_6s_6ns_6_2_1_U2.top_sub_6s_6ns_6_2_1_Adder_1_U.u2.s ;
wire [15:0] tmp_13_fu_872_p3;
wire tmp_6_fu_672_p3;
wire tmp_7_fu_679_p3;
wire [5:0] trunc_ln851_1_fu_478_p1;
wire trunc_ln851_2_fu_393_p1;
wire [2:0] trunc_ln851_3_fu_789_p1;
wire [7:0] trunc_ln851_4_fu_889_p0;
wire [6:0] trunc_ln851_4_fu_889_p1;
wire [7:0] trunc_ln851_5_fu_954_p0;
wire [4:0] trunc_ln851_5_fu_954_p1;
wire [7:0] trunc_ln851_fu_448_p0;
wire [2:0] trunc_ln851_fu_448_p1;
wire [3:0] ush_fu_262_p3;
wire xor_ln340_fu_713_p2;
wire xor_ln365_1_fu_692_p2;
wire xor_ln365_fu_686_p2;
wire xor_ln785_1_fu_750_p2;
wire xor_ln785_fu_587_p2;
wire xor_ln786_1_fu_633_p2;
wire xor_ln786_fu_618_p2;
wire [15:0] zext_ln1367_fu_313_p1;
wire [15:0] zext_ln1494_fu_372_p1;


assign _0070_ = icmp_ln851_3_reg_1474 & ap_CS_fsm[25];
assign _0071_ = icmp_ln851_4_reg_1511 & ap_CS_fsm[30];
assign _0072_ = icmp_ln851_2_reg_1422 & ap_CS_fsm[20];
assign _0073_ = _0082_ & ap_CS_fsm[9];
assign _0074_ = ap_CS_fsm[15] & _0083_;
assign _0075_ = ap_CS_fsm[11] & _0084_;
assign _0076_ = _0085_ & ap_CS_fsm[15];
assign _0077_ = ap_CS_fsm[8] & p_Result_14_reg_1147;
assign _0078_ = isNeg_reg_1033 & ap_CS_fsm[9];
assign _0079_ = ap_CS_fsm[15] & p_Result_14_reg_1147;
assign _0080_ = _0086_ & ap_CS_fsm[0];
assign _0081_ = ap_start & ap_CS_fsm[0];
assign and_ln340_1_fu_730_p2 = or_ln786_reg_1314 & or_ln340_reg_1320;
assign and_ln340_fu_718_p2 = xor_ln340_fu_713_p2 & or_ln786_reg_1314;
assign and_ln785_1_fu_734_p2 = xor_ln785_reg_1298 & and_ln786_reg_1326;
assign and_ln785_fu_760_p2 = or_ln785_1_fu_755_p2 & and_ln786_reg_1326;
assign and_ln786_fu_638_p2 = xor_ln786_1_fu_633_p2 & p_Result_12_reg_1248;
assign overflow_fu_614_p2 = xor_ln785_reg_1298 & or_ln785_reg_1292;
assign sel_tmp11_fu_744_p2 = xor_ln365_1_fu_692_p2 & or_ln785_2_fu_738_p2;
assign xor_ln340_fu_713_p2 = ~ or_ln340_reg_1320;
assign xor_ln785_1_fu_750_p2 = ~ or_ln785_reg_1292;
assign xor_ln786_1_fu_633_p2 = ~ icmp_ln786_reg_1276;
assign xor_ln786_fu_618_p2 = ~ p_Result_12_reg_1248;
assign xor_ln365_1_fu_692_p2 = ~ xor_ln365_fu_686_p2;
assign xor_ln785_fu_587_p2 = ~ p_Result_11_reg_1233;
assign p_Val2_3_fu_698_p2 = ~ p_Val2_2_reg_1240[6:0];
assign _0082_ = ~ isNeg_reg_1033;
assign _0083_ = ~ p_Result_14_reg_1147;
assign _0084_ = ~ icmp_ln851_reg_1167;
assign _0085_ = ~ sel_tmp11_reg_1352;
assign _0086_ = ~ ap_start;
assign _0087_ = ! trunc_ln851_1_reg_1211;
assign _0088_ = ! op_1[2:0];
always @(posedge \add_10ns_10s_10_2_1_U18.top_add_10ns_10s_10_2_1_Adder_12_U.clk )
\add_10ns_10s_10_2_1_U18.top_add_10ns_10s_10_2_1_Adder_12_U.bin_s1  <= _0090_;
always @(posedge \add_10ns_10s_10_2_1_U18.top_add_10ns_10s_10_2_1_Adder_12_U.clk )
\add_10ns_10s_10_2_1_U18.top_add_10ns_10s_10_2_1_Adder_12_U.ain_s1  <= _0089_;
always @(posedge \add_10ns_10s_10_2_1_U18.top_add_10ns_10s_10_2_1_Adder_12_U.clk )
\add_10ns_10s_10_2_1_U18.top_add_10ns_10s_10_2_1_Adder_12_U.sum_s1  <= _0092_;
always @(posedge \add_10ns_10s_10_2_1_U18.top_add_10ns_10s_10_2_1_Adder_12_U.clk )
\add_10ns_10s_10_2_1_U18.top_add_10ns_10s_10_2_1_Adder_12_U.carry_s1  <= _0091_;
assign _0090_ = \add_10ns_10s_10_2_1_U18.top_add_10ns_10s_10_2_1_Adder_12_U.ce  ? \add_10ns_10s_10_2_1_U18.top_add_10ns_10s_10_2_1_Adder_12_U.b [9:5] : \add_10ns_10s_10_2_1_U18.top_add_10ns_10s_10_2_1_Adder_12_U.bin_s1 ;
assign _0089_ = \add_10ns_10s_10_2_1_U18.top_add_10ns_10s_10_2_1_Adder_12_U.ce  ? \add_10ns_10s_10_2_1_U18.top_add_10ns_10s_10_2_1_Adder_12_U.a [9:5] : \add_10ns_10s_10_2_1_U18.top_add_10ns_10s_10_2_1_Adder_12_U.ain_s1 ;
assign _0091_ = \add_10ns_10s_10_2_1_U18.top_add_10ns_10s_10_2_1_Adder_12_U.ce  ? \add_10ns_10s_10_2_1_U18.top_add_10ns_10s_10_2_1_Adder_12_U.facout_s1  : \add_10ns_10s_10_2_1_U18.top_add_10ns_10s_10_2_1_Adder_12_U.carry_s1 ;
assign _0092_ = \add_10ns_10s_10_2_1_U18.top_add_10ns_10s_10_2_1_Adder_12_U.ce  ? \add_10ns_10s_10_2_1_U18.top_add_10ns_10s_10_2_1_Adder_12_U.fas_s1  : \add_10ns_10s_10_2_1_U18.top_add_10ns_10s_10_2_1_Adder_12_U.sum_s1 ;
assign _0093_ = \add_10ns_10s_10_2_1_U18.top_add_10ns_10s_10_2_1_Adder_12_U.u1.a  + \add_10ns_10s_10_2_1_U18.top_add_10ns_10s_10_2_1_Adder_12_U.u1.b ;
assign { \add_10ns_10s_10_2_1_U18.top_add_10ns_10s_10_2_1_Adder_12_U.u1.cout , \add_10ns_10s_10_2_1_U18.top_add_10ns_10s_10_2_1_Adder_12_U.u1.s  } = _0093_ + \add_10ns_10s_10_2_1_U18.top_add_10ns_10s_10_2_1_Adder_12_U.u1.cin ;
assign _0094_ = \add_10ns_10s_10_2_1_U18.top_add_10ns_10s_10_2_1_Adder_12_U.u2.a  + \add_10ns_10s_10_2_1_U18.top_add_10ns_10s_10_2_1_Adder_12_U.u2.b ;
assign { \add_10ns_10s_10_2_1_U18.top_add_10ns_10s_10_2_1_Adder_12_U.u2.cout , \add_10ns_10s_10_2_1_U18.top_add_10ns_10s_10_2_1_Adder_12_U.u2.s  } = _0094_ + \add_10ns_10s_10_2_1_U18.top_add_10ns_10s_10_2_1_Adder_12_U.u2.cin ;
always @(posedge \add_11s_11s_11_2_1_U17.top_add_11s_11s_11_2_1_Adder_11_U.clk )
\add_11s_11s_11_2_1_U17.top_add_11s_11s_11_2_1_Adder_11_U.bin_s1  <= _0096_;
always @(posedge \add_11s_11s_11_2_1_U17.top_add_11s_11s_11_2_1_Adder_11_U.clk )
\add_11s_11s_11_2_1_U17.top_add_11s_11s_11_2_1_Adder_11_U.ain_s1  <= _0095_;
always @(posedge \add_11s_11s_11_2_1_U17.top_add_11s_11s_11_2_1_Adder_11_U.clk )
\add_11s_11s_11_2_1_U17.top_add_11s_11s_11_2_1_Adder_11_U.sum_s1  <= _0098_;
always @(posedge \add_11s_11s_11_2_1_U17.top_add_11s_11s_11_2_1_Adder_11_U.clk )
\add_11s_11s_11_2_1_U17.top_add_11s_11s_11_2_1_Adder_11_U.carry_s1  <= _0097_;
assign _0096_ = \add_11s_11s_11_2_1_U17.top_add_11s_11s_11_2_1_Adder_11_U.ce  ? \add_11s_11s_11_2_1_U17.top_add_11s_11s_11_2_1_Adder_11_U.b [10:5] : \add_11s_11s_11_2_1_U17.top_add_11s_11s_11_2_1_Adder_11_U.bin_s1 ;
assign _0095_ = \add_11s_11s_11_2_1_U17.top_add_11s_11s_11_2_1_Adder_11_U.ce  ? \add_11s_11s_11_2_1_U17.top_add_11s_11s_11_2_1_Adder_11_U.a [10:5] : \add_11s_11s_11_2_1_U17.top_add_11s_11s_11_2_1_Adder_11_U.ain_s1 ;
assign _0097_ = \add_11s_11s_11_2_1_U17.top_add_11s_11s_11_2_1_Adder_11_U.ce  ? \add_11s_11s_11_2_1_U17.top_add_11s_11s_11_2_1_Adder_11_U.facout_s1  : \add_11s_11s_11_2_1_U17.top_add_11s_11s_11_2_1_Adder_11_U.carry_s1 ;
assign _0098_ = \add_11s_11s_11_2_1_U17.top_add_11s_11s_11_2_1_Adder_11_U.ce  ? \add_11s_11s_11_2_1_U17.top_add_11s_11s_11_2_1_Adder_11_U.fas_s1  : \add_11s_11s_11_2_1_U17.top_add_11s_11s_11_2_1_Adder_11_U.sum_s1 ;
assign _0099_ = \add_11s_11s_11_2_1_U17.top_add_11s_11s_11_2_1_Adder_11_U.u1.a  + \add_11s_11s_11_2_1_U17.top_add_11s_11s_11_2_1_Adder_11_U.u1.b ;
assign { \add_11s_11s_11_2_1_U17.top_add_11s_11s_11_2_1_Adder_11_U.u1.cout , \add_11s_11s_11_2_1_U17.top_add_11s_11s_11_2_1_Adder_11_U.u1.s  } = _0099_ + \add_11s_11s_11_2_1_U17.top_add_11s_11s_11_2_1_Adder_11_U.u1.cin ;
assign _0100_ = \add_11s_11s_11_2_1_U17.top_add_11s_11s_11_2_1_Adder_11_U.u2.a  + \add_11s_11s_11_2_1_U17.top_add_11s_11s_11_2_1_Adder_11_U.u2.b ;
assign { \add_11s_11s_11_2_1_U17.top_add_11s_11s_11_2_1_Adder_11_U.u2.cout , \add_11s_11s_11_2_1_U17.top_add_11s_11s_11_2_1_Adder_11_U.u2.s  } = _0100_ + \add_11s_11s_11_2_1_U17.top_add_11s_11s_11_2_1_Adder_11_U.u2.cin ;
always @(posedge \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.clk )
\add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.bin_s1  <= _0102_;
always @(posedge \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.clk )
\add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.ain_s1  <= _0101_;
always @(posedge \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.clk )
\add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.sum_s1  <= _0104_;
always @(posedge \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.clk )
\add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.carry_s1  <= _0103_;
assign _0102_ = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.ce  ? \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.b [31:16] : \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.bin_s1 ;
assign _0101_ = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.ce  ? \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.a [31:16] : \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.ain_s1 ;
assign _0103_ = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.ce  ? \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.facout_s1  : \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.carry_s1 ;
assign _0104_ = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.ce  ? \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.fas_s1  : \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.sum_s1 ;
assign _0105_ = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.a  + \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.b ;
assign { \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.cout , \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.s  } = _0105_ + \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.cin ;
assign _0106_ = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.a  + \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.b ;
assign { \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.cout , \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.s  } = _0106_ + \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.cin ;
always @(posedge \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.clk )
\add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.bin_s1  <= _0108_;
always @(posedge \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.clk )
\add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.ain_s1  <= _0107_;
always @(posedge \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.clk )
\add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.sum_s1  <= _0110_;
always @(posedge \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.clk )
\add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.carry_s1  <= _0109_;
assign _0108_ = \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.ce  ? \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.b [31:16] : \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.bin_s1 ;
assign _0107_ = \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.ce  ? \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.a [31:16] : \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.ain_s1 ;
assign _0109_ = \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.ce  ? \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.facout_s1  : \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.carry_s1 ;
assign _0110_ = \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.ce  ? \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.fas_s1  : \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.sum_s1 ;
assign _0111_ = \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.a  + \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.b ;
assign { \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.cout , \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.s  } = _0111_ + \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.cin ;
assign _0112_ = \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.a  + \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.b ;
assign { \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.cout , \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.s  } = _0112_ + \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.cin ;
always @(posedge \add_32ns_32s_32_2_1_U24.top_add_32ns_32s_32_2_1_Adder_17_U.clk )
\add_32ns_32s_32_2_1_U24.top_add_32ns_32s_32_2_1_Adder_17_U.bin_s1  <= _0114_;
always @(posedge \add_32ns_32s_32_2_1_U24.top_add_32ns_32s_32_2_1_Adder_17_U.clk )
\add_32ns_32s_32_2_1_U24.top_add_32ns_32s_32_2_1_Adder_17_U.ain_s1  <= _0113_;
always @(posedge \add_32ns_32s_32_2_1_U24.top_add_32ns_32s_32_2_1_Adder_17_U.clk )
\add_32ns_32s_32_2_1_U24.top_add_32ns_32s_32_2_1_Adder_17_U.sum_s1  <= _0116_;
always @(posedge \add_32ns_32s_32_2_1_U24.top_add_32ns_32s_32_2_1_Adder_17_U.clk )
\add_32ns_32s_32_2_1_U24.top_add_32ns_32s_32_2_1_Adder_17_U.carry_s1  <= _0115_;
assign _0114_ = \add_32ns_32s_32_2_1_U24.top_add_32ns_32s_32_2_1_Adder_17_U.ce  ? \add_32ns_32s_32_2_1_U24.top_add_32ns_32s_32_2_1_Adder_17_U.b [31:16] : \add_32ns_32s_32_2_1_U24.top_add_32ns_32s_32_2_1_Adder_17_U.bin_s1 ;
assign _0113_ = \add_32ns_32s_32_2_1_U24.top_add_32ns_32s_32_2_1_Adder_17_U.ce  ? \add_32ns_32s_32_2_1_U24.top_add_32ns_32s_32_2_1_Adder_17_U.a [31:16] : \add_32ns_32s_32_2_1_U24.top_add_32ns_32s_32_2_1_Adder_17_U.ain_s1 ;
assign _0115_ = \add_32ns_32s_32_2_1_U24.top_add_32ns_32s_32_2_1_Adder_17_U.ce  ? \add_32ns_32s_32_2_1_U24.top_add_32ns_32s_32_2_1_Adder_17_U.facout_s1  : \add_32ns_32s_32_2_1_U24.top_add_32ns_32s_32_2_1_Adder_17_U.carry_s1 ;
assign _0116_ = \add_32ns_32s_32_2_1_U24.top_add_32ns_32s_32_2_1_Adder_17_U.ce  ? \add_32ns_32s_32_2_1_U24.top_add_32ns_32s_32_2_1_Adder_17_U.fas_s1  : \add_32ns_32s_32_2_1_U24.top_add_32ns_32s_32_2_1_Adder_17_U.sum_s1 ;
assign _0117_ = \add_32ns_32s_32_2_1_U24.top_add_32ns_32s_32_2_1_Adder_17_U.u1.a  + \add_32ns_32s_32_2_1_U24.top_add_32ns_32s_32_2_1_Adder_17_U.u1.b ;
assign { \add_32ns_32s_32_2_1_U24.top_add_32ns_32s_32_2_1_Adder_17_U.u1.cout , \add_32ns_32s_32_2_1_U24.top_add_32ns_32s_32_2_1_Adder_17_U.u1.s  } = _0117_ + \add_32ns_32s_32_2_1_U24.top_add_32ns_32s_32_2_1_Adder_17_U.u1.cin ;
assign _0118_ = \add_32ns_32s_32_2_1_U24.top_add_32ns_32s_32_2_1_Adder_17_U.u2.a  + \add_32ns_32s_32_2_1_U24.top_add_32ns_32s_32_2_1_Adder_17_U.u2.b ;
assign { \add_32ns_32s_32_2_1_U24.top_add_32ns_32s_32_2_1_Adder_17_U.u2.cout , \add_32ns_32s_32_2_1_U24.top_add_32ns_32s_32_2_1_Adder_17_U.u2.s  } = _0118_ + \add_32ns_32s_32_2_1_U24.top_add_32ns_32s_32_2_1_Adder_17_U.u2.cin ;
always @(posedge \add_32ns_32s_32_2_1_U25.top_add_32ns_32s_32_2_1_Adder_17_U.clk )
\add_32ns_32s_32_2_1_U25.top_add_32ns_32s_32_2_1_Adder_17_U.bin_s1  <= _0120_;
always @(posedge \add_32ns_32s_32_2_1_U25.top_add_32ns_32s_32_2_1_Adder_17_U.clk )
\add_32ns_32s_32_2_1_U25.top_add_32ns_32s_32_2_1_Adder_17_U.ain_s1  <= _0119_;
always @(posedge \add_32ns_32s_32_2_1_U25.top_add_32ns_32s_32_2_1_Adder_17_U.clk )
\add_32ns_32s_32_2_1_U25.top_add_32ns_32s_32_2_1_Adder_17_U.sum_s1  <= _0122_;
always @(posedge \add_32ns_32s_32_2_1_U25.top_add_32ns_32s_32_2_1_Adder_17_U.clk )
\add_32ns_32s_32_2_1_U25.top_add_32ns_32s_32_2_1_Adder_17_U.carry_s1  <= _0121_;
assign _0120_ = \add_32ns_32s_32_2_1_U25.top_add_32ns_32s_32_2_1_Adder_17_U.ce  ? \add_32ns_32s_32_2_1_U25.top_add_32ns_32s_32_2_1_Adder_17_U.b [31:16] : \add_32ns_32s_32_2_1_U25.top_add_32ns_32s_32_2_1_Adder_17_U.bin_s1 ;
assign _0119_ = \add_32ns_32s_32_2_1_U25.top_add_32ns_32s_32_2_1_Adder_17_U.ce  ? \add_32ns_32s_32_2_1_U25.top_add_32ns_32s_32_2_1_Adder_17_U.a [31:16] : \add_32ns_32s_32_2_1_U25.top_add_32ns_32s_32_2_1_Adder_17_U.ain_s1 ;
assign _0121_ = \add_32ns_32s_32_2_1_U25.top_add_32ns_32s_32_2_1_Adder_17_U.ce  ? \add_32ns_32s_32_2_1_U25.top_add_32ns_32s_32_2_1_Adder_17_U.facout_s1  : \add_32ns_32s_32_2_1_U25.top_add_32ns_32s_32_2_1_Adder_17_U.carry_s1 ;
assign _0122_ = \add_32ns_32s_32_2_1_U25.top_add_32ns_32s_32_2_1_Adder_17_U.ce  ? \add_32ns_32s_32_2_1_U25.top_add_32ns_32s_32_2_1_Adder_17_U.fas_s1  : \add_32ns_32s_32_2_1_U25.top_add_32ns_32s_32_2_1_Adder_17_U.sum_s1 ;
assign _0123_ = \add_32ns_32s_32_2_1_U25.top_add_32ns_32s_32_2_1_Adder_17_U.u1.a  + \add_32ns_32s_32_2_1_U25.top_add_32ns_32s_32_2_1_Adder_17_U.u1.b ;
assign { \add_32ns_32s_32_2_1_U25.top_add_32ns_32s_32_2_1_Adder_17_U.u1.cout , \add_32ns_32s_32_2_1_U25.top_add_32ns_32s_32_2_1_Adder_17_U.u1.s  } = _0123_ + \add_32ns_32s_32_2_1_U25.top_add_32ns_32s_32_2_1_Adder_17_U.u1.cin ;
assign _0124_ = \add_32ns_32s_32_2_1_U25.top_add_32ns_32s_32_2_1_Adder_17_U.u2.a  + \add_32ns_32s_32_2_1_U25.top_add_32ns_32s_32_2_1_Adder_17_U.u2.b ;
assign { \add_32ns_32s_32_2_1_U25.top_add_32ns_32s_32_2_1_Adder_17_U.u2.cout , \add_32ns_32s_32_2_1_U25.top_add_32ns_32s_32_2_1_Adder_17_U.u2.s  } = _0124_ + \add_32ns_32s_32_2_1_U25.top_add_32ns_32s_32_2_1_Adder_17_U.u2.cin ;
always @(posedge \add_32s_32ns_32_2_1_U26.top_add_32s_32ns_32_2_1_Adder_18_U.clk )
\add_32s_32ns_32_2_1_U26.top_add_32s_32ns_32_2_1_Adder_18_U.bin_s1  <= _0126_;
always @(posedge \add_32s_32ns_32_2_1_U26.top_add_32s_32ns_32_2_1_Adder_18_U.clk )
\add_32s_32ns_32_2_1_U26.top_add_32s_32ns_32_2_1_Adder_18_U.ain_s1  <= _0125_;
always @(posedge \add_32s_32ns_32_2_1_U26.top_add_32s_32ns_32_2_1_Adder_18_U.clk )
\add_32s_32ns_32_2_1_U26.top_add_32s_32ns_32_2_1_Adder_18_U.sum_s1  <= _0128_;
always @(posedge \add_32s_32ns_32_2_1_U26.top_add_32s_32ns_32_2_1_Adder_18_U.clk )
\add_32s_32ns_32_2_1_U26.top_add_32s_32ns_32_2_1_Adder_18_U.carry_s1  <= _0127_;
assign _0126_ = \add_32s_32ns_32_2_1_U26.top_add_32s_32ns_32_2_1_Adder_18_U.ce  ? \add_32s_32ns_32_2_1_U26.top_add_32s_32ns_32_2_1_Adder_18_U.b [31:16] : \add_32s_32ns_32_2_1_U26.top_add_32s_32ns_32_2_1_Adder_18_U.bin_s1 ;
assign _0125_ = \add_32s_32ns_32_2_1_U26.top_add_32s_32ns_32_2_1_Adder_18_U.ce  ? \add_32s_32ns_32_2_1_U26.top_add_32s_32ns_32_2_1_Adder_18_U.a [31:16] : \add_32s_32ns_32_2_1_U26.top_add_32s_32ns_32_2_1_Adder_18_U.ain_s1 ;
assign _0127_ = \add_32s_32ns_32_2_1_U26.top_add_32s_32ns_32_2_1_Adder_18_U.ce  ? \add_32s_32ns_32_2_1_U26.top_add_32s_32ns_32_2_1_Adder_18_U.facout_s1  : \add_32s_32ns_32_2_1_U26.top_add_32s_32ns_32_2_1_Adder_18_U.carry_s1 ;
assign _0128_ = \add_32s_32ns_32_2_1_U26.top_add_32s_32ns_32_2_1_Adder_18_U.ce  ? \add_32s_32ns_32_2_1_U26.top_add_32s_32ns_32_2_1_Adder_18_U.fas_s1  : \add_32s_32ns_32_2_1_U26.top_add_32s_32ns_32_2_1_Adder_18_U.sum_s1 ;
assign _0129_ = \add_32s_32ns_32_2_1_U26.top_add_32s_32ns_32_2_1_Adder_18_U.u1.a  + \add_32s_32ns_32_2_1_U26.top_add_32s_32ns_32_2_1_Adder_18_U.u1.b ;
assign { \add_32s_32ns_32_2_1_U26.top_add_32s_32ns_32_2_1_Adder_18_U.u1.cout , \add_32s_32ns_32_2_1_U26.top_add_32s_32ns_32_2_1_Adder_18_U.u1.s  } = _0129_ + \add_32s_32ns_32_2_1_U26.top_add_32s_32ns_32_2_1_Adder_18_U.u1.cin ;
assign _0130_ = \add_32s_32ns_32_2_1_U26.top_add_32s_32ns_32_2_1_Adder_18_U.u2.a  + \add_32s_32ns_32_2_1_U26.top_add_32s_32ns_32_2_1_Adder_18_U.u2.b ;
assign { \add_32s_32ns_32_2_1_U26.top_add_32s_32ns_32_2_1_Adder_18_U.u2.cout , \add_32s_32ns_32_2_1_U26.top_add_32s_32ns_32_2_1_Adder_18_U.u2.s  } = _0130_ + \add_32s_32ns_32_2_1_U26.top_add_32s_32ns_32_2_1_Adder_18_U.u2.cin ;
always @(posedge \add_38s_38s_38_2_1_U22.top_add_38s_38s_38_2_1_Adder_16_U.clk )
\add_38s_38s_38_2_1_U22.top_add_38s_38s_38_2_1_Adder_16_U.bin_s1  <= _0132_;
always @(posedge \add_38s_38s_38_2_1_U22.top_add_38s_38s_38_2_1_Adder_16_U.clk )
\add_38s_38s_38_2_1_U22.top_add_38s_38s_38_2_1_Adder_16_U.ain_s1  <= _0131_;
always @(posedge \add_38s_38s_38_2_1_U22.top_add_38s_38s_38_2_1_Adder_16_U.clk )
\add_38s_38s_38_2_1_U22.top_add_38s_38s_38_2_1_Adder_16_U.sum_s1  <= _0134_;
always @(posedge \add_38s_38s_38_2_1_U22.top_add_38s_38s_38_2_1_Adder_16_U.clk )
\add_38s_38s_38_2_1_U22.top_add_38s_38s_38_2_1_Adder_16_U.carry_s1  <= _0133_;
assign _0132_ = \add_38s_38s_38_2_1_U22.top_add_38s_38s_38_2_1_Adder_16_U.ce  ? \add_38s_38s_38_2_1_U22.top_add_38s_38s_38_2_1_Adder_16_U.b [37:19] : \add_38s_38s_38_2_1_U22.top_add_38s_38s_38_2_1_Adder_16_U.bin_s1 ;
assign _0131_ = \add_38s_38s_38_2_1_U22.top_add_38s_38s_38_2_1_Adder_16_U.ce  ? \add_38s_38s_38_2_1_U22.top_add_38s_38s_38_2_1_Adder_16_U.a [37:19] : \add_38s_38s_38_2_1_U22.top_add_38s_38s_38_2_1_Adder_16_U.ain_s1 ;
assign _0133_ = \add_38s_38s_38_2_1_U22.top_add_38s_38s_38_2_1_Adder_16_U.ce  ? \add_38s_38s_38_2_1_U22.top_add_38s_38s_38_2_1_Adder_16_U.facout_s1  : \add_38s_38s_38_2_1_U22.top_add_38s_38s_38_2_1_Adder_16_U.carry_s1 ;
assign _0134_ = \add_38s_38s_38_2_1_U22.top_add_38s_38s_38_2_1_Adder_16_U.ce  ? \add_38s_38s_38_2_1_U22.top_add_38s_38s_38_2_1_Adder_16_U.fas_s1  : \add_38s_38s_38_2_1_U22.top_add_38s_38s_38_2_1_Adder_16_U.sum_s1 ;
assign _0135_ = \add_38s_38s_38_2_1_U22.top_add_38s_38s_38_2_1_Adder_16_U.u1.a  + \add_38s_38s_38_2_1_U22.top_add_38s_38s_38_2_1_Adder_16_U.u1.b ;
assign { \add_38s_38s_38_2_1_U22.top_add_38s_38s_38_2_1_Adder_16_U.u1.cout , \add_38s_38s_38_2_1_U22.top_add_38s_38s_38_2_1_Adder_16_U.u1.s  } = _0135_ + \add_38s_38s_38_2_1_U22.top_add_38s_38s_38_2_1_Adder_16_U.u1.cin ;
assign _0136_ = \add_38s_38s_38_2_1_U22.top_add_38s_38s_38_2_1_Adder_16_U.u2.a  + \add_38s_38s_38_2_1_U22.top_add_38s_38s_38_2_1_Adder_16_U.u2.b ;
assign { \add_38s_38s_38_2_1_U22.top_add_38s_38s_38_2_1_Adder_16_U.u2.cout , \add_38s_38s_38_2_1_U22.top_add_38s_38s_38_2_1_Adder_16_U.u2.s  } = _0136_ + \add_38s_38s_38_2_1_U22.top_add_38s_38s_38_2_1_Adder_16_U.u2.cin ;
always @(posedge \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_9_U.clk )
\add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_9_U.bin_s1  <= _0138_;
always @(posedge \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_9_U.clk )
\add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_9_U.ain_s1  <= _0137_;
always @(posedge \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_9_U.clk )
\add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_9_U.sum_s1  <= _0140_;
always @(posedge \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_9_U.clk )
\add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_9_U.carry_s1  <= _0139_;
assign _0138_ = \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_9_U.ce  ? \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_9_U.b [2:1] : \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_9_U.bin_s1 ;
assign _0137_ = \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_9_U.ce  ? \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_9_U.a [2:1] : \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_9_U.ain_s1 ;
assign _0139_ = \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_9_U.ce  ? \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_9_U.facout_s1  : \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_9_U.carry_s1 ;
assign _0140_ = \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_9_U.ce  ? \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_9_U.fas_s1  : \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_9_U.sum_s1 ;
assign _0141_ = \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_9_U.u1.a  + \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_9_U.u1.b ;
assign { \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_9_U.u1.cout , \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_9_U.u1.s  } = _0141_ + \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_9_U.u1.cin ;
assign _0142_ = \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_9_U.u2.a  + \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_9_U.u2.b ;
assign { \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_9_U.u2.cout , \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_9_U.u2.s  } = _0142_ + \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_9_U.u2.cin ;
always @(posedge \add_3s_3s_3_2_1_U6.top_add_3s_3s_3_2_1_Adder_2_U.clk )
\add_3s_3s_3_2_1_U6.top_add_3s_3s_3_2_1_Adder_2_U.bin_s1  <= _0144_;
always @(posedge \add_3s_3s_3_2_1_U6.top_add_3s_3s_3_2_1_Adder_2_U.clk )
\add_3s_3s_3_2_1_U6.top_add_3s_3s_3_2_1_Adder_2_U.ain_s1  <= _0143_;
always @(posedge \add_3s_3s_3_2_1_U6.top_add_3s_3s_3_2_1_Adder_2_U.clk )
\add_3s_3s_3_2_1_U6.top_add_3s_3s_3_2_1_Adder_2_U.sum_s1  <= _0146_;
always @(posedge \add_3s_3s_3_2_1_U6.top_add_3s_3s_3_2_1_Adder_2_U.clk )
\add_3s_3s_3_2_1_U6.top_add_3s_3s_3_2_1_Adder_2_U.carry_s1  <= _0145_;
assign _0144_ = \add_3s_3s_3_2_1_U6.top_add_3s_3s_3_2_1_Adder_2_U.ce  ? \add_3s_3s_3_2_1_U6.top_add_3s_3s_3_2_1_Adder_2_U.b [2:1] : \add_3s_3s_3_2_1_U6.top_add_3s_3s_3_2_1_Adder_2_U.bin_s1 ;
assign _0143_ = \add_3s_3s_3_2_1_U6.top_add_3s_3s_3_2_1_Adder_2_U.ce  ? \add_3s_3s_3_2_1_U6.top_add_3s_3s_3_2_1_Adder_2_U.a [2:1] : \add_3s_3s_3_2_1_U6.top_add_3s_3s_3_2_1_Adder_2_U.ain_s1 ;
assign _0145_ = \add_3s_3s_3_2_1_U6.top_add_3s_3s_3_2_1_Adder_2_U.ce  ? \add_3s_3s_3_2_1_U6.top_add_3s_3s_3_2_1_Adder_2_U.facout_s1  : \add_3s_3s_3_2_1_U6.top_add_3s_3s_3_2_1_Adder_2_U.carry_s1 ;
assign _0146_ = \add_3s_3s_3_2_1_U6.top_add_3s_3s_3_2_1_Adder_2_U.ce  ? \add_3s_3s_3_2_1_U6.top_add_3s_3s_3_2_1_Adder_2_U.fas_s1  : \add_3s_3s_3_2_1_U6.top_add_3s_3s_3_2_1_Adder_2_U.sum_s1 ;
assign _0147_ = \add_3s_3s_3_2_1_U6.top_add_3s_3s_3_2_1_Adder_2_U.u1.a  + \add_3s_3s_3_2_1_U6.top_add_3s_3s_3_2_1_Adder_2_U.u1.b ;
assign { \add_3s_3s_3_2_1_U6.top_add_3s_3s_3_2_1_Adder_2_U.u1.cout , \add_3s_3s_3_2_1_U6.top_add_3s_3s_3_2_1_Adder_2_U.u1.s  } = _0147_ + \add_3s_3s_3_2_1_U6.top_add_3s_3s_3_2_1_Adder_2_U.u1.cin ;
assign _0148_ = \add_3s_3s_3_2_1_U6.top_add_3s_3s_3_2_1_Adder_2_U.u2.a  + \add_3s_3s_3_2_1_U6.top_add_3s_3s_3_2_1_Adder_2_U.u2.b ;
assign { \add_3s_3s_3_2_1_U6.top_add_3s_3s_3_2_1_Adder_2_U.u2.cout , \add_3s_3s_3_2_1_U6.top_add_3s_3s_3_2_1_Adder_2_U.u2.s  } = _0148_ + \add_3s_3s_3_2_1_U6.top_add_3s_3s_3_2_1_Adder_2_U.u2.cin ;
always @(posedge \add_40s_40s_40_2_1_U20.top_add_40s_40s_40_2_1_Adder_14_U.clk )
\add_40s_40s_40_2_1_U20.top_add_40s_40s_40_2_1_Adder_14_U.bin_s1  <= _0150_;
always @(posedge \add_40s_40s_40_2_1_U20.top_add_40s_40s_40_2_1_Adder_14_U.clk )
\add_40s_40s_40_2_1_U20.top_add_40s_40s_40_2_1_Adder_14_U.ain_s1  <= _0149_;
always @(posedge \add_40s_40s_40_2_1_U20.top_add_40s_40s_40_2_1_Adder_14_U.clk )
\add_40s_40s_40_2_1_U20.top_add_40s_40s_40_2_1_Adder_14_U.sum_s1  <= _0152_;
always @(posedge \add_40s_40s_40_2_1_U20.top_add_40s_40s_40_2_1_Adder_14_U.clk )
\add_40s_40s_40_2_1_U20.top_add_40s_40s_40_2_1_Adder_14_U.carry_s1  <= _0151_;
assign _0150_ = \add_40s_40s_40_2_1_U20.top_add_40s_40s_40_2_1_Adder_14_U.ce  ? \add_40s_40s_40_2_1_U20.top_add_40s_40s_40_2_1_Adder_14_U.b [39:20] : \add_40s_40s_40_2_1_U20.top_add_40s_40s_40_2_1_Adder_14_U.bin_s1 ;
assign _0149_ = \add_40s_40s_40_2_1_U20.top_add_40s_40s_40_2_1_Adder_14_U.ce  ? \add_40s_40s_40_2_1_U20.top_add_40s_40s_40_2_1_Adder_14_U.a [39:20] : \add_40s_40s_40_2_1_U20.top_add_40s_40s_40_2_1_Adder_14_U.ain_s1 ;
assign _0151_ = \add_40s_40s_40_2_1_U20.top_add_40s_40s_40_2_1_Adder_14_U.ce  ? \add_40s_40s_40_2_1_U20.top_add_40s_40s_40_2_1_Adder_14_U.facout_s1  : \add_40s_40s_40_2_1_U20.top_add_40s_40s_40_2_1_Adder_14_U.carry_s1 ;
assign _0152_ = \add_40s_40s_40_2_1_U20.top_add_40s_40s_40_2_1_Adder_14_U.ce  ? \add_40s_40s_40_2_1_U20.top_add_40s_40s_40_2_1_Adder_14_U.fas_s1  : \add_40s_40s_40_2_1_U20.top_add_40s_40s_40_2_1_Adder_14_U.sum_s1 ;
assign _0153_ = \add_40s_40s_40_2_1_U20.top_add_40s_40s_40_2_1_Adder_14_U.u1.a  + \add_40s_40s_40_2_1_U20.top_add_40s_40s_40_2_1_Adder_14_U.u1.b ;
assign { \add_40s_40s_40_2_1_U20.top_add_40s_40s_40_2_1_Adder_14_U.u1.cout , \add_40s_40s_40_2_1_U20.top_add_40s_40s_40_2_1_Adder_14_U.u1.s  } = _0153_ + \add_40s_40s_40_2_1_U20.top_add_40s_40s_40_2_1_Adder_14_U.u1.cin ;
assign _0154_ = \add_40s_40s_40_2_1_U20.top_add_40s_40s_40_2_1_Adder_14_U.u2.a  + \add_40s_40s_40_2_1_U20.top_add_40s_40s_40_2_1_Adder_14_U.u2.b ;
assign { \add_40s_40s_40_2_1_U20.top_add_40s_40s_40_2_1_Adder_14_U.u2.cout , \add_40s_40s_40_2_1_U20.top_add_40s_40s_40_2_1_Adder_14_U.u2.s  } = _0154_ + \add_40s_40s_40_2_1_U20.top_add_40s_40s_40_2_1_Adder_14_U.u2.cin ;
always @(posedge \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_7_U.clk )
\add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_7_U.bin_s1  <= _0156_;
always @(posedge \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_7_U.clk )
\add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_7_U.ain_s1  <= _0155_;
always @(posedge \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_7_U.clk )
\add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_7_U.sum_s1  <= _0158_;
always @(posedge \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_7_U.clk )
\add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_7_U.carry_s1  <= _0157_;
assign _0156_ = \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_7_U.ce  ? \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_7_U.b [3:2] : \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_7_U.bin_s1 ;
assign _0155_ = \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_7_U.ce  ? \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_7_U.a [3:2] : \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_7_U.ain_s1 ;
assign _0157_ = \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_7_U.ce  ? \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_7_U.facout_s1  : \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_7_U.carry_s1 ;
assign _0158_ = \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_7_U.ce  ? \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_7_U.fas_s1  : \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_7_U.sum_s1 ;
assign _0159_ = \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_7_U.u1.a  + \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_7_U.u1.b ;
assign { \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_7_U.u1.cout , \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_7_U.u1.s  } = _0159_ + \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_7_U.u1.cin ;
assign _0160_ = \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_7_U.u2.a  + \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_7_U.u2.b ;
assign { \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_7_U.u2.cout , \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_7_U.u2.s  } = _0160_ + \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_7_U.u2.cin ;
always @(posedge \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_3_U.clk )
\add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_3_U.bin_s1  <= _0162_;
always @(posedge \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_3_U.clk )
\add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_3_U.ain_s1  <= _0161_;
always @(posedge \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_3_U.clk )
\add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_3_U.sum_s1  <= _0164_;
always @(posedge \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_3_U.clk )
\add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_3_U.carry_s1  <= _0163_;
assign _0162_ = \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_3_U.ce  ? \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_3_U.b [4:2] : \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_3_U.bin_s1 ;
assign _0161_ = \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_3_U.ce  ? \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_3_U.a [4:2] : \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_3_U.ain_s1 ;
assign _0163_ = \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_3_U.ce  ? \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_3_U.facout_s1  : \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_3_U.carry_s1 ;
assign _0164_ = \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_3_U.ce  ? \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_3_U.fas_s1  : \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_3_U.sum_s1 ;
assign _0165_ = \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_3_U.u1.a  + \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_3_U.u1.b ;
assign { \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_3_U.u1.cout , \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_3_U.u1.s  } = _0165_ + \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_3_U.u1.cin ;
assign _0166_ = \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_3_U.u2.a  + \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_3_U.u2.b ;
assign { \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_3_U.u2.cout , \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_3_U.u2.s  } = _0166_ + \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_3_U.u2.cin ;
always @(posedge \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_6_U.clk )
\add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_6_U.bin_s1  <= _0168_;
always @(posedge \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_6_U.clk )
\add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_6_U.ain_s1  <= _0167_;
always @(posedge \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_6_U.clk )
\add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_6_U.sum_s1  <= _0170_;
always @(posedge \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_6_U.clk )
\add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_6_U.carry_s1  <= _0169_;
assign _0168_ = \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_6_U.ce  ? \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_6_U.b [5:3] : \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_6_U.bin_s1 ;
assign _0167_ = \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_6_U.ce  ? \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_6_U.a [5:3] : \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_6_U.ain_s1 ;
assign _0169_ = \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_6_U.ce  ? \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_6_U.facout_s1  : \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_6_U.carry_s1 ;
assign _0170_ = \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_6_U.ce  ? \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_6_U.fas_s1  : \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_6_U.sum_s1 ;
assign _0171_ = \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_6_U.u1.a  + \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_6_U.u1.b ;
assign { \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_6_U.u1.cout , \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_6_U.u1.s  } = _0171_ + \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_6_U.u1.cin ;
assign _0172_ = \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_6_U.u2.a  + \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_6_U.u2.b ;
assign { \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_6_U.u2.cout , \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_6_U.u2.s  } = _0172_ + \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_6_U.u2.cin ;
always @(posedge \add_7ns_7ns_7_2_1_U16.top_add_7ns_7ns_7_2_1_Adder_10_U.clk )
\add_7ns_7ns_7_2_1_U16.top_add_7ns_7ns_7_2_1_Adder_10_U.bin_s1  <= _0174_;
always @(posedge \add_7ns_7ns_7_2_1_U16.top_add_7ns_7ns_7_2_1_Adder_10_U.clk )
\add_7ns_7ns_7_2_1_U16.top_add_7ns_7ns_7_2_1_Adder_10_U.ain_s1  <= _0173_;
always @(posedge \add_7ns_7ns_7_2_1_U16.top_add_7ns_7ns_7_2_1_Adder_10_U.clk )
\add_7ns_7ns_7_2_1_U16.top_add_7ns_7ns_7_2_1_Adder_10_U.sum_s1  <= _0176_;
always @(posedge \add_7ns_7ns_7_2_1_U16.top_add_7ns_7ns_7_2_1_Adder_10_U.clk )
\add_7ns_7ns_7_2_1_U16.top_add_7ns_7ns_7_2_1_Adder_10_U.carry_s1  <= _0175_;
assign _0174_ = \add_7ns_7ns_7_2_1_U16.top_add_7ns_7ns_7_2_1_Adder_10_U.ce  ? \add_7ns_7ns_7_2_1_U16.top_add_7ns_7ns_7_2_1_Adder_10_U.b [6:3] : \add_7ns_7ns_7_2_1_U16.top_add_7ns_7ns_7_2_1_Adder_10_U.bin_s1 ;
assign _0173_ = \add_7ns_7ns_7_2_1_U16.top_add_7ns_7ns_7_2_1_Adder_10_U.ce  ? \add_7ns_7ns_7_2_1_U16.top_add_7ns_7ns_7_2_1_Adder_10_U.a [6:3] : \add_7ns_7ns_7_2_1_U16.top_add_7ns_7ns_7_2_1_Adder_10_U.ain_s1 ;
assign _0175_ = \add_7ns_7ns_7_2_1_U16.top_add_7ns_7ns_7_2_1_Adder_10_U.ce  ? \add_7ns_7ns_7_2_1_U16.top_add_7ns_7ns_7_2_1_Adder_10_U.facout_s1  : \add_7ns_7ns_7_2_1_U16.top_add_7ns_7ns_7_2_1_Adder_10_U.carry_s1 ;
assign _0176_ = \add_7ns_7ns_7_2_1_U16.top_add_7ns_7ns_7_2_1_Adder_10_U.ce  ? \add_7ns_7ns_7_2_1_U16.top_add_7ns_7ns_7_2_1_Adder_10_U.fas_s1  : \add_7ns_7ns_7_2_1_U16.top_add_7ns_7ns_7_2_1_Adder_10_U.sum_s1 ;
assign _0177_ = \add_7ns_7ns_7_2_1_U16.top_add_7ns_7ns_7_2_1_Adder_10_U.u1.a  + \add_7ns_7ns_7_2_1_U16.top_add_7ns_7ns_7_2_1_Adder_10_U.u1.b ;
assign { \add_7ns_7ns_7_2_1_U16.top_add_7ns_7ns_7_2_1_Adder_10_U.u1.cout , \add_7ns_7ns_7_2_1_U16.top_add_7ns_7ns_7_2_1_Adder_10_U.u1.s  } = _0177_ + \add_7ns_7ns_7_2_1_U16.top_add_7ns_7ns_7_2_1_Adder_10_U.u1.cin ;
assign _0178_ = \add_7ns_7ns_7_2_1_U16.top_add_7ns_7ns_7_2_1_Adder_10_U.u2.a  + \add_7ns_7ns_7_2_1_U16.top_add_7ns_7ns_7_2_1_Adder_10_U.u2.b ;
assign { \add_7ns_7ns_7_2_1_U16.top_add_7ns_7ns_7_2_1_Adder_10_U.u2.cout , \add_7ns_7ns_7_2_1_U16.top_add_7ns_7ns_7_2_1_Adder_10_U.u2.s  } = _0178_ + \add_7ns_7ns_7_2_1_U16.top_add_7ns_7ns_7_2_1_Adder_10_U.u2.cin ;
always @(posedge \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_8_U.clk )
\add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_8_U.bin_s1  <= _0180_;
always @(posedge \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_8_U.clk )
\add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_8_U.ain_s1  <= _0179_;
always @(posedge \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_8_U.clk )
\add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_8_U.sum_s1  <= _0182_;
always @(posedge \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_8_U.clk )
\add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_8_U.carry_s1  <= _0181_;
assign _0180_ = \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_8_U.ce  ? \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_8_U.b [6:3] : \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_8_U.bin_s1 ;
assign _0179_ = \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_8_U.ce  ? \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_8_U.a [6:3] : \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_8_U.ain_s1 ;
assign _0181_ = \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_8_U.ce  ? \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_8_U.facout_s1  : \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_8_U.carry_s1 ;
assign _0182_ = \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_8_U.ce  ? \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_8_U.fas_s1  : \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_8_U.sum_s1 ;
assign _0183_ = \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_8_U.u1.a  + \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_8_U.u1.b ;
assign { \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_8_U.u1.cout , \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_8_U.u1.s  } = _0183_ + \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_8_U.u1.cin ;
assign _0184_ = \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_8_U.u2.a  + \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_8_U.u2.b ;
assign { \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_8_U.u2.cout , \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_8_U.u2.s  } = _0184_ + \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_8_U.u2.cin ;
always @(posedge \add_9ns_9s_9_2_1_U9.top_add_9ns_9s_9_2_1_Adder_5_U.clk )
\add_9ns_9s_9_2_1_U9.top_add_9ns_9s_9_2_1_Adder_5_U.bin_s1  <= _0186_;
always @(posedge \add_9ns_9s_9_2_1_U9.top_add_9ns_9s_9_2_1_Adder_5_U.clk )
\add_9ns_9s_9_2_1_U9.top_add_9ns_9s_9_2_1_Adder_5_U.ain_s1  <= _0185_;
always @(posedge \add_9ns_9s_9_2_1_U9.top_add_9ns_9s_9_2_1_Adder_5_U.clk )
\add_9ns_9s_9_2_1_U9.top_add_9ns_9s_9_2_1_Adder_5_U.sum_s1  <= _0188_;
always @(posedge \add_9ns_9s_9_2_1_U9.top_add_9ns_9s_9_2_1_Adder_5_U.clk )
\add_9ns_9s_9_2_1_U9.top_add_9ns_9s_9_2_1_Adder_5_U.carry_s1  <= _0187_;
assign _0186_ = \add_9ns_9s_9_2_1_U9.top_add_9ns_9s_9_2_1_Adder_5_U.ce  ? \add_9ns_9s_9_2_1_U9.top_add_9ns_9s_9_2_1_Adder_5_U.b [8:4] : \add_9ns_9s_9_2_1_U9.top_add_9ns_9s_9_2_1_Adder_5_U.bin_s1 ;
assign _0185_ = \add_9ns_9s_9_2_1_U9.top_add_9ns_9s_9_2_1_Adder_5_U.ce  ? \add_9ns_9s_9_2_1_U9.top_add_9ns_9s_9_2_1_Adder_5_U.a [8:4] : \add_9ns_9s_9_2_1_U9.top_add_9ns_9s_9_2_1_Adder_5_U.ain_s1 ;
assign _0187_ = \add_9ns_9s_9_2_1_U9.top_add_9ns_9s_9_2_1_Adder_5_U.ce  ? \add_9ns_9s_9_2_1_U9.top_add_9ns_9s_9_2_1_Adder_5_U.facout_s1  : \add_9ns_9s_9_2_1_U9.top_add_9ns_9s_9_2_1_Adder_5_U.carry_s1 ;
assign _0188_ = \add_9ns_9s_9_2_1_U9.top_add_9ns_9s_9_2_1_Adder_5_U.ce  ? \add_9ns_9s_9_2_1_U9.top_add_9ns_9s_9_2_1_Adder_5_U.fas_s1  : \add_9ns_9s_9_2_1_U9.top_add_9ns_9s_9_2_1_Adder_5_U.sum_s1 ;
assign _0189_ = \add_9ns_9s_9_2_1_U9.top_add_9ns_9s_9_2_1_Adder_5_U.u1.a  + \add_9ns_9s_9_2_1_U9.top_add_9ns_9s_9_2_1_Adder_5_U.u1.b ;
assign { \add_9ns_9s_9_2_1_U9.top_add_9ns_9s_9_2_1_Adder_5_U.u1.cout , \add_9ns_9s_9_2_1_U9.top_add_9ns_9s_9_2_1_Adder_5_U.u1.s  } = _0189_ + \add_9ns_9s_9_2_1_U9.top_add_9ns_9s_9_2_1_Adder_5_U.u1.cin ;
assign _0190_ = \add_9ns_9s_9_2_1_U9.top_add_9ns_9s_9_2_1_Adder_5_U.u2.a  + \add_9ns_9s_9_2_1_U9.top_add_9ns_9s_9_2_1_Adder_5_U.u2.b ;
assign { \add_9ns_9s_9_2_1_U9.top_add_9ns_9s_9_2_1_Adder_5_U.u2.cout , \add_9ns_9s_9_2_1_U9.top_add_9ns_9s_9_2_1_Adder_5_U.u2.s  } = _0190_ + \add_9ns_9s_9_2_1_U9.top_add_9ns_9s_9_2_1_Adder_5_U.u2.cin ;
always @(posedge \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_13_U.clk )
\add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_13_U.bin_s1  <= _0192_;
always @(posedge \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_13_U.clk )
\add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_13_U.ain_s1  <= _0191_;
always @(posedge \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_13_U.clk )
\add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_13_U.sum_s1  <= _0194_;
always @(posedge \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_13_U.clk )
\add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_13_U.carry_s1  <= _0193_;
assign _0192_ = \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_13_U.ce  ? \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_13_U.b [8:4] : \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_13_U.bin_s1 ;
assign _0191_ = \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_13_U.ce  ? \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_13_U.a [8:4] : \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_13_U.ain_s1 ;
assign _0193_ = \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_13_U.ce  ? \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_13_U.facout_s1  : \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_13_U.carry_s1 ;
assign _0194_ = \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_13_U.ce  ? \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_13_U.fas_s1  : \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_13_U.sum_s1 ;
assign _0195_ = \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_13_U.u1.a  + \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_13_U.u1.b ;
assign { \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_13_U.u1.cout , \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_13_U.u1.s  } = _0195_ + \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_13_U.u1.cin ;
assign _0196_ = \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_13_U.u2.a  + \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_13_U.u2.b ;
assign { \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_13_U.u2.cout , \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_13_U.u2.s  } = _0196_ + \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_13_U.u2.cin ;
always @(posedge \ashr_16s_4ns_16_7_1_U4.clk )
\ashr_16s_4ns_16_7_1_U4.dout_array[5]  <= _0208_;
always @(posedge \ashr_16s_4ns_16_7_1_U4.clk )
\ashr_16s_4ns_16_7_1_U4.din1_cast_array[5]  <= _0202_;
always @(posedge \ashr_16s_4ns_16_7_1_U4.clk )
\ashr_16s_4ns_16_7_1_U4.dout_array[4]  <= _0207_;
always @(posedge \ashr_16s_4ns_16_7_1_U4.clk )
\ashr_16s_4ns_16_7_1_U4.din1_cast_array[4]  <= _0201_;
always @(posedge \ashr_16s_4ns_16_7_1_U4.clk )
\ashr_16s_4ns_16_7_1_U4.dout_array[3]  <= _0206_;
always @(posedge \ashr_16s_4ns_16_7_1_U4.clk )
\ashr_16s_4ns_16_7_1_U4.din1_cast_array[3]  <= _0200_;
always @(posedge \ashr_16s_4ns_16_7_1_U4.clk )
\ashr_16s_4ns_16_7_1_U4.dout_array[2]  <= _0205_;
always @(posedge \ashr_16s_4ns_16_7_1_U4.clk )
\ashr_16s_4ns_16_7_1_U4.din1_cast_array[2]  <= _0199_;
always @(posedge \ashr_16s_4ns_16_7_1_U4.clk )
\ashr_16s_4ns_16_7_1_U4.dout_array[1]  <= _0204_;
always @(posedge \ashr_16s_4ns_16_7_1_U4.clk )
\ashr_16s_4ns_16_7_1_U4.din1_cast_array[1]  <= _0198_;
always @(posedge \ashr_16s_4ns_16_7_1_U4.clk )
\ashr_16s_4ns_16_7_1_U4.dout_array[0]  <= _0203_;
always @(posedge \ashr_16s_4ns_16_7_1_U4.clk )
\ashr_16s_4ns_16_7_1_U4.din1_cast_array[0]  <= _0197_;
assign _0209_ = \ashr_16s_4ns_16_7_1_U4.ce  ? \ashr_16s_4ns_16_7_1_U4.din1_cast_array[4]  : \ashr_16s_4ns_16_7_1_U4.din1_cast_array[5] ;
assign _0202_ = \ashr_16s_4ns_16_7_1_U4.reset  ? 4'h0 : _0209_;
assign _0210_ = \ashr_16s_4ns_16_7_1_U4.ce  ? _0223_ : \ashr_16s_4ns_16_7_1_U4.dout_array[5] ;
assign _0208_ = \ashr_16s_4ns_16_7_1_U4.reset  ? 16'h0000 : _0210_;
assign _0211_ = \ashr_16s_4ns_16_7_1_U4.ce  ? \ashr_16s_4ns_16_7_1_U4.din1_cast_array[3]  : \ashr_16s_4ns_16_7_1_U4.din1_cast_array[4] ;
assign _0201_ = \ashr_16s_4ns_16_7_1_U4.reset  ? 4'h0 : _0211_;
assign _0212_ = \ashr_16s_4ns_16_7_1_U4.ce  ? _0222_ : \ashr_16s_4ns_16_7_1_U4.dout_array[4] ;
assign _0207_ = \ashr_16s_4ns_16_7_1_U4.reset  ? 16'h0000 : _0212_;
assign _0213_ = \ashr_16s_4ns_16_7_1_U4.ce  ? \ashr_16s_4ns_16_7_1_U4.din1_cast_array[2]  : \ashr_16s_4ns_16_7_1_U4.din1_cast_array[3] ;
assign _0200_ = \ashr_16s_4ns_16_7_1_U4.reset  ? 4'h0 : _0213_;
assign _0214_ = \ashr_16s_4ns_16_7_1_U4.ce  ? _0221_ : \ashr_16s_4ns_16_7_1_U4.dout_array[3] ;
assign _0206_ = \ashr_16s_4ns_16_7_1_U4.reset  ? 16'h0000 : _0214_;
assign _0215_ = \ashr_16s_4ns_16_7_1_U4.ce  ? \ashr_16s_4ns_16_7_1_U4.din1_cast_array[1]  : \ashr_16s_4ns_16_7_1_U4.din1_cast_array[2] ;
assign _0199_ = \ashr_16s_4ns_16_7_1_U4.reset  ? 4'h0 : _0215_;
assign _0216_ = \ashr_16s_4ns_16_7_1_U4.ce  ? \ashr_16s_4ns_16_7_1_U4.dout_array[1]  : \ashr_16s_4ns_16_7_1_U4.dout_array[2] ;
assign _0205_ = \ashr_16s_4ns_16_7_1_U4.reset  ? 16'h0000 : _0216_;
assign _0217_ = \ashr_16s_4ns_16_7_1_U4.ce  ? \ashr_16s_4ns_16_7_1_U4.din1_cast_array[0]  : \ashr_16s_4ns_16_7_1_U4.din1_cast_array[1] ;
assign _0198_ = \ashr_16s_4ns_16_7_1_U4.reset  ? 4'h0 : _0217_;
assign _0218_ = \ashr_16s_4ns_16_7_1_U4.ce  ? \ashr_16s_4ns_16_7_1_U4.dout_array[0]  : \ashr_16s_4ns_16_7_1_U4.dout_array[1] ;
assign _0204_ = \ashr_16s_4ns_16_7_1_U4.reset  ? 16'h0000 : _0218_;
assign _0219_ = \ashr_16s_4ns_16_7_1_U4.ce  ? \ashr_16s_4ns_16_7_1_U4.din1 [3:0] : \ashr_16s_4ns_16_7_1_U4.din1_cast_array[0] ;
assign _0197_ = \ashr_16s_4ns_16_7_1_U4.reset  ? 4'h0 : _0219_;
assign _0220_ = \ashr_16s_4ns_16_7_1_U4.ce  ? \ashr_16s_4ns_16_7_1_U4.din0  : \ashr_16s_4ns_16_7_1_U4.dout_array[0] ;
assign _0203_ = \ashr_16s_4ns_16_7_1_U4.reset  ? 16'h0000 : _0220_;
assign _0221_ = $signed(\ashr_16s_4ns_16_7_1_U4.dout_array[2] ) >>> { \ashr_16s_4ns_16_7_1_U4.din1_cast_array[2] [3], 3'h0 };
assign _0222_ = $signed(\ashr_16s_4ns_16_7_1_U4.dout_array[3] ) >>> { \ashr_16s_4ns_16_7_1_U4.din1_cast_array[3] [2], 2'h0 };
assign _0223_ = $signed(\ashr_16s_4ns_16_7_1_U4.dout_array[4] ) >>> { \ashr_16s_4ns_16_7_1_U4.din1_cast_array[4] [1], 1'h0 };
assign \ashr_16s_4ns_16_7_1_U4.dout  = $signed(\ashr_16s_4ns_16_7_1_U4.dout_array[5] ) >>> \ashr_16s_4ns_16_7_1_U4.din1_cast_array[5] [0];
always @(posedge \ashr_8ns_8s_8_7_1_U11.clk )
\ashr_8ns_8s_8_7_1_U11.dout_array[5]  <= _0235_;
always @(posedge \ashr_8ns_8s_8_7_1_U11.clk )
\ashr_8ns_8s_8_7_1_U11.din1_cast_array[5]  <= _0229_;
always @(posedge \ashr_8ns_8s_8_7_1_U11.clk )
\ashr_8ns_8s_8_7_1_U11.dout_array[4]  <= _0234_;
always @(posedge \ashr_8ns_8s_8_7_1_U11.clk )
\ashr_8ns_8s_8_7_1_U11.din1_cast_array[4]  <= _0228_;
always @(posedge \ashr_8ns_8s_8_7_1_U11.clk )
\ashr_8ns_8s_8_7_1_U11.dout_array[3]  <= _0233_;
always @(posedge \ashr_8ns_8s_8_7_1_U11.clk )
\ashr_8ns_8s_8_7_1_U11.din1_cast_array[3]  <= _0227_;
always @(posedge \ashr_8ns_8s_8_7_1_U11.clk )
\ashr_8ns_8s_8_7_1_U11.dout_array[2]  <= _0232_;
always @(posedge \ashr_8ns_8s_8_7_1_U11.clk )
\ashr_8ns_8s_8_7_1_U11.din1_cast_array[2]  <= _0226_;
always @(posedge \ashr_8ns_8s_8_7_1_U11.clk )
\ashr_8ns_8s_8_7_1_U11.dout_array[1]  <= _0231_;
always @(posedge \ashr_8ns_8s_8_7_1_U11.clk )
\ashr_8ns_8s_8_7_1_U11.din1_cast_array[1]  <= _0225_;
always @(posedge \ashr_8ns_8s_8_7_1_U11.clk )
\ashr_8ns_8s_8_7_1_U11.dout_array[0]  <= _0230_;
always @(posedge \ashr_8ns_8s_8_7_1_U11.clk )
\ashr_8ns_8s_8_7_1_U11.din1_cast_array[0]  <= _0224_;
assign _0236_ = \ashr_8ns_8s_8_7_1_U11.ce  ? \ashr_8ns_8s_8_7_1_U11.din1_cast_array[4]  : \ashr_8ns_8s_8_7_1_U11.din1_cast_array[5] ;
assign _0229_ = \ashr_8ns_8s_8_7_1_U11.reset  ? 8'h00 : _0236_;
assign _0237_ = \ashr_8ns_8s_8_7_1_U11.ce  ? _0250_ : \ashr_8ns_8s_8_7_1_U11.dout_array[5] ;
assign _0235_ = \ashr_8ns_8s_8_7_1_U11.reset  ? 8'h00 : _0237_;
assign _0238_ = \ashr_8ns_8s_8_7_1_U11.ce  ? \ashr_8ns_8s_8_7_1_U11.din1_cast_array[3]  : \ashr_8ns_8s_8_7_1_U11.din1_cast_array[4] ;
assign _0228_ = \ashr_8ns_8s_8_7_1_U11.reset  ? 8'h00 : _0238_;
assign _0239_ = \ashr_8ns_8s_8_7_1_U11.ce  ? _0249_ : \ashr_8ns_8s_8_7_1_U11.dout_array[4] ;
assign _0234_ = \ashr_8ns_8s_8_7_1_U11.reset  ? 8'h00 : _0239_;
assign _0240_ = \ashr_8ns_8s_8_7_1_U11.ce  ? \ashr_8ns_8s_8_7_1_U11.din1_cast_array[2]  : \ashr_8ns_8s_8_7_1_U11.din1_cast_array[3] ;
assign _0227_ = \ashr_8ns_8s_8_7_1_U11.reset  ? 8'h00 : _0240_;
assign _0241_ = \ashr_8ns_8s_8_7_1_U11.ce  ? _0248_ : \ashr_8ns_8s_8_7_1_U11.dout_array[3] ;
assign _0233_ = \ashr_8ns_8s_8_7_1_U11.reset  ? 8'h00 : _0241_;
assign _0242_ = \ashr_8ns_8s_8_7_1_U11.ce  ? \ashr_8ns_8s_8_7_1_U11.din1_cast_array[1]  : \ashr_8ns_8s_8_7_1_U11.din1_cast_array[2] ;
assign _0226_ = \ashr_8ns_8s_8_7_1_U11.reset  ? 8'h00 : _0242_;
assign _0243_ = \ashr_8ns_8s_8_7_1_U11.ce  ? \ashr_8ns_8s_8_7_1_U11.dout_array[1]  : \ashr_8ns_8s_8_7_1_U11.dout_array[2] ;
assign _0232_ = \ashr_8ns_8s_8_7_1_U11.reset  ? 8'h00 : _0243_;
assign _0244_ = \ashr_8ns_8s_8_7_1_U11.ce  ? \ashr_8ns_8s_8_7_1_U11.din1_cast_array[0]  : \ashr_8ns_8s_8_7_1_U11.din1_cast_array[1] ;
assign _0225_ = \ashr_8ns_8s_8_7_1_U11.reset  ? 8'h00 : _0244_;
assign _0245_ = \ashr_8ns_8s_8_7_1_U11.ce  ? \ashr_8ns_8s_8_7_1_U11.dout_array[0]  : \ashr_8ns_8s_8_7_1_U11.dout_array[1] ;
assign _0231_ = \ashr_8ns_8s_8_7_1_U11.reset  ? 8'h00 : _0245_;
assign _0246_ = \ashr_8ns_8s_8_7_1_U11.ce  ? \ashr_8ns_8s_8_7_1_U11.din1  : \ashr_8ns_8s_8_7_1_U11.din1_cast_array[0] ;
assign _0224_ = \ashr_8ns_8s_8_7_1_U11.reset  ? 8'h00 : _0246_;
assign _0247_ = \ashr_8ns_8s_8_7_1_U11.ce  ? \ashr_8ns_8s_8_7_1_U11.din0  : \ashr_8ns_8s_8_7_1_U11.dout_array[0] ;
assign _0230_ = \ashr_8ns_8s_8_7_1_U11.reset  ? 8'h00 : _0247_;
assign _0248_ = $signed(\ashr_8ns_8s_8_7_1_U11.dout_array[2] ) >>> { \ashr_8ns_8s_8_7_1_U11.din1_cast_array[2] [7:6], 6'h00 };
assign _0249_ = $signed(\ashr_8ns_8s_8_7_1_U11.dout_array[3] ) >>> { \ashr_8ns_8s_8_7_1_U11.din1_cast_array[3] [5:4], 4'h0 };
assign _0250_ = $signed(\ashr_8ns_8s_8_7_1_U11.dout_array[4] ) >>> { \ashr_8ns_8s_8_7_1_U11.din1_cast_array[4] [3:2], 2'h0 };
assign \ashr_8ns_8s_8_7_1_U11.dout  = $signed(\ashr_8ns_8s_8_7_1_U11.dout_array[5] ) >>> \ashr_8ns_8s_8_7_1_U11.din1_cast_array[5] [1:0];
assign \mul_16s_2s_18_7_1_U5.top_mul_16s_2s_18_7_1_Mul_DSP_0_U.tmp_product  = $signed(\mul_16s_2s_18_7_1_U5.top_mul_16s_2s_18_7_1_Mul_DSP_0_U.a_reg0 ) * $signed(\mul_16s_2s_18_7_1_U5.top_mul_16s_2s_18_7_1_Mul_DSP_0_U.b_reg0 );
always @(posedge \mul_16s_2s_18_7_1_U5.top_mul_16s_2s_18_7_1_Mul_DSP_0_U.clk )
\mul_16s_2s_18_7_1_U5.top_mul_16s_2s_18_7_1_Mul_DSP_0_U.a_reg0  <= _0251_;
always @(posedge \mul_16s_2s_18_7_1_U5.top_mul_16s_2s_18_7_1_Mul_DSP_0_U.clk )
\mul_16s_2s_18_7_1_U5.top_mul_16s_2s_18_7_1_Mul_DSP_0_U.b_reg0  <= _0252_;
always @(posedge \mul_16s_2s_18_7_1_U5.top_mul_16s_2s_18_7_1_Mul_DSP_0_U.clk )
\mul_16s_2s_18_7_1_U5.top_mul_16s_2s_18_7_1_Mul_DSP_0_U.buff0  <= _0253_;
always @(posedge \mul_16s_2s_18_7_1_U5.top_mul_16s_2s_18_7_1_Mul_DSP_0_U.clk )
\mul_16s_2s_18_7_1_U5.top_mul_16s_2s_18_7_1_Mul_DSP_0_U.buff1  <= _0254_;
always @(posedge \mul_16s_2s_18_7_1_U5.top_mul_16s_2s_18_7_1_Mul_DSP_0_U.clk )
\mul_16s_2s_18_7_1_U5.top_mul_16s_2s_18_7_1_Mul_DSP_0_U.buff2  <= _0255_;
always @(posedge \mul_16s_2s_18_7_1_U5.top_mul_16s_2s_18_7_1_Mul_DSP_0_U.clk )
\mul_16s_2s_18_7_1_U5.top_mul_16s_2s_18_7_1_Mul_DSP_0_U.buff3  <= _0256_;
always @(posedge \mul_16s_2s_18_7_1_U5.top_mul_16s_2s_18_7_1_Mul_DSP_0_U.clk )
\mul_16s_2s_18_7_1_U5.top_mul_16s_2s_18_7_1_Mul_DSP_0_U.buff4  <= _0257_;
assign _0257_ = \mul_16s_2s_18_7_1_U5.top_mul_16s_2s_18_7_1_Mul_DSP_0_U.ce  ? \mul_16s_2s_18_7_1_U5.top_mul_16s_2s_18_7_1_Mul_DSP_0_U.buff3  : \mul_16s_2s_18_7_1_U5.top_mul_16s_2s_18_7_1_Mul_DSP_0_U.buff4 ;
assign _0256_ = \mul_16s_2s_18_7_1_U5.top_mul_16s_2s_18_7_1_Mul_DSP_0_U.ce  ? \mul_16s_2s_18_7_1_U5.top_mul_16s_2s_18_7_1_Mul_DSP_0_U.buff2  : \mul_16s_2s_18_7_1_U5.top_mul_16s_2s_18_7_1_Mul_DSP_0_U.buff3 ;
assign _0255_ = \mul_16s_2s_18_7_1_U5.top_mul_16s_2s_18_7_1_Mul_DSP_0_U.ce  ? \mul_16s_2s_18_7_1_U5.top_mul_16s_2s_18_7_1_Mul_DSP_0_U.buff1  : \mul_16s_2s_18_7_1_U5.top_mul_16s_2s_18_7_1_Mul_DSP_0_U.buff2 ;
assign _0254_ = \mul_16s_2s_18_7_1_U5.top_mul_16s_2s_18_7_1_Mul_DSP_0_U.ce  ? \mul_16s_2s_18_7_1_U5.top_mul_16s_2s_18_7_1_Mul_DSP_0_U.buff0  : \mul_16s_2s_18_7_1_U5.top_mul_16s_2s_18_7_1_Mul_DSP_0_U.buff1 ;
assign _0253_ = \mul_16s_2s_18_7_1_U5.top_mul_16s_2s_18_7_1_Mul_DSP_0_U.ce  ? \mul_16s_2s_18_7_1_U5.top_mul_16s_2s_18_7_1_Mul_DSP_0_U.tmp_product  : \mul_16s_2s_18_7_1_U5.top_mul_16s_2s_18_7_1_Mul_DSP_0_U.buff0 ;
assign _0252_ = \mul_16s_2s_18_7_1_U5.top_mul_16s_2s_18_7_1_Mul_DSP_0_U.ce  ? \mul_16s_2s_18_7_1_U5.top_mul_16s_2s_18_7_1_Mul_DSP_0_U.b  : \mul_16s_2s_18_7_1_U5.top_mul_16s_2s_18_7_1_Mul_DSP_0_U.b_reg0 ;
assign _0251_ = \mul_16s_2s_18_7_1_U5.top_mul_16s_2s_18_7_1_Mul_DSP_0_U.ce  ? \mul_16s_2s_18_7_1_U5.top_mul_16s_2s_18_7_1_Mul_DSP_0_U.a  : \mul_16s_2s_18_7_1_U5.top_mul_16s_2s_18_7_1_Mul_DSP_0_U.a_reg0 ;
always @(posedge \shl_16s_4ns_16_7_1_U3.clk )
\shl_16s_4ns_16_7_1_U3.dout_array[5]  <= _0269_;
always @(posedge \shl_16s_4ns_16_7_1_U3.clk )
\shl_16s_4ns_16_7_1_U3.din1_cast_array[5]  <= _0263_;
always @(posedge \shl_16s_4ns_16_7_1_U3.clk )
\shl_16s_4ns_16_7_1_U3.dout_array[4]  <= _0268_;
always @(posedge \shl_16s_4ns_16_7_1_U3.clk )
\shl_16s_4ns_16_7_1_U3.din1_cast_array[4]  <= _0262_;
always @(posedge \shl_16s_4ns_16_7_1_U3.clk )
\shl_16s_4ns_16_7_1_U3.dout_array[3]  <= _0267_;
always @(posedge \shl_16s_4ns_16_7_1_U3.clk )
\shl_16s_4ns_16_7_1_U3.din1_cast_array[3]  <= _0261_;
always @(posedge \shl_16s_4ns_16_7_1_U3.clk )
\shl_16s_4ns_16_7_1_U3.dout_array[2]  <= _0266_;
always @(posedge \shl_16s_4ns_16_7_1_U3.clk )
\shl_16s_4ns_16_7_1_U3.din1_cast_array[2]  <= _0260_;
always @(posedge \shl_16s_4ns_16_7_1_U3.clk )
\shl_16s_4ns_16_7_1_U3.dout_array[1]  <= _0265_;
always @(posedge \shl_16s_4ns_16_7_1_U3.clk )
\shl_16s_4ns_16_7_1_U3.din1_cast_array[1]  <= _0259_;
always @(posedge \shl_16s_4ns_16_7_1_U3.clk )
\shl_16s_4ns_16_7_1_U3.dout_array[0]  <= _0264_;
always @(posedge \shl_16s_4ns_16_7_1_U3.clk )
\shl_16s_4ns_16_7_1_U3.din1_cast_array[0]  <= _0258_;
assign _0270_ = \shl_16s_4ns_16_7_1_U3.ce  ? \shl_16s_4ns_16_7_1_U3.din1_cast_array[4]  : \shl_16s_4ns_16_7_1_U3.din1_cast_array[5] ;
assign _0263_ = \shl_16s_4ns_16_7_1_U3.reset  ? 4'h0 : _0270_;
assign _0271_ = \shl_16s_4ns_16_7_1_U3.ce  ? _0284_ : \shl_16s_4ns_16_7_1_U3.dout_array[5] ;
assign _0269_ = \shl_16s_4ns_16_7_1_U3.reset  ? 16'h0000 : _0271_;
assign _0272_ = \shl_16s_4ns_16_7_1_U3.ce  ? \shl_16s_4ns_16_7_1_U3.din1_cast_array[3]  : \shl_16s_4ns_16_7_1_U3.din1_cast_array[4] ;
assign _0262_ = \shl_16s_4ns_16_7_1_U3.reset  ? 4'h0 : _0272_;
assign _0273_ = \shl_16s_4ns_16_7_1_U3.ce  ? _0283_ : \shl_16s_4ns_16_7_1_U3.dout_array[4] ;
assign _0268_ = \shl_16s_4ns_16_7_1_U3.reset  ? 16'h0000 : _0273_;
assign _0274_ = \shl_16s_4ns_16_7_1_U3.ce  ? \shl_16s_4ns_16_7_1_U3.din1_cast_array[2]  : \shl_16s_4ns_16_7_1_U3.din1_cast_array[3] ;
assign _0261_ = \shl_16s_4ns_16_7_1_U3.reset  ? 4'h0 : _0274_;
assign _0275_ = \shl_16s_4ns_16_7_1_U3.ce  ? _0282_ : \shl_16s_4ns_16_7_1_U3.dout_array[3] ;
assign _0267_ = \shl_16s_4ns_16_7_1_U3.reset  ? 16'h0000 : _0275_;
assign _0276_ = \shl_16s_4ns_16_7_1_U3.ce  ? \shl_16s_4ns_16_7_1_U3.din1_cast_array[1]  : \shl_16s_4ns_16_7_1_U3.din1_cast_array[2] ;
assign _0260_ = \shl_16s_4ns_16_7_1_U3.reset  ? 4'h0 : _0276_;
assign _0277_ = \shl_16s_4ns_16_7_1_U3.ce  ? \shl_16s_4ns_16_7_1_U3.dout_array[1]  : \shl_16s_4ns_16_7_1_U3.dout_array[2] ;
assign _0266_ = \shl_16s_4ns_16_7_1_U3.reset  ? 16'h0000 : _0277_;
assign _0278_ = \shl_16s_4ns_16_7_1_U3.ce  ? \shl_16s_4ns_16_7_1_U3.din1_cast_array[0]  : \shl_16s_4ns_16_7_1_U3.din1_cast_array[1] ;
assign _0259_ = \shl_16s_4ns_16_7_1_U3.reset  ? 4'h0 : _0278_;
assign _0279_ = \shl_16s_4ns_16_7_1_U3.ce  ? \shl_16s_4ns_16_7_1_U3.dout_array[0]  : \shl_16s_4ns_16_7_1_U3.dout_array[1] ;
assign _0265_ = \shl_16s_4ns_16_7_1_U3.reset  ? 16'h0000 : _0279_;
assign _0280_ = \shl_16s_4ns_16_7_1_U3.ce  ? \shl_16s_4ns_16_7_1_U3.din1 [3:0] : \shl_16s_4ns_16_7_1_U3.din1_cast_array[0] ;
assign _0258_ = \shl_16s_4ns_16_7_1_U3.reset  ? 4'h0 : _0280_;
assign _0281_ = \shl_16s_4ns_16_7_1_U3.ce  ? \shl_16s_4ns_16_7_1_U3.din0  : \shl_16s_4ns_16_7_1_U3.dout_array[0] ;
assign _0264_ = \shl_16s_4ns_16_7_1_U3.reset  ? 16'h0000 : _0281_;
assign _0282_ = \shl_16s_4ns_16_7_1_U3.dout_array[2]  << { \shl_16s_4ns_16_7_1_U3.din1_cast_array[2] [3], 3'h0 };
assign _0283_ = \shl_16s_4ns_16_7_1_U3.dout_array[3]  << { \shl_16s_4ns_16_7_1_U3.din1_cast_array[3] [2], 2'h0 };
assign _0284_ = \shl_16s_4ns_16_7_1_U3.dout_array[4]  << { \shl_16s_4ns_16_7_1_U3.din1_cast_array[4] [1], 1'h0 };
assign \shl_16s_4ns_16_7_1_U3.dout  = \shl_16s_4ns_16_7_1_U3.dout_array[5]  << \shl_16s_4ns_16_7_1_U3.din1_cast_array[5] [0];
always @(posedge \shl_8ns_8s_8_7_1_U10.clk )
\shl_8ns_8s_8_7_1_U10.dout_array[5]  <= _0296_;
always @(posedge \shl_8ns_8s_8_7_1_U10.clk )
\shl_8ns_8s_8_7_1_U10.din1_cast_array[5]  <= _0290_;
always @(posedge \shl_8ns_8s_8_7_1_U10.clk )
\shl_8ns_8s_8_7_1_U10.dout_array[4]  <= _0295_;
always @(posedge \shl_8ns_8s_8_7_1_U10.clk )
\shl_8ns_8s_8_7_1_U10.din1_cast_array[4]  <= _0289_;
always @(posedge \shl_8ns_8s_8_7_1_U10.clk )
\shl_8ns_8s_8_7_1_U10.dout_array[3]  <= _0294_;
always @(posedge \shl_8ns_8s_8_7_1_U10.clk )
\shl_8ns_8s_8_7_1_U10.din1_cast_array[3]  <= _0288_;
always @(posedge \shl_8ns_8s_8_7_1_U10.clk )
\shl_8ns_8s_8_7_1_U10.dout_array[2]  <= _0293_;
always @(posedge \shl_8ns_8s_8_7_1_U10.clk )
\shl_8ns_8s_8_7_1_U10.din1_cast_array[2]  <= _0287_;
always @(posedge \shl_8ns_8s_8_7_1_U10.clk )
\shl_8ns_8s_8_7_1_U10.dout_array[1]  <= _0292_;
always @(posedge \shl_8ns_8s_8_7_1_U10.clk )
\shl_8ns_8s_8_7_1_U10.din1_cast_array[1]  <= _0286_;
always @(posedge \shl_8ns_8s_8_7_1_U10.clk )
\shl_8ns_8s_8_7_1_U10.dout_array[0]  <= _0291_;
always @(posedge \shl_8ns_8s_8_7_1_U10.clk )
\shl_8ns_8s_8_7_1_U10.din1_cast_array[0]  <= _0285_;
assign _0286_ = \shl_8ns_8s_8_7_1_U10.reset  ? 8'h00 : _0308_;
assign _0297_ = \shl_8ns_8s_8_7_1_U10.ce  ? \shl_8ns_8s_8_7_1_U10.dout_array[0]  : \shl_8ns_8s_8_7_1_U10.dout_array[1] ;
assign _0292_ = \shl_8ns_8s_8_7_1_U10.reset  ? 8'h00 : _0297_;
assign _0298_ = \shl_8ns_8s_8_7_1_U10.ce  ? \shl_8ns_8s_8_7_1_U10.din1  : \shl_8ns_8s_8_7_1_U10.din1_cast_array[0] ;
assign _0285_ = \shl_8ns_8s_8_7_1_U10.reset  ? 8'h00 : _0298_;
assign _0299_ = \shl_8ns_8s_8_7_1_U10.ce  ? \shl_8ns_8s_8_7_1_U10.din0  : \shl_8ns_8s_8_7_1_U10.dout_array[0] ;
assign _0291_ = \shl_8ns_8s_8_7_1_U10.reset  ? 8'h00 : _0299_;
assign _0300_ = \shl_8ns_8s_8_7_1_U10.ce  ? \shl_8ns_8s_8_7_1_U10.din1_cast_array[4]  : \shl_8ns_8s_8_7_1_U10.din1_cast_array[5] ;
assign _0290_ = \shl_8ns_8s_8_7_1_U10.reset  ? 8'h00 : _0300_;
assign _0301_ = \shl_8ns_8s_8_7_1_U10.ce  ? _0311_ : \shl_8ns_8s_8_7_1_U10.dout_array[5] ;
assign _0296_ = \shl_8ns_8s_8_7_1_U10.reset  ? 8'h00 : _0301_;
assign _0302_ = \shl_8ns_8s_8_7_1_U10.ce  ? \shl_8ns_8s_8_7_1_U10.din1_cast_array[3]  : \shl_8ns_8s_8_7_1_U10.din1_cast_array[4] ;
assign _0289_ = \shl_8ns_8s_8_7_1_U10.reset  ? 8'h00 : _0302_;
assign _0303_ = \shl_8ns_8s_8_7_1_U10.ce  ? _0310_ : \shl_8ns_8s_8_7_1_U10.dout_array[4] ;
assign _0295_ = \shl_8ns_8s_8_7_1_U10.reset  ? 8'h00 : _0303_;
assign _0304_ = \shl_8ns_8s_8_7_1_U10.ce  ? \shl_8ns_8s_8_7_1_U10.din1_cast_array[2]  : \shl_8ns_8s_8_7_1_U10.din1_cast_array[3] ;
assign _0288_ = \shl_8ns_8s_8_7_1_U10.reset  ? 8'h00 : _0304_;
assign _0305_ = \shl_8ns_8s_8_7_1_U10.ce  ? _0309_ : \shl_8ns_8s_8_7_1_U10.dout_array[3] ;
assign _0294_ = \shl_8ns_8s_8_7_1_U10.reset  ? 8'h00 : _0305_;
assign _0306_ = \shl_8ns_8s_8_7_1_U10.ce  ? \shl_8ns_8s_8_7_1_U10.din1_cast_array[1]  : \shl_8ns_8s_8_7_1_U10.din1_cast_array[2] ;
assign _0287_ = \shl_8ns_8s_8_7_1_U10.reset  ? 8'h00 : _0306_;
assign _0307_ = \shl_8ns_8s_8_7_1_U10.ce  ? \shl_8ns_8s_8_7_1_U10.dout_array[1]  : \shl_8ns_8s_8_7_1_U10.dout_array[2] ;
assign _0293_ = \shl_8ns_8s_8_7_1_U10.reset  ? 8'h00 : _0307_;
assign _0308_ = \shl_8ns_8s_8_7_1_U10.ce  ? \shl_8ns_8s_8_7_1_U10.din1_cast_array[0]  : \shl_8ns_8s_8_7_1_U10.din1_cast_array[1] ;
assign _0309_ = \shl_8ns_8s_8_7_1_U10.dout_array[2]  << { \shl_8ns_8s_8_7_1_U10.din1_cast_array[2] [7:6], 6'h00 };
assign _0310_ = \shl_8ns_8s_8_7_1_U10.dout_array[3]  << { \shl_8ns_8s_8_7_1_U10.din1_cast_array[3] [5:4], 4'h0 };
assign _0311_ = \shl_8ns_8s_8_7_1_U10.dout_array[4]  << { \shl_8ns_8s_8_7_1_U10.din1_cast_array[4] [3:2], 2'h0 };
assign \shl_8ns_8s_8_7_1_U10.dout  = \shl_8ns_8s_8_7_1_U10.dout_array[5]  << \shl_8ns_8s_8_7_1_U10.din1_cast_array[5] [1:0];
assign \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.bin_s0  = ~ \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.b ;
always @(posedge \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.clk )
\sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.bin_s1  <= _0313_;
always @(posedge \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.clk )
\sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.ain_s1  <= _0312_;
always @(posedge \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.clk )
\sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.sum_s1  <= _0315_;
always @(posedge \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.clk )
\sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.carry_s1  <= _0314_;
assign _0313_ = \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.ce  ? \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.bin_s0 [3:2] : \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.bin_s1 ;
assign _0312_ = \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.ce  ? \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.a [3:2] : \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.ain_s1 ;
assign _0314_ = \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.ce  ? \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.facout_s1  : \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.carry_s1 ;
assign _0315_ = \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.ce  ? \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.fas_s1  : \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.sum_s1 ;
assign _0316_ = \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.u1.a  + \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.u1.b ;
assign { \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.u1.cout , \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.u1.s  } = _0316_ + \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.u1.cin ;
assign _0317_ = \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.u2.a  + \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.u2.b ;
assign { \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.u2.cout , \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.u2.s  } = _0317_ + \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.u2.cin ;
assign \sub_6ns_6s_6_2_1_U8.top_sub_6ns_6s_6_2_1_Adder_4_U.bin_s0  = ~ \sub_6ns_6s_6_2_1_U8.top_sub_6ns_6s_6_2_1_Adder_4_U.b ;
always @(posedge \sub_6ns_6s_6_2_1_U8.top_sub_6ns_6s_6_2_1_Adder_4_U.clk )
\sub_6ns_6s_6_2_1_U8.top_sub_6ns_6s_6_2_1_Adder_4_U.bin_s1  <= _0319_;
always @(posedge \sub_6ns_6s_6_2_1_U8.top_sub_6ns_6s_6_2_1_Adder_4_U.clk )
\sub_6ns_6s_6_2_1_U8.top_sub_6ns_6s_6_2_1_Adder_4_U.ain_s1  <= _0318_;
always @(posedge \sub_6ns_6s_6_2_1_U8.top_sub_6ns_6s_6_2_1_Adder_4_U.clk )
\sub_6ns_6s_6_2_1_U8.top_sub_6ns_6s_6_2_1_Adder_4_U.sum_s1  <= _0321_;
always @(posedge \sub_6ns_6s_6_2_1_U8.top_sub_6ns_6s_6_2_1_Adder_4_U.clk )
\sub_6ns_6s_6_2_1_U8.top_sub_6ns_6s_6_2_1_Adder_4_U.carry_s1  <= _0320_;
assign _0319_ = \sub_6ns_6s_6_2_1_U8.top_sub_6ns_6s_6_2_1_Adder_4_U.ce  ? \sub_6ns_6s_6_2_1_U8.top_sub_6ns_6s_6_2_1_Adder_4_U.bin_s0 [5:3] : \sub_6ns_6s_6_2_1_U8.top_sub_6ns_6s_6_2_1_Adder_4_U.bin_s1 ;
assign _0318_ = \sub_6ns_6s_6_2_1_U8.top_sub_6ns_6s_6_2_1_Adder_4_U.ce  ? \sub_6ns_6s_6_2_1_U8.top_sub_6ns_6s_6_2_1_Adder_4_U.a [5:3] : \sub_6ns_6s_6_2_1_U8.top_sub_6ns_6s_6_2_1_Adder_4_U.ain_s1 ;
assign _0320_ = \sub_6ns_6s_6_2_1_U8.top_sub_6ns_6s_6_2_1_Adder_4_U.ce  ? \sub_6ns_6s_6_2_1_U8.top_sub_6ns_6s_6_2_1_Adder_4_U.facout_s1  : \sub_6ns_6s_6_2_1_U8.top_sub_6ns_6s_6_2_1_Adder_4_U.carry_s1 ;
assign _0321_ = \sub_6ns_6s_6_2_1_U8.top_sub_6ns_6s_6_2_1_Adder_4_U.ce  ? \sub_6ns_6s_6_2_1_U8.top_sub_6ns_6s_6_2_1_Adder_4_U.fas_s1  : \sub_6ns_6s_6_2_1_U8.top_sub_6ns_6s_6_2_1_Adder_4_U.sum_s1 ;
assign _0322_ = \sub_6ns_6s_6_2_1_U8.top_sub_6ns_6s_6_2_1_Adder_4_U.u1.a  + \sub_6ns_6s_6_2_1_U8.top_sub_6ns_6s_6_2_1_Adder_4_U.u1.b ;
assign { \sub_6ns_6s_6_2_1_U8.top_sub_6ns_6s_6_2_1_Adder_4_U.u1.cout , \sub_6ns_6s_6_2_1_U8.top_sub_6ns_6s_6_2_1_Adder_4_U.u1.s  } = _0322_ + \sub_6ns_6s_6_2_1_U8.top_sub_6ns_6s_6_2_1_Adder_4_U.u1.cin ;
assign _0323_ = \sub_6ns_6s_6_2_1_U8.top_sub_6ns_6s_6_2_1_Adder_4_U.u2.a  + \sub_6ns_6s_6_2_1_U8.top_sub_6ns_6s_6_2_1_Adder_4_U.u2.b ;
assign { \sub_6ns_6s_6_2_1_U8.top_sub_6ns_6s_6_2_1_Adder_4_U.u2.cout , \sub_6ns_6s_6_2_1_U8.top_sub_6ns_6s_6_2_1_Adder_4_U.u2.s  } = _0323_ + \sub_6ns_6s_6_2_1_U8.top_sub_6ns_6s_6_2_1_Adder_4_U.u2.cin ;
assign \sub_6s_6ns_6_2_1_U2.top_sub_6s_6ns_6_2_1_Adder_1_U.bin_s0  = ~ \sub_6s_6ns_6_2_1_U2.top_sub_6s_6ns_6_2_1_Adder_1_U.b ;
always @(posedge \sub_6s_6ns_6_2_1_U2.top_sub_6s_6ns_6_2_1_Adder_1_U.clk )
\sub_6s_6ns_6_2_1_U2.top_sub_6s_6ns_6_2_1_Adder_1_U.bin_s1  <= _0325_;
always @(posedge \sub_6s_6ns_6_2_1_U2.top_sub_6s_6ns_6_2_1_Adder_1_U.clk )
\sub_6s_6ns_6_2_1_U2.top_sub_6s_6ns_6_2_1_Adder_1_U.ain_s1  <= _0324_;
always @(posedge \sub_6s_6ns_6_2_1_U2.top_sub_6s_6ns_6_2_1_Adder_1_U.clk )
\sub_6s_6ns_6_2_1_U2.top_sub_6s_6ns_6_2_1_Adder_1_U.sum_s1  <= _0327_;
always @(posedge \sub_6s_6ns_6_2_1_U2.top_sub_6s_6ns_6_2_1_Adder_1_U.clk )
\sub_6s_6ns_6_2_1_U2.top_sub_6s_6ns_6_2_1_Adder_1_U.carry_s1  <= _0326_;
assign _0325_ = \sub_6s_6ns_6_2_1_U2.top_sub_6s_6ns_6_2_1_Adder_1_U.ce  ? \sub_6s_6ns_6_2_1_U2.top_sub_6s_6ns_6_2_1_Adder_1_U.bin_s0 [5:3] : \sub_6s_6ns_6_2_1_U2.top_sub_6s_6ns_6_2_1_Adder_1_U.bin_s1 ;
assign _0324_ = \sub_6s_6ns_6_2_1_U2.top_sub_6s_6ns_6_2_1_Adder_1_U.ce  ? \sub_6s_6ns_6_2_1_U2.top_sub_6s_6ns_6_2_1_Adder_1_U.a [5:3] : \sub_6s_6ns_6_2_1_U2.top_sub_6s_6ns_6_2_1_Adder_1_U.ain_s1 ;
assign _0326_ = \sub_6s_6ns_6_2_1_U2.top_sub_6s_6ns_6_2_1_Adder_1_U.ce  ? \sub_6s_6ns_6_2_1_U2.top_sub_6s_6ns_6_2_1_Adder_1_U.facout_s1  : \sub_6s_6ns_6_2_1_U2.top_sub_6s_6ns_6_2_1_Adder_1_U.carry_s1 ;
assign _0327_ = \sub_6s_6ns_6_2_1_U2.top_sub_6s_6ns_6_2_1_Adder_1_U.ce  ? \sub_6s_6ns_6_2_1_U2.top_sub_6s_6ns_6_2_1_Adder_1_U.fas_s1  : \sub_6s_6ns_6_2_1_U2.top_sub_6s_6ns_6_2_1_Adder_1_U.sum_s1 ;
assign _0328_ = \sub_6s_6ns_6_2_1_U2.top_sub_6s_6ns_6_2_1_Adder_1_U.u1.a  + \sub_6s_6ns_6_2_1_U2.top_sub_6s_6ns_6_2_1_Adder_1_U.u1.b ;
assign { \sub_6s_6ns_6_2_1_U2.top_sub_6s_6ns_6_2_1_Adder_1_U.u1.cout , \sub_6s_6ns_6_2_1_U2.top_sub_6s_6ns_6_2_1_Adder_1_U.u1.s  } = _0328_ + \sub_6s_6ns_6_2_1_U2.top_sub_6s_6ns_6_2_1_Adder_1_U.u1.cin ;
assign _0329_ = \sub_6s_6ns_6_2_1_U2.top_sub_6s_6ns_6_2_1_Adder_1_U.u2.a  + \sub_6s_6ns_6_2_1_U2.top_sub_6s_6ns_6_2_1_Adder_1_U.u2.b ;
assign { \sub_6s_6ns_6_2_1_U2.top_sub_6s_6ns_6_2_1_Adder_1_U.u2.cout , \sub_6s_6ns_6_2_1_U2.top_sub_6s_6ns_6_2_1_Adder_1_U.u2.s  } = _0329_ + \sub_6s_6ns_6_2_1_U2.top_sub_6s_6ns_6_2_1_Adder_1_U.u2.cin ;
assign _0330_ = $signed({ 1'h0, icmp_ln1499_reg_1082, 6'h00 }) < $signed(op_4);
assign _0331_ = $signed(op_8) < $signed(op_5);
assign _0332_ = $signed({ op_3, 6'h00 }) != $signed(op_4);
assign _0333_ = | p_Result_s_18_reg_1255;
assign _0334_ = p_Result_s_18_reg_1255 != 5'h1f;
assign _0335_ = | trunc_ln851_3_reg_1402;
assign _0336_ = | op_13[6:0];
assign _0337_ = | op_15[4:0];
assign or_ln340_fu_628_p2 = p_Result_11_reg_1233 | overflow_fu_614_p2;
assign or_ln785_1_fu_755_p2 = xor_ln785_1_fu_750_p2 | p_Result_11_reg_1233;
assign or_ln785_2_fu_738_p2 = and_ln785_1_fu_734_p2 | and_ln340_1_fu_730_p2;
assign or_ln785_fu_583_p2 = p_Result_12_reg_1248 | icmp_ln768_reg_1271;
assign or_ln786_fu_623_p2 = xor_ln786_fu_618_p2 | icmp_ln786_reg_1276;
always @(posedge ap_clk)
ush_reg_1054 <= _0067_;
always @(posedge ap_clk)
sub_ln1367_reg_1044 <= _0063_;
always @(posedge ap_clk)
signbit_reg_1049 <= _0062_;
always @(posedge ap_clk)
shl_ln781_reg_1372 <= _0061_;
always @(posedge ap_clk)
shl_ln1299_reg_1189 <= _0060_;
always @(posedge ap_clk)
sh_V_1_reg_1172 <= _0059_;
always @(posedge ap_clk)
sext_ln850_reg_1447 <= _0058_;
always @(posedge ap_clk)
select_ln785_reg_1367 <= _0057_;
always @(posedge ap_clk)
select_ln353_reg_1459 <= _0056_;
always @(posedge ap_clk)
select_ln353_1_reg_1496 <= _0055_;
always @(posedge ap_clk)
ret_V_8_reg_1136 <= _0050_;
always @(posedge ap_clk)
ret_V_2_reg_1266 <= _0046_;
always @(posedge ap_clk)
ret_V_26_reg_1553 <= _0045_;
always @(posedge ap_clk)
ret_V_25_reg_1543 <= _0044_;
always @(posedge ap_clk)
ret_V_24_reg_1533 <= _0042_;
always @(posedge ap_clk)
ret_V_23_reg_1516 <= _0041_;
always @(posedge ap_clk)
ret_V_25_cast_reg_1521 <= _0043_;
always @(posedge ap_clk)
ret_V_22_reg_1479 <= _0039_;
always @(posedge ap_clk)
ret_V_23_cast_reg_1484 <= _0040_;
always @(posedge ap_clk)
ret_V_16_reg_1177 <= _0033_;
always @(posedge ap_clk)
ret_V_reg_1182 <= _0051_;
always @(posedge ap_clk)
r_V_1_reg_1199 <= _0030_;
always @(posedge ap_clk)
ret_V_3_cast_reg_1204 <= _0047_;
always @(posedge ap_clk)
trunc_ln851_1_reg_1211 <= _0065_;
always @(posedge ap_clk)
ret_V_20_reg_1141 <= _0037_;
always @(posedge ap_clk)
p_Result_14_reg_1147 <= _0027_;
always @(posedge ap_clk)
ret_V_17_reg_1287 <= _0034_;
always @(posedge ap_clk)
or_ln785_reg_1292 <= _0023_;
always @(posedge ap_clk)
xor_ln785_reg_1298 <= _0068_;
always @(posedge ap_clk)
ret_V_18_reg_1304 <= _0035_;
always @(posedge ap_clk)
op_12_V_reg_1387 <= _0020_;
always @(posedge ap_clk)
r_reg_1392 <= _0032_;
always @(posedge ap_clk)
op_23_V_reg_1397 <= _0021_;
always @(posedge ap_clk)
trunc_ln851_3_reg_1402 <= _0066_;
always @(posedge ap_clk)
isNeg_reg_1033 <= _0019_;
always @(posedge ap_clk)
icmp_ln851_reg_1167 <= _0018_;
always @(posedge ap_clk)
icmp_ln851_4_reg_1511 <= _0017_;
always @(posedge ap_clk)
icmp_ln851_3_reg_1474 <= _0016_;
always @(posedge ap_clk)
icmp_ln851_2_reg_1422 <= _0015_;
always @(posedge ap_clk)
r_V_reg_1226 <= _0031_;
always @(posedge ap_clk)
p_Result_11_reg_1233 <= _0025_;
always @(posedge ap_clk)
p_Val2_2_reg_1240 <= _0029_;
always @(posedge ap_clk)
p_Result_12_reg_1248 <= _0026_;
always @(posedge ap_clk)
p_Result_s_18_reg_1255 <= _0028_;
always @(posedge ap_clk)
icmp_ln851_1_reg_1261 <= _0014_;
always @(posedge ap_clk)
icmp_ln768_reg_1271 <= _0012_;
always @(posedge ap_clk)
icmp_ln786_reg_1276 <= _0013_;
always @(posedge ap_clk)
ret_V_4_reg_1282 <= _0048_;
always @(posedge ap_clk)
icmp_ln1499_reg_1082 <= _0011_;
always @(posedge ap_clk)
ret_V_19_reg_1113 <= _0036_;
always @(posedge ap_clk)
ret_V_7_reg_1119 <= _0049_;
always @(posedge ap_clk)
ret_reg_1126 <= _0052_;
always @(posedge ap_clk)
icmp_ln1494_reg_1131 <= _0010_;
always @(posedge ap_clk)
ashr_ln799_reg_1377 <= _0009_;
always @(posedge ap_clk)
ashr_ln1333_reg_1194 <= _0008_;
always @(posedge ap_clk)
or_ln786_reg_1314 <= _0024_;
always @(posedge ap_clk)
or_ln340_reg_1320 <= _0022_;
always @(posedge ap_clk)
and_ln786_reg_1326 <= _0006_;
always @(posedge ap_clk)
ret_V_21_reg_1432 <= _0038_;
always @(posedge ap_clk)
tmp_reg_1437 <= _0064_;
always @(posedge ap_clk)
add_ln69_3_reg_1442 <= _0004_;
always @(posedge ap_clk)
select_ln340_reg_1347 <= _0054_;
always @(posedge ap_clk)
sel_tmp11_reg_1352 <= _0053_;
always @(posedge ap_clk)
add_ln69_reg_1357 <= _0005_;
always @(posedge ap_clk)
add_ln69_1_reg_1362 <= _0003_;
always @(posedge ap_clk)
add_ln691_reg_1454 <= _0002_;
always @(posedge ap_clk)
add_ln691_2_reg_1528 <= _0001_;
always @(posedge ap_clk)
add_ln691_1_reg_1491 <= _0000_;
always @(posedge ap_clk)
ap_CS_fsm <= _0007_;
assign _0069_ = _0081_ ? 2'h2 : 2'h1;
assign _0338_ = ap_CS_fsm == 1'h1;
function [37:0] _0923_;
input [37:0] a;
input [1443:0] b;
input [37:0] s;
case (s)
38'b00000000000000000000000000000000000001:
_0923_ = b[37:0];
38'b00000000000000000000000000000000000010:
_0923_ = b[75:38];
38'b00000000000000000000000000000000000100:
_0923_ = b[113:76];
38'b00000000000000000000000000000000001000:
_0923_ = b[151:114];
38'b00000000000000000000000000000000010000:
_0923_ = b[189:152];
38'b00000000000000000000000000000000100000:
_0923_ = b[227:190];
38'b00000000000000000000000000000001000000:
_0923_ = b[265:228];
38'b00000000000000000000000000000010000000:
_0923_ = b[303:266];
38'b00000000000000000000000000000100000000:
_0923_ = b[341:304];
38'b00000000000000000000000000001000000000:
_0923_ = b[379:342];
38'b00000000000000000000000000010000000000:
_0923_ = b[417:380];
38'b00000000000000000000000000100000000000:
_0923_ = b[455:418];
38'b00000000000000000000000001000000000000:
_0923_ = b[493:456];
38'b00000000000000000000000010000000000000:
_0923_ = b[531:494];
38'b00000000000000000000000100000000000000:
_0923_ = b[569:532];
38'b00000000000000000000001000000000000000:
_0923_ = b[607:570];
38'b00000000000000000000010000000000000000:
_0923_ = b[645:608];
38'b00000000000000000000100000000000000000:
_0923_ = b[683:646];
38'b00000000000000000001000000000000000000:
_0923_ = b[721:684];
38'b00000000000000000010000000000000000000:
_0923_ = b[759:722];
38'b00000000000000000100000000000000000000:
_0923_ = b[797:760];
38'b00000000000000001000000000000000000000:
_0923_ = b[835:798];
38'b00000000000000010000000000000000000000:
_0923_ = b[873:836];
38'b00000000000000100000000000000000000000:
_0923_ = b[911:874];
38'b00000000000001000000000000000000000000:
_0923_ = b[949:912];
38'b00000000000010000000000000000000000000:
_0923_ = b[987:950];
38'b00000000000100000000000000000000000000:
_0923_ = b[1025:988];
38'b00000000001000000000000000000000000000:
_0923_ = b[1063:1026];
38'b00000000010000000000000000000000000000:
_0923_ = b[1101:1064];
38'b00000000100000000000000000000000000000:
_0923_ = b[1139:1102];
38'b00000001000000000000000000000000000000:
_0923_ = b[1177:1140];
38'b00000010000000000000000000000000000000:
_0923_ = b[1215:1178];
38'b00000100000000000000000000000000000000:
_0923_ = b[1253:1216];
38'b00001000000000000000000000000000000000:
_0923_ = b[1291:1254];
38'b00010000000000000000000000000000000000:
_0923_ = b[1329:1292];
38'b00100000000000000000000000000000000000:
_0923_ = b[1367:1330];
38'b01000000000000000000000000000000000000:
_0923_ = b[1405:1368];
38'b10000000000000000000000000000000000000:
_0923_ = b[1443:1406];
38'b00000000000000000000000000000000000000:
_0923_ = a;
default:
_0923_ = 38'bx;
endcase
endfunction
assign ap_NS_fsm = _0923_(38'hxxxxxxxxxx, { 36'h000000000, _0069_, 1406'h0000000004000000002000000001000000000800000000400000000200000000100000000080000000040000000020000000010000000008000000004000000002000000001000000000800000000400000000200000000100000000080000000040000000020000000010000000008000000004000000002000000001000000000800000000400000000200000000100000000080000000040000000020000000010000000008000000000000000001 }, { _0338_, _0375_, _0374_, _0373_, _0372_, _0371_, _0370_, _0369_, _0368_, _0367_, _0366_, _0365_, _0364_, _0363_, _0362_, _0361_, _0360_, _0359_, _0358_, _0357_, _0356_, _0355_, _0354_, _0353_, _0352_, _0351_, _0350_, _0349_, _0348_, _0347_, _0346_, _0345_, _0344_, _0343_, _0342_, _0341_, _0340_, _0339_ });
assign _0339_ = ap_CS_fsm == 38'h2000000000;
assign _0340_ = ap_CS_fsm == 37'h1000000000;
assign _0341_ = ap_CS_fsm == 36'h800000000;
assign _0342_ = ap_CS_fsm == 35'h400000000;
assign _0343_ = ap_CS_fsm == 34'h200000000;
assign _0344_ = ap_CS_fsm == 33'h100000000;
assign _0345_ = ap_CS_fsm == 32'd2147483648;
assign _0346_ = ap_CS_fsm == 31'h40000000;
assign _0347_ = ap_CS_fsm == 30'h20000000;
assign _0348_ = ap_CS_fsm == 29'h10000000;
assign _0349_ = ap_CS_fsm == 28'h8000000;
assign _0350_ = ap_CS_fsm == 27'h4000000;
assign _0351_ = ap_CS_fsm == 26'h2000000;
assign _0352_ = ap_CS_fsm == 25'h1000000;
assign _0353_ = ap_CS_fsm == 24'h800000;
assign _0354_ = ap_CS_fsm == 23'h400000;
assign _0355_ = ap_CS_fsm == 22'h200000;
assign _0356_ = ap_CS_fsm == 21'h100000;
assign _0357_ = ap_CS_fsm == 20'h80000;
assign _0358_ = ap_CS_fsm == 19'h40000;
assign _0359_ = ap_CS_fsm == 18'h20000;
assign _0360_ = ap_CS_fsm == 17'h10000;
assign _0361_ = ap_CS_fsm == 16'h8000;
assign _0362_ = ap_CS_fsm == 15'h4000;
assign _0363_ = ap_CS_fsm == 14'h2000;
assign _0364_ = ap_CS_fsm == 13'h1000;
assign _0365_ = ap_CS_fsm == 12'h800;
assign _0366_ = ap_CS_fsm == 11'h400;
assign _0367_ = ap_CS_fsm == 10'h200;
assign _0368_ = ap_CS_fsm == 9'h100;
assign _0369_ = ap_CS_fsm == 8'h80;
assign _0370_ = ap_CS_fsm == 7'h40;
assign _0371_ = ap_CS_fsm == 6'h20;
assign _0372_ = ap_CS_fsm == 5'h10;
assign _0373_ = ap_CS_fsm == 4'h8;
assign _0374_ = ap_CS_fsm == 3'h4;
assign _0375_ = ap_CS_fsm == 2'h2;
assign op_30_ap_vld = ap_CS_fsm[37] ? 1'h1 : 1'h0;
assign ap_idle = _0080_ ? 1'h1 : 1'h0;
assign _0067_ = ap_CS_fsm[2] ? ush_fu_262_p3 : ush_reg_1054;
assign _0062_ = ap_CS_fsm[1] ? signbit_fu_257_p2 : signbit_reg_1049;
assign _0063_ = ap_CS_fsm[1] ? grp_fu_247_p2 : sub_ln1367_reg_1044;
assign _0061_ = _0079_ ? grp_fu_485_p2 : shl_ln781_reg_1372;
assign _0060_ = _0078_ ? grp_fu_316_p2 : shl_ln1299_reg_1189;
assign _0059_ = _0077_ ? grp_fu_420_p2 : sh_V_1_reg_1172;
assign _0058_ = ap_CS_fsm[19] ? { tmp_reg_1437[7], tmp_reg_1437 } : sext_ln850_reg_1447;
assign _0057_ = _0076_ ? select_ln785_fu_765_p3 : select_ln785_reg_1367;
assign _0056_ = ap_CS_fsm[21] ? select_ln353_fu_861_p3 : select_ln353_reg_1459;
assign _0055_ = ap_CS_fsm[26] ? select_ln353_1_fu_926_p3 : select_ln353_1_reg_1496;
assign _0050_ = ap_CS_fsm[5] ? grp_fu_381_p2 : ret_V_8_reg_1136;
assign _0046_ = _0075_ ? grp_fu_498_p2 : ret_V_2_reg_1266;
assign _0045_ = ap_CS_fsm[35] ? grp_fu_1011_p2 : ret_V_26_reg_1553;
assign _0044_ = ap_CS_fsm[33] ? grp_fu_1002_p2 : ret_V_25_reg_1543;
assign _0042_ = ap_CS_fsm[31] ? ret_V_24_fu_991_p3 : ret_V_24_reg_1533;
assign _0043_ = ap_CS_fsm[28] ? grp_fu_948_p2[36:5] : ret_V_25_cast_reg_1521;
assign _0041_ = ap_CS_fsm[28] ? grp_fu_948_p2 : ret_V_23_reg_1516;
assign _0040_ = ap_CS_fsm[23] ? grp_fu_883_p2[38:7] : ret_V_23_cast_reg_1484;
assign _0039_ = ap_CS_fsm[23] ? grp_fu_883_p2 : ret_V_22_reg_1479;
assign _0065_ = ap_CS_fsm[9] ? grp_fu_336_p2[5:0] : trunc_ln851_1_reg_1211;
assign _0047_ = ap_CS_fsm[9] ? grp_fu_336_p2[9:6] : ret_V_3_cast_reg_1204;
assign _0030_ = ap_CS_fsm[9] ? grp_fu_336_p2 : r_V_1_reg_1199;
assign _0051_ = ap_CS_fsm[9] ? grp_fu_442_p2[8:3] : ret_V_reg_1182;
assign _0033_ = ap_CS_fsm[9] ? grp_fu_442_p2 : ret_V_16_reg_1177;
assign _0027_ = ap_CS_fsm[6] ? ret_V_20_fu_402_p3[4] : p_Result_14_reg_1147;
assign _0037_ = ap_CS_fsm[6] ? ret_V_20_fu_402_p3 : ret_V_20_reg_1141;
assign _0035_ = ap_CS_fsm[12] ? ret_V_18_fu_604_p3 : ret_V_18_reg_1304;
assign _0068_ = ap_CS_fsm[12] ? xor_ln785_fu_587_p2 : xor_ln785_reg_1298;
assign _0023_ = ap_CS_fsm[12] ? or_ln785_fu_583_p2 : or_ln785_reg_1292;
assign _0034_ = ap_CS_fsm[12] ? ret_V_17_fu_576_p3 : ret_V_17_reg_1287;
assign _0066_ = ap_CS_fsm[16] ? op_12_V_fu_779_p3[2:0] : trunc_ln851_3_reg_1402;
assign _0021_ = ap_CS_fsm[16] ? grp_fu_774_p2 : op_23_V_reg_1397;
assign _0032_ = ap_CS_fsm[16] ? r_fu_784_p3 : r_reg_1392;
assign _0020_ = ap_CS_fsm[16] ? op_12_V_fu_779_p3 : op_12_V_reg_1387;
assign _0019_ = ap_CS_fsm[0] ? op_5[3] : isNeg_reg_1033;
assign _0018_ = ap_CS_fsm[8] ? icmp_ln851_fu_452_p2 : icmp_ln851_reg_1167;
assign _0017_ = ap_CS_fsm[27] ? icmp_ln851_4_fu_958_p2 : icmp_ln851_4_reg_1511;
assign _0016_ = ap_CS_fsm[22] ? icmp_ln851_3_fu_893_p2 : icmp_ln851_3_reg_1474;
assign _0015_ = ap_CS_fsm[17] ? icmp_ln851_2_fu_816_p2 : icmp_ln851_2_reg_1422;
assign _0014_ = ap_CS_fsm[10] ? icmp_ln851_1_fu_544_p2 : icmp_ln851_1_reg_1261;
assign _0028_ = ap_CS_fsm[10] ? r_V_fu_503_p3[15:11] : p_Result_s_18_reg_1255;
assign _0026_ = ap_CS_fsm[10] ? r_V_fu_503_p3[10] : p_Result_12_reg_1248;
assign _0029_ = ap_CS_fsm[10] ? r_V_fu_503_p3[10:3] : p_Val2_2_reg_1240;
assign _0025_ = ap_CS_fsm[10] ? r_V_fu_503_p3[15] : p_Result_11_reg_1233;
assign _0031_ = ap_CS_fsm[10] ? r_V_fu_503_p3 : r_V_reg_1226;
assign _0048_ = ap_CS_fsm[11] ? grp_fu_549_p2 : ret_V_4_reg_1282;
assign _0013_ = ap_CS_fsm[11] ? icmp_ln786_fu_559_p2 : icmp_ln786_reg_1276;
assign _0012_ = ap_CS_fsm[11] ? icmp_ln768_fu_554_p2 : icmp_ln768_reg_1271;
assign _0049_ = ap_CS_fsm[3] ? grp_fu_289_p2[5:1] : ret_V_7_reg_1119;
assign _0036_ = ap_CS_fsm[3] ? grp_fu_289_p2 : ret_V_19_reg_1113;
assign _0011_ = ap_CS_fsm[3] ? icmp_ln1499_fu_307_p2 : icmp_ln1499_reg_1082;
assign _0010_ = ap_CS_fsm[4] ? icmp_ln1494_fu_376_p2 : icmp_ln1494_reg_1131;
assign _0052_ = ap_CS_fsm[4] ? grp_fu_349_p2 : ret_reg_1126;
assign _0009_ = _0074_ ? grp_fu_493_p2 : ashr_ln799_reg_1377;
assign _0008_ = _0073_ ? grp_fu_322_p2 : ashr_ln1333_reg_1194;
assign _0006_ = ap_CS_fsm[13] ? and_ln786_fu_638_p2 : and_ln786_reg_1326;
assign _0022_ = ap_CS_fsm[13] ? or_ln340_fu_628_p2 : or_ln340_reg_1320;
assign _0024_ = ap_CS_fsm[13] ? or_ln786_fu_623_p2 : or_ln786_reg_1314;
assign _0004_ = ap_CS_fsm[18] ? grp_fu_824_p2 : add_ln69_3_reg_1442;
assign _0064_ = ap_CS_fsm[18] ? grp_fu_810_p2[10:3] : tmp_reg_1437;
assign _0038_ = ap_CS_fsm[18] ? grp_fu_810_p2 : ret_V_21_reg_1432;
assign _0003_ = ap_CS_fsm[14] ? grp_fu_659_p2 : add_ln69_1_reg_1362;
assign _0005_ = ap_CS_fsm[14] ? grp_fu_653_p2 : add_ln69_reg_1357;
assign _0053_ = ap_CS_fsm[14] ? sel_tmp11_fu_744_p2 : sel_tmp11_reg_1352;
assign _0054_ = ap_CS_fsm[14] ? select_ln340_fu_723_p3 : select_ln340_reg_1347;
assign _0002_ = _0072_ ? grp_fu_843_p2 : add_ln691_reg_1454;
assign _0001_ = _0071_ ? grp_fu_974_p2 : add_ln691_2_reg_1528;
assign _0000_ = _0070_ ? grp_fu_909_p2 : add_ln691_1_reg_1491;
assign _0007_ = ap_rst ? 38'h0000000001 : ap_NS_fsm;
assign icmp_ln1494_fu_376_p2 = _0330_ ? 1'h1 : 1'h0;
assign icmp_ln1499_fu_307_p2 = _0332_ ? 1'h1 : 1'h0;
assign icmp_ln768_fu_554_p2 = _0333_ ? 1'h1 : 1'h0;
assign icmp_ln786_fu_559_p2 = _0334_ ? 1'h1 : 1'h0;
assign icmp_ln851_1_fu_544_p2 = _0087_ ? 1'h1 : 1'h0;
assign icmp_ln851_2_fu_816_p2 = _0335_ ? 1'h1 : 1'h0;
assign icmp_ln851_3_fu_893_p2 = _0336_ ? 1'h1 : 1'h0;
assign icmp_ln851_4_fu_958_p2 = _0337_ ? 1'h1 : 1'h0;
assign icmp_ln851_fu_452_p2 = _0088_ ? 1'h1 : 1'h0;
assign op_12_V_fu_779_p3 = sel_tmp11_reg_1352 ? p_Val2_2_reg_1240 : select_ln785_reg_1367;
assign r_V_fu_503_p3 = isNeg_reg_1033 ? shl_ln1299_reg_1189 : ashr_ln1333_reg_1194;
assign r_fu_784_p3 = p_Result_14_reg_1147 ? shl_ln781_reg_1372 : ashr_ln799_reg_1377;
assign ret_V_17_fu_576_p3 = ret_V_16_reg_1177[8] ? select_ln850_fu_571_p3 : ret_V_reg_1182;
assign ret_V_18_fu_604_p3 = r_V_1_reg_1199[17] ? select_ln850_1_fu_599_p3 : ret_V_3_cast_reg_1204;
assign ret_V_20_fu_402_p3 = ret_V_19_reg_1113[5] ? select_ln850_2_fu_396_p3 : ret_V_7_reg_1119;
assign ret_V_24_fu_991_p3 = ret_V_23_reg_1516[37] ? select_ln850_5_fu_986_p3 : ret_V_25_cast_reg_1521;
assign select_ln340_fu_723_p3 = and_ln340_fu_718_p2 ? p_Val2_2_reg_1240 : { r_V_reg_1226[11], p_Val2_3_fu_698_p2 };
assign select_ln353_1_fu_926_p3 = ret_V_22_reg_1479[39] ? select_ln850_7_fu_921_p3 : ret_V_23_cast_reg_1484;
assign select_ln353_fu_861_p3 = ret_V_21_reg_1432[10] ? select_ln850_6_fu_856_p3 : sext_ln850_reg_1447;
assign select_ln785_fu_765_p3 = and_ln785_fu_760_p2 ? p_Val2_2_reg_1240 : select_ln340_reg_1347;
assign select_ln850_1_fu_599_p3 = icmp_ln851_1_reg_1261 ? ret_V_3_cast_reg_1204 : ret_V_4_reg_1282;
assign select_ln850_2_fu_396_p3 = ret_V_19_reg_1113[0] ? ret_V_8_reg_1136 : ret_V_7_reg_1119;
assign select_ln850_5_fu_986_p3 = icmp_ln851_4_reg_1511 ? add_ln691_2_reg_1528 : ret_V_25_cast_reg_1521;
assign select_ln850_6_fu_856_p3 = icmp_ln851_2_reg_1422 ? add_ln691_reg_1454 : sext_ln850_reg_1447;
assign select_ln850_7_fu_921_p3 = icmp_ln851_3_reg_1474 ? add_ln691_1_reg_1491 : ret_V_23_cast_reg_1484;
assign select_ln850_fu_571_p3 = icmp_ln851_reg_1167 ? ret_V_reg_1182 : ret_V_2_reg_1266;
assign signbit_fu_257_p2 = _0331_ ? 1'h1 : 1'h0;
assign ush_fu_262_p3 = isNeg_reg_1033 ? sub_ln1367_reg_1044 : op_5;
assign xor_ln365_fu_686_p2 = r_V_reg_1226[10] ^ r_V_reg_1226[11];
assign ap_CS_fsm_state1 = ap_CS_fsm[0];
assign ap_CS_fsm_state10 = ap_CS_fsm[9];
assign ap_CS_fsm_state11 = ap_CS_fsm[10];
assign ap_CS_fsm_state12 = ap_CS_fsm[11];
assign ap_CS_fsm_state13 = ap_CS_fsm[12];
assign ap_CS_fsm_state14 = ap_CS_fsm[13];
assign ap_CS_fsm_state15 = ap_CS_fsm[14];
assign ap_CS_fsm_state16 = ap_CS_fsm[15];
assign ap_CS_fsm_state17 = ap_CS_fsm[16];
assign ap_CS_fsm_state18 = ap_CS_fsm[17];
assign ap_CS_fsm_state19 = ap_CS_fsm[18];
assign ap_CS_fsm_state2 = ap_CS_fsm[1];
assign ap_CS_fsm_state20 = ap_CS_fsm[19];
assign ap_CS_fsm_state21 = ap_CS_fsm[20];
assign ap_CS_fsm_state22 = ap_CS_fsm[21];
assign ap_CS_fsm_state23 = ap_CS_fsm[22];
assign ap_CS_fsm_state24 = ap_CS_fsm[23];
assign ap_CS_fsm_state25 = ap_CS_fsm[24];
assign ap_CS_fsm_state26 = ap_CS_fsm[25];
assign ap_CS_fsm_state27 = ap_CS_fsm[26];
assign ap_CS_fsm_state28 = ap_CS_fsm[27];
assign ap_CS_fsm_state29 = ap_CS_fsm[28];
assign ap_CS_fsm_state3 = ap_CS_fsm[2];
assign ap_CS_fsm_state30 = ap_CS_fsm[29];
assign ap_CS_fsm_state31 = ap_CS_fsm[30];
assign ap_CS_fsm_state32 = ap_CS_fsm[31];
assign ap_CS_fsm_state33 = ap_CS_fsm[32];
assign ap_CS_fsm_state34 = ap_CS_fsm[33];
assign ap_CS_fsm_state35 = ap_CS_fsm[34];
assign ap_CS_fsm_state36 = ap_CS_fsm[35];
assign ap_CS_fsm_state37 = ap_CS_fsm[36];
assign ap_CS_fsm_state38 = ap_CS_fsm[37];
assign ap_CS_fsm_state4 = ap_CS_fsm[3];
assign ap_CS_fsm_state5 = ap_CS_fsm[4];
assign ap_CS_fsm_state6 = ap_CS_fsm[5];
assign ap_CS_fsm_state7 = ap_CS_fsm[6];
assign ap_CS_fsm_state8 = ap_CS_fsm[7];
assign ap_CS_fsm_state9 = ap_CS_fsm[8];
assign ap_done = op_30_ap_vld;
assign ap_ready = op_30_ap_vld;
assign grp_fu_1002_p1 = { op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16 };
assign grp_fu_1011_p1 = { op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17 };
assign grp_fu_1019_p0 = { add_ln69_3_reg_1442[9], add_ln69_3_reg_1442[9], add_ln69_3_reg_1442[9], add_ln69_3_reg_1442[9], add_ln69_3_reg_1442[9], add_ln69_3_reg_1442[9], add_ln69_3_reg_1442[9], add_ln69_3_reg_1442[9], add_ln69_3_reg_1442[9], add_ln69_3_reg_1442[9], add_ln69_3_reg_1442[9], add_ln69_3_reg_1442[9], add_ln69_3_reg_1442[9], add_ln69_3_reg_1442[9], add_ln69_3_reg_1442[9], add_ln69_3_reg_1442[9], add_ln69_3_reg_1442[9], add_ln69_3_reg_1442[9], add_ln69_3_reg_1442[9], add_ln69_3_reg_1442[9], add_ln69_3_reg_1442[9], add_ln69_3_reg_1442[9], add_ln69_3_reg_1442 };
assign grp_fu_289_p0 = { op_5[3], op_5, 1'h0 };
assign grp_fu_289_p1 = { 4'h0, signbit_reg_1049, 1'h0 };
assign grp_fu_349_p0 = { op_8[1], op_8 };
assign grp_fu_349_p1 = { op_7[1], op_7 };
assign grp_fu_420_p1 = { ret_V_20_reg_1141[4], ret_V_20_reg_1141 };
assign grp_fu_442_p0 = { 4'h0, op_0, 3'h0 };
assign grp_fu_442_p1 = { op_1[7], op_1 };
assign grp_fu_485_p1 = { sh_V_1_reg_1172[5], sh_V_1_reg_1172[5], sh_V_1_reg_1172 };
assign grp_fu_493_p1 = { ret_V_20_reg_1141[4], ret_V_20_reg_1141[4], ret_V_20_reg_1141[4], ret_V_20_reg_1141 };
assign grp_fu_653_p0 = { ret_V_17_reg_1287[5], ret_V_17_reg_1287 };
assign grp_fu_653_p1 = { 3'h0, ret_V_18_reg_1304 };
assign grp_fu_659_p0 = { 1'h0, op_2 };
assign grp_fu_659_p1 = { 2'h0, icmp_ln1494_reg_1131 };
assign grp_fu_774_p0 = { 4'h0, add_ln69_1_reg_1362 };
assign grp_fu_810_p0 = { op_23_V_reg_1397[6], op_23_V_reg_1397, 3'h0 };
assign grp_fu_810_p1 = { op_12_V_reg_1387[7], op_12_V_reg_1387[7], op_12_V_reg_1387[7], op_12_V_reg_1387 };
assign grp_fu_824_p0 = { 2'h0, r_reg_1392 };
assign grp_fu_824_p1 = { ret_reg_1126[2], ret_reg_1126[2], ret_reg_1126[2], ret_reg_1126[2], ret_reg_1126[2], ret_reg_1126[2], ret_reg_1126[2], ret_reg_1126 };
assign grp_fu_843_p0 = { tmp_reg_1437[7], tmp_reg_1437 };
assign grp_fu_883_p0 = { select_ln353_reg_1459[8], select_ln353_reg_1459[8], select_ln353_reg_1459[8], select_ln353_reg_1459[8], select_ln353_reg_1459[8], select_ln353_reg_1459[8], select_ln353_reg_1459[8], select_ln353_reg_1459[8], select_ln353_reg_1459[8], select_ln353_reg_1459[8], select_ln353_reg_1459[8], select_ln353_reg_1459[8], select_ln353_reg_1459[8], select_ln353_reg_1459[8], select_ln353_reg_1459[8], select_ln353_reg_1459[8], select_ln353_reg_1459[8], select_ln353_reg_1459[8], select_ln353_reg_1459[8], select_ln353_reg_1459[8], select_ln353_reg_1459[8], select_ln353_reg_1459[8], select_ln353_reg_1459[8], select_ln353_reg_1459[8], select_ln353_reg_1459, 7'h00 };
assign grp_fu_883_p1 = { op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13 };
assign grp_fu_948_p0 = { select_ln353_1_reg_1496[31], select_ln353_1_reg_1496, 5'h00 };
assign grp_fu_948_p1 = { op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15 };
assign icmp_ln1494_fu_376_p1 = op_4;
assign icmp_ln1499_fu_307_p1 = op_4;
assign lhs_V_fu_274_p3 = { op_5, 1'h0 };
assign lhs_fu_426_p3 = { op_0, 3'h0 };
assign op_30 = grp_fu_1019_p2;
assign op_9_V_fu_267_p3 = { signbit_reg_1049, 1'h0 };
assign p_Result_10_fu_979_p3 = ret_V_23_reg_1516[37];
assign p_Result_13_fu_665_p3 = r_V_reg_1226[11];
assign p_Result_4_fu_703_p4 = { r_V_reg_1226[11], p_Val2_3_fu_698_p2 };
assign p_Result_5_fu_592_p3 = r_V_1_reg_1199[17];
assign p_Result_6_fu_386_p3 = ret_V_19_reg_1113[5];
assign p_Result_8_fu_849_p3 = ret_V_21_reg_1432[10];
assign p_Result_9_fu_914_p3 = ret_V_22_reg_1479[39];
assign p_Result_s_fu_564_p3 = ret_V_16_reg_1177[8];
assign rhs_2_fu_799_p3 = { op_23_V_reg_1397, 3'h0 };
assign rhs_3_fu_937_p3 = { select_ln353_1_reg_1496, 5'h00 };
assign sext_ln1499_fu_303_p1 = { op_3[7], op_3[7], op_3, 6'h00 };
assign sext_ln215_1_fu_346_p0 = op_8;
assign sext_ln215_fu_342_p0 = op_7;
assign sext_ln703_1_fu_868_p0 = op_13;
assign sext_ln703_2_fu_933_p0 = op_15;
assign sext_ln703_fu_438_p0 = op_1;
assign sext_ln850_fu_840_p1 = { tmp_reg_1437[7], tmp_reg_1437 };
assign sext_ln886_fu_253_p0 = op_8;
assign sext_ln886_fu_253_p1 = { op_8[1], op_8[1], op_8 };
assign shl_ln728_2_fu_365_p3 = { icmp_ln1499_reg_1082, 6'h00 };
assign shl_ln_fu_295_p3 = { op_3, 6'h00 };
assign tmp_13_fu_872_p3 = { select_ln353_reg_1459, 7'h00 };
assign tmp_6_fu_672_p3 = r_V_reg_1226[11];
assign tmp_7_fu_679_p3 = r_V_reg_1226[10];
assign trunc_ln851_1_fu_478_p1 = grp_fu_336_p2[5:0];
assign trunc_ln851_2_fu_393_p1 = ret_V_19_reg_1113[0];
assign trunc_ln851_3_fu_789_p1 = op_12_V_fu_779_p3[2:0];
assign trunc_ln851_4_fu_889_p0 = op_13;
assign trunc_ln851_4_fu_889_p1 = op_13[6:0];
assign trunc_ln851_5_fu_954_p0 = op_15;
assign trunc_ln851_5_fu_954_p1 = op_15[4:0];
assign trunc_ln851_fu_448_p0 = op_1;
assign trunc_ln851_fu_448_p1 = op_1[2:0];
assign zext_ln1367_fu_313_p1 = { 12'h000, ush_reg_1054 };
assign zext_ln1494_fu_372_p1 = { 9'h000, icmp_ln1499_reg_1082, 6'h00 };
assign \sub_6s_6ns_6_2_1_U2.top_sub_6s_6ns_6_2_1_Adder_1_U.ain_s0  = \sub_6s_6ns_6_2_1_U2.top_sub_6s_6ns_6_2_1_Adder_1_U.a ;
assign \sub_6s_6ns_6_2_1_U2.top_sub_6s_6ns_6_2_1_Adder_1_U.s  = { \sub_6s_6ns_6_2_1_U2.top_sub_6s_6ns_6_2_1_Adder_1_U.fas_s2 , \sub_6s_6ns_6_2_1_U2.top_sub_6s_6ns_6_2_1_Adder_1_U.sum_s1  };
assign \sub_6s_6ns_6_2_1_U2.top_sub_6s_6ns_6_2_1_Adder_1_U.u2.a  = \sub_6s_6ns_6_2_1_U2.top_sub_6s_6ns_6_2_1_Adder_1_U.ain_s1 ;
assign \sub_6s_6ns_6_2_1_U2.top_sub_6s_6ns_6_2_1_Adder_1_U.u2.b  = \sub_6s_6ns_6_2_1_U2.top_sub_6s_6ns_6_2_1_Adder_1_U.bin_s1 ;
assign \sub_6s_6ns_6_2_1_U2.top_sub_6s_6ns_6_2_1_Adder_1_U.u2.cin  = \sub_6s_6ns_6_2_1_U2.top_sub_6s_6ns_6_2_1_Adder_1_U.carry_s1 ;
assign \sub_6s_6ns_6_2_1_U2.top_sub_6s_6ns_6_2_1_Adder_1_U.facout_s2  = \sub_6s_6ns_6_2_1_U2.top_sub_6s_6ns_6_2_1_Adder_1_U.u2.cout ;
assign \sub_6s_6ns_6_2_1_U2.top_sub_6s_6ns_6_2_1_Adder_1_U.fas_s2  = \sub_6s_6ns_6_2_1_U2.top_sub_6s_6ns_6_2_1_Adder_1_U.u2.s ;
assign \sub_6s_6ns_6_2_1_U2.top_sub_6s_6ns_6_2_1_Adder_1_U.u1.a  = \sub_6s_6ns_6_2_1_U2.top_sub_6s_6ns_6_2_1_Adder_1_U.a [2:0];
assign \sub_6s_6ns_6_2_1_U2.top_sub_6s_6ns_6_2_1_Adder_1_U.u1.b  = \sub_6s_6ns_6_2_1_U2.top_sub_6s_6ns_6_2_1_Adder_1_U.bin_s0 [2:0];
assign \sub_6s_6ns_6_2_1_U2.top_sub_6s_6ns_6_2_1_Adder_1_U.u1.cin  = 1'h1;
assign \sub_6s_6ns_6_2_1_U2.top_sub_6s_6ns_6_2_1_Adder_1_U.facout_s1  = \sub_6s_6ns_6_2_1_U2.top_sub_6s_6ns_6_2_1_Adder_1_U.u1.cout ;
assign \sub_6s_6ns_6_2_1_U2.top_sub_6s_6ns_6_2_1_Adder_1_U.fas_s1  = \sub_6s_6ns_6_2_1_U2.top_sub_6s_6ns_6_2_1_Adder_1_U.u1.s ;
assign \sub_6s_6ns_6_2_1_U2.top_sub_6s_6ns_6_2_1_Adder_1_U.a  = \sub_6s_6ns_6_2_1_U2.din0 ;
assign \sub_6s_6ns_6_2_1_U2.top_sub_6s_6ns_6_2_1_Adder_1_U.b  = \sub_6s_6ns_6_2_1_U2.din1 ;
assign \sub_6s_6ns_6_2_1_U2.top_sub_6s_6ns_6_2_1_Adder_1_U.ce  = \sub_6s_6ns_6_2_1_U2.ce ;
assign \sub_6s_6ns_6_2_1_U2.top_sub_6s_6ns_6_2_1_Adder_1_U.clk  = \sub_6s_6ns_6_2_1_U2.clk ;
assign \sub_6s_6ns_6_2_1_U2.top_sub_6s_6ns_6_2_1_Adder_1_U.reset  = \sub_6s_6ns_6_2_1_U2.reset ;
assign \sub_6s_6ns_6_2_1_U2.dout  = \sub_6s_6ns_6_2_1_U2.top_sub_6s_6ns_6_2_1_Adder_1_U.s ;
assign \sub_6s_6ns_6_2_1_U2.ce  = 1'h1;
assign \sub_6s_6ns_6_2_1_U2.clk  = ap_clk;
assign \sub_6s_6ns_6_2_1_U2.din0  = { op_5[3], op_5, 1'h0 };
assign \sub_6s_6ns_6_2_1_U2.din1  = { 4'h0, signbit_reg_1049, 1'h0 };
assign grp_fu_289_p2 = \sub_6s_6ns_6_2_1_U2.dout ;
assign \sub_6s_6ns_6_2_1_U2.reset  = ap_rst;
assign \sub_6ns_6s_6_2_1_U8.top_sub_6ns_6s_6_2_1_Adder_4_U.ain_s0  = \sub_6ns_6s_6_2_1_U8.top_sub_6ns_6s_6_2_1_Adder_4_U.a ;
assign \sub_6ns_6s_6_2_1_U8.top_sub_6ns_6s_6_2_1_Adder_4_U.s  = { \sub_6ns_6s_6_2_1_U8.top_sub_6ns_6s_6_2_1_Adder_4_U.fas_s2 , \sub_6ns_6s_6_2_1_U8.top_sub_6ns_6s_6_2_1_Adder_4_U.sum_s1  };
assign \sub_6ns_6s_6_2_1_U8.top_sub_6ns_6s_6_2_1_Adder_4_U.u2.a  = \sub_6ns_6s_6_2_1_U8.top_sub_6ns_6s_6_2_1_Adder_4_U.ain_s1 ;
assign \sub_6ns_6s_6_2_1_U8.top_sub_6ns_6s_6_2_1_Adder_4_U.u2.b  = \sub_6ns_6s_6_2_1_U8.top_sub_6ns_6s_6_2_1_Adder_4_U.bin_s1 ;
assign \sub_6ns_6s_6_2_1_U8.top_sub_6ns_6s_6_2_1_Adder_4_U.u2.cin  = \sub_6ns_6s_6_2_1_U8.top_sub_6ns_6s_6_2_1_Adder_4_U.carry_s1 ;
assign \sub_6ns_6s_6_2_1_U8.top_sub_6ns_6s_6_2_1_Adder_4_U.facout_s2  = \sub_6ns_6s_6_2_1_U8.top_sub_6ns_6s_6_2_1_Adder_4_U.u2.cout ;
assign \sub_6ns_6s_6_2_1_U8.top_sub_6ns_6s_6_2_1_Adder_4_U.fas_s2  = \sub_6ns_6s_6_2_1_U8.top_sub_6ns_6s_6_2_1_Adder_4_U.u2.s ;
assign \sub_6ns_6s_6_2_1_U8.top_sub_6ns_6s_6_2_1_Adder_4_U.u1.a  = \sub_6ns_6s_6_2_1_U8.top_sub_6ns_6s_6_2_1_Adder_4_U.a [2:0];
assign \sub_6ns_6s_6_2_1_U8.top_sub_6ns_6s_6_2_1_Adder_4_U.u1.b  = \sub_6ns_6s_6_2_1_U8.top_sub_6ns_6s_6_2_1_Adder_4_U.bin_s0 [2:0];
assign \sub_6ns_6s_6_2_1_U8.top_sub_6ns_6s_6_2_1_Adder_4_U.u1.cin  = 1'h1;
assign \sub_6ns_6s_6_2_1_U8.top_sub_6ns_6s_6_2_1_Adder_4_U.facout_s1  = \sub_6ns_6s_6_2_1_U8.top_sub_6ns_6s_6_2_1_Adder_4_U.u1.cout ;
assign \sub_6ns_6s_6_2_1_U8.top_sub_6ns_6s_6_2_1_Adder_4_U.fas_s1  = \sub_6ns_6s_6_2_1_U8.top_sub_6ns_6s_6_2_1_Adder_4_U.u1.s ;
assign \sub_6ns_6s_6_2_1_U8.top_sub_6ns_6s_6_2_1_Adder_4_U.a  = \sub_6ns_6s_6_2_1_U8.din0 ;
assign \sub_6ns_6s_6_2_1_U8.top_sub_6ns_6s_6_2_1_Adder_4_U.b  = \sub_6ns_6s_6_2_1_U8.din1 ;
assign \sub_6ns_6s_6_2_1_U8.top_sub_6ns_6s_6_2_1_Adder_4_U.ce  = \sub_6ns_6s_6_2_1_U8.ce ;
assign \sub_6ns_6s_6_2_1_U8.top_sub_6ns_6s_6_2_1_Adder_4_U.clk  = \sub_6ns_6s_6_2_1_U8.clk ;
assign \sub_6ns_6s_6_2_1_U8.top_sub_6ns_6s_6_2_1_Adder_4_U.reset  = \sub_6ns_6s_6_2_1_U8.reset ;
assign \sub_6ns_6s_6_2_1_U8.dout  = \sub_6ns_6s_6_2_1_U8.top_sub_6ns_6s_6_2_1_Adder_4_U.s ;
assign \sub_6ns_6s_6_2_1_U8.ce  = 1'h1;
assign \sub_6ns_6s_6_2_1_U8.clk  = ap_clk;
assign \sub_6ns_6s_6_2_1_U8.din0  = 6'h00;
assign \sub_6ns_6s_6_2_1_U8.din1  = { ret_V_20_reg_1141[4], ret_V_20_reg_1141 };
assign grp_fu_420_p2 = \sub_6ns_6s_6_2_1_U8.dout ;
assign \sub_6ns_6s_6_2_1_U8.reset  = ap_rst;
assign \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.ain_s0  = \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.a ;
assign \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.s  = { \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.fas_s2 , \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.sum_s1  };
assign \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.u2.a  = \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.ain_s1 ;
assign \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.u2.b  = \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.bin_s1 ;
assign \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.u2.cin  = \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.carry_s1 ;
assign \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.facout_s2  = \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.u2.cout ;
assign \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.fas_s2  = \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.u2.s ;
assign \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.u1.a  = \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.a [1:0];
assign \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.u1.b  = \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.bin_s0 [1:0];
assign \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.u1.cin  = 1'h1;
assign \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.facout_s1  = \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.u1.cout ;
assign \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.fas_s1  = \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.u1.s ;
assign \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.a  = \sub_4ns_4ns_4_2_1_U1.din0 ;
assign \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.b  = \sub_4ns_4ns_4_2_1_U1.din1 ;
assign \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.ce  = \sub_4ns_4ns_4_2_1_U1.ce ;
assign \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.clk  = \sub_4ns_4ns_4_2_1_U1.clk ;
assign \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.reset  = \sub_4ns_4ns_4_2_1_U1.reset ;
assign \sub_4ns_4ns_4_2_1_U1.dout  = \sub_4ns_4ns_4_2_1_U1.top_sub_4ns_4ns_4_2_1_Adder_0_U.s ;
assign \sub_4ns_4ns_4_2_1_U1.ce  = 1'h1;
assign \sub_4ns_4ns_4_2_1_U1.clk  = ap_clk;
assign \sub_4ns_4ns_4_2_1_U1.din0  = 4'h0;
assign \sub_4ns_4ns_4_2_1_U1.din1  = op_5;
assign grp_fu_247_p2 = \sub_4ns_4ns_4_2_1_U1.dout ;
assign \sub_4ns_4ns_4_2_1_U1.reset  = ap_rst;
assign \shl_8ns_8s_8_7_1_U10.din1_cast  = \shl_8ns_8s_8_7_1_U10.din1 ;
assign \shl_8ns_8s_8_7_1_U10.din1_mask  = 8'h03;
assign \shl_8ns_8s_8_7_1_U10.ce  = 1'h1;
assign \shl_8ns_8s_8_7_1_U10.clk  = ap_clk;
assign \shl_8ns_8s_8_7_1_U10.din0  = op_3;
assign \shl_8ns_8s_8_7_1_U10.din1  = { sh_V_1_reg_1172[5], sh_V_1_reg_1172[5], sh_V_1_reg_1172 };
assign grp_fu_485_p2 = \shl_8ns_8s_8_7_1_U10.dout ;
assign \shl_8ns_8s_8_7_1_U10.reset  = ap_rst;
assign \shl_16s_4ns_16_7_1_U3.din1_cast  = \shl_16s_4ns_16_7_1_U3.din1 [3:0];
assign \shl_16s_4ns_16_7_1_U3.din1_mask  = 4'h1;
assign \shl_16s_4ns_16_7_1_U3.ce  = 1'h1;
assign \shl_16s_4ns_16_7_1_U3.clk  = ap_clk;
assign \shl_16s_4ns_16_7_1_U3.din0  = op_4;
assign \shl_16s_4ns_16_7_1_U3.din1  = { 12'h000, ush_reg_1054 };
assign grp_fu_316_p2 = \shl_16s_4ns_16_7_1_U3.dout ;
assign \shl_16s_4ns_16_7_1_U3.reset  = ap_rst;
assign \mul_16s_2s_18_7_1_U5.top_mul_16s_2s_18_7_1_Mul_DSP_0_U.p  = \mul_16s_2s_18_7_1_U5.top_mul_16s_2s_18_7_1_Mul_DSP_0_U.buff4 ;
assign \mul_16s_2s_18_7_1_U5.top_mul_16s_2s_18_7_1_Mul_DSP_0_U.a  = \mul_16s_2s_18_7_1_U5.din0 ;
assign \mul_16s_2s_18_7_1_U5.top_mul_16s_2s_18_7_1_Mul_DSP_0_U.b  = \mul_16s_2s_18_7_1_U5.din1 ;
assign \mul_16s_2s_18_7_1_U5.top_mul_16s_2s_18_7_1_Mul_DSP_0_U.ce  = \mul_16s_2s_18_7_1_U5.ce ;
assign \mul_16s_2s_18_7_1_U5.top_mul_16s_2s_18_7_1_Mul_DSP_0_U.clk  = \mul_16s_2s_18_7_1_U5.clk ;
assign \mul_16s_2s_18_7_1_U5.dout  = \mul_16s_2s_18_7_1_U5.top_mul_16s_2s_18_7_1_Mul_DSP_0_U.p ;
assign \mul_16s_2s_18_7_1_U5.ce  = 1'h1;
assign \mul_16s_2s_18_7_1_U5.clk  = ap_clk;
assign \mul_16s_2s_18_7_1_U5.din0  = op_4;
assign \mul_16s_2s_18_7_1_U5.din1  = op_7;
assign grp_fu_336_p2 = \mul_16s_2s_18_7_1_U5.dout ;
assign \mul_16s_2s_18_7_1_U5.reset  = ap_rst;
assign \ashr_8ns_8s_8_7_1_U11.din1_cast  = \ashr_8ns_8s_8_7_1_U11.din1 ;
assign \ashr_8ns_8s_8_7_1_U11.din1_mask  = 8'h03;
assign \ashr_8ns_8s_8_7_1_U11.ce  = 1'h1;
assign \ashr_8ns_8s_8_7_1_U11.clk  = ap_clk;
assign \ashr_8ns_8s_8_7_1_U11.din0  = op_3;
assign \ashr_8ns_8s_8_7_1_U11.din1  = { ret_V_20_reg_1141[4], ret_V_20_reg_1141[4], ret_V_20_reg_1141[4], ret_V_20_reg_1141 };
assign grp_fu_493_p2 = \ashr_8ns_8s_8_7_1_U11.dout ;
assign \ashr_8ns_8s_8_7_1_U11.reset  = ap_rst;
assign \ashr_16s_4ns_16_7_1_U4.din1_cast  = \ashr_16s_4ns_16_7_1_U4.din1 [3:0];
assign \ashr_16s_4ns_16_7_1_U4.din1_mask  = 4'h1;
assign \ashr_16s_4ns_16_7_1_U4.ce  = 1'h1;
assign \ashr_16s_4ns_16_7_1_U4.clk  = ap_clk;
assign \ashr_16s_4ns_16_7_1_U4.din0  = op_4;
assign \ashr_16s_4ns_16_7_1_U4.din1  = { 12'h000, ush_reg_1054 };
assign grp_fu_322_p2 = \ashr_16s_4ns_16_7_1_U4.dout ;
assign \ashr_16s_4ns_16_7_1_U4.reset  = ap_rst;
assign \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_13_U.ain_s0  = \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_13_U.a ;
assign \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_13_U.bin_s0  = \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_13_U.b ;
assign \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_13_U.s  = { \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_13_U.fas_s2 , \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_13_U.sum_s1  };
assign \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_13_U.u2.a  = \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_13_U.ain_s1 ;
assign \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_13_U.u2.b  = \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_13_U.bin_s1 ;
assign \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_13_U.u2.cin  = \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_13_U.carry_s1 ;
assign \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_13_U.facout_s2  = \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_13_U.u2.cout ;
assign \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_13_U.fas_s2  = \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_13_U.u2.s ;
assign \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_13_U.u1.a  = \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_13_U.a [3:0];
assign \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_13_U.u1.b  = \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_13_U.b [3:0];
assign \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_13_U.u1.cin  = 1'h0;
assign \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_13_U.facout_s1  = \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_13_U.u1.cout ;
assign \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_13_U.fas_s1  = \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_13_U.u1.s ;
assign \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_13_U.a  = \add_9s_9ns_9_2_1_U19.din0 ;
assign \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_13_U.b  = \add_9s_9ns_9_2_1_U19.din1 ;
assign \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_13_U.ce  = \add_9s_9ns_9_2_1_U19.ce ;
assign \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_13_U.clk  = \add_9s_9ns_9_2_1_U19.clk ;
assign \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_13_U.reset  = \add_9s_9ns_9_2_1_U19.reset ;
assign \add_9s_9ns_9_2_1_U19.dout  = \add_9s_9ns_9_2_1_U19.top_add_9s_9ns_9_2_1_Adder_13_U.s ;
assign \add_9s_9ns_9_2_1_U19.ce  = 1'h1;
assign \add_9s_9ns_9_2_1_U19.clk  = ap_clk;
assign \add_9s_9ns_9_2_1_U19.din0  = { tmp_reg_1437[7], tmp_reg_1437 };
assign \add_9s_9ns_9_2_1_U19.din1  = 9'h001;
assign grp_fu_843_p2 = \add_9s_9ns_9_2_1_U19.dout ;
assign \add_9s_9ns_9_2_1_U19.reset  = ap_rst;
assign \add_9ns_9s_9_2_1_U9.top_add_9ns_9s_9_2_1_Adder_5_U.ain_s0  = \add_9ns_9s_9_2_1_U9.top_add_9ns_9s_9_2_1_Adder_5_U.a ;
assign \add_9ns_9s_9_2_1_U9.top_add_9ns_9s_9_2_1_Adder_5_U.bin_s0  = \add_9ns_9s_9_2_1_U9.top_add_9ns_9s_9_2_1_Adder_5_U.b ;
assign \add_9ns_9s_9_2_1_U9.top_add_9ns_9s_9_2_1_Adder_5_U.s  = { \add_9ns_9s_9_2_1_U9.top_add_9ns_9s_9_2_1_Adder_5_U.fas_s2 , \add_9ns_9s_9_2_1_U9.top_add_9ns_9s_9_2_1_Adder_5_U.sum_s1  };
assign \add_9ns_9s_9_2_1_U9.top_add_9ns_9s_9_2_1_Adder_5_U.u2.a  = \add_9ns_9s_9_2_1_U9.top_add_9ns_9s_9_2_1_Adder_5_U.ain_s1 ;
assign \add_9ns_9s_9_2_1_U9.top_add_9ns_9s_9_2_1_Adder_5_U.u2.b  = \add_9ns_9s_9_2_1_U9.top_add_9ns_9s_9_2_1_Adder_5_U.bin_s1 ;
assign \add_9ns_9s_9_2_1_U9.top_add_9ns_9s_9_2_1_Adder_5_U.u2.cin  = \add_9ns_9s_9_2_1_U9.top_add_9ns_9s_9_2_1_Adder_5_U.carry_s1 ;
assign \add_9ns_9s_9_2_1_U9.top_add_9ns_9s_9_2_1_Adder_5_U.facout_s2  = \add_9ns_9s_9_2_1_U9.top_add_9ns_9s_9_2_1_Adder_5_U.u2.cout ;
assign \add_9ns_9s_9_2_1_U9.top_add_9ns_9s_9_2_1_Adder_5_U.fas_s2  = \add_9ns_9s_9_2_1_U9.top_add_9ns_9s_9_2_1_Adder_5_U.u2.s ;
assign \add_9ns_9s_9_2_1_U9.top_add_9ns_9s_9_2_1_Adder_5_U.u1.a  = \add_9ns_9s_9_2_1_U9.top_add_9ns_9s_9_2_1_Adder_5_U.a [3:0];
assign \add_9ns_9s_9_2_1_U9.top_add_9ns_9s_9_2_1_Adder_5_U.u1.b  = \add_9ns_9s_9_2_1_U9.top_add_9ns_9s_9_2_1_Adder_5_U.b [3:0];
assign \add_9ns_9s_9_2_1_U9.top_add_9ns_9s_9_2_1_Adder_5_U.u1.cin  = 1'h0;
assign \add_9ns_9s_9_2_1_U9.top_add_9ns_9s_9_2_1_Adder_5_U.facout_s1  = \add_9ns_9s_9_2_1_U9.top_add_9ns_9s_9_2_1_Adder_5_U.u1.cout ;
assign \add_9ns_9s_9_2_1_U9.top_add_9ns_9s_9_2_1_Adder_5_U.fas_s1  = \add_9ns_9s_9_2_1_U9.top_add_9ns_9s_9_2_1_Adder_5_U.u1.s ;
assign \add_9ns_9s_9_2_1_U9.top_add_9ns_9s_9_2_1_Adder_5_U.a  = \add_9ns_9s_9_2_1_U9.din0 ;
assign \add_9ns_9s_9_2_1_U9.top_add_9ns_9s_9_2_1_Adder_5_U.b  = \add_9ns_9s_9_2_1_U9.din1 ;
assign \add_9ns_9s_9_2_1_U9.top_add_9ns_9s_9_2_1_Adder_5_U.ce  = \add_9ns_9s_9_2_1_U9.ce ;
assign \add_9ns_9s_9_2_1_U9.top_add_9ns_9s_9_2_1_Adder_5_U.clk  = \add_9ns_9s_9_2_1_U9.clk ;
assign \add_9ns_9s_9_2_1_U9.top_add_9ns_9s_9_2_1_Adder_5_U.reset  = \add_9ns_9s_9_2_1_U9.reset ;
assign \add_9ns_9s_9_2_1_U9.dout  = \add_9ns_9s_9_2_1_U9.top_add_9ns_9s_9_2_1_Adder_5_U.s ;
assign \add_9ns_9s_9_2_1_U9.ce  = 1'h1;
assign \add_9ns_9s_9_2_1_U9.clk  = ap_clk;
assign \add_9ns_9s_9_2_1_U9.din0  = { 4'h0, op_0, 3'h0 };
assign \add_9ns_9s_9_2_1_U9.din1  = { op_1[7], op_1 };
assign grp_fu_442_p2 = \add_9ns_9s_9_2_1_U9.dout ;
assign \add_9ns_9s_9_2_1_U9.reset  = ap_rst;
assign \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_8_U.ain_s0  = \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_8_U.a ;
assign \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_8_U.bin_s0  = \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_8_U.b ;
assign \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_8_U.s  = { \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_8_U.fas_s2 , \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_8_U.sum_s1  };
assign \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_8_U.u2.a  = \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_8_U.ain_s1 ;
assign \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_8_U.u2.b  = \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_8_U.bin_s1 ;
assign \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_8_U.u2.cin  = \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_8_U.carry_s1 ;
assign \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_8_U.facout_s2  = \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_8_U.u2.cout ;
assign \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_8_U.fas_s2  = \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_8_U.u2.s ;
assign \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_8_U.u1.a  = \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_8_U.a [2:0];
assign \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_8_U.u1.b  = \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_8_U.b [2:0];
assign \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_8_U.u1.cin  = 1'h0;
assign \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_8_U.facout_s1  = \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_8_U.u1.cout ;
assign \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_8_U.fas_s1  = \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_8_U.u1.s ;
assign \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_8_U.a  = \add_7s_7ns_7_2_1_U14.din0 ;
assign \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_8_U.b  = \add_7s_7ns_7_2_1_U14.din1 ;
assign \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_8_U.ce  = \add_7s_7ns_7_2_1_U14.ce ;
assign \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_8_U.clk  = \add_7s_7ns_7_2_1_U14.clk ;
assign \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_8_U.reset  = \add_7s_7ns_7_2_1_U14.reset ;
assign \add_7s_7ns_7_2_1_U14.dout  = \add_7s_7ns_7_2_1_U14.top_add_7s_7ns_7_2_1_Adder_8_U.s ;
assign \add_7s_7ns_7_2_1_U14.ce  = 1'h1;
assign \add_7s_7ns_7_2_1_U14.clk  = ap_clk;
assign \add_7s_7ns_7_2_1_U14.din0  = { ret_V_17_reg_1287[5], ret_V_17_reg_1287 };
assign \add_7s_7ns_7_2_1_U14.din1  = { 3'h0, ret_V_18_reg_1304 };
assign grp_fu_653_p2 = \add_7s_7ns_7_2_1_U14.dout ;
assign \add_7s_7ns_7_2_1_U14.reset  = ap_rst;
assign \add_7ns_7ns_7_2_1_U16.top_add_7ns_7ns_7_2_1_Adder_10_U.ain_s0  = \add_7ns_7ns_7_2_1_U16.top_add_7ns_7ns_7_2_1_Adder_10_U.a ;
assign \add_7ns_7ns_7_2_1_U16.top_add_7ns_7ns_7_2_1_Adder_10_U.bin_s0  = \add_7ns_7ns_7_2_1_U16.top_add_7ns_7ns_7_2_1_Adder_10_U.b ;
assign \add_7ns_7ns_7_2_1_U16.top_add_7ns_7ns_7_2_1_Adder_10_U.s  = { \add_7ns_7ns_7_2_1_U16.top_add_7ns_7ns_7_2_1_Adder_10_U.fas_s2 , \add_7ns_7ns_7_2_1_U16.top_add_7ns_7ns_7_2_1_Adder_10_U.sum_s1  };
assign \add_7ns_7ns_7_2_1_U16.top_add_7ns_7ns_7_2_1_Adder_10_U.u2.a  = \add_7ns_7ns_7_2_1_U16.top_add_7ns_7ns_7_2_1_Adder_10_U.ain_s1 ;
assign \add_7ns_7ns_7_2_1_U16.top_add_7ns_7ns_7_2_1_Adder_10_U.u2.b  = \add_7ns_7ns_7_2_1_U16.top_add_7ns_7ns_7_2_1_Adder_10_U.bin_s1 ;
assign \add_7ns_7ns_7_2_1_U16.top_add_7ns_7ns_7_2_1_Adder_10_U.u2.cin  = \add_7ns_7ns_7_2_1_U16.top_add_7ns_7ns_7_2_1_Adder_10_U.carry_s1 ;
assign \add_7ns_7ns_7_2_1_U16.top_add_7ns_7ns_7_2_1_Adder_10_U.facout_s2  = \add_7ns_7ns_7_2_1_U16.top_add_7ns_7ns_7_2_1_Adder_10_U.u2.cout ;
assign \add_7ns_7ns_7_2_1_U16.top_add_7ns_7ns_7_2_1_Adder_10_U.fas_s2  = \add_7ns_7ns_7_2_1_U16.top_add_7ns_7ns_7_2_1_Adder_10_U.u2.s ;
assign \add_7ns_7ns_7_2_1_U16.top_add_7ns_7ns_7_2_1_Adder_10_U.u1.a  = \add_7ns_7ns_7_2_1_U16.top_add_7ns_7ns_7_2_1_Adder_10_U.a [2:0];
assign \add_7ns_7ns_7_2_1_U16.top_add_7ns_7ns_7_2_1_Adder_10_U.u1.b  = \add_7ns_7ns_7_2_1_U16.top_add_7ns_7ns_7_2_1_Adder_10_U.b [2:0];
assign \add_7ns_7ns_7_2_1_U16.top_add_7ns_7ns_7_2_1_Adder_10_U.u1.cin  = 1'h0;
assign \add_7ns_7ns_7_2_1_U16.top_add_7ns_7ns_7_2_1_Adder_10_U.facout_s1  = \add_7ns_7ns_7_2_1_U16.top_add_7ns_7ns_7_2_1_Adder_10_U.u1.cout ;
assign \add_7ns_7ns_7_2_1_U16.top_add_7ns_7ns_7_2_1_Adder_10_U.fas_s1  = \add_7ns_7ns_7_2_1_U16.top_add_7ns_7ns_7_2_1_Adder_10_U.u1.s ;
assign \add_7ns_7ns_7_2_1_U16.top_add_7ns_7ns_7_2_1_Adder_10_U.a  = \add_7ns_7ns_7_2_1_U16.din0 ;
assign \add_7ns_7ns_7_2_1_U16.top_add_7ns_7ns_7_2_1_Adder_10_U.b  = \add_7ns_7ns_7_2_1_U16.din1 ;
assign \add_7ns_7ns_7_2_1_U16.top_add_7ns_7ns_7_2_1_Adder_10_U.ce  = \add_7ns_7ns_7_2_1_U16.ce ;
assign \add_7ns_7ns_7_2_1_U16.top_add_7ns_7ns_7_2_1_Adder_10_U.clk  = \add_7ns_7ns_7_2_1_U16.clk ;
assign \add_7ns_7ns_7_2_1_U16.top_add_7ns_7ns_7_2_1_Adder_10_U.reset  = \add_7ns_7ns_7_2_1_U16.reset ;
assign \add_7ns_7ns_7_2_1_U16.dout  = \add_7ns_7ns_7_2_1_U16.top_add_7ns_7ns_7_2_1_Adder_10_U.s ;
assign \add_7ns_7ns_7_2_1_U16.ce  = 1'h1;
assign \add_7ns_7ns_7_2_1_U16.clk  = ap_clk;
assign \add_7ns_7ns_7_2_1_U16.din0  = { 4'h0, add_ln69_1_reg_1362 };
assign \add_7ns_7ns_7_2_1_U16.din1  = add_ln69_reg_1357;
assign grp_fu_774_p2 = \add_7ns_7ns_7_2_1_U16.dout ;
assign \add_7ns_7ns_7_2_1_U16.reset  = ap_rst;
assign \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_6_U.ain_s0  = \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_6_U.a ;
assign \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_6_U.bin_s0  = \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_6_U.b ;
assign \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_6_U.s  = { \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_6_U.fas_s2 , \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_6_U.sum_s1  };
assign \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_6_U.u2.a  = \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_6_U.ain_s1 ;
assign \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_6_U.u2.b  = \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_6_U.bin_s1 ;
assign \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_6_U.u2.cin  = \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_6_U.carry_s1 ;
assign \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_6_U.facout_s2  = \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_6_U.u2.cout ;
assign \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_6_U.fas_s2  = \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_6_U.u2.s ;
assign \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_6_U.u1.a  = \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_6_U.a [2:0];
assign \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_6_U.u1.b  = \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_6_U.b [2:0];
assign \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_6_U.u1.cin  = 1'h0;
assign \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_6_U.facout_s1  = \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_6_U.u1.cout ;
assign \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_6_U.fas_s1  = \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_6_U.u1.s ;
assign \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_6_U.a  = \add_6ns_6ns_6_2_1_U12.din0 ;
assign \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_6_U.b  = \add_6ns_6ns_6_2_1_U12.din1 ;
assign \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_6_U.ce  = \add_6ns_6ns_6_2_1_U12.ce ;
assign \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_6_U.clk  = \add_6ns_6ns_6_2_1_U12.clk ;
assign \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_6_U.reset  = \add_6ns_6ns_6_2_1_U12.reset ;
assign \add_6ns_6ns_6_2_1_U12.dout  = \add_6ns_6ns_6_2_1_U12.top_add_6ns_6ns_6_2_1_Adder_6_U.s ;
assign \add_6ns_6ns_6_2_1_U12.ce  = 1'h1;
assign \add_6ns_6ns_6_2_1_U12.clk  = ap_clk;
assign \add_6ns_6ns_6_2_1_U12.din0  = ret_V_reg_1182;
assign \add_6ns_6ns_6_2_1_U12.din1  = 6'h01;
assign grp_fu_498_p2 = \add_6ns_6ns_6_2_1_U12.dout ;
assign \add_6ns_6ns_6_2_1_U12.reset  = ap_rst;
assign \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_3_U.ain_s0  = \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_3_U.a ;
assign \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_3_U.bin_s0  = \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_3_U.b ;
assign \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_3_U.s  = { \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_3_U.fas_s2 , \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_3_U.sum_s1  };
assign \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_3_U.u2.a  = \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_3_U.ain_s1 ;
assign \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_3_U.u2.b  = \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_3_U.bin_s1 ;
assign \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_3_U.u2.cin  = \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_3_U.carry_s1 ;
assign \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_3_U.facout_s2  = \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_3_U.u2.cout ;
assign \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_3_U.fas_s2  = \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_3_U.u2.s ;
assign \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_3_U.u1.a  = \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_3_U.a [1:0];
assign \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_3_U.u1.b  = \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_3_U.b [1:0];
assign \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_3_U.u1.cin  = 1'h0;
assign \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_3_U.facout_s1  = \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_3_U.u1.cout ;
assign \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_3_U.fas_s1  = \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_3_U.u1.s ;
assign \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_3_U.a  = \add_5ns_5ns_5_2_1_U7.din0 ;
assign \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_3_U.b  = \add_5ns_5ns_5_2_1_U7.din1 ;
assign \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_3_U.ce  = \add_5ns_5ns_5_2_1_U7.ce ;
assign \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_3_U.clk  = \add_5ns_5ns_5_2_1_U7.clk ;
assign \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_3_U.reset  = \add_5ns_5ns_5_2_1_U7.reset ;
assign \add_5ns_5ns_5_2_1_U7.dout  = \add_5ns_5ns_5_2_1_U7.top_add_5ns_5ns_5_2_1_Adder_3_U.s ;
assign \add_5ns_5ns_5_2_1_U7.ce  = 1'h1;
assign \add_5ns_5ns_5_2_1_U7.clk  = ap_clk;
assign \add_5ns_5ns_5_2_1_U7.din0  = ret_V_7_reg_1119;
assign \add_5ns_5ns_5_2_1_U7.din1  = 5'h01;
assign grp_fu_381_p2 = \add_5ns_5ns_5_2_1_U7.dout ;
assign \add_5ns_5ns_5_2_1_U7.reset  = ap_rst;
assign \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_7_U.ain_s0  = \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_7_U.a ;
assign \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_7_U.bin_s0  = \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_7_U.b ;
assign \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_7_U.s  = { \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_7_U.fas_s2 , \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_7_U.sum_s1  };
assign \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_7_U.u2.a  = \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_7_U.ain_s1 ;
assign \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_7_U.u2.b  = \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_7_U.bin_s1 ;
assign \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_7_U.u2.cin  = \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_7_U.carry_s1 ;
assign \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_7_U.facout_s2  = \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_7_U.u2.cout ;
assign \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_7_U.fas_s2  = \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_7_U.u2.s ;
assign \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_7_U.u1.a  = \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_7_U.a [1:0];
assign \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_7_U.u1.b  = \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_7_U.b [1:0];
assign \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_7_U.u1.cin  = 1'h0;
assign \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_7_U.facout_s1  = \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_7_U.u1.cout ;
assign \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_7_U.fas_s1  = \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_7_U.u1.s ;
assign \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_7_U.a  = \add_4ns_4ns_4_2_1_U13.din0 ;
assign \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_7_U.b  = \add_4ns_4ns_4_2_1_U13.din1 ;
assign \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_7_U.ce  = \add_4ns_4ns_4_2_1_U13.ce ;
assign \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_7_U.clk  = \add_4ns_4ns_4_2_1_U13.clk ;
assign \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_7_U.reset  = \add_4ns_4ns_4_2_1_U13.reset ;
assign \add_4ns_4ns_4_2_1_U13.dout  = \add_4ns_4ns_4_2_1_U13.top_add_4ns_4ns_4_2_1_Adder_7_U.s ;
assign \add_4ns_4ns_4_2_1_U13.ce  = 1'h1;
assign \add_4ns_4ns_4_2_1_U13.clk  = ap_clk;
assign \add_4ns_4ns_4_2_1_U13.din0  = ret_V_3_cast_reg_1204;
assign \add_4ns_4ns_4_2_1_U13.din1  = 4'h1;
assign grp_fu_549_p2 = \add_4ns_4ns_4_2_1_U13.dout ;
assign \add_4ns_4ns_4_2_1_U13.reset  = ap_rst;
assign \add_40s_40s_40_2_1_U20.top_add_40s_40s_40_2_1_Adder_14_U.ain_s0  = \add_40s_40s_40_2_1_U20.top_add_40s_40s_40_2_1_Adder_14_U.a ;
assign \add_40s_40s_40_2_1_U20.top_add_40s_40s_40_2_1_Adder_14_U.bin_s0  = \add_40s_40s_40_2_1_U20.top_add_40s_40s_40_2_1_Adder_14_U.b ;
assign \add_40s_40s_40_2_1_U20.top_add_40s_40s_40_2_1_Adder_14_U.s  = { \add_40s_40s_40_2_1_U20.top_add_40s_40s_40_2_1_Adder_14_U.fas_s2 , \add_40s_40s_40_2_1_U20.top_add_40s_40s_40_2_1_Adder_14_U.sum_s1  };
assign \add_40s_40s_40_2_1_U20.top_add_40s_40s_40_2_1_Adder_14_U.u2.a  = \add_40s_40s_40_2_1_U20.top_add_40s_40s_40_2_1_Adder_14_U.ain_s1 ;
assign \add_40s_40s_40_2_1_U20.top_add_40s_40s_40_2_1_Adder_14_U.u2.b  = \add_40s_40s_40_2_1_U20.top_add_40s_40s_40_2_1_Adder_14_U.bin_s1 ;
assign \add_40s_40s_40_2_1_U20.top_add_40s_40s_40_2_1_Adder_14_U.u2.cin  = \add_40s_40s_40_2_1_U20.top_add_40s_40s_40_2_1_Adder_14_U.carry_s1 ;
assign \add_40s_40s_40_2_1_U20.top_add_40s_40s_40_2_1_Adder_14_U.facout_s2  = \add_40s_40s_40_2_1_U20.top_add_40s_40s_40_2_1_Adder_14_U.u2.cout ;
assign \add_40s_40s_40_2_1_U20.top_add_40s_40s_40_2_1_Adder_14_U.fas_s2  = \add_40s_40s_40_2_1_U20.top_add_40s_40s_40_2_1_Adder_14_U.u2.s ;
assign \add_40s_40s_40_2_1_U20.top_add_40s_40s_40_2_1_Adder_14_U.u1.a  = \add_40s_40s_40_2_1_U20.top_add_40s_40s_40_2_1_Adder_14_U.a [19:0];
assign \add_40s_40s_40_2_1_U20.top_add_40s_40s_40_2_1_Adder_14_U.u1.b  = \add_40s_40s_40_2_1_U20.top_add_40s_40s_40_2_1_Adder_14_U.b [19:0];
assign \add_40s_40s_40_2_1_U20.top_add_40s_40s_40_2_1_Adder_14_U.u1.cin  = 1'h0;
assign \add_40s_40s_40_2_1_U20.top_add_40s_40s_40_2_1_Adder_14_U.facout_s1  = \add_40s_40s_40_2_1_U20.top_add_40s_40s_40_2_1_Adder_14_U.u1.cout ;
assign \add_40s_40s_40_2_1_U20.top_add_40s_40s_40_2_1_Adder_14_U.fas_s1  = \add_40s_40s_40_2_1_U20.top_add_40s_40s_40_2_1_Adder_14_U.u1.s ;
assign \add_40s_40s_40_2_1_U20.top_add_40s_40s_40_2_1_Adder_14_U.a  = \add_40s_40s_40_2_1_U20.din0 ;
assign \add_40s_40s_40_2_1_U20.top_add_40s_40s_40_2_1_Adder_14_U.b  = \add_40s_40s_40_2_1_U20.din1 ;
assign \add_40s_40s_40_2_1_U20.top_add_40s_40s_40_2_1_Adder_14_U.ce  = \add_40s_40s_40_2_1_U20.ce ;
assign \add_40s_40s_40_2_1_U20.top_add_40s_40s_40_2_1_Adder_14_U.clk  = \add_40s_40s_40_2_1_U20.clk ;
assign \add_40s_40s_40_2_1_U20.top_add_40s_40s_40_2_1_Adder_14_U.reset  = \add_40s_40s_40_2_1_U20.reset ;
assign \add_40s_40s_40_2_1_U20.dout  = \add_40s_40s_40_2_1_U20.top_add_40s_40s_40_2_1_Adder_14_U.s ;
assign \add_40s_40s_40_2_1_U20.ce  = 1'h1;
assign \add_40s_40s_40_2_1_U20.clk  = ap_clk;
assign \add_40s_40s_40_2_1_U20.din0  = { select_ln353_reg_1459[8], select_ln353_reg_1459[8], select_ln353_reg_1459[8], select_ln353_reg_1459[8], select_ln353_reg_1459[8], select_ln353_reg_1459[8], select_ln353_reg_1459[8], select_ln353_reg_1459[8], select_ln353_reg_1459[8], select_ln353_reg_1459[8], select_ln353_reg_1459[8], select_ln353_reg_1459[8], select_ln353_reg_1459[8], select_ln353_reg_1459[8], select_ln353_reg_1459[8], select_ln353_reg_1459[8], select_ln353_reg_1459[8], select_ln353_reg_1459[8], select_ln353_reg_1459[8], select_ln353_reg_1459[8], select_ln353_reg_1459[8], select_ln353_reg_1459[8], select_ln353_reg_1459[8], select_ln353_reg_1459[8], select_ln353_reg_1459, 7'h00 };
assign \add_40s_40s_40_2_1_U20.din1  = { op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13 };
assign grp_fu_883_p2 = \add_40s_40s_40_2_1_U20.dout ;
assign \add_40s_40s_40_2_1_U20.reset  = ap_rst;
assign \add_3s_3s_3_2_1_U6.top_add_3s_3s_3_2_1_Adder_2_U.ain_s0  = \add_3s_3s_3_2_1_U6.top_add_3s_3s_3_2_1_Adder_2_U.a ;
assign \add_3s_3s_3_2_1_U6.top_add_3s_3s_3_2_1_Adder_2_U.bin_s0  = \add_3s_3s_3_2_1_U6.top_add_3s_3s_3_2_1_Adder_2_U.b ;
assign \add_3s_3s_3_2_1_U6.top_add_3s_3s_3_2_1_Adder_2_U.s  = { \add_3s_3s_3_2_1_U6.top_add_3s_3s_3_2_1_Adder_2_U.fas_s2 , \add_3s_3s_3_2_1_U6.top_add_3s_3s_3_2_1_Adder_2_U.sum_s1  };
assign \add_3s_3s_3_2_1_U6.top_add_3s_3s_3_2_1_Adder_2_U.u2.a  = \add_3s_3s_3_2_1_U6.top_add_3s_3s_3_2_1_Adder_2_U.ain_s1 ;
assign \add_3s_3s_3_2_1_U6.top_add_3s_3s_3_2_1_Adder_2_U.u2.b  = \add_3s_3s_3_2_1_U6.top_add_3s_3s_3_2_1_Adder_2_U.bin_s1 ;
assign \add_3s_3s_3_2_1_U6.top_add_3s_3s_3_2_1_Adder_2_U.u2.cin  = \add_3s_3s_3_2_1_U6.top_add_3s_3s_3_2_1_Adder_2_U.carry_s1 ;
assign \add_3s_3s_3_2_1_U6.top_add_3s_3s_3_2_1_Adder_2_U.facout_s2  = \add_3s_3s_3_2_1_U6.top_add_3s_3s_3_2_1_Adder_2_U.u2.cout ;
assign \add_3s_3s_3_2_1_U6.top_add_3s_3s_3_2_1_Adder_2_U.fas_s2  = \add_3s_3s_3_2_1_U6.top_add_3s_3s_3_2_1_Adder_2_U.u2.s ;
assign \add_3s_3s_3_2_1_U6.top_add_3s_3s_3_2_1_Adder_2_U.u1.a  = \add_3s_3s_3_2_1_U6.top_add_3s_3s_3_2_1_Adder_2_U.a [0];
assign \add_3s_3s_3_2_1_U6.top_add_3s_3s_3_2_1_Adder_2_U.u1.b  = \add_3s_3s_3_2_1_U6.top_add_3s_3s_3_2_1_Adder_2_U.b [0];
assign \add_3s_3s_3_2_1_U6.top_add_3s_3s_3_2_1_Adder_2_U.u1.cin  = 1'h0;
assign \add_3s_3s_3_2_1_U6.top_add_3s_3s_3_2_1_Adder_2_U.facout_s1  = \add_3s_3s_3_2_1_U6.top_add_3s_3s_3_2_1_Adder_2_U.u1.cout ;
assign \add_3s_3s_3_2_1_U6.top_add_3s_3s_3_2_1_Adder_2_U.fas_s1  = \add_3s_3s_3_2_1_U6.top_add_3s_3s_3_2_1_Adder_2_U.u1.s ;
assign \add_3s_3s_3_2_1_U6.top_add_3s_3s_3_2_1_Adder_2_U.a  = \add_3s_3s_3_2_1_U6.din0 ;
assign \add_3s_3s_3_2_1_U6.top_add_3s_3s_3_2_1_Adder_2_U.b  = \add_3s_3s_3_2_1_U6.din1 ;
assign \add_3s_3s_3_2_1_U6.top_add_3s_3s_3_2_1_Adder_2_U.ce  = \add_3s_3s_3_2_1_U6.ce ;
assign \add_3s_3s_3_2_1_U6.top_add_3s_3s_3_2_1_Adder_2_U.clk  = \add_3s_3s_3_2_1_U6.clk ;
assign \add_3s_3s_3_2_1_U6.top_add_3s_3s_3_2_1_Adder_2_U.reset  = \add_3s_3s_3_2_1_U6.reset ;
assign \add_3s_3s_3_2_1_U6.dout  = \add_3s_3s_3_2_1_U6.top_add_3s_3s_3_2_1_Adder_2_U.s ;
assign \add_3s_3s_3_2_1_U6.ce  = 1'h1;
assign \add_3s_3s_3_2_1_U6.clk  = ap_clk;
assign \add_3s_3s_3_2_1_U6.din0  = { op_8[1], op_8 };
assign \add_3s_3s_3_2_1_U6.din1  = { op_7[1], op_7 };
assign grp_fu_349_p2 = \add_3s_3s_3_2_1_U6.dout ;
assign \add_3s_3s_3_2_1_U6.reset  = ap_rst;
assign \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_9_U.ain_s0  = \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_9_U.a ;
assign \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_9_U.bin_s0  = \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_9_U.b ;
assign \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_9_U.s  = { \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_9_U.fas_s2 , \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_9_U.sum_s1  };
assign \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_9_U.u2.a  = \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_9_U.ain_s1 ;
assign \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_9_U.u2.b  = \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_9_U.bin_s1 ;
assign \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_9_U.u2.cin  = \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_9_U.carry_s1 ;
assign \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_9_U.facout_s2  = \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_9_U.u2.cout ;
assign \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_9_U.fas_s2  = \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_9_U.u2.s ;
assign \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_9_U.u1.a  = \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_9_U.a [0];
assign \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_9_U.u1.b  = \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_9_U.b [0];
assign \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_9_U.u1.cin  = 1'h0;
assign \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_9_U.facout_s1  = \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_9_U.u1.cout ;
assign \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_9_U.fas_s1  = \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_9_U.u1.s ;
assign \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_9_U.a  = \add_3ns_3ns_3_2_1_U15.din0 ;
assign \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_9_U.b  = \add_3ns_3ns_3_2_1_U15.din1 ;
assign \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_9_U.ce  = \add_3ns_3ns_3_2_1_U15.ce ;
assign \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_9_U.clk  = \add_3ns_3ns_3_2_1_U15.clk ;
assign \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_9_U.reset  = \add_3ns_3ns_3_2_1_U15.reset ;
assign \add_3ns_3ns_3_2_1_U15.dout  = \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_9_U.s ;
assign \add_3ns_3ns_3_2_1_U15.ce  = 1'h1;
assign \add_3ns_3ns_3_2_1_U15.clk  = ap_clk;
assign \add_3ns_3ns_3_2_1_U15.din0  = { 1'h0, op_2 };
assign \add_3ns_3ns_3_2_1_U15.din1  = { 2'h0, icmp_ln1494_reg_1131 };
assign grp_fu_659_p2 = \add_3ns_3ns_3_2_1_U15.dout ;
assign \add_3ns_3ns_3_2_1_U15.reset  = ap_rst;
assign \add_38s_38s_38_2_1_U22.top_add_38s_38s_38_2_1_Adder_16_U.ain_s0  = \add_38s_38s_38_2_1_U22.top_add_38s_38s_38_2_1_Adder_16_U.a ;
assign \add_38s_38s_38_2_1_U22.top_add_38s_38s_38_2_1_Adder_16_U.bin_s0  = \add_38s_38s_38_2_1_U22.top_add_38s_38s_38_2_1_Adder_16_U.b ;
assign \add_38s_38s_38_2_1_U22.top_add_38s_38s_38_2_1_Adder_16_U.s  = { \add_38s_38s_38_2_1_U22.top_add_38s_38s_38_2_1_Adder_16_U.fas_s2 , \add_38s_38s_38_2_1_U22.top_add_38s_38s_38_2_1_Adder_16_U.sum_s1  };
assign \add_38s_38s_38_2_1_U22.top_add_38s_38s_38_2_1_Adder_16_U.u2.a  = \add_38s_38s_38_2_1_U22.top_add_38s_38s_38_2_1_Adder_16_U.ain_s1 ;
assign \add_38s_38s_38_2_1_U22.top_add_38s_38s_38_2_1_Adder_16_U.u2.b  = \add_38s_38s_38_2_1_U22.top_add_38s_38s_38_2_1_Adder_16_U.bin_s1 ;
assign \add_38s_38s_38_2_1_U22.top_add_38s_38s_38_2_1_Adder_16_U.u2.cin  = \add_38s_38s_38_2_1_U22.top_add_38s_38s_38_2_1_Adder_16_U.carry_s1 ;
assign \add_38s_38s_38_2_1_U22.top_add_38s_38s_38_2_1_Adder_16_U.facout_s2  = \add_38s_38s_38_2_1_U22.top_add_38s_38s_38_2_1_Adder_16_U.u2.cout ;
assign \add_38s_38s_38_2_1_U22.top_add_38s_38s_38_2_1_Adder_16_U.fas_s2  = \add_38s_38s_38_2_1_U22.top_add_38s_38s_38_2_1_Adder_16_U.u2.s ;
assign \add_38s_38s_38_2_1_U22.top_add_38s_38s_38_2_1_Adder_16_U.u1.a  = \add_38s_38s_38_2_1_U22.top_add_38s_38s_38_2_1_Adder_16_U.a [18:0];
assign \add_38s_38s_38_2_1_U22.top_add_38s_38s_38_2_1_Adder_16_U.u1.b  = \add_38s_38s_38_2_1_U22.top_add_38s_38s_38_2_1_Adder_16_U.b [18:0];
assign \add_38s_38s_38_2_1_U22.top_add_38s_38s_38_2_1_Adder_16_U.u1.cin  = 1'h0;
assign \add_38s_38s_38_2_1_U22.top_add_38s_38s_38_2_1_Adder_16_U.facout_s1  = \add_38s_38s_38_2_1_U22.top_add_38s_38s_38_2_1_Adder_16_U.u1.cout ;
assign \add_38s_38s_38_2_1_U22.top_add_38s_38s_38_2_1_Adder_16_U.fas_s1  = \add_38s_38s_38_2_1_U22.top_add_38s_38s_38_2_1_Adder_16_U.u1.s ;
assign \add_38s_38s_38_2_1_U22.top_add_38s_38s_38_2_1_Adder_16_U.a  = \add_38s_38s_38_2_1_U22.din0 ;
assign \add_38s_38s_38_2_1_U22.top_add_38s_38s_38_2_1_Adder_16_U.b  = \add_38s_38s_38_2_1_U22.din1 ;
assign \add_38s_38s_38_2_1_U22.top_add_38s_38s_38_2_1_Adder_16_U.ce  = \add_38s_38s_38_2_1_U22.ce ;
assign \add_38s_38s_38_2_1_U22.top_add_38s_38s_38_2_1_Adder_16_U.clk  = \add_38s_38s_38_2_1_U22.clk ;
assign \add_38s_38s_38_2_1_U22.top_add_38s_38s_38_2_1_Adder_16_U.reset  = \add_38s_38s_38_2_1_U22.reset ;
assign \add_38s_38s_38_2_1_U22.dout  = \add_38s_38s_38_2_1_U22.top_add_38s_38s_38_2_1_Adder_16_U.s ;
assign \add_38s_38s_38_2_1_U22.ce  = 1'h1;
assign \add_38s_38s_38_2_1_U22.clk  = ap_clk;
assign \add_38s_38s_38_2_1_U22.din0  = { select_ln353_1_reg_1496[31], select_ln353_1_reg_1496, 5'h00 };
assign \add_38s_38s_38_2_1_U22.din1  = { op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15 };
assign grp_fu_948_p2 = \add_38s_38s_38_2_1_U22.dout ;
assign \add_38s_38s_38_2_1_U22.reset  = ap_rst;
assign \add_32s_32ns_32_2_1_U26.top_add_32s_32ns_32_2_1_Adder_18_U.ain_s0  = \add_32s_32ns_32_2_1_U26.top_add_32s_32ns_32_2_1_Adder_18_U.a ;
assign \add_32s_32ns_32_2_1_U26.top_add_32s_32ns_32_2_1_Adder_18_U.bin_s0  = \add_32s_32ns_32_2_1_U26.top_add_32s_32ns_32_2_1_Adder_18_U.b ;
assign \add_32s_32ns_32_2_1_U26.top_add_32s_32ns_32_2_1_Adder_18_U.s  = { \add_32s_32ns_32_2_1_U26.top_add_32s_32ns_32_2_1_Adder_18_U.fas_s2 , \add_32s_32ns_32_2_1_U26.top_add_32s_32ns_32_2_1_Adder_18_U.sum_s1  };
assign \add_32s_32ns_32_2_1_U26.top_add_32s_32ns_32_2_1_Adder_18_U.u2.a  = \add_32s_32ns_32_2_1_U26.top_add_32s_32ns_32_2_1_Adder_18_U.ain_s1 ;
assign \add_32s_32ns_32_2_1_U26.top_add_32s_32ns_32_2_1_Adder_18_U.u2.b  = \add_32s_32ns_32_2_1_U26.top_add_32s_32ns_32_2_1_Adder_18_U.bin_s1 ;
assign \add_32s_32ns_32_2_1_U26.top_add_32s_32ns_32_2_1_Adder_18_U.u2.cin  = \add_32s_32ns_32_2_1_U26.top_add_32s_32ns_32_2_1_Adder_18_U.carry_s1 ;
assign \add_32s_32ns_32_2_1_U26.top_add_32s_32ns_32_2_1_Adder_18_U.facout_s2  = \add_32s_32ns_32_2_1_U26.top_add_32s_32ns_32_2_1_Adder_18_U.u2.cout ;
assign \add_32s_32ns_32_2_1_U26.top_add_32s_32ns_32_2_1_Adder_18_U.fas_s2  = \add_32s_32ns_32_2_1_U26.top_add_32s_32ns_32_2_1_Adder_18_U.u2.s ;
assign \add_32s_32ns_32_2_1_U26.top_add_32s_32ns_32_2_1_Adder_18_U.u1.a  = \add_32s_32ns_32_2_1_U26.top_add_32s_32ns_32_2_1_Adder_18_U.a [15:0];
assign \add_32s_32ns_32_2_1_U26.top_add_32s_32ns_32_2_1_Adder_18_U.u1.b  = \add_32s_32ns_32_2_1_U26.top_add_32s_32ns_32_2_1_Adder_18_U.b [15:0];
assign \add_32s_32ns_32_2_1_U26.top_add_32s_32ns_32_2_1_Adder_18_U.u1.cin  = 1'h0;
assign \add_32s_32ns_32_2_1_U26.top_add_32s_32ns_32_2_1_Adder_18_U.facout_s1  = \add_32s_32ns_32_2_1_U26.top_add_32s_32ns_32_2_1_Adder_18_U.u1.cout ;
assign \add_32s_32ns_32_2_1_U26.top_add_32s_32ns_32_2_1_Adder_18_U.fas_s1  = \add_32s_32ns_32_2_1_U26.top_add_32s_32ns_32_2_1_Adder_18_U.u1.s ;
assign \add_32s_32ns_32_2_1_U26.top_add_32s_32ns_32_2_1_Adder_18_U.a  = \add_32s_32ns_32_2_1_U26.din0 ;
assign \add_32s_32ns_32_2_1_U26.top_add_32s_32ns_32_2_1_Adder_18_U.b  = \add_32s_32ns_32_2_1_U26.din1 ;
assign \add_32s_32ns_32_2_1_U26.top_add_32s_32ns_32_2_1_Adder_18_U.ce  = \add_32s_32ns_32_2_1_U26.ce ;
assign \add_32s_32ns_32_2_1_U26.top_add_32s_32ns_32_2_1_Adder_18_U.clk  = \add_32s_32ns_32_2_1_U26.clk ;
assign \add_32s_32ns_32_2_1_U26.top_add_32s_32ns_32_2_1_Adder_18_U.reset  = \add_32s_32ns_32_2_1_U26.reset ;
assign \add_32s_32ns_32_2_1_U26.dout  = \add_32s_32ns_32_2_1_U26.top_add_32s_32ns_32_2_1_Adder_18_U.s ;
assign \add_32s_32ns_32_2_1_U26.ce  = 1'h1;
assign \add_32s_32ns_32_2_1_U26.clk  = ap_clk;
assign \add_32s_32ns_32_2_1_U26.din0  = { add_ln69_3_reg_1442[9], add_ln69_3_reg_1442[9], add_ln69_3_reg_1442[9], add_ln69_3_reg_1442[9], add_ln69_3_reg_1442[9], add_ln69_3_reg_1442[9], add_ln69_3_reg_1442[9], add_ln69_3_reg_1442[9], add_ln69_3_reg_1442[9], add_ln69_3_reg_1442[9], add_ln69_3_reg_1442[9], add_ln69_3_reg_1442[9], add_ln69_3_reg_1442[9], add_ln69_3_reg_1442[9], add_ln69_3_reg_1442[9], add_ln69_3_reg_1442[9], add_ln69_3_reg_1442[9], add_ln69_3_reg_1442[9], add_ln69_3_reg_1442[9], add_ln69_3_reg_1442[9], add_ln69_3_reg_1442[9], add_ln69_3_reg_1442[9], add_ln69_3_reg_1442 };
assign \add_32s_32ns_32_2_1_U26.din1  = ret_V_26_reg_1553;
assign grp_fu_1019_p2 = \add_32s_32ns_32_2_1_U26.dout ;
assign \add_32s_32ns_32_2_1_U26.reset  = ap_rst;
assign \add_32ns_32s_32_2_1_U25.top_add_32ns_32s_32_2_1_Adder_17_U.ain_s0  = \add_32ns_32s_32_2_1_U25.top_add_32ns_32s_32_2_1_Adder_17_U.a ;
assign \add_32ns_32s_32_2_1_U25.top_add_32ns_32s_32_2_1_Adder_17_U.bin_s0  = \add_32ns_32s_32_2_1_U25.top_add_32ns_32s_32_2_1_Adder_17_U.b ;
assign \add_32ns_32s_32_2_1_U25.top_add_32ns_32s_32_2_1_Adder_17_U.s  = { \add_32ns_32s_32_2_1_U25.top_add_32ns_32s_32_2_1_Adder_17_U.fas_s2 , \add_32ns_32s_32_2_1_U25.top_add_32ns_32s_32_2_1_Adder_17_U.sum_s1  };
assign \add_32ns_32s_32_2_1_U25.top_add_32ns_32s_32_2_1_Adder_17_U.u2.a  = \add_32ns_32s_32_2_1_U25.top_add_32ns_32s_32_2_1_Adder_17_U.ain_s1 ;
assign \add_32ns_32s_32_2_1_U25.top_add_32ns_32s_32_2_1_Adder_17_U.u2.b  = \add_32ns_32s_32_2_1_U25.top_add_32ns_32s_32_2_1_Adder_17_U.bin_s1 ;
assign \add_32ns_32s_32_2_1_U25.top_add_32ns_32s_32_2_1_Adder_17_U.u2.cin  = \add_32ns_32s_32_2_1_U25.top_add_32ns_32s_32_2_1_Adder_17_U.carry_s1 ;
assign \add_32ns_32s_32_2_1_U25.top_add_32ns_32s_32_2_1_Adder_17_U.facout_s2  = \add_32ns_32s_32_2_1_U25.top_add_32ns_32s_32_2_1_Adder_17_U.u2.cout ;
assign \add_32ns_32s_32_2_1_U25.top_add_32ns_32s_32_2_1_Adder_17_U.fas_s2  = \add_32ns_32s_32_2_1_U25.top_add_32ns_32s_32_2_1_Adder_17_U.u2.s ;
assign \add_32ns_32s_32_2_1_U25.top_add_32ns_32s_32_2_1_Adder_17_U.u1.a  = \add_32ns_32s_32_2_1_U25.top_add_32ns_32s_32_2_1_Adder_17_U.a [15:0];
assign \add_32ns_32s_32_2_1_U25.top_add_32ns_32s_32_2_1_Adder_17_U.u1.b  = \add_32ns_32s_32_2_1_U25.top_add_32ns_32s_32_2_1_Adder_17_U.b [15:0];
assign \add_32ns_32s_32_2_1_U25.top_add_32ns_32s_32_2_1_Adder_17_U.u1.cin  = 1'h0;
assign \add_32ns_32s_32_2_1_U25.top_add_32ns_32s_32_2_1_Adder_17_U.facout_s1  = \add_32ns_32s_32_2_1_U25.top_add_32ns_32s_32_2_1_Adder_17_U.u1.cout ;
assign \add_32ns_32s_32_2_1_U25.top_add_32ns_32s_32_2_1_Adder_17_U.fas_s1  = \add_32ns_32s_32_2_1_U25.top_add_32ns_32s_32_2_1_Adder_17_U.u1.s ;
assign \add_32ns_32s_32_2_1_U25.top_add_32ns_32s_32_2_1_Adder_17_U.a  = \add_32ns_32s_32_2_1_U25.din0 ;
assign \add_32ns_32s_32_2_1_U25.top_add_32ns_32s_32_2_1_Adder_17_U.b  = \add_32ns_32s_32_2_1_U25.din1 ;
assign \add_32ns_32s_32_2_1_U25.top_add_32ns_32s_32_2_1_Adder_17_U.ce  = \add_32ns_32s_32_2_1_U25.ce ;
assign \add_32ns_32s_32_2_1_U25.top_add_32ns_32s_32_2_1_Adder_17_U.clk  = \add_32ns_32s_32_2_1_U25.clk ;
assign \add_32ns_32s_32_2_1_U25.top_add_32ns_32s_32_2_1_Adder_17_U.reset  = \add_32ns_32s_32_2_1_U25.reset ;
assign \add_32ns_32s_32_2_1_U25.dout  = \add_32ns_32s_32_2_1_U25.top_add_32ns_32s_32_2_1_Adder_17_U.s ;
assign \add_32ns_32s_32_2_1_U25.ce  = 1'h1;
assign \add_32ns_32s_32_2_1_U25.clk  = ap_clk;
assign \add_32ns_32s_32_2_1_U25.din0  = ret_V_25_reg_1543;
assign \add_32ns_32s_32_2_1_U25.din1  = { op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17 };
assign grp_fu_1011_p2 = \add_32ns_32s_32_2_1_U25.dout ;
assign \add_32ns_32s_32_2_1_U25.reset  = ap_rst;
assign \add_32ns_32s_32_2_1_U24.top_add_32ns_32s_32_2_1_Adder_17_U.ain_s0  = \add_32ns_32s_32_2_1_U24.top_add_32ns_32s_32_2_1_Adder_17_U.a ;
assign \add_32ns_32s_32_2_1_U24.top_add_32ns_32s_32_2_1_Adder_17_U.bin_s0  = \add_32ns_32s_32_2_1_U24.top_add_32ns_32s_32_2_1_Adder_17_U.b ;
assign \add_32ns_32s_32_2_1_U24.top_add_32ns_32s_32_2_1_Adder_17_U.s  = { \add_32ns_32s_32_2_1_U24.top_add_32ns_32s_32_2_1_Adder_17_U.fas_s2 , \add_32ns_32s_32_2_1_U24.top_add_32ns_32s_32_2_1_Adder_17_U.sum_s1  };
assign \add_32ns_32s_32_2_1_U24.top_add_32ns_32s_32_2_1_Adder_17_U.u2.a  = \add_32ns_32s_32_2_1_U24.top_add_32ns_32s_32_2_1_Adder_17_U.ain_s1 ;
assign \add_32ns_32s_32_2_1_U24.top_add_32ns_32s_32_2_1_Adder_17_U.u2.b  = \add_32ns_32s_32_2_1_U24.top_add_32ns_32s_32_2_1_Adder_17_U.bin_s1 ;
assign \add_32ns_32s_32_2_1_U24.top_add_32ns_32s_32_2_1_Adder_17_U.u2.cin  = \add_32ns_32s_32_2_1_U24.top_add_32ns_32s_32_2_1_Adder_17_U.carry_s1 ;
assign \add_32ns_32s_32_2_1_U24.top_add_32ns_32s_32_2_1_Adder_17_U.facout_s2  = \add_32ns_32s_32_2_1_U24.top_add_32ns_32s_32_2_1_Adder_17_U.u2.cout ;
assign \add_32ns_32s_32_2_1_U24.top_add_32ns_32s_32_2_1_Adder_17_U.fas_s2  = \add_32ns_32s_32_2_1_U24.top_add_32ns_32s_32_2_1_Adder_17_U.u2.s ;
assign \add_32ns_32s_32_2_1_U24.top_add_32ns_32s_32_2_1_Adder_17_U.u1.a  = \add_32ns_32s_32_2_1_U24.top_add_32ns_32s_32_2_1_Adder_17_U.a [15:0];
assign \add_32ns_32s_32_2_1_U24.top_add_32ns_32s_32_2_1_Adder_17_U.u1.b  = \add_32ns_32s_32_2_1_U24.top_add_32ns_32s_32_2_1_Adder_17_U.b [15:0];
assign \add_32ns_32s_32_2_1_U24.top_add_32ns_32s_32_2_1_Adder_17_U.u1.cin  = 1'h0;
assign \add_32ns_32s_32_2_1_U24.top_add_32ns_32s_32_2_1_Adder_17_U.facout_s1  = \add_32ns_32s_32_2_1_U24.top_add_32ns_32s_32_2_1_Adder_17_U.u1.cout ;
assign \add_32ns_32s_32_2_1_U24.top_add_32ns_32s_32_2_1_Adder_17_U.fas_s1  = \add_32ns_32s_32_2_1_U24.top_add_32ns_32s_32_2_1_Adder_17_U.u1.s ;
assign \add_32ns_32s_32_2_1_U24.top_add_32ns_32s_32_2_1_Adder_17_U.a  = \add_32ns_32s_32_2_1_U24.din0 ;
assign \add_32ns_32s_32_2_1_U24.top_add_32ns_32s_32_2_1_Adder_17_U.b  = \add_32ns_32s_32_2_1_U24.din1 ;
assign \add_32ns_32s_32_2_1_U24.top_add_32ns_32s_32_2_1_Adder_17_U.ce  = \add_32ns_32s_32_2_1_U24.ce ;
assign \add_32ns_32s_32_2_1_U24.top_add_32ns_32s_32_2_1_Adder_17_U.clk  = \add_32ns_32s_32_2_1_U24.clk ;
assign \add_32ns_32s_32_2_1_U24.top_add_32ns_32s_32_2_1_Adder_17_U.reset  = \add_32ns_32s_32_2_1_U24.reset ;
assign \add_32ns_32s_32_2_1_U24.dout  = \add_32ns_32s_32_2_1_U24.top_add_32ns_32s_32_2_1_Adder_17_U.s ;
assign \add_32ns_32s_32_2_1_U24.ce  = 1'h1;
assign \add_32ns_32s_32_2_1_U24.clk  = ap_clk;
assign \add_32ns_32s_32_2_1_U24.din0  = ret_V_24_reg_1533;
assign \add_32ns_32s_32_2_1_U24.din1  = { op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16 };
assign grp_fu_1002_p2 = \add_32ns_32s_32_2_1_U24.dout ;
assign \add_32ns_32s_32_2_1_U24.reset  = ap_rst;
assign \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.ain_s0  = \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.a ;
assign \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.bin_s0  = \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.b ;
assign \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.s  = { \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.fas_s2 , \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.sum_s1  };
assign \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.a  = \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.ain_s1 ;
assign \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.b  = \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.bin_s1 ;
assign \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.cin  = \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.carry_s1 ;
assign \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.facout_s2  = \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.cout ;
assign \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.fas_s2  = \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.s ;
assign \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.a  = \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.a [15:0];
assign \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.b  = \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.b [15:0];
assign \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.cin  = 1'h0;
assign \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.facout_s1  = \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.cout ;
assign \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.fas_s1  = \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.s ;
assign \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.a  = \add_32ns_32ns_32_2_1_U23.din0 ;
assign \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.b  = \add_32ns_32ns_32_2_1_U23.din1 ;
assign \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.ce  = \add_32ns_32ns_32_2_1_U23.ce ;
assign \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.clk  = \add_32ns_32ns_32_2_1_U23.clk ;
assign \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.reset  = \add_32ns_32ns_32_2_1_U23.reset ;
assign \add_32ns_32ns_32_2_1_U23.dout  = \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_15_U.s ;
assign \add_32ns_32ns_32_2_1_U23.ce  = 1'h1;
assign \add_32ns_32ns_32_2_1_U23.clk  = ap_clk;
assign \add_32ns_32ns_32_2_1_U23.din0  = ret_V_25_cast_reg_1521;
assign \add_32ns_32ns_32_2_1_U23.din1  = 32'd1;
assign grp_fu_974_p2 = \add_32ns_32ns_32_2_1_U23.dout ;
assign \add_32ns_32ns_32_2_1_U23.reset  = ap_rst;
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.ain_s0  = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.a ;
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.bin_s0  = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.b ;
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.s  = { \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.fas_s2 , \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.sum_s1  };
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.a  = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.ain_s1 ;
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.b  = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.bin_s1 ;
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.cin  = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.carry_s1 ;
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.facout_s2  = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.cout ;
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.fas_s2  = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.u2.s ;
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.a  = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.a [15:0];
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.b  = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.b [15:0];
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.cin  = 1'h0;
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.facout_s1  = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.cout ;
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.fas_s1  = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.u1.s ;
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.a  = \add_32ns_32ns_32_2_1_U21.din0 ;
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.b  = \add_32ns_32ns_32_2_1_U21.din1 ;
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.ce  = \add_32ns_32ns_32_2_1_U21.ce ;
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.clk  = \add_32ns_32ns_32_2_1_U21.clk ;
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.reset  = \add_32ns_32ns_32_2_1_U21.reset ;
assign \add_32ns_32ns_32_2_1_U21.dout  = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_15_U.s ;
assign \add_32ns_32ns_32_2_1_U21.ce  = 1'h1;
assign \add_32ns_32ns_32_2_1_U21.clk  = ap_clk;
assign \add_32ns_32ns_32_2_1_U21.din0  = ret_V_23_cast_reg_1484;
assign \add_32ns_32ns_32_2_1_U21.din1  = 32'd1;
assign grp_fu_909_p2 = \add_32ns_32ns_32_2_1_U21.dout ;
assign \add_32ns_32ns_32_2_1_U21.reset  = ap_rst;
assign \add_11s_11s_11_2_1_U17.top_add_11s_11s_11_2_1_Adder_11_U.ain_s0  = \add_11s_11s_11_2_1_U17.top_add_11s_11s_11_2_1_Adder_11_U.a ;
assign \add_11s_11s_11_2_1_U17.top_add_11s_11s_11_2_1_Adder_11_U.bin_s0  = \add_11s_11s_11_2_1_U17.top_add_11s_11s_11_2_1_Adder_11_U.b ;
assign \add_11s_11s_11_2_1_U17.top_add_11s_11s_11_2_1_Adder_11_U.s  = { \add_11s_11s_11_2_1_U17.top_add_11s_11s_11_2_1_Adder_11_U.fas_s2 , \add_11s_11s_11_2_1_U17.top_add_11s_11s_11_2_1_Adder_11_U.sum_s1  };
assign \add_11s_11s_11_2_1_U17.top_add_11s_11s_11_2_1_Adder_11_U.u2.a  = \add_11s_11s_11_2_1_U17.top_add_11s_11s_11_2_1_Adder_11_U.ain_s1 ;
assign \add_11s_11s_11_2_1_U17.top_add_11s_11s_11_2_1_Adder_11_U.u2.b  = \add_11s_11s_11_2_1_U17.top_add_11s_11s_11_2_1_Adder_11_U.bin_s1 ;
assign \add_11s_11s_11_2_1_U17.top_add_11s_11s_11_2_1_Adder_11_U.u2.cin  = \add_11s_11s_11_2_1_U17.top_add_11s_11s_11_2_1_Adder_11_U.carry_s1 ;
assign \add_11s_11s_11_2_1_U17.top_add_11s_11s_11_2_1_Adder_11_U.facout_s2  = \add_11s_11s_11_2_1_U17.top_add_11s_11s_11_2_1_Adder_11_U.u2.cout ;
assign \add_11s_11s_11_2_1_U17.top_add_11s_11s_11_2_1_Adder_11_U.fas_s2  = \add_11s_11s_11_2_1_U17.top_add_11s_11s_11_2_1_Adder_11_U.u2.s ;
assign \add_11s_11s_11_2_1_U17.top_add_11s_11s_11_2_1_Adder_11_U.u1.a  = \add_11s_11s_11_2_1_U17.top_add_11s_11s_11_2_1_Adder_11_U.a [4:0];
assign \add_11s_11s_11_2_1_U17.top_add_11s_11s_11_2_1_Adder_11_U.u1.b  = \add_11s_11s_11_2_1_U17.top_add_11s_11s_11_2_1_Adder_11_U.b [4:0];
assign \add_11s_11s_11_2_1_U17.top_add_11s_11s_11_2_1_Adder_11_U.u1.cin  = 1'h0;
assign \add_11s_11s_11_2_1_U17.top_add_11s_11s_11_2_1_Adder_11_U.facout_s1  = \add_11s_11s_11_2_1_U17.top_add_11s_11s_11_2_1_Adder_11_U.u1.cout ;
assign \add_11s_11s_11_2_1_U17.top_add_11s_11s_11_2_1_Adder_11_U.fas_s1  = \add_11s_11s_11_2_1_U17.top_add_11s_11s_11_2_1_Adder_11_U.u1.s ;
assign \add_11s_11s_11_2_1_U17.top_add_11s_11s_11_2_1_Adder_11_U.a  = \add_11s_11s_11_2_1_U17.din0 ;
assign \add_11s_11s_11_2_1_U17.top_add_11s_11s_11_2_1_Adder_11_U.b  = \add_11s_11s_11_2_1_U17.din1 ;
assign \add_11s_11s_11_2_1_U17.top_add_11s_11s_11_2_1_Adder_11_U.ce  = \add_11s_11s_11_2_1_U17.ce ;
assign \add_11s_11s_11_2_1_U17.top_add_11s_11s_11_2_1_Adder_11_U.clk  = \add_11s_11s_11_2_1_U17.clk ;
assign \add_11s_11s_11_2_1_U17.top_add_11s_11s_11_2_1_Adder_11_U.reset  = \add_11s_11s_11_2_1_U17.reset ;
assign \add_11s_11s_11_2_1_U17.dout  = \add_11s_11s_11_2_1_U17.top_add_11s_11s_11_2_1_Adder_11_U.s ;
assign \add_11s_11s_11_2_1_U17.ce  = 1'h1;
assign \add_11s_11s_11_2_1_U17.clk  = ap_clk;
assign \add_11s_11s_11_2_1_U17.din0  = { op_23_V_reg_1397[6], op_23_V_reg_1397, 3'h0 };
assign \add_11s_11s_11_2_1_U17.din1  = { op_12_V_reg_1387[7], op_12_V_reg_1387[7], op_12_V_reg_1387[7], op_12_V_reg_1387 };
assign grp_fu_810_p2 = \add_11s_11s_11_2_1_U17.dout ;
assign \add_11s_11s_11_2_1_U17.reset  = ap_rst;
assign \add_10ns_10s_10_2_1_U18.top_add_10ns_10s_10_2_1_Adder_12_U.ain_s0  = \add_10ns_10s_10_2_1_U18.top_add_10ns_10s_10_2_1_Adder_12_U.a ;
assign \add_10ns_10s_10_2_1_U18.top_add_10ns_10s_10_2_1_Adder_12_U.bin_s0  = \add_10ns_10s_10_2_1_U18.top_add_10ns_10s_10_2_1_Adder_12_U.b ;
assign \add_10ns_10s_10_2_1_U18.top_add_10ns_10s_10_2_1_Adder_12_U.s  = { \add_10ns_10s_10_2_1_U18.top_add_10ns_10s_10_2_1_Adder_12_U.fas_s2 , \add_10ns_10s_10_2_1_U18.top_add_10ns_10s_10_2_1_Adder_12_U.sum_s1  };
assign \add_10ns_10s_10_2_1_U18.top_add_10ns_10s_10_2_1_Adder_12_U.u2.a  = \add_10ns_10s_10_2_1_U18.top_add_10ns_10s_10_2_1_Adder_12_U.ain_s1 ;
assign \add_10ns_10s_10_2_1_U18.top_add_10ns_10s_10_2_1_Adder_12_U.u2.b  = \add_10ns_10s_10_2_1_U18.top_add_10ns_10s_10_2_1_Adder_12_U.bin_s1 ;
assign \add_10ns_10s_10_2_1_U18.top_add_10ns_10s_10_2_1_Adder_12_U.u2.cin  = \add_10ns_10s_10_2_1_U18.top_add_10ns_10s_10_2_1_Adder_12_U.carry_s1 ;
assign \add_10ns_10s_10_2_1_U18.top_add_10ns_10s_10_2_1_Adder_12_U.facout_s2  = \add_10ns_10s_10_2_1_U18.top_add_10ns_10s_10_2_1_Adder_12_U.u2.cout ;
assign \add_10ns_10s_10_2_1_U18.top_add_10ns_10s_10_2_1_Adder_12_U.fas_s2  = \add_10ns_10s_10_2_1_U18.top_add_10ns_10s_10_2_1_Adder_12_U.u2.s ;
assign \add_10ns_10s_10_2_1_U18.top_add_10ns_10s_10_2_1_Adder_12_U.u1.a  = \add_10ns_10s_10_2_1_U18.top_add_10ns_10s_10_2_1_Adder_12_U.a [4:0];
assign \add_10ns_10s_10_2_1_U18.top_add_10ns_10s_10_2_1_Adder_12_U.u1.b  = \add_10ns_10s_10_2_1_U18.top_add_10ns_10s_10_2_1_Adder_12_U.b [4:0];
assign \add_10ns_10s_10_2_1_U18.top_add_10ns_10s_10_2_1_Adder_12_U.u1.cin  = 1'h0;
assign \add_10ns_10s_10_2_1_U18.top_add_10ns_10s_10_2_1_Adder_12_U.facout_s1  = \add_10ns_10s_10_2_1_U18.top_add_10ns_10s_10_2_1_Adder_12_U.u1.cout ;
assign \add_10ns_10s_10_2_1_U18.top_add_10ns_10s_10_2_1_Adder_12_U.fas_s1  = \add_10ns_10s_10_2_1_U18.top_add_10ns_10s_10_2_1_Adder_12_U.u1.s ;
assign \add_10ns_10s_10_2_1_U18.top_add_10ns_10s_10_2_1_Adder_12_U.a  = \add_10ns_10s_10_2_1_U18.din0 ;
assign \add_10ns_10s_10_2_1_U18.top_add_10ns_10s_10_2_1_Adder_12_U.b  = \add_10ns_10s_10_2_1_U18.din1 ;
assign \add_10ns_10s_10_2_1_U18.top_add_10ns_10s_10_2_1_Adder_12_U.ce  = \add_10ns_10s_10_2_1_U18.ce ;
assign \add_10ns_10s_10_2_1_U18.top_add_10ns_10s_10_2_1_Adder_12_U.clk  = \add_10ns_10s_10_2_1_U18.clk ;
assign \add_10ns_10s_10_2_1_U18.top_add_10ns_10s_10_2_1_Adder_12_U.reset  = \add_10ns_10s_10_2_1_U18.reset ;
assign \add_10ns_10s_10_2_1_U18.dout  = \add_10ns_10s_10_2_1_U18.top_add_10ns_10s_10_2_1_Adder_12_U.s ;
assign \add_10ns_10s_10_2_1_U18.ce  = 1'h1;
assign \add_10ns_10s_10_2_1_U18.clk  = ap_clk;
assign \add_10ns_10s_10_2_1_U18.din0  = { 2'h0, r_reg_1392 };
assign \add_10ns_10s_10_2_1_U18.din1  = { ret_reg_1126[2], ret_reg_1126[2], ret_reg_1126[2], ret_reg_1126[2], ret_reg_1126[2], ret_reg_1126[2], ret_reg_1126[2], ret_reg_1126 };
assign grp_fu_824_p2 = \add_10ns_10s_10_2_1_U18.dout ;
assign \add_10ns_10s_10_2_1_U18.reset  = ap_rst;
endmodule


// Machine B:
// Processed by function `add_clk_enable_signal` in `verilog_tricks.py`.
// Processed by function `remove_reset_signal` in `verilog_tricks.py`.
module top_B (
  ap_clk,
  ap_start,
  ap_done,
  ap_idle,
  ap_ready,
  op_0,
  op_1,
  op_2,
  op_3,
  op_4,
  op_5,
  op_7,
  op_8,
  op_13,
  op_15,
  op_16,
  op_17,
  op_30,
  op_30_ap_vld,
clk_enable
);
input clk_enable;


input ap_clk;
wire ap_rst;
assign ap_rst = op_30_ap_vld;
input ap_start;
input [1:0] op_0;
input [7:0] op_1;
input [7:0] op_13;
input [7:0] op_15;
input [3:0] op_16;
input [3:0] op_17;
input [1:0] op_2;
input [7:0] op_3;
input [15:0] op_4;
input [3:0] op_5;
input [1:0] op_7;
input [1:0] op_8;
output ap_done;
output ap_idle;
output ap_ready;
output [31:0] op_30;
output op_30_ap_vld;


reg [9:0] add_ln69_3_reg_1182;
reg [5:0] ap_CS_fsm = 6'h01;
reg icmp_ln1494_reg_1155;
reg icmp_ln851_1_reg_1145;
reg icmp_ln851_3_reg_1199;
reg icmp_ln851_4_reg_1216;
reg [7:0] op_12_V_reg_1167;
reg [6:0] op_23_V_reg_1172;
reg p_Result_11_reg_1105;
reg p_Result_12_reg_1120;
reg [4:0] p_Result_s_18_reg_1127;
reg [7:0] p_Val2_2_reg_1112;
reg [17:0] r_V_1_reg_1133;
reg [15:0] r_V_reg_1098;
reg [5:0] ret_V_17_reg_1093;
reg [4:0] ret_V_20_reg_1160;
reg [39:0] ret_V_22_reg_1187;
reg [31:0] ret_V_23_cast_reg_1192;
reg [37:0] ret_V_23_reg_1204;
reg [31:0] ret_V_25_cast_reg_1209;
reg [31:0] ret_V_25_reg_1221;
reg [3:0] ret_V_3_cast_reg_1138;
reg [2:0] ret_reg_1150;
reg [2:0] trunc_ln851_3_reg_1177;
wire [9:0] _000_;
wire [5:0] _001_;
wire _002_;
wire _003_;
wire _004_;
wire _005_;
wire [7:0] _006_;
wire [6:0] _007_;
wire _008_;
wire _009_;
wire [4:0] _010_;
wire [7:0] _011_;
wire [17:0] _012_;
wire [15:0] _013_;
wire [5:0] _014_;
wire [4:0] _015_;
wire [39:0] _016_;
wire [31:0] _017_;
wire [37:0] _018_;
wire [31:0] _019_;
wire [31:0] _020_;
wire [3:0] _021_;
wire [2:0] _022_;
wire [2:0] _023_;
wire [1:0] _024_;
wire _025_;
wire _026_;
wire _027_;
wire _028_;
wire _029_;
wire _030_;
wire _031_;
wire _032_;
wire _033_;
wire _034_;
wire _035_;
wire _036_;
wire _037_;
wire _038_;
wire _039_;
wire _040_;
wire _041_;
wire _042_;
wire _043_;
wire [31:0] add_ln691_1_fu_973_p2;
wire [31:0] add_ln691_2_fu_1040_p2;
wire [8:0] add_ln691_fu_902_p2;
wire [2:0] add_ln69_1_fu_825_p2;
wire [9:0] add_ln69_3_fu_849_p2;
wire [6:0] add_ln69_fu_819_p2;
wire and_ln340_1_fu_708_p2;
wire and_ln340_fu_660_p2;
wire and_ln785_1_fu_714_p2;
wire and_ln785_fu_695_p2;
wire and_ln786_fu_679_p2;
wire ap_CS_fsm_state1;
wire ap_CS_fsm_state2;
wire ap_CS_fsm_state3;
wire ap_CS_fsm_state4;
wire ap_CS_fsm_state5;
wire ap_CS_fsm_state6;
wire [5:0] ap_NS_fsm;
wire ap_clk;
wire ap_done;
wire ap_idle;
wire ap_ready;
wire ap_rst;
wire ap_start;
wire [15:0] ashr_ln1333_fu_361_p0;
wire [15:0] ashr_ln1333_fu_361_p2;
wire [7:0] ashr_ln799_fu_803_p2;
wire [15:0] icmp_ln1494_fu_489_p1;
wire icmp_ln1494_fu_489_p2;
wire [15:0] icmp_ln1499_fu_323_p1;
wire icmp_ln1499_fu_323_p2;
wire icmp_ln768_fu_571_p2;
wire icmp_ln786_fu_597_p2;
wire icmp_ln851_1_fu_439_p2;
wire icmp_ln851_2_fu_897_p2;
wire icmp_ln851_3_fu_960_p2;
wire icmp_ln851_4_fu_1027_p2;
wire icmp_ln851_fu_283_p2;
wire isNeg_fu_329_p3;
wire [4:0] lhs_V_fu_495_p3;
wire [4:0] lhs_fu_239_p3;
wire [15:0] \mul_16s_2s_18_1_1_U1.din0 ;
wire [1:0] \mul_16s_2s_18_1_1_U1.din1 ;
wire [17:0] \mul_16s_2s_18_1_1_U1.dout ;
wire [15:0] \mul_16s_2s_18_1_1_U1.top_mul_16s_2s_18_1_1_Multiplier_0_U.a ;
wire [1:0] \mul_16s_2s_18_1_1_U1.top_mul_16s_2s_18_1_1_Multiplier_0_U.b ;
wire [17:0] \mul_16s_2s_18_1_1_U1.top_mul_16s_2s_18_1_1_Multiplier_0_U.p ;
wire [1:0] op_0;
wire [7:0] op_1;
wire [7:0] op_12_V_fu_732_p3;
wire [7:0] op_13;
wire [7:0] op_15;
wire [3:0] op_16;
wire [3:0] op_17;
wire [1:0] op_2;
wire [6:0] op_23_V_fu_835_p2;
wire [7:0] op_3;
wire [31:0] op_30;
wire op_30_ap_vld;
wire [15:0] op_4;
wire [3:0] op_5;
wire [1:0] op_7;
wire [1:0] op_8;
wire [1:0] op_9_V_fu_455_p3;
wire or_ln340_fu_608_p2;
wire or_ln785_1_fu_690_p2;
wire or_ln785_2_fu_720_p2;
wire or_ln785_fu_576_p2;
wire or_ln786_fu_602_p2;
wire overflow_fu_586_p2;
wire p_Result_10_fu_1033_p3;
wire p_Result_13_fu_564_p3;
wire p_Result_14_fu_778_p3;
wire [7:0] p_Result_4_fu_644_p4;
wire p_Result_5_fu_739_p3;
wire p_Result_6_fu_527_p3;
wire p_Result_8_fu_889_p3;
wire p_Result_9_fu_966_p3;
wire p_Result_s_fu_271_p3;
wire [6:0] p_Val2_3_fu_639_p2;
wire [17:0] r_V_1_fu_419_p2;
wire [15:0] r_V_fu_367_p3;
wire [7:0] r_fu_808_p3;
wire [8:0] ret_V_16_fu_255_p2;
wire [5:0] ret_V_17_fu_303_p3;
wire [3:0] ret_V_18_fu_757_p3;
wire [5:0] ret_V_19_fu_511_p2;
wire [4:0] ret_V_20_fu_553_p3;
wire [10:0] ret_V_21_fu_869_p2;
wire [39:0] ret_V_22_fu_940_p2;
wire [37:0] ret_V_23_fu_1007_p2;
wire [31:0] ret_V_24_fu_1051_p3;
wire [31:0] ret_V_25_fu_1062_p2;
wire [31:0] ret_V_26_fu_1072_p2;
wire [5:0] ret_V_2_fu_289_p2;
wire [3:0] ret_V_4_fu_746_p2;
wire [4:0] ret_V_7_fu_517_p4;
wire [4:0] ret_V_8_fu_539_p2;
wire [5:0] ret_V_fu_261_p4;
wire [2:0] ret_fu_471_p2;
wire [9:0] rhs_2_fu_858_p3;
wire [36:0] rhs_3_fu_995_p3;
wire sel_tmp11_fu_726_p2;
wire [7:0] select_ln340_fu_666_p3;
wire [31:0] select_ln353_1_fu_988_p3;
wire [8:0] select_ln353_fu_920_p3;
wire [7:0] select_ln785_fu_701_p3;
wire [3:0] select_ln850_1_fu_751_p3;
wire [4:0] select_ln850_2_fu_545_p3;
wire [31:0] select_ln850_5_fu_1045_p3;
wire [8:0] select_ln850_6_fu_912_p3;
wire [31:0] select_ln850_7_fu_982_p3;
wire [5:0] select_ln850_fu_295_p3;
wire [10:0] sext_ln1192_1_fu_865_p1;
wire [39:0] sext_ln1192_2_fu_936_p1;
wire [37:0] sext_ln1192_3_fu_1003_p1;
wire [31:0] sext_ln1192_4_fu_1058_p1;
wire [31:0] sext_ln1192_5_fu_1068_p1;
wire [10:0] sext_ln1192_fu_855_p1;
wire [5:0] sext_ln1193_fu_503_p1;
wire [15:0] sext_ln1499_fu_319_p1;
wire [5:0] sext_ln17_fu_771_p1;
wire [9:0] sext_ln18_fu_764_p1;
wire [6:0] sext_ln20_fu_561_p1;
wire [1:0] sext_ln215_1_fu_467_p0;
wire [2:0] sext_ln215_1_fu_467_p1;
wire [1:0] sext_ln215_fu_463_p0;
wire [2:0] sext_ln215_fu_463_p1;
wire [7:0] sext_ln546_1_fu_800_p1;
wire [7:0] sext_ln546_fu_791_p1;
wire [31:0] sext_ln69_fu_1077_p1;
wire [7:0] sext_ln703_1_fu_908_p0;
wire [39:0] sext_ln703_1_fu_908_p1;
wire [7:0] sext_ln703_2_fu_978_p0;
wire [37:0] sext_ln703_2_fu_978_p1;
wire [7:0] sext_ln703_fu_251_p0;
wire [8:0] sext_ln703_fu_251_p1;
wire [8:0] sext_ln850_fu_885_p1;
wire [1:0] sext_ln886_fu_445_p0;
wire [3:0] sext_ln886_fu_445_p1;
wire [5:0] sh_V_1_fu_785_p2;
wire [15:0] shl_ln1299_fu_355_p0;
wire [15:0] shl_ln1299_fu_355_p2;
wire [6:0] shl_ln728_2_fu_477_p3;
wire [7:0] shl_ln781_fu_795_p2;
wire [13:0] shl_ln_fu_311_p3;
wire signbit_fu_449_p2;
wire [3:0] sub_ln1367_fu_337_p2;
wire [15:0] tmp_13_fu_928_p3;
wire tmp_6_fu_613_p3;
wire tmp_7_fu_620_p3;
wire [7:0] tmp_fu_875_p4;
wire [5:0] trunc_ln851_1_fu_435_p1;
wire trunc_ln851_2_fu_535_p1;
wire [2:0] trunc_ln851_3_fu_841_p1;
wire [7:0] trunc_ln851_4_fu_956_p0;
wire [6:0] trunc_ln851_4_fu_956_p1;
wire [7:0] trunc_ln851_5_fu_1023_p0;
wire [4:0] trunc_ln851_5_fu_1023_p1;
wire [7:0] trunc_ln851_fu_279_p0;
wire [2:0] trunc_ln851_fu_279_p1;
wire [3:0] ush_fu_343_p3;
wire xor_ln340_fu_654_p2;
wire xor_ln365_1_fu_633_p2;
wire xor_ln365_fu_627_p2;
wire xor_ln785_1_fu_684_p2;
wire xor_ln785_fu_581_p2;
wire xor_ln786_1_fu_673_p2;
wire xor_ln786_fu_592_p2;
wire [8:0] zext_ln1192_fu_247_p1;
wire [15:0] zext_ln1367_fu_351_p1;
wire [15:0] zext_ln1494_fu_485_p1;
wire [6:0] zext_ln69_1_fu_831_p1;
wire [9:0] zext_ln69_2_fu_845_p1;
wire [2:0] zext_ln69_fu_816_p1;
wire [5:0] zext_ln703_fu_507_p1;
wire [2:0] zext_ln727_fu_767_p1;
wire [6:0] zext_ln787_fu_774_p1;


assign add_ln691_1_fu_973_p2 = ret_V_23_cast_reg_1192 + 1'h1;
assign add_ln691_2_fu_1040_p2 = ret_V_25_cast_reg_1209 + 1'h1;
assign add_ln691_fu_902_p2 = $signed(ret_V_21_fu_869_p2[10:3]) + $signed(2'h1);
assign add_ln69_1_fu_825_p2 = op_2 + icmp_ln1494_reg_1155;
assign add_ln69_3_fu_849_p2 = $signed({ 1'h0, r_fu_808_p3 }) + $signed(ret_reg_1150);
assign add_ln69_fu_819_p2 = $signed(ret_V_17_reg_1093) + $signed({ 1'h0, ret_V_18_fu_757_p3 });
assign op_23_V_fu_835_p2 = add_ln69_1_fu_825_p2 + add_ln69_fu_819_p2;
assign op_30 = $signed(add_ln69_3_reg_1182) + $signed(ret_V_26_fu_1072_p2);
assign ret_V_16_fu_255_p2 = $signed({ 1'h0, op_0, 3'h0 }) + $signed(op_1);
assign ret_V_21_fu_869_p2 = $signed({ op_23_V_reg_1172, 3'h0 }) + $signed(op_12_V_reg_1167);
assign { ret_V_22_fu_940_p2[39], ret_V_22_fu_940_p2[15:0] } = $signed({ select_ln353_fu_920_p3, 7'h00 }) + $signed(op_13);
assign ret_V_23_fu_1007_p2 = $signed({ select_ln353_1_fu_988_p3, 5'h00 }) + $signed(op_15);
assign ret_V_25_fu_1062_p2 = $signed(ret_V_24_fu_1051_p3) + $signed(op_16);
assign ret_V_26_fu_1072_p2 = $signed(ret_V_25_reg_1221) + $signed(op_17);
assign ret_V_2_fu_289_p2 = ret_V_16_fu_255_p2[8:3] + 1'h1;
assign ret_V_4_fu_746_p2 = ret_V_3_cast_reg_1138 + 1'h1;
assign ret_V_8_fu_539_p2 = ret_V_19_fu_511_p2[5:1] + 1'h1;
assign ret_fu_471_p2 = $signed(op_8) + $signed(op_7);
assign _025_ = ap_CS_fsm[0] & _027_;
assign _026_ = ap_CS_fsm[0] & ap_start;
assign and_ln340_1_fu_708_p2 = or_ln786_fu_602_p2 & or_ln340_fu_608_p2;
assign and_ln340_fu_660_p2 = xor_ln340_fu_654_p2 & or_ln786_fu_602_p2;
assign and_ln785_1_fu_714_p2 = xor_ln785_fu_581_p2 & and_ln786_fu_679_p2;
assign and_ln785_fu_695_p2 = or_ln785_1_fu_690_p2 & and_ln786_fu_679_p2;
assign and_ln786_fu_679_p2 = xor_ln786_1_fu_673_p2 & p_Result_12_reg_1120;
assign overflow_fu_586_p2 = xor_ln785_fu_581_p2 & or_ln785_fu_576_p2;
assign sel_tmp11_fu_726_p2 = xor_ln365_1_fu_633_p2 & or_ln785_2_fu_720_p2;
assign xor_ln785_fu_581_p2 = ~ p_Result_11_reg_1105;
assign xor_ln786_fu_592_p2 = ~ p_Result_12_reg_1120;
assign xor_ln340_fu_654_p2 = ~ or_ln340_fu_608_p2;
assign xor_ln786_1_fu_673_p2 = ~ icmp_ln786_fu_597_p2;
assign xor_ln785_1_fu_684_p2 = ~ or_ln785_fu_576_p2;
assign xor_ln365_1_fu_633_p2 = ~ xor_ln365_fu_627_p2;
assign p_Val2_3_fu_639_p2 = ~ p_Val2_2_reg_1112[6:0];
assign _027_ = ~ ap_start;
assign _028_ = ! r_V_1_fu_419_p2[5:0];
assign _029_ = ! op_1[2:0];
assign \mul_16s_2s_18_1_1_U1.top_mul_16s_2s_18_1_1_Multiplier_0_U.p  = $signed(\mul_16s_2s_18_1_1_U1.top_mul_16s_2s_18_1_1_Multiplier_0_U.a ) * $signed(\mul_16s_2s_18_1_1_U1.top_mul_16s_2s_18_1_1_Multiplier_0_U.b );
assign _030_ = $signed({ 1'h0, icmp_ln1499_fu_323_p2, 6'h00 }) < $signed(op_4);
assign _031_ = $signed(op_8) < $signed(op_5);
assign _032_ = $signed({ op_3, 6'h00 }) != $signed(op_4);
assign _033_ = | p_Result_s_18_reg_1127;
assign _034_ = p_Result_s_18_reg_1127 != 5'h1f;
assign _035_ = | trunc_ln851_3_reg_1177;
assign _036_ = | op_13[6:0];
assign _037_ = | op_15[4:0];
assign or_ln340_fu_608_p2 = p_Result_11_reg_1105 | overflow_fu_586_p2;
assign or_ln785_1_fu_690_p2 = xor_ln785_1_fu_684_p2 | p_Result_11_reg_1105;
assign or_ln785_2_fu_720_p2 = and_ln785_1_fu_714_p2 | and_ln340_1_fu_708_p2;
assign or_ln785_fu_576_p2 = p_Result_12_reg_1120 | icmp_ln768_fu_571_p2;
assign or_ln786_fu_602_p2 = xor_ln786_fu_592_p2 | icmp_ln786_fu_597_p2;
always @(posedge ap_clk)
ret_V_25_reg_1221 <= _020_;
always @(posedge ap_clk)
ret_V_23_reg_1204 <= _018_;
always @(posedge ap_clk)
ret_V_25_cast_reg_1209 <= _019_;
always @(posedge ap_clk)
icmp_ln851_4_reg_1216 <= _005_;
always @(posedge ap_clk)
ret_V_22_reg_1187 <= _016_;
always @(posedge ap_clk)
ret_V_23_cast_reg_1192 <= _017_;
always @(posedge ap_clk)
icmp_ln851_3_reg_1199 <= _004_;
always @(posedge ap_clk)
ret_V_17_reg_1093 <= _014_;
always @(posedge ap_clk)
r_V_reg_1098 <= _013_;
always @(posedge ap_clk)
p_Result_11_reg_1105 <= _008_;
always @(posedge ap_clk)
p_Val2_2_reg_1112 <= _011_;
always @(posedge ap_clk)
p_Result_12_reg_1120 <= _009_;
always @(posedge ap_clk)
p_Result_s_18_reg_1127 <= _010_;
always @(posedge ap_clk)
r_V_1_reg_1133 <= _012_;
always @(posedge ap_clk)
ret_V_3_cast_reg_1138 <= _021_;
always @(posedge ap_clk)
icmp_ln851_1_reg_1145 <= _003_;
always @(posedge ap_clk)
ret_reg_1150 <= _022_;
always @(posedge ap_clk)
icmp_ln1494_reg_1155 <= _002_;
always @(posedge ap_clk)
ret_V_20_reg_1160 <= _015_;
always @(posedge ap_clk)
op_12_V_reg_1167 <= _006_;
always @(posedge ap_clk)
op_23_V_reg_1172 <= _007_;
always @(posedge ap_clk)
trunc_ln851_3_reg_1177 <= _023_;
always @(posedge ap_clk)
add_ln69_3_reg_1182 <= _000_;
always @(posedge ap_clk)
ap_CS_fsm <= _001_;
assign _024_ = _026_ ? 2'h2 : 2'h1;
assign _038_ = ap_CS_fsm == 1'h1;
function [5:0] _121_;
input [5:0] a;
input [35:0] b;
input [5:0] s;
case (s)
6'b000001:
_121_ = b[5:0];
6'b000010:
_121_ = b[11:6];
6'b000100:
_121_ = b[17:12];
6'b001000:
_121_ = b[23:18];
6'b010000:
_121_ = b[29:24];
6'b100000:
_121_ = b[35:30];
6'b000000:
_121_ = a;
default:
_121_ = 6'bx;
endcase
endfunction
assign ap_NS_fsm = _121_(6'hxx, { 4'h0, _024_, 30'h04210801 }, { _038_, _043_, _042_, _041_, _040_, _039_ });
assign _039_ = ap_CS_fsm == 6'h20;
assign _040_ = ap_CS_fsm == 5'h10;
assign _041_ = ap_CS_fsm == 4'h8;
assign _042_ = ap_CS_fsm == 3'h4;
assign _043_ = ap_CS_fsm == 2'h2;
assign op_30_ap_vld = ap_CS_fsm[5] ? 1'h1 : 1'h0;
assign ap_idle = _025_ ? 1'h1 : 1'h0;
assign _020_ = ap_CS_fsm[4] ? ret_V_25_fu_1062_p2 : ret_V_25_reg_1221;
assign _005_ = ap_CS_fsm[3] ? icmp_ln851_4_fu_1027_p2 : icmp_ln851_4_reg_1216;
assign _019_ = ap_CS_fsm[3] ? ret_V_23_fu_1007_p2[36:5] : ret_V_25_cast_reg_1209;
assign _018_ = ap_CS_fsm[3] ? ret_V_23_fu_1007_p2 : ret_V_23_reg_1204;
assign _004_ = ap_CS_fsm[2] ? icmp_ln851_3_fu_960_p2 : icmp_ln851_3_reg_1199;
assign _017_ = ap_CS_fsm[2] ? { ret_V_22_fu_940_p2[39], ret_V_22_fu_940_p2[39], ret_V_22_fu_940_p2[39], ret_V_22_fu_940_p2[39], ret_V_22_fu_940_p2[39], ret_V_22_fu_940_p2[39], ret_V_22_fu_940_p2[39], ret_V_22_fu_940_p2[39], ret_V_22_fu_940_p2[39], ret_V_22_fu_940_p2[39], ret_V_22_fu_940_p2[39], ret_V_22_fu_940_p2[39], ret_V_22_fu_940_p2[39], ret_V_22_fu_940_p2[39], ret_V_22_fu_940_p2[39], ret_V_22_fu_940_p2[39], ret_V_22_fu_940_p2[39], ret_V_22_fu_940_p2[39], ret_V_22_fu_940_p2[39], ret_V_22_fu_940_p2[39], ret_V_22_fu_940_p2[39], ret_V_22_fu_940_p2[39], ret_V_22_fu_940_p2[39], ret_V_22_fu_940_p2[15:7] } : ret_V_23_cast_reg_1192;
assign _016_ = ap_CS_fsm[2] ? { ret_V_22_fu_940_p2[39], ret_V_22_fu_940_p2[39], ret_V_22_fu_940_p2[39], ret_V_22_fu_940_p2[39], ret_V_22_fu_940_p2[39], ret_V_22_fu_940_p2[39], ret_V_22_fu_940_p2[39], ret_V_22_fu_940_p2[39], ret_V_22_fu_940_p2[39], ret_V_22_fu_940_p2[39], ret_V_22_fu_940_p2[39], ret_V_22_fu_940_p2[39], ret_V_22_fu_940_p2[39], ret_V_22_fu_940_p2[39], ret_V_22_fu_940_p2[39], ret_V_22_fu_940_p2[39], ret_V_22_fu_940_p2[39], ret_V_22_fu_940_p2[39], ret_V_22_fu_940_p2[39], ret_V_22_fu_940_p2[39], ret_V_22_fu_940_p2[39], ret_V_22_fu_940_p2[39], ret_V_22_fu_940_p2[39], ret_V_22_fu_940_p2[39], ret_V_22_fu_940_p2[15:0] } : ret_V_22_reg_1187;
assign _015_ = ap_CS_fsm[0] ? ret_V_20_fu_553_p3 : ret_V_20_reg_1160;
assign _002_ = ap_CS_fsm[0] ? icmp_ln1494_fu_489_p2 : icmp_ln1494_reg_1155;
assign _022_ = ap_CS_fsm[0] ? ret_fu_471_p2 : ret_reg_1150;
assign _003_ = ap_CS_fsm[0] ? icmp_ln851_1_fu_439_p2 : icmp_ln851_1_reg_1145;
assign _021_ = ap_CS_fsm[0] ? r_V_1_fu_419_p2[9:6] : ret_V_3_cast_reg_1138;
assign _012_ = ap_CS_fsm[0] ? r_V_1_fu_419_p2 : r_V_1_reg_1133;
assign _010_ = ap_CS_fsm[0] ? r_V_fu_367_p3[15:11] : p_Result_s_18_reg_1127;
assign _009_ = ap_CS_fsm[0] ? r_V_fu_367_p3[10] : p_Result_12_reg_1120;
assign _011_ = ap_CS_fsm[0] ? r_V_fu_367_p3[10:3] : p_Val2_2_reg_1112;
assign _008_ = ap_CS_fsm[0] ? r_V_fu_367_p3[15] : p_Result_11_reg_1105;
assign _013_ = ap_CS_fsm[0] ? r_V_fu_367_p3 : r_V_reg_1098;
assign _014_ = ap_CS_fsm[0] ? ret_V_17_fu_303_p3 : ret_V_17_reg_1093;
assign _000_ = ap_CS_fsm[1] ? add_ln69_3_fu_849_p2 : add_ln69_3_reg_1182;
assign _023_ = ap_CS_fsm[1] ? op_12_V_fu_732_p3[2:0] : trunc_ln851_3_reg_1177;
assign _007_ = ap_CS_fsm[1] ? op_23_V_fu_835_p2 : op_23_V_reg_1172;
assign _006_ = ap_CS_fsm[1] ? op_12_V_fu_732_p3 : op_12_V_reg_1167;
assign _001_ = ap_rst ? 6'h01 : ap_NS_fsm;
assign shl_ln1299_fu_355_p2 = $signed(op_4) << ush_fu_343_p3;
assign shl_ln781_fu_795_p2 = op_3 << { sh_V_1_fu_785_p2[5], sh_V_1_fu_785_p2[5], sh_V_1_fu_785_p2 };
assign ashr_ln1333_fu_361_p2 = $signed(op_4) >>> ush_fu_343_p3;
assign ashr_ln799_fu_803_p2 = $signed(op_3) >>> { ret_V_20_reg_1160[4], ret_V_20_reg_1160[4], ret_V_20_reg_1160[4], ret_V_20_reg_1160 };
assign ret_V_19_fu_511_p2 = $signed({ op_5, 1'h0 }) - $signed({ 1'h0, signbit_fu_449_p2, 1'h0 });
assign sh_V_1_fu_785_p2 = $signed(1'h0) - $signed(ret_V_20_reg_1160);
assign sub_ln1367_fu_337_p2 = 1'h0 - op_5;
assign icmp_ln1494_fu_489_p2 = _030_ ? 1'h1 : 1'h0;
assign icmp_ln1499_fu_323_p2 = _032_ ? 1'h1 : 1'h0;
assign icmp_ln768_fu_571_p2 = _033_ ? 1'h1 : 1'h0;
assign icmp_ln786_fu_597_p2 = _034_ ? 1'h1 : 1'h0;
assign icmp_ln851_1_fu_439_p2 = _028_ ? 1'h1 : 1'h0;
assign icmp_ln851_2_fu_897_p2 = _035_ ? 1'h1 : 1'h0;
assign icmp_ln851_3_fu_960_p2 = _036_ ? 1'h1 : 1'h0;
assign icmp_ln851_4_fu_1027_p2 = _037_ ? 1'h1 : 1'h0;
assign icmp_ln851_fu_283_p2 = _029_ ? 1'h1 : 1'h0;
assign op_12_V_fu_732_p3 = sel_tmp11_fu_726_p2 ? p_Val2_2_reg_1112 : select_ln785_fu_701_p3;
assign r_V_fu_367_p3 = op_5[3] ? shl_ln1299_fu_355_p2 : ashr_ln1333_fu_361_p2;
assign r_fu_808_p3 = ret_V_20_reg_1160[4] ? shl_ln781_fu_795_p2 : ashr_ln799_fu_803_p2;
assign ret_V_17_fu_303_p3 = ret_V_16_fu_255_p2[8] ? select_ln850_fu_295_p3 : { 1'h0, ret_V_16_fu_255_p2[7:3] };
assign ret_V_18_fu_757_p3 = r_V_1_reg_1133[17] ? select_ln850_1_fu_751_p3 : ret_V_3_cast_reg_1138;
assign ret_V_20_fu_553_p3 = ret_V_19_fu_511_p2[5] ? select_ln850_2_fu_545_p3 : { 1'h0, ret_V_19_fu_511_p2[4:1] };
assign ret_V_24_fu_1051_p3 = ret_V_23_reg_1204[37] ? select_ln850_5_fu_1045_p3 : ret_V_25_cast_reg_1209;
assign select_ln340_fu_666_p3 = and_ln340_fu_660_p2 ? p_Val2_2_reg_1112 : { r_V_reg_1098[11], p_Val2_3_fu_639_p2 };
assign select_ln353_1_fu_988_p3 = ret_V_22_reg_1187[39] ? select_ln850_7_fu_982_p3 : ret_V_23_cast_reg_1192;
assign select_ln353_fu_920_p3 = ret_V_21_fu_869_p2[10] ? select_ln850_6_fu_912_p3 : { 2'h0, ret_V_21_fu_869_p2[9:3] };
assign select_ln785_fu_701_p3 = and_ln785_fu_695_p2 ? p_Val2_2_reg_1112 : select_ln340_fu_666_p3;
assign select_ln850_1_fu_751_p3 = icmp_ln851_1_reg_1145 ? ret_V_3_cast_reg_1138 : ret_V_4_fu_746_p2;
assign select_ln850_2_fu_545_p3 = ret_V_19_fu_511_p2[0] ? ret_V_8_fu_539_p2 : { 1'h1, ret_V_19_fu_511_p2[4:1] };
assign select_ln850_5_fu_1045_p3 = icmp_ln851_4_reg_1216 ? add_ln691_2_fu_1040_p2 : ret_V_25_cast_reg_1209;
assign select_ln850_6_fu_912_p3 = icmp_ln851_2_fu_897_p2 ? add_ln691_fu_902_p2 : { 2'h3, ret_V_21_fu_869_p2[9:3] };
assign select_ln850_7_fu_982_p3 = icmp_ln851_3_reg_1199 ? add_ln691_1_fu_973_p2 : ret_V_23_cast_reg_1192;
assign select_ln850_fu_295_p3 = icmp_ln851_fu_283_p2 ? { 1'h1, ret_V_16_fu_255_p2[7:3] } : ret_V_2_fu_289_p2;
assign signbit_fu_449_p2 = _031_ ? 1'h1 : 1'h0;
assign ush_fu_343_p3 = op_5[3] ? sub_ln1367_fu_337_p2 : { 1'h0, op_5[2:0] };
assign xor_ln365_fu_627_p2 = r_V_reg_1098[10] ^ r_V_reg_1098[11];
assign ap_CS_fsm_state1 = ap_CS_fsm[0];
assign ap_CS_fsm_state2 = ap_CS_fsm[1];
assign ap_CS_fsm_state3 = ap_CS_fsm[2];
assign ap_CS_fsm_state4 = ap_CS_fsm[3];
assign ap_CS_fsm_state5 = ap_CS_fsm[4];
assign ap_CS_fsm_state6 = ap_CS_fsm[5];
assign ap_done = op_30_ap_vld;
assign ap_ready = op_30_ap_vld;
assign ashr_ln1333_fu_361_p0 = op_4;
assign icmp_ln1494_fu_489_p1 = op_4;
assign icmp_ln1499_fu_323_p1 = op_4;
assign isNeg_fu_329_p3 = op_5[3];
assign lhs_V_fu_495_p3 = { op_5, 1'h0 };
assign lhs_fu_239_p3 = { op_0, 3'h0 };
assign op_9_V_fu_455_p3 = { signbit_fu_449_p2, 1'h0 };
assign p_Result_10_fu_1033_p3 = ret_V_23_reg_1204[37];
assign p_Result_13_fu_564_p3 = r_V_reg_1098[11];
assign p_Result_14_fu_778_p3 = ret_V_20_reg_1160[4];
assign p_Result_4_fu_644_p4 = { r_V_reg_1098[11], p_Val2_3_fu_639_p2 };
assign p_Result_5_fu_739_p3 = r_V_1_reg_1133[17];
assign p_Result_6_fu_527_p3 = ret_V_19_fu_511_p2[5];
assign p_Result_8_fu_889_p3 = ret_V_21_fu_869_p2[10];
assign p_Result_9_fu_966_p3 = ret_V_22_reg_1187[39];
assign p_Result_s_fu_271_p3 = ret_V_16_fu_255_p2[8];
assign ret_V_22_fu_940_p2[38:16] = { ret_V_22_fu_940_p2[39], ret_V_22_fu_940_p2[39], ret_V_22_fu_940_p2[39], ret_V_22_fu_940_p2[39], ret_V_22_fu_940_p2[39], ret_V_22_fu_940_p2[39], ret_V_22_fu_940_p2[39], ret_V_22_fu_940_p2[39], ret_V_22_fu_940_p2[39], ret_V_22_fu_940_p2[39], ret_V_22_fu_940_p2[39], ret_V_22_fu_940_p2[39], ret_V_22_fu_940_p2[39], ret_V_22_fu_940_p2[39], ret_V_22_fu_940_p2[39], ret_V_22_fu_940_p2[39], ret_V_22_fu_940_p2[39], ret_V_22_fu_940_p2[39], ret_V_22_fu_940_p2[39], ret_V_22_fu_940_p2[39], ret_V_22_fu_940_p2[39], ret_V_22_fu_940_p2[39], ret_V_22_fu_940_p2[39] };
assign ret_V_7_fu_517_p4 = ret_V_19_fu_511_p2[5:1];
assign ret_V_fu_261_p4 = ret_V_16_fu_255_p2[8:3];
assign rhs_2_fu_858_p3 = { op_23_V_reg_1172, 3'h0 };
assign rhs_3_fu_995_p3 = { select_ln353_1_fu_988_p3, 5'h00 };
assign sext_ln1192_1_fu_865_p1 = { op_23_V_reg_1172[6], op_23_V_reg_1172, 3'h0 };
assign sext_ln1192_2_fu_936_p1 = { select_ln353_fu_920_p3[8], select_ln353_fu_920_p3[8], select_ln353_fu_920_p3[8], select_ln353_fu_920_p3[8], select_ln353_fu_920_p3[8], select_ln353_fu_920_p3[8], select_ln353_fu_920_p3[8], select_ln353_fu_920_p3[8], select_ln353_fu_920_p3[8], select_ln353_fu_920_p3[8], select_ln353_fu_920_p3[8], select_ln353_fu_920_p3[8], select_ln353_fu_920_p3[8], select_ln353_fu_920_p3[8], select_ln353_fu_920_p3[8], select_ln353_fu_920_p3[8], select_ln353_fu_920_p3[8], select_ln353_fu_920_p3[8], select_ln353_fu_920_p3[8], select_ln353_fu_920_p3[8], select_ln353_fu_920_p3[8], select_ln353_fu_920_p3[8], select_ln353_fu_920_p3[8], select_ln353_fu_920_p3[8], select_ln353_fu_920_p3, 7'h00 };
assign sext_ln1192_3_fu_1003_p1 = { select_ln353_1_fu_988_p3[31], select_ln353_1_fu_988_p3, 5'h00 };
assign sext_ln1192_4_fu_1058_p1 = { op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16 };
assign sext_ln1192_5_fu_1068_p1 = { op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17 };
assign sext_ln1192_fu_855_p1 = { op_12_V_reg_1167[7], op_12_V_reg_1167[7], op_12_V_reg_1167[7], op_12_V_reg_1167 };
assign sext_ln1193_fu_503_p1 = { op_5[3], op_5, 1'h0 };
assign sext_ln1499_fu_319_p1 = { op_3[7], op_3[7], op_3, 6'h00 };
assign sext_ln17_fu_771_p1 = { ret_V_20_reg_1160[4], ret_V_20_reg_1160 };
assign sext_ln18_fu_764_p1 = { ret_reg_1150[2], ret_reg_1150[2], ret_reg_1150[2], ret_reg_1150[2], ret_reg_1150[2], ret_reg_1150[2], ret_reg_1150[2], ret_reg_1150 };
assign sext_ln20_fu_561_p1 = { ret_V_17_reg_1093[5], ret_V_17_reg_1093 };
assign sext_ln215_1_fu_467_p0 = op_8;
assign sext_ln215_1_fu_467_p1 = { op_8[1], op_8 };
assign sext_ln215_fu_463_p0 = op_7;
assign sext_ln215_fu_463_p1 = { op_7[1], op_7 };
assign sext_ln546_1_fu_800_p1 = { ret_V_20_reg_1160[4], ret_V_20_reg_1160[4], ret_V_20_reg_1160[4], ret_V_20_reg_1160 };
assign sext_ln546_fu_791_p1 = { sh_V_1_fu_785_p2[5], sh_V_1_fu_785_p2[5], sh_V_1_fu_785_p2 };
assign sext_ln69_fu_1077_p1 = { add_ln69_3_reg_1182[9], add_ln69_3_reg_1182[9], add_ln69_3_reg_1182[9], add_ln69_3_reg_1182[9], add_ln69_3_reg_1182[9], add_ln69_3_reg_1182[9], add_ln69_3_reg_1182[9], add_ln69_3_reg_1182[9], add_ln69_3_reg_1182[9], add_ln69_3_reg_1182[9], add_ln69_3_reg_1182[9], add_ln69_3_reg_1182[9], add_ln69_3_reg_1182[9], add_ln69_3_reg_1182[9], add_ln69_3_reg_1182[9], add_ln69_3_reg_1182[9], add_ln69_3_reg_1182[9], add_ln69_3_reg_1182[9], add_ln69_3_reg_1182[9], add_ln69_3_reg_1182[9], add_ln69_3_reg_1182[9], add_ln69_3_reg_1182[9], add_ln69_3_reg_1182 };
assign sext_ln703_1_fu_908_p0 = op_13;
assign sext_ln703_1_fu_908_p1 = { op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13 };
assign sext_ln703_2_fu_978_p0 = op_15;
assign sext_ln703_2_fu_978_p1 = { op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15[7], op_15 };
assign sext_ln703_fu_251_p0 = op_1;
assign sext_ln703_fu_251_p1 = { op_1[7], op_1 };
assign sext_ln850_fu_885_p1 = { ret_V_21_fu_869_p2[10], ret_V_21_fu_869_p2[10:3] };
assign sext_ln886_fu_445_p0 = op_8;
assign sext_ln886_fu_445_p1 = { op_8[1], op_8[1], op_8 };
assign shl_ln1299_fu_355_p0 = op_4;
assign shl_ln728_2_fu_477_p3 = { icmp_ln1499_fu_323_p2, 6'h00 };
assign shl_ln_fu_311_p3 = { op_3, 6'h00 };
assign tmp_13_fu_928_p3 = { select_ln353_fu_920_p3, 7'h00 };
assign tmp_6_fu_613_p3 = r_V_reg_1098[11];
assign tmp_7_fu_620_p3 = r_V_reg_1098[10];
assign tmp_fu_875_p4 = ret_V_21_fu_869_p2[10:3];
assign trunc_ln851_1_fu_435_p1 = r_V_1_fu_419_p2[5:0];
assign trunc_ln851_2_fu_535_p1 = ret_V_19_fu_511_p2[0];
assign trunc_ln851_3_fu_841_p1 = op_12_V_fu_732_p3[2:0];
assign trunc_ln851_4_fu_956_p0 = op_13;
assign trunc_ln851_4_fu_956_p1 = op_13[6:0];
assign trunc_ln851_5_fu_1023_p0 = op_15;
assign trunc_ln851_5_fu_1023_p1 = op_15[4:0];
assign trunc_ln851_fu_279_p0 = op_1;
assign trunc_ln851_fu_279_p1 = op_1[2:0];
assign zext_ln1192_fu_247_p1 = { 4'h0, op_0, 3'h0 };
assign zext_ln1367_fu_351_p1 = { 12'h000, ush_fu_343_p3 };
assign zext_ln1494_fu_485_p1 = { 9'h000, icmp_ln1499_fu_323_p2, 6'h00 };
assign zext_ln69_1_fu_831_p1 = { 4'h0, add_ln69_1_fu_825_p2 };
assign zext_ln69_2_fu_845_p1 = { 2'h0, r_fu_808_p3 };
assign zext_ln69_fu_816_p1 = { 2'h0, icmp_ln1494_reg_1155 };
assign zext_ln703_fu_507_p1 = { 4'h0, signbit_fu_449_p2, 1'h0 };
assign zext_ln727_fu_767_p1 = { 1'h0, op_2 };
assign zext_ln787_fu_774_p1 = { 3'h0, ret_V_18_fu_757_p3 };
assign \mul_16s_2s_18_1_1_U1.top_mul_16s_2s_18_1_1_Multiplier_0_U.a  = \mul_16s_2s_18_1_1_U1.din0 ;
assign \mul_16s_2s_18_1_1_U1.top_mul_16s_2s_18_1_1_Multiplier_0_U.b  = \mul_16s_2s_18_1_1_U1.din1 ;
assign \mul_16s_2s_18_1_1_U1.dout  = \mul_16s_2s_18_1_1_U1.top_mul_16s_2s_18_1_1_Multiplier_0_U.p ;
assign \mul_16s_2s_18_1_1_U1.din0  = op_4;
assign \mul_16s_2s_18_1_1_U1.din1  = op_7;
assign r_V_1_fu_419_p2 = \mul_16s_2s_18_1_1_U1.dout ;
endmodule


// Product machine:
module top_A_times_top_B (ap_start, op_0, op_1, op_13, op_15, op_16, op_17, op_2, op_3, op_4, op_5, op_7, op_8, ap_clk, unsafe_signal);
input ap_start;
input [1:0] op_0;
input [7:0] op_1;
input [7:0] op_13;
input [7:0] op_15;
input [3:0] op_16;
input [3:0] op_17;
input [1:0] op_2;
input [7:0] op_3;
input [15:0] op_4;
input [3:0] op_5;
input [1:0] op_7;
input [1:0] op_8;
input ap_clk;
output unsafe_signal;
reg _setup;
initial _setup = 1'b0;
always @ (posedge ap_clk) _setup <= 1'b1;
reg ap_start_internal;
always @ (posedge ap_clk) if (!_setup) ap_start_internal <= ap_start;
reg [1:0] op_0_internal;
always @ (posedge ap_clk) if (!_setup) op_0_internal <= op_0;
reg [7:0] op_1_internal;
always @ (posedge ap_clk) if (!_setup) op_1_internal <= op_1;
reg [7:0] op_13_internal;
always @ (posedge ap_clk) if (!_setup) op_13_internal <= op_13;
reg [7:0] op_15_internal;
always @ (posedge ap_clk) if (!_setup) op_15_internal <= op_15;
reg [3:0] op_16_internal;
always @ (posedge ap_clk) if (!_setup) op_16_internal <= op_16;
reg [3:0] op_17_internal;
always @ (posedge ap_clk) if (!_setup) op_17_internal <= op_17;
reg [1:0] op_2_internal;
always @ (posedge ap_clk) if (!_setup) op_2_internal <= op_2;
reg [7:0] op_3_internal;
always @ (posedge ap_clk) if (!_setup) op_3_internal <= op_3;
reg [15:0] op_4_internal;
always @ (posedge ap_clk) if (!_setup) op_4_internal <= op_4;
reg [3:0] op_5_internal;
always @ (posedge ap_clk) if (!_setup) op_5_internal <= op_5;
reg [1:0] op_7_internal;
always @ (posedge ap_clk) if (!_setup) op_7_internal <= op_7;
reg [1:0] op_8_internal;
always @ (posedge ap_clk) if (!_setup) op_8_internal <= op_8;
wire ap_done_A;
wire ap_done_B;
wire ap_done_eq;
assign ap_done_eq = ap_done_A == ap_done_B;
wire ap_idle_A;
wire ap_idle_B;
wire ap_idle_eq;
assign ap_idle_eq = ap_idle_A == ap_idle_B;
wire ap_ready_A;
wire ap_ready_B;
wire ap_ready_eq;
assign ap_ready_eq = ap_ready_A == ap_ready_B;
wire [31:0] op_30_A;
wire [31:0] op_30_B;
wire op_30_eq;
assign op_30_eq = op_30_A == op_30_B;
wire op_30_ap_vld_A;
wire op_30_ap_vld_B;
wire clk_enable_A;
wire clk_enable_B;
assign clk_enable_A = _setup & (~op_30_ap_vld_A | op_30_ap_vld_B);
assign clk_enable_B = _setup;
wire divergent;
assign divergent = ~(ap_done_eq & ap_idle_eq & ap_ready_eq & op_30_eq);
assign unsafe_signal = op_30_ap_vld_A & op_30_ap_vld_B & divergent;
top_A instance_A (
    .ap_clk(ap_clk),
    .clk_enable(clk_enable_A),
    .ap_start(ap_start_internal),
    .op_0(op_0_internal),
    .op_1(op_1_internal),
    .op_13(op_13_internal),
    .op_15(op_15_internal),
    .op_16(op_16_internal),
    .op_17(op_17_internal),
    .op_2(op_2_internal),
    .op_3(op_3_internal),
    .op_4(op_4_internal),
    .op_5(op_5_internal),
    .op_7(op_7_internal),
    .op_8(op_8_internal),
    .ap_done(ap_done_A),
    .ap_idle(ap_idle_A),
    .ap_ready(ap_ready_A),
    .op_30(op_30_A),
    .op_30_ap_vld(op_30_ap_vld_A)
);
top_B instance_B (
    .ap_clk(ap_clk),
    .clk_enable(clk_enable_B),
    .ap_start(ap_start_internal),
    .op_0(op_0_internal),
    .op_1(op_1_internal),
    .op_13(op_13_internal),
    .op_15(op_15_internal),
    .op_16(op_16_internal),
    .op_17(op_17_internal),
    .op_2(op_2_internal),
    .op_3(op_3_internal),
    .op_4(op_4_internal),
    .op_5(op_5_internal),
    .op_7(op_7_internal),
    .op_8(op_8_internal),
    .ap_done(ap_done_B),
    .ap_idle(ap_idle_B),
    .ap_ready(ap_ready_B),
    .op_30(op_30_B),
    .op_30_ap_vld(op_30_ap_vld_B)
);
endmodule
