// Processed by function `construct_kairos` in `verilog_tricks.py`.
// Machine A:
// Processed by function `add_clk_enable_signal` in `verilog_tricks.py`.
// Processed by function `remove_reset_signal` in `verilog_tricks.py`.
module top_A (
  ap_clk,
  ap_start,
  ap_done,
  ap_idle,
  ap_ready,
  op_0,
  op_1,
  op_2,
  op_3,
  op_7,
  op_8,
  op_13,
  op_16,
  op_17,
  op_29,
  op_29_ap_vld,
clk_enable
);
input clk_enable;


input ap_clk;
wire ap_rst;
assign ap_rst = op_29_ap_vld;
input ap_start;
input [7:0] op_0;
input op_1;
input [31:0] op_13;
input [7:0] op_16;
input [7:0] op_17;
input [3:0] op_2;
input [31:0] op_3;
input [3:0] op_7;
input [31:0] op_8;
output ap_done;
output ap_idle;
output ap_ready;
output [31:0] op_29;
output op_29_ap_vld;


reg [31:0] add_ln691_3_reg_1222;
reg [31:0] add_ln691_4_reg_1253;
reg and_ln786_1_reg_1146;
reg [8:0] ap_CS_fsm = 9'h001;
reg [9:0] empty_reg_1056;
reg icmp_ln851_2_reg_1168;
reg icmp_ln851_3_reg_1196;
reg icmp_ln851_4_reg_1217;
reg icmp_ln851_5_reg_1248;
reg icmp_ln851_reg_1115;
reg icmp_ln878_reg_1068;
reg [2:0] op_10_V_reg_1125;
reg [3:0] op_18_V_reg_1227;
reg [31:0] op_25_V_reg_1201;
reg or_ln785_1_reg_1136;
reg p_Result_13_reg_1074;
reg p_Result_14_reg_1091;
reg [24:0] p_Result_s_20_reg_1098;
reg [15:0] p_Val2_3_reg_1130;
reg [8:0] ret_V_16_reg_1104;
reg [1:0] ret_V_18_reg_1061;
reg [39:0] ret_V_19_reg_1156;
reg [52:0] ret_V_21_reg_1184;
reg [31:0] ret_V_22_cast_reg_1189;
reg [37:0] ret_V_23_reg_1206;
reg [31:0] ret_V_24_cast_reg_1211;
reg [38:0] ret_V_24_reg_1237;
reg [31:0] ret_V_26_cast_reg_1242;
reg [3:0] ret_V_2_reg_1120;
reg [31:0] ret_V_8_cast_reg_1161;
reg [3:0] ret_V_reg_1109;
reg sel_tmp18_reg_1151;
reg [15:0] select_ln340_1_reg_1141;
reg [31:0] tmp_2_reg_1178;
reg tmp_3_reg_1080;
reg [8:0] trunc_ln1346_reg_1086;
reg [3:0] trunc_ln2_reg_1232;
reg [32:0] _118_;
wire [31:0] _000_;
wire [31:0] _001_;
wire _002_;
wire [8:0] _003_;
wire [9:0] _004_;
wire _005_;
wire _006_;
wire _007_;
wire _008_;
wire _009_;
wire _010_;
wire [1:0] _011_;
wire [3:0] _012_;
wire [31:0] _013_;
wire _014_;
wire _015_;
wire _016_;
wire [24:0] _017_;
wire [8:0] _018_;
wire [8:0] _019_;
wire [1:0] _020_;
wire [39:0] _021_;
wire [32:0] _022_;
wire [52:0] _023_;
wire [31:0] _024_;
wire [37:0] _025_;
wire [31:0] _026_;
wire [38:0] _027_;
wire [31:0] _028_;
wire [3:0] _029_;
wire [31:0] _030_;
wire [3:0] _031_;
wire _032_;
wire [15:0] _033_;
wire [31:0] _034_;
wire _035_;
wire [8:0] _036_;
wire [3:0] _037_;
wire [1:0] _038_;
wire _039_;
wire _040_;
wire _041_;
wire _042_;
wire _043_;
wire _044_;
wire _045_;
wire _046_;
wire _047_;
wire _048_;
wire _049_;
wire _050_;
wire _051_;
wire _052_;
wire _053_;
wire _054_;
wire _055_;
wire _056_;
wire _057_;
wire _058_;
wire _059_;
wire [9:0] add_ln1346_1_fu_428_p2;
wire [31:0] add_ln691_2_fu_834_p2;
wire [31:0] add_ln691_3_fu_903_p2;
wire [31:0] add_ln691_4_fu_1012_p2;
wire [31:0] add_ln691_fu_711_p2;
wire [8:0] add_ln731_fu_433_p2;
wire [31:0] add_ln850_fu_764_p2;
wire and_ln340_1_fu_582_p2;
wire and_ln340_fu_556_p2;
wire and_ln785_1_fu_588_p2;
wire and_ln785_fu_645_p2;
wire and_ln786_1_fu_576_p2;
wire and_ln786_fu_405_p2;
wire ap_CS_fsm_state1;
wire ap_CS_fsm_state2;
wire ap_CS_fsm_state3;
wire ap_CS_fsm_state4;
wire ap_CS_fsm_state5;
wire ap_CS_fsm_state6;
wire ap_CS_fsm_state7;
wire ap_CS_fsm_state8;
wire ap_CS_fsm_state9;
wire [8:0] ap_NS_fsm;
wire ap_clk;
wire ap_done;
wire ap_idle;
wire ap_ready;
wire ap_rst;
wire ap_start;
wire [9:0] empty_fu_231_p1;
wire icmp_ln768_fu_462_p2;
wire icmp_ln786_fu_490_p2;
wire icmp_ln851_1_fu_257_p2;
wire icmp_ln851_2_fu_698_p2;
wire icmp_ln851_3_fu_812_p2;
wire icmp_ln851_4_fu_897_p2;
wire icmp_ln851_5_fu_1006_p2;
wire icmp_ln851_fu_379_p2;
wire icmp_ln878_fu_289_p2;
wire [7:0] op_0;
wire op_1;
wire [2:0] op_10_V_fu_417_p3;
wire [15:0] op_11_V_fu_656_p3;
wire [31:0] op_13;
wire [4:0] op_14_V_fu_915_p3;
wire [7:0] op_16;
wire [7:0] op_17;
wire [3:0] op_18_V_fu_926_p2;
wire [3:0] op_2;
wire [31:0] op_21_V_fu_629_p2;
wire [31:0] op_25_V_fu_856_p2;
wire [31:0] op_28_V_fu_1040_p2;
wire [31:0] op_29;
wire op_29_ap_vld;
wire [31:0] op_3;
wire [3:0] op_7;
wire [31:0] op_8;
wire or_ln340_fu_501_p2;
wire or_ln785_1_fu_467_p2;
wire or_ln785_2_fu_640_p2;
wire or_ln785_3_fu_594_p2;
wire or_ln785_fu_401_p2;
wire or_ln786_fu_495_p2;
wire overflow_fu_478_p2;
wire p_Result_10_fu_827_p3;
wire p_Result_11_fu_951_p3;
wire p_Result_12_fu_1018_p3;
wire p_Result_15_fu_446_p3;
wire p_Result_16_fu_454_p3;
wire p_Result_1_fu_245_p3;
wire [15:0] p_Result_7_fu_540_p4;
wire p_Result_8_fu_704_p3;
wire p_Result_9_fu_757_p3;
wire p_Result_s_fu_606_p3;
wire [2:0] p_Val2_1_fu_394_p3;
wire [15:0] p_Val2_3_fu_438_p3;
wire [14:0] p_Val2_4_fu_534_p2;
wire [3:0] r_2_fu_909_p2;
wire [1:0] r_fu_821_p2;
wire [8:0] ret_V_16_fu_359_p2;
wire [3:0] ret_V_17_fu_618_p3;
wire [1:0] ret_V_18_fu_277_p3;
wire [39:0] ret_V_19_fu_678_p2;
wire [33:0] ret_V_20_fu_741_p2;
wire [33:0] ret_V_20_reg_1173;
wire [52:0] ret_V_21_fu_792_p2;
wire [31:0] ret_V_22_fu_845_p3;
wire [37:0] ret_V_23_fu_877_p2;
wire [31:0] ret_V_24_cast_fu_883_p4;
wire [38:0] ret_V_24_fu_986_p2;
wire [31:0] ret_V_25_fu_1030_p3;
wire [31:0] ret_V_26_cast_fu_992_p4;
wire [3:0] ret_V_2_fu_385_p2;
wire [1:0] ret_V_3_fu_235_p4;
wire [1:0] ret_V_5_fu_263_p2;
wire [4:0] ret_V_7_fu_935_p2;
wire [3:0] ret_V_fu_365_p4;
wire [33:0] ret_fu_323_p2;
wire [38:0] rhs_3_fu_666_p3;
wire [32:0] rhs_4_fu_729_p3;
wire [51:0] rhs_5_fu_780_p3;
wire [36:0] rhs_7_fu_866_p3;
wire [37:0] rhs_8_fu_974_p3;
wire sel_tmp18_fu_600_p2;
wire select_ln1192_fu_351_p0;
wire [8:0] select_ln1192_fu_351_p3;
wire [15:0] select_ln340_1_fu_562_p3;
wire [2:0] select_ln340_fu_409_p3;
wire [31:0] select_ln353_2_fu_967_p3;
wire [31:0] select_ln353_fu_722_p3;
wire [15:0] select_ln785_fu_650_p3;
wire [1:0] select_ln850_1_fu_269_p3;
wire [31:0] select_ln850_4_fu_839_p3;
wire [31:0] select_ln850_5_fu_716_p3;
wire [31:0] select_ln850_6_fu_1025_p3;
wire [31:0] select_ln850_7_fu_773_p3;
wire [31:0] select_ln850_8_fu_962_p3;
wire [3:0] select_ln850_fu_613_p3;
wire [33:0] sext_ln1192_1_fu_737_p1;
wire [52:0] sext_ln1192_2_fu_788_p1;
wire [37:0] sext_ln1192_3_fu_873_p1;
wire [38:0] sext_ln1192_4_fu_982_p1;
wire [31:0] sext_ln1192_5_fu_1046_p1;
wire [39:0] sext_ln1192_fu_674_p1;
wire [4:0] sext_ln1194_fu_932_p1;
wire [8:0] sext_ln1346_fu_425_p1;
wire [33:0] sext_ln215_fu_315_p1;
wire [31:0] sext_ln353_fu_625_p1;
wire [31:0] sext_ln69_fu_1037_p1;
wire [39:0] sext_ln703_1_fu_662_p1;
wire [31:0] sext_ln703_2_fu_769_p0;
wire [52:0] sext_ln703_2_fu_769_p1;
wire [7:0] sext_ln703_3_fu_862_p0;
wire [37:0] sext_ln703_3_fu_862_p1;
wire [7:0] sext_ln703_4_fu_958_p0;
wire [38:0] sext_ln703_4_fu_958_p1;
wire [8:0] sext_ln703_fu_347_p1;
wire [31:0] sext_ln870_fu_285_p1;
wire [9:0] sext_ln878_fu_391_p1;
wire tmp_7_fu_506_p3;
wire tmp_8_fu_514_p3;
wire [8:0] trunc_ln1346_fu_319_p1;
wire [1:0] trunc_ln851_1_fu_253_p1;
wire [6:0] trunc_ln851_2_fu_694_p1;
wire [31:0] trunc_ln851_3_fu_808_p0;
wire [19:0] trunc_ln851_3_fu_808_p1;
wire [7:0] trunc_ln851_4_fu_893_p0;
wire [4:0] trunc_ln851_4_fu_893_p1;
wire [7:0] trunc_ln851_5_fu_1002_p0;
wire [5:0] trunc_ln851_5_fu_1002_p1;
wire [4:0] trunc_ln851_fu_375_p1;
wire xor_ln340_fu_550_p2;
wire xor_ln365_1_fu_528_p2;
wire xor_ln365_fu_522_p2;
wire xor_ln785_1_fu_635_p2;
wire xor_ln785_fu_473_p2;
wire xor_ln786_1_fu_570_p2;
wire xor_ln786_fu_484_p2;
wire [33:0] zext_ln215_fu_311_p1;
wire [31:0] zext_ln69_1_fu_852_p1;
wire [3:0] zext_ln69_fu_923_p1;
wire [1:0] zext_ln799_fu_818_p1;


assign add_ln1346_1_fu_428_p2 = $signed(empty_reg_1056) + $signed(ret_V_18_reg_1061);
assign add_ln691_2_fu_834_p2 = ret_V_22_cast_reg_1189 + 1'h1;
assign add_ln691_3_fu_903_p2 = ret_V_23_fu_877_p2[36:5] + 1'h1;
assign add_ln691_4_fu_1012_p2 = ret_V_24_fu_986_p2[37:6] + 1'h1;
assign add_ln691_fu_711_p2 = ret_V_8_cast_reg_1161 + 1'h1;
assign add_ln731_fu_433_p2 = $signed(trunc_ln1346_reg_1086) + $signed(ret_V_18_reg_1061);
assign add_ln850_fu_764_p2 = tmp_2_reg_1178 + 1'h1;
assign op_18_V_fu_926_p2 = icmp_ln878_reg_1068 + op_7;
assign op_21_V_fu_629_p2 = $signed(ret_V_17_fu_618_p3) + $signed(op_8);
assign op_25_V_fu_856_p2 = ret_V_22_fu_845_p3 + r_fu_821_p2;
assign op_28_V_fu_1040_p2 = $signed(ret_V_25_fu_1030_p3) + $signed(op_18_V_reg_1227);
assign op_29 = $signed(op_28_V_fu_1040_p2) + $signed(trunc_ln2_reg_1232);
assign ret_V_16_fu_359_p2 = $signed(select_ln1192_fu_351_p3) + $signed(op_0);
assign ret_V_19_fu_678_p2 = $signed({ op_21_V_fu_629_p2, 7'h00 }) + $signed(op_11_V_fu_656_p3);
assign ret_V_20_fu_741_p2 = $signed({ select_ln353_fu_722_p3, 1'h0 }) + $signed(1'h1);
assign ret_V_21_fu_792_p2 = $signed({ select_ln850_7_fu_773_p3, 20'h00000 }) + $signed(op_13);
assign ret_V_23_fu_877_p2 = $signed({ op_25_V_reg_1201, 5'h00 }) + $signed(op_16);
assign ret_V_24_fu_986_p2 = $signed({ select_ln353_2_fu_967_p3, 6'h00 }) + $signed(op_17);
assign ret_V_2_fu_385_p2 = ret_V_16_fu_359_p2[8:5] + 1'h1;
assign ret_V_5_fu_263_p2 = op_2[3:2] + 1'h1;
assign ret_fu_323_p2 = $signed({ 1'h0, op_3 }) + $signed(ret_V_18_fu_277_p3);
assign _039_ = ap_CS_fsm[0] & _041_;
assign _040_ = ap_CS_fsm[0] & ap_start;
assign and_ln340_1_fu_582_p2 = or_ln786_fu_495_p2 & or_ln340_fu_501_p2;
assign and_ln340_fu_556_p2 = xor_ln340_fu_550_p2 & or_ln786_fu_495_p2;
assign and_ln785_1_fu_588_p2 = xor_ln785_fu_473_p2 & and_ln786_1_fu_576_p2;
assign and_ln785_fu_645_p2 = or_ln785_2_fu_640_p2 & and_ln786_1_reg_1146;
assign and_ln786_1_fu_576_p2 = xor_ln786_1_fu_570_p2 & add_ln731_fu_433_p2[8];
assign and_ln786_fu_405_p2 = tmp_3_reg_1080 & p_Result_13_reg_1074;
assign overflow_fu_478_p2 = xor_ln785_fu_473_p2 & or_ln785_1_fu_467_p2;
assign ret_V_7_fu_935_p2 = { op_10_V_reg_1125[2], op_10_V_reg_1125[2], op_10_V_reg_1125 } & { r_2_fu_909_p2, 1'h0 };
assign sel_tmp18_fu_600_p2 = xor_ln365_1_fu_528_p2 & or_ln785_3_fu_594_p2;
assign xor_ln785_fu_473_p2 = ~ p_Result_14_reg_1091;
assign xor_ln786_fu_484_p2 = ~ add_ln731_fu_433_p2[8];
assign xor_ln340_fu_550_p2 = ~ or_ln340_fu_501_p2;
assign xor_ln786_1_fu_570_p2 = ~ icmp_ln786_fu_490_p2;
assign xor_ln785_1_fu_635_p2 = ~ or_ln785_1_reg_1136;
assign xor_ln365_1_fu_528_p2 = ~ xor_ln365_fu_522_p2;
assign p_Val2_4_fu_534_p2 = ~ { add_ln731_fu_433_p2[7:0], 7'h00 };
assign r_2_fu_909_p2 = ~ op_7;
assign _041_ = ~ ap_start;
assign _042_ = ! op_2[1:0];
assign _043_ = ! ret_V_16_fu_359_p2[4:0];
assign _044_ = { ret_V_18_fu_277_p3[1], ret_V_18_fu_277_p3[1], ret_V_18_fu_277_p3[1], ret_V_18_fu_277_p3[1], ret_V_18_fu_277_p3[1], ret_V_18_fu_277_p3[1], ret_V_18_fu_277_p3[1], ret_V_18_fu_277_p3[1], ret_V_18_fu_277_p3[1], ret_V_18_fu_277_p3[1], ret_V_18_fu_277_p3[1], ret_V_18_fu_277_p3[1], ret_V_18_fu_277_p3[1], ret_V_18_fu_277_p3[1], ret_V_18_fu_277_p3[1], ret_V_18_fu_277_p3[1], ret_V_18_fu_277_p3[1], ret_V_18_fu_277_p3[1], ret_V_18_fu_277_p3[1], ret_V_18_fu_277_p3[1], ret_V_18_fu_277_p3[1], ret_V_18_fu_277_p3[1], ret_V_18_fu_277_p3[1], ret_V_18_fu_277_p3[1], ret_V_18_fu_277_p3[1], ret_V_18_fu_277_p3[1], ret_V_18_fu_277_p3[1], ret_V_18_fu_277_p3[1], ret_V_18_fu_277_p3[1], ret_V_18_fu_277_p3[1], ret_V_18_fu_277_p3 } > op_3;
assign _045_ = | p_Result_s_20_reg_1098;
assign _046_ = p_Result_s_20_reg_1098 != 25'h1ffffff;
assign _047_ = | op_11_V_fu_656_p3[6:0];
assign _048_ = | op_13[19:0];
assign _049_ = | op_16[4:0];
assign _050_ = | op_17[5:0];
assign or_ln340_fu_501_p2 = p_Result_14_reg_1091 | overflow_fu_478_p2;
assign or_ln785_1_fu_467_p2 = add_ln731_fu_433_p2[8] | icmp_ln768_fu_462_p2;
assign or_ln785_2_fu_640_p2 = xor_ln785_1_fu_635_p2 | p_Result_14_reg_1091;
assign or_ln785_3_fu_594_p2 = and_ln785_1_fu_588_p2 | and_ln340_1_fu_582_p2;
assign or_ln785_fu_401_p2 = tmp_3_reg_1080 | p_Result_13_reg_1074;
assign or_ln786_fu_495_p2 = xor_ln786_fu_484_p2 | icmp_ln786_fu_490_p2;
always @(posedge ap_clk)
op_10_V_reg_1125[0] <= 1'h0;
always @(posedge ap_clk)
p_Val2_3_reg_1130[6:0] <= 7'h00;
always @(posedge ap_clk)
_118_ <= _022_;
assign ret_V_20_reg_1173[33:1] = _118_;
always @(posedge ap_clk)
tmp_2_reg_1178 <= _034_;
always @(posedge ap_clk)
op_25_V_reg_1201 <= _013_;
always @(posedge ap_clk)
ret_V_21_reg_1184 <= _023_;
always @(posedge ap_clk)
ret_V_22_cast_reg_1189 <= _024_;
always @(posedge ap_clk)
icmp_ln851_3_reg_1196 <= _006_;
always @(posedge ap_clk)
ret_V_19_reg_1156 <= _021_;
always @(posedge ap_clk)
ret_V_8_cast_reg_1161 <= _030_;
always @(posedge ap_clk)
icmp_ln851_2_reg_1168 <= _005_;
always @(posedge ap_clk)
empty_reg_1056 <= _004_;
always @(posedge ap_clk)
ret_V_18_reg_1061 <= _020_;
always @(posedge ap_clk)
icmp_ln878_reg_1068 <= _010_;
always @(posedge ap_clk)
p_Result_13_reg_1074 <= _015_;
always @(posedge ap_clk)
tmp_3_reg_1080 <= _035_;
always @(posedge ap_clk)
trunc_ln1346_reg_1086 <= _036_;
always @(posedge ap_clk)
p_Result_14_reg_1091 <= _016_;
always @(posedge ap_clk)
p_Result_s_20_reg_1098 <= _017_;
always @(posedge ap_clk)
ret_V_16_reg_1104 <= _019_;
always @(posedge ap_clk)
ret_V_reg_1109 <= _031_;
always @(posedge ap_clk)
icmp_ln851_reg_1115 <= _009_;
always @(posedge ap_clk)
ret_V_2_reg_1120 <= _029_;
always @(posedge ap_clk)
op_10_V_reg_1125[2:1] <= _011_;
always @(posedge ap_clk)
p_Val2_3_reg_1130[15:7] <= _018_;
always @(posedge ap_clk)
or_ln785_1_reg_1136 <= _014_;
always @(posedge ap_clk)
select_ln340_1_reg_1141 <= _033_;
always @(posedge ap_clk)
and_ln786_1_reg_1146 <= _002_;
always @(posedge ap_clk)
sel_tmp18_reg_1151 <= _032_;
always @(posedge ap_clk)
op_18_V_reg_1227 <= _012_;
always @(posedge ap_clk)
trunc_ln2_reg_1232 <= _037_;
always @(posedge ap_clk)
ret_V_24_reg_1237 <= _027_;
always @(posedge ap_clk)
ret_V_26_cast_reg_1242 <= _028_;
always @(posedge ap_clk)
icmp_ln851_5_reg_1248 <= _008_;
always @(posedge ap_clk)
add_ln691_4_reg_1253 <= _001_;
always @(posedge ap_clk)
ret_V_23_reg_1206 <= _025_;
always @(posedge ap_clk)
ret_V_24_cast_reg_1211 <= _026_;
always @(posedge ap_clk)
icmp_ln851_4_reg_1217 <= _007_;
always @(posedge ap_clk)
add_ln691_3_reg_1222 <= _000_;
always @(posedge ap_clk)
ap_CS_fsm <= _003_;
assign _038_ = _040_ ? 2'h2 : 2'h1;
assign _051_ = ap_CS_fsm == 1'h1;
function [8:0] _158_;
input [8:0] a;
input [80:0] b;
input [8:0] s;
case (s)
9'b000000001:
_158_ = b[8:0];
9'b000000010:
_158_ = b[17:9];
9'b000000100:
_158_ = b[26:18];
9'b000001000:
_158_ = b[35:27];
9'b000010000:
_158_ = b[44:36];
9'b000100000:
_158_ = b[53:45];
9'b001000000:
_158_ = b[62:54];
9'b010000000:
_158_ = b[71:63];
9'b100000000:
_158_ = b[80:72];
9'b000000000:
_158_ = a;
default:
_158_ = 9'bx;
endcase
endfunction
assign ap_NS_fsm = _158_(9'hxxx, { 7'h00, _038_, 72'h020202020202020001 }, { _051_, _059_, _058_, _057_, _056_, _055_, _054_, _053_, _052_ });
assign _052_ = ap_CS_fsm == 9'h100;
assign _053_ = ap_CS_fsm == 8'h80;
assign _054_ = ap_CS_fsm == 7'h40;
assign _055_ = ap_CS_fsm == 6'h20;
assign _056_ = ap_CS_fsm == 5'h10;
assign _057_ = ap_CS_fsm == 4'h8;
assign _058_ = ap_CS_fsm == 3'h4;
assign _059_ = ap_CS_fsm == 2'h2;
assign op_29_ap_vld = ap_CS_fsm[8] ? 1'h1 : 1'h0;
assign ap_idle = _039_ ? 1'h1 : 1'h0;
assign _034_ = ap_CS_fsm[3] ? ret_V_20_fu_741_p2[32:1] : tmp_2_reg_1178;
assign _022_ = ap_CS_fsm[3] ? ret_V_20_fu_741_p2[33:1] : ret_V_20_reg_1173[33:1];
assign _013_ = ap_CS_fsm[5] ? op_25_V_fu_856_p2 : op_25_V_reg_1201;
assign _006_ = ap_CS_fsm[4] ? icmp_ln851_3_fu_812_p2 : icmp_ln851_3_reg_1196;
assign _024_ = ap_CS_fsm[4] ? ret_V_21_fu_792_p2[51:20] : ret_V_22_cast_reg_1189;
assign _023_ = ap_CS_fsm[4] ? ret_V_21_fu_792_p2 : ret_V_21_reg_1184;
assign _005_ = ap_CS_fsm[2] ? icmp_ln851_2_fu_698_p2 : icmp_ln851_2_reg_1168;
assign _030_ = ap_CS_fsm[2] ? ret_V_19_fu_678_p2[38:7] : ret_V_8_cast_reg_1161;
assign _021_ = ap_CS_fsm[2] ? ret_V_19_fu_678_p2 : ret_V_19_reg_1156;
assign _017_ = ap_CS_fsm[0] ? ret_fu_323_p2[33:9] : p_Result_s_20_reg_1098;
assign _016_ = ap_CS_fsm[0] ? ret_fu_323_p2[33] : p_Result_14_reg_1091;
assign _036_ = ap_CS_fsm[0] ? op_3[8:0] : trunc_ln1346_reg_1086;
assign _035_ = ap_CS_fsm[0] ? ret_V_18_fu_277_p3[1] : tmp_3_reg_1080;
assign _015_ = ap_CS_fsm[0] ? ret_V_18_fu_277_p3[1] : p_Result_13_reg_1074;
assign _010_ = ap_CS_fsm[0] ? icmp_ln878_fu_289_p2 : icmp_ln878_reg_1068;
assign _020_ = ap_CS_fsm[0] ? ret_V_18_fu_277_p3 : ret_V_18_reg_1061;
assign _004_ = ap_CS_fsm[0] ? op_3[9:0] : empty_reg_1056;
assign _032_ = ap_CS_fsm[1] ? sel_tmp18_fu_600_p2 : sel_tmp18_reg_1151;
assign _002_ = ap_CS_fsm[1] ? and_ln786_1_fu_576_p2 : and_ln786_1_reg_1146;
assign _033_ = ap_CS_fsm[1] ? select_ln340_1_fu_562_p3 : select_ln340_1_reg_1141;
assign _014_ = ap_CS_fsm[1] ? or_ln785_1_fu_467_p2 : or_ln785_1_reg_1136;
assign _018_ = ap_CS_fsm[1] ? add_ln731_fu_433_p2 : p_Val2_3_reg_1130[15:7];
assign _011_ = ap_CS_fsm[1] ? op_10_V_fu_417_p3[2:1] : op_10_V_reg_1125[2:1];
assign _029_ = ap_CS_fsm[1] ? ret_V_2_fu_385_p2 : ret_V_2_reg_1120;
assign _009_ = ap_CS_fsm[1] ? icmp_ln851_fu_379_p2 : icmp_ln851_reg_1115;
assign _031_ = ap_CS_fsm[1] ? ret_V_16_fu_359_p2[8:5] : ret_V_reg_1109;
assign _019_ = ap_CS_fsm[1] ? ret_V_16_fu_359_p2 : ret_V_16_reg_1104;
assign _001_ = ap_CS_fsm[7] ? add_ln691_4_fu_1012_p2 : add_ln691_4_reg_1253;
assign _008_ = ap_CS_fsm[7] ? icmp_ln851_5_fu_1006_p2 : icmp_ln851_5_reg_1248;
assign _028_ = ap_CS_fsm[7] ? ret_V_24_fu_986_p2[37:6] : ret_V_26_cast_reg_1242;
assign _027_ = ap_CS_fsm[7] ? ret_V_24_fu_986_p2 : ret_V_24_reg_1237;
assign _037_ = ap_CS_fsm[7] ? ret_V_7_fu_935_p2[4:1] : trunc_ln2_reg_1232;
assign _012_ = ap_CS_fsm[7] ? op_18_V_fu_926_p2 : op_18_V_reg_1227;
assign _000_ = ap_CS_fsm[6] ? add_ln691_3_fu_903_p2 : add_ln691_3_reg_1222;
assign _007_ = ap_CS_fsm[6] ? icmp_ln851_4_fu_897_p2 : icmp_ln851_4_reg_1217;
assign _026_ = ap_CS_fsm[6] ? ret_V_23_fu_877_p2[36:5] : ret_V_24_cast_reg_1211;
assign _025_ = ap_CS_fsm[6] ? ret_V_23_fu_877_p2 : ret_V_23_reg_1206;
assign _003_ = ap_rst ? 9'h001 : ap_NS_fsm;
assign r_fu_821_p2 = icmp_ln878_reg_1068 >> icmp_ln878_reg_1068;
assign icmp_ln768_fu_462_p2 = _045_ ? 1'h1 : 1'h0;
assign icmp_ln786_fu_490_p2 = _046_ ? 1'h1 : 1'h0;
assign icmp_ln851_1_fu_257_p2 = _042_ ? 1'h1 : 1'h0;
assign icmp_ln851_2_fu_698_p2 = _047_ ? 1'h1 : 1'h0;
assign icmp_ln851_3_fu_812_p2 = _048_ ? 1'h1 : 1'h0;
assign icmp_ln851_4_fu_897_p2 = _049_ ? 1'h1 : 1'h0;
assign icmp_ln851_5_fu_1006_p2 = _050_ ? 1'h1 : 1'h0;
assign icmp_ln851_fu_379_p2 = _043_ ? 1'h1 : 1'h0;
assign icmp_ln878_fu_289_p2 = _044_ ? 1'h1 : 1'h0;
assign op_10_V_fu_417_p3 = and_ln786_fu_405_p2 ? { ret_V_18_reg_1061, 1'h0 } : select_ln340_fu_409_p3;
assign op_11_V_fu_656_p3 = sel_tmp18_reg_1151 ? p_Val2_3_reg_1130 : select_ln785_fu_650_p3;
assign ret_V_17_fu_618_p3 = ret_V_16_reg_1104[8] ? select_ln850_fu_613_p3 : ret_V_reg_1109;
assign ret_V_18_fu_277_p3 = op_2[3] ? select_ln850_1_fu_269_p3 : { 1'h0, op_2[2] };
assign ret_V_22_fu_845_p3 = ret_V_21_reg_1184[52] ? select_ln850_4_fu_839_p3 : ret_V_22_cast_reg_1189;
assign ret_V_25_fu_1030_p3 = ret_V_24_reg_1237[38] ? select_ln850_6_fu_1025_p3 : ret_V_26_cast_reg_1242;
assign select_ln1192_fu_351_p3 = op_1 ? 9'h1e0 : 9'h000;
assign select_ln340_1_fu_562_p3 = and_ln340_fu_556_p2 ? { add_ln731_fu_433_p2, 7'h00 } : { add_ln1346_1_fu_428_p2[9], p_Val2_4_fu_534_p2 };
assign select_ln340_fu_409_p3 = or_ln785_fu_401_p2 ? 3'h0 : { ret_V_18_reg_1061, 1'h0 };
assign select_ln353_2_fu_967_p3 = ret_V_23_reg_1206[37] ? select_ln850_8_fu_962_p3 : ret_V_24_cast_reg_1211;
assign select_ln353_fu_722_p3 = ret_V_19_reg_1156[39] ? select_ln850_5_fu_716_p3 : ret_V_8_cast_reg_1161;
assign select_ln785_fu_650_p3 = and_ln785_fu_645_p2 ? p_Val2_3_reg_1130 : select_ln340_1_reg_1141;
assign select_ln850_1_fu_269_p3 = icmp_ln851_1_fu_257_p2 ? { 1'h1, op_2[2] } : ret_V_5_fu_263_p2;
assign select_ln850_4_fu_839_p3 = icmp_ln851_3_reg_1196 ? add_ln691_2_fu_834_p2 : ret_V_22_cast_reg_1189;
assign select_ln850_5_fu_716_p3 = icmp_ln851_2_reg_1168 ? add_ln691_fu_711_p2 : ret_V_8_cast_reg_1161;
assign select_ln850_6_fu_1025_p3 = icmp_ln851_5_reg_1248 ? add_ln691_4_reg_1253 : ret_V_26_cast_reg_1242;
assign select_ln850_7_fu_773_p3 = ret_V_20_reg_1173[33] ? add_ln850_fu_764_p2 : tmp_2_reg_1178;
assign select_ln850_8_fu_962_p3 = icmp_ln851_4_reg_1217 ? add_ln691_3_reg_1222 : ret_V_24_cast_reg_1211;
assign select_ln850_fu_613_p3 = icmp_ln851_reg_1115 ? ret_V_reg_1109 : ret_V_2_reg_1120;
assign xor_ln365_fu_522_p2 = add_ln731_fu_433_p2[8] ^ add_ln1346_1_fu_428_p2[9];
assign ap_CS_fsm_state1 = ap_CS_fsm[0];
assign ap_CS_fsm_state2 = ap_CS_fsm[1];
assign ap_CS_fsm_state3 = ap_CS_fsm[2];
assign ap_CS_fsm_state4 = ap_CS_fsm[3];
assign ap_CS_fsm_state5 = ap_CS_fsm[4];
assign ap_CS_fsm_state6 = ap_CS_fsm[5];
assign ap_CS_fsm_state7 = ap_CS_fsm[6];
assign ap_CS_fsm_state8 = ap_CS_fsm[7];
assign ap_CS_fsm_state9 = ap_CS_fsm[8];
assign ap_done = op_29_ap_vld;
assign ap_ready = op_29_ap_vld;
assign empty_fu_231_p1 = op_3[9:0];
assign op_14_V_fu_915_p3 = { r_2_fu_909_p2, 1'h0 };
assign p_Result_10_fu_827_p3 = ret_V_21_reg_1184[52];
assign p_Result_11_fu_951_p3 = ret_V_23_reg_1206[37];
assign p_Result_12_fu_1018_p3 = ret_V_24_reg_1237[38];
assign p_Result_15_fu_446_p3 = add_ln731_fu_433_p2[8];
assign p_Result_16_fu_454_p3 = add_ln1346_1_fu_428_p2[9];
assign p_Result_1_fu_245_p3 = op_2[3];
assign p_Result_7_fu_540_p4 = { add_ln1346_1_fu_428_p2[9], p_Val2_4_fu_534_p2 };
assign p_Result_8_fu_704_p3 = ret_V_19_reg_1156[39];
assign p_Result_9_fu_757_p3 = ret_V_20_reg_1173[33];
assign p_Result_s_fu_606_p3 = ret_V_16_reg_1104[8];
assign p_Val2_1_fu_394_p3 = { ret_V_18_reg_1061, 1'h0 };
assign p_Val2_3_fu_438_p3 = { add_ln731_fu_433_p2, 7'h00 };
assign ret_V_24_cast_fu_883_p4 = ret_V_23_fu_877_p2[36:5];
assign ret_V_26_cast_fu_992_p4 = ret_V_24_fu_986_p2[37:6];
assign ret_V_3_fu_235_p4 = op_2[3:2];
assign ret_V_fu_365_p4 = ret_V_16_fu_359_p2[8:5];
assign rhs_3_fu_666_p3 = { op_21_V_fu_629_p2, 7'h00 };
assign rhs_4_fu_729_p3 = { select_ln353_fu_722_p3, 1'h0 };
assign rhs_5_fu_780_p3 = { select_ln850_7_fu_773_p3, 20'h00000 };
assign rhs_7_fu_866_p3 = { op_25_V_reg_1201, 5'h00 };
assign rhs_8_fu_974_p3 = { select_ln353_2_fu_967_p3, 6'h00 };
assign select_ln1192_fu_351_p0 = op_1;
assign sext_ln1192_1_fu_737_p1 = { select_ln353_fu_722_p3[31], select_ln353_fu_722_p3, 1'h0 };
assign sext_ln1192_2_fu_788_p1 = { select_ln850_7_fu_773_p3[31], select_ln850_7_fu_773_p3, 20'h00000 };
assign sext_ln1192_3_fu_873_p1 = { op_25_V_reg_1201[31], op_25_V_reg_1201, 5'h00 };
assign sext_ln1192_4_fu_982_p1 = { select_ln353_2_fu_967_p3[31], select_ln353_2_fu_967_p3, 6'h00 };
assign sext_ln1192_5_fu_1046_p1 = { trunc_ln2_reg_1232[3], trunc_ln2_reg_1232[3], trunc_ln2_reg_1232[3], trunc_ln2_reg_1232[3], trunc_ln2_reg_1232[3], trunc_ln2_reg_1232[3], trunc_ln2_reg_1232[3], trunc_ln2_reg_1232[3], trunc_ln2_reg_1232[3], trunc_ln2_reg_1232[3], trunc_ln2_reg_1232[3], trunc_ln2_reg_1232[3], trunc_ln2_reg_1232[3], trunc_ln2_reg_1232[3], trunc_ln2_reg_1232[3], trunc_ln2_reg_1232[3], trunc_ln2_reg_1232[3], trunc_ln2_reg_1232[3], trunc_ln2_reg_1232[3], trunc_ln2_reg_1232[3], trunc_ln2_reg_1232[3], trunc_ln2_reg_1232[3], trunc_ln2_reg_1232[3], trunc_ln2_reg_1232[3], trunc_ln2_reg_1232[3], trunc_ln2_reg_1232[3], trunc_ln2_reg_1232[3], trunc_ln2_reg_1232[3], trunc_ln2_reg_1232 };
assign sext_ln1192_fu_674_p1 = { op_21_V_fu_629_p2[31], op_21_V_fu_629_p2, 7'h00 };
assign sext_ln1194_fu_932_p1 = { op_10_V_reg_1125[2], op_10_V_reg_1125[2], op_10_V_reg_1125 };
assign sext_ln1346_fu_425_p1 = { ret_V_18_reg_1061[1], ret_V_18_reg_1061[1], ret_V_18_reg_1061[1], ret_V_18_reg_1061[1], ret_V_18_reg_1061[1], ret_V_18_reg_1061[1], ret_V_18_reg_1061[1], ret_V_18_reg_1061 };
assign sext_ln215_fu_315_p1 = { ret_V_18_fu_277_p3[1], ret_V_18_fu_277_p3[1], ret_V_18_fu_277_p3[1], ret_V_18_fu_277_p3[1], ret_V_18_fu_277_p3[1], ret_V_18_fu_277_p3[1], ret_V_18_fu_277_p3[1], ret_V_18_fu_277_p3[1], ret_V_18_fu_277_p3[1], ret_V_18_fu_277_p3[1], ret_V_18_fu_277_p3[1], ret_V_18_fu_277_p3[1], ret_V_18_fu_277_p3[1], ret_V_18_fu_277_p3[1], ret_V_18_fu_277_p3[1], ret_V_18_fu_277_p3[1], ret_V_18_fu_277_p3[1], ret_V_18_fu_277_p3[1], ret_V_18_fu_277_p3[1], ret_V_18_fu_277_p3[1], ret_V_18_fu_277_p3[1], ret_V_18_fu_277_p3[1], ret_V_18_fu_277_p3[1], ret_V_18_fu_277_p3[1], ret_V_18_fu_277_p3[1], ret_V_18_fu_277_p3[1], ret_V_18_fu_277_p3[1], ret_V_18_fu_277_p3[1], ret_V_18_fu_277_p3[1], ret_V_18_fu_277_p3[1], ret_V_18_fu_277_p3[1], ret_V_18_fu_277_p3[1], ret_V_18_fu_277_p3 };
assign sext_ln353_fu_625_p1 = { ret_V_17_fu_618_p3[3], ret_V_17_fu_618_p3[3], ret_V_17_fu_618_p3[3], ret_V_17_fu_618_p3[3], ret_V_17_fu_618_p3[3], ret_V_17_fu_618_p3[3], ret_V_17_fu_618_p3[3], ret_V_17_fu_618_p3[3], ret_V_17_fu_618_p3[3], ret_V_17_fu_618_p3[3], ret_V_17_fu_618_p3[3], ret_V_17_fu_618_p3[3], ret_V_17_fu_618_p3[3], ret_V_17_fu_618_p3[3], ret_V_17_fu_618_p3[3], ret_V_17_fu_618_p3[3], ret_V_17_fu_618_p3[3], ret_V_17_fu_618_p3[3], ret_V_17_fu_618_p3[3], ret_V_17_fu_618_p3[3], ret_V_17_fu_618_p3[3], ret_V_17_fu_618_p3[3], ret_V_17_fu_618_p3[3], ret_V_17_fu_618_p3[3], ret_V_17_fu_618_p3[3], ret_V_17_fu_618_p3[3], ret_V_17_fu_618_p3[3], ret_V_17_fu_618_p3[3], ret_V_17_fu_618_p3 };
assign sext_ln69_fu_1037_p1 = { op_18_V_reg_1227[3], op_18_V_reg_1227[3], op_18_V_reg_1227[3], op_18_V_reg_1227[3], op_18_V_reg_1227[3], op_18_V_reg_1227[3], op_18_V_reg_1227[3], op_18_V_reg_1227[3], op_18_V_reg_1227[3], op_18_V_reg_1227[3], op_18_V_reg_1227[3], op_18_V_reg_1227[3], op_18_V_reg_1227[3], op_18_V_reg_1227[3], op_18_V_reg_1227[3], op_18_V_reg_1227[3], op_18_V_reg_1227[3], op_18_V_reg_1227[3], op_18_V_reg_1227[3], op_18_V_reg_1227[3], op_18_V_reg_1227[3], op_18_V_reg_1227[3], op_18_V_reg_1227[3], op_18_V_reg_1227[3], op_18_V_reg_1227[3], op_18_V_reg_1227[3], op_18_V_reg_1227[3], op_18_V_reg_1227[3], op_18_V_reg_1227 };
assign sext_ln703_1_fu_662_p1 = { op_11_V_fu_656_p3[15], op_11_V_fu_656_p3[15], op_11_V_fu_656_p3[15], op_11_V_fu_656_p3[15], op_11_V_fu_656_p3[15], op_11_V_fu_656_p3[15], op_11_V_fu_656_p3[15], op_11_V_fu_656_p3[15], op_11_V_fu_656_p3[15], op_11_V_fu_656_p3[15], op_11_V_fu_656_p3[15], op_11_V_fu_656_p3[15], op_11_V_fu_656_p3[15], op_11_V_fu_656_p3[15], op_11_V_fu_656_p3[15], op_11_V_fu_656_p3[15], op_11_V_fu_656_p3[15], op_11_V_fu_656_p3[15], op_11_V_fu_656_p3[15], op_11_V_fu_656_p3[15], op_11_V_fu_656_p3[15], op_11_V_fu_656_p3[15], op_11_V_fu_656_p3[15], op_11_V_fu_656_p3[15], op_11_V_fu_656_p3 };
assign sext_ln703_2_fu_769_p0 = op_13;
assign sext_ln703_2_fu_769_p1 = { op_13[31], op_13[31], op_13[31], op_13[31], op_13[31], op_13[31], op_13[31], op_13[31], op_13[31], op_13[31], op_13[31], op_13[31], op_13[31], op_13[31], op_13[31], op_13[31], op_13[31], op_13[31], op_13[31], op_13[31], op_13[31], op_13 };
assign sext_ln703_3_fu_862_p0 = op_16;
assign sext_ln703_3_fu_862_p1 = { op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16 };
assign sext_ln703_4_fu_958_p0 = op_17;
assign sext_ln703_4_fu_958_p1 = { op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17 };
assign sext_ln703_fu_347_p1 = { op_0[7], op_0 };
assign sext_ln870_fu_285_p1 = { ret_V_18_fu_277_p3[1], ret_V_18_fu_277_p3[1], ret_V_18_fu_277_p3[1], ret_V_18_fu_277_p3[1], ret_V_18_fu_277_p3[1], ret_V_18_fu_277_p3[1], ret_V_18_fu_277_p3[1], ret_V_18_fu_277_p3[1], ret_V_18_fu_277_p3[1], ret_V_18_fu_277_p3[1], ret_V_18_fu_277_p3[1], ret_V_18_fu_277_p3[1], ret_V_18_fu_277_p3[1], ret_V_18_fu_277_p3[1], ret_V_18_fu_277_p3[1], ret_V_18_fu_277_p3[1], ret_V_18_fu_277_p3[1], ret_V_18_fu_277_p3[1], ret_V_18_fu_277_p3[1], ret_V_18_fu_277_p3[1], ret_V_18_fu_277_p3[1], ret_V_18_fu_277_p3[1], ret_V_18_fu_277_p3[1], ret_V_18_fu_277_p3[1], ret_V_18_fu_277_p3[1], ret_V_18_fu_277_p3[1], ret_V_18_fu_277_p3[1], ret_V_18_fu_277_p3[1], ret_V_18_fu_277_p3[1], ret_V_18_fu_277_p3[1], ret_V_18_fu_277_p3 };
assign sext_ln878_fu_391_p1 = { ret_V_18_reg_1061[1], ret_V_18_reg_1061[1], ret_V_18_reg_1061[1], ret_V_18_reg_1061[1], ret_V_18_reg_1061[1], ret_V_18_reg_1061[1], ret_V_18_reg_1061[1], ret_V_18_reg_1061[1], ret_V_18_reg_1061 };
assign tmp_7_fu_506_p3 = add_ln1346_1_fu_428_p2[9];
assign tmp_8_fu_514_p3 = add_ln731_fu_433_p2[8];
assign trunc_ln1346_fu_319_p1 = op_3[8:0];
assign trunc_ln851_1_fu_253_p1 = op_2[1:0];
assign trunc_ln851_2_fu_694_p1 = op_11_V_fu_656_p3[6:0];
assign trunc_ln851_3_fu_808_p0 = op_13;
assign trunc_ln851_3_fu_808_p1 = op_13[19:0];
assign trunc_ln851_4_fu_893_p0 = op_16;
assign trunc_ln851_4_fu_893_p1 = op_16[4:0];
assign trunc_ln851_5_fu_1002_p0 = op_17;
assign trunc_ln851_5_fu_1002_p1 = op_17[5:0];
assign trunc_ln851_fu_375_p1 = ret_V_16_fu_359_p2[4:0];
assign zext_ln215_fu_311_p1 = { 2'h0, op_3 };
assign zext_ln69_1_fu_852_p1 = { 30'h00000000, r_fu_821_p2 };
assign zext_ln69_fu_923_p1 = { 3'h0, icmp_ln878_reg_1068 };
assign zext_ln799_fu_818_p1 = { 1'h0, icmp_ln878_reg_1068 };
endmodule


// Machine B:
// Processed by function `add_clk_enable_signal` in `verilog_tricks.py`.
// Processed by function `remove_reset_signal` in `verilog_tricks.py`.
module top_B (
  ap_clk,
  ap_start,
  ap_done,
  ap_idle,
  ap_ready,
  op_0,
  op_1,
  op_2,
  op_3,
  op_7,
  op_8,
  op_13,
  op_16,
  op_17,
  op_29,
  op_29_ap_vld,
clk_enable
);
input clk_enable;


input ap_clk;
wire ap_rst;
assign ap_rst = op_29_ap_vld;
input ap_start;
input [7:0] op_0;
input op_1;
input [31:0] op_13;
input [7:0] op_16;
input [7:0] op_17;
input [3:0] op_2;
input [31:0] op_3;
input [3:0] op_7;
input [31:0] op_8;
output ap_done;
output ap_idle;
output ap_ready;
output [31:0] op_29;
output op_29_ap_vld;


reg [15:0] \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s1 ;
reg \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.carry_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.sum_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s1 ;
reg \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_7_U.carry_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_7_U.sum_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s1 ;
reg \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.carry_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.sum_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s1 ;
reg \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.carry_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.sum_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s1 ;
reg \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.carry_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.sum_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s1 ;
reg \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.carry_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.sum_s1 ;
reg [15:0] \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_12_U.ain_s1 ;
reg [15:0] \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_12_U.bin_s1 ;
reg \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_12_U.carry_s1 ;
reg [15:0] \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_12_U.sum_s1 ;
reg [15:0] \add_32ns_32s_32_2_1_U21.top_add_32ns_32s_32_2_1_Adder_12_U.ain_s1 ;
reg [15:0] \add_32ns_32s_32_2_1_U21.top_add_32ns_32s_32_2_1_Adder_12_U.bin_s1 ;
reg \add_32ns_32s_32_2_1_U21.top_add_32ns_32s_32_2_1_Adder_12_U.carry_s1 ;
reg [15:0] \add_32ns_32s_32_2_1_U21.top_add_32ns_32s_32_2_1_Adder_12_U.sum_s1 ;
reg [15:0] \add_32s_32ns_32_2_1_U7.top_add_32s_32ns_32_2_1_Adder_5_U.ain_s1 ;
reg [15:0] \add_32s_32ns_32_2_1_U7.top_add_32s_32ns_32_2_1_Adder_5_U.bin_s1 ;
reg \add_32s_32ns_32_2_1_U7.top_add_32s_32ns_32_2_1_Adder_5_U.carry_s1 ;
reg [15:0] \add_32s_32ns_32_2_1_U7.top_add_32s_32ns_32_2_1_Adder_5_U.sum_s1 ;
reg [16:0] \add_34ns_34s_34_2_1_U2.top_add_34ns_34s_34_2_1_Adder_1_U.ain_s1 ;
reg [16:0] \add_34ns_34s_34_2_1_U2.top_add_34ns_34s_34_2_1_Adder_1_U.bin_s1 ;
reg \add_34ns_34s_34_2_1_U2.top_add_34ns_34s_34_2_1_Adder_1_U.carry_s1 ;
reg [16:0] \add_34ns_34s_34_2_1_U2.top_add_34ns_34s_34_2_1_Adder_1_U.sum_s1 ;
reg [16:0] \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_8_U.ain_s1 ;
reg [16:0] \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_8_U.bin_s1 ;
reg \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_8_U.carry_s1 ;
reg [16:0] \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_8_U.sum_s1 ;
reg [18:0] \add_38s_38s_38_2_1_U15.top_add_38s_38s_38_2_1_Adder_10_U.ain_s1 ;
reg [18:0] \add_38s_38s_38_2_1_U15.top_add_38s_38s_38_2_1_Adder_10_U.bin_s1 ;
reg \add_38s_38s_38_2_1_U15.top_add_38s_38s_38_2_1_Adder_10_U.carry_s1 ;
reg [18:0] \add_38s_38s_38_2_1_U15.top_add_38s_38s_38_2_1_Adder_10_U.sum_s1 ;
reg [19:0] \add_39s_39s_39_2_1_U17.top_add_39s_39s_39_2_1_Adder_11_U.ain_s1 ;
reg [19:0] \add_39s_39s_39_2_1_U17.top_add_39s_39s_39_2_1_Adder_11_U.bin_s1 ;
reg \add_39s_39s_39_2_1_U17.top_add_39s_39s_39_2_1_Adder_11_U.carry_s1 ;
reg [18:0] \add_39s_39s_39_2_1_U17.top_add_39s_39s_39_2_1_Adder_11_U.sum_s1 ;
reg [19:0] \add_40s_40s_40_2_1_U8.top_add_40s_40s_40_2_1_Adder_6_U.ain_s1 ;
reg [19:0] \add_40s_40s_40_2_1_U8.top_add_40s_40s_40_2_1_Adder_6_U.bin_s1 ;
reg \add_40s_40s_40_2_1_U8.top_add_40s_40s_40_2_1_Adder_6_U.carry_s1 ;
reg [19:0] \add_40s_40s_40_2_1_U8.top_add_40s_40s_40_2_1_Adder_6_U.sum_s1 ;
reg [26:0] \add_53s_53s_53_2_1_U12.top_add_53s_53s_53_2_1_Adder_9_U.ain_s1 ;
reg [26:0] \add_53s_53s_53_2_1_U12.top_add_53s_53s_53_2_1_Adder_9_U.bin_s1 ;
reg \add_53s_53s_53_2_1_U12.top_add_53s_53s_53_2_1_Adder_9_U.carry_s1 ;
reg [25:0] \add_53s_53s_53_2_1_U12.top_add_53s_53s_53_2_1_Adder_9_U.sum_s1 ;
reg [9:0] add_ln1346_1_reg_1129;
reg [31:0] add_ln691_2_reg_1322;
reg [31:0] add_ln691_3_reg_1374;
reg [31:0] add_ln691_4_reg_1411;
reg [31:0] add_ln691_reg_1259;
reg [8:0] add_ln731_reg_1135;
reg [31:0] add_ln850_reg_1285;
reg and_ln786_1_reg_1186;
reg [38:0] ap_CS_fsm = 39'h0000000001;
reg [9:0] empty_reg_1058;
reg icmp_ln768_reg_1148;
reg icmp_ln786_reg_1153;
reg icmp_ln851_1_reg_1027;
reg icmp_ln851_2_reg_1242;
reg icmp_ln851_3_reg_1305;
reg icmp_ln851_4_reg_1357;
reg icmp_ln851_5_reg_1394;
reg icmp_ln851_reg_1114;
reg icmp_ln878_reg_1063;
reg [2:0] op_10_V_reg_1124;
reg [15:0] op_11_V_reg_1222;
reg [3:0] op_18_V_reg_1416;
reg [31:0] op_21_V_reg_1217;
reg [31:0] op_25_V_reg_1342;
reg [31:0] op_28_V_reg_1436;
reg or_ln340_reg_1180;
reg or_ln785_1_reg_1164;
reg or_ln786_reg_1174;
reg p_Result_13_reg_1046;
reg p_Result_14_reg_1101;
reg p_Result_15_reg_1141;
reg p_Result_9_reg_1274;
reg [24:0] p_Result_s_20_reg_1108;
reg [15:0] p_Val2_3_reg_1202;
reg [1:0] r_reg_1327;
reg [8:0] ret_V_16_reg_1084;
reg [3:0] ret_V_17_reg_1159;
reg [1:0] ret_V_18_reg_1037;
reg [39:0] ret_V_19_reg_1247;
reg [52:0] ret_V_21_reg_1310;
reg [31:0] ret_V_22_cast_reg_1315;
reg [31:0] ret_V_22_reg_1332;
reg [37:0] ret_V_23_reg_1362;
reg [31:0] ret_V_24_cast_reg_1367;
reg [38:0] ret_V_24_reg_1399;
reg [31:0] ret_V_25_reg_1426;
reg [31:0] ret_V_26_cast_reg_1404;
reg [3:0] ret_V_2_reg_1119;
reg [1:0] ret_V_3_reg_1021;
reg [1:0] ret_V_5_reg_1032;
reg [31:0] ret_V_8_cast_reg_1252;
reg [3:0] ret_V_reg_1089;
reg sel_tmp18_reg_1212;
reg [31:0] select_ln353_2_reg_1379;
reg [31:0] select_ln353_reg_1264;
reg [15:0] select_ln785_reg_1207;
reg [31:0] select_ln850_7_reg_1290;
reg [31:0] tmp_2_reg_1279;
reg tmp_3_reg_1052;
reg [8:0] trunc_ln1346_reg_1079;
reg [3:0] trunc_ln2_reg_1421;
reg [6:0] trunc_ln851_2_reg_1227;
reg [4:0] trunc_ln851_reg_1096;
reg xor_ln785_reg_1169;
wire [9:0] _000_;
wire [31:0] _001_;
wire [31:0] _002_;
wire [31:0] _003_;
wire [31:0] _004_;
wire [8:0] _005_;
wire [31:0] _006_;
wire _007_;
wire [38:0] _008_;
wire [9:0] _009_;
wire _010_;
wire _011_;
wire _012_;
wire _013_;
wire _014_;
wire _015_;
wire _016_;
wire _017_;
wire _018_;
wire [1:0] _019_;
wire [15:0] _020_;
wire [3:0] _021_;
wire [31:0] _022_;
wire [31:0] _023_;
wire [31:0] _024_;
wire _025_;
wire _026_;
wire _027_;
wire _028_;
wire _029_;
wire _030_;
wire _031_;
wire [24:0] _032_;
wire [8:0] _033_;
wire [1:0] _034_;
wire [8:0] _035_;
wire [3:0] _036_;
wire [1:0] _037_;
wire [39:0] _038_;
wire [52:0] _039_;
wire [31:0] _040_;
wire [31:0] _041_;
wire [37:0] _042_;
wire [31:0] _043_;
wire [38:0] _044_;
wire [31:0] _045_;
wire [31:0] _046_;
wire [3:0] _047_;
wire [1:0] _048_;
wire [1:0] _049_;
wire [31:0] _050_;
wire [3:0] _051_;
wire _052_;
wire [31:0] _053_;
wire [31:0] _054_;
wire [15:0] _055_;
wire [31:0] _056_;
wire [31:0] _057_;
wire _058_;
wire [8:0] _059_;
wire [3:0] _060_;
wire [6:0] _061_;
wire [4:0] _062_;
wire _063_;
wire [1:0] _064_;
wire _065_;
wire _066_;
wire _067_;
wire _068_;
wire _069_;
wire _070_;
wire _071_;
wire _072_;
wire _073_;
wire _074_;
wire [15:0] _075_;
wire [15:0] _076_;
wire _077_;
wire [15:0] _078_;
wire [16:0] _079_;
wire [16:0] _080_;
wire [15:0] _081_;
wire [15:0] _082_;
wire _083_;
wire [15:0] _084_;
wire [16:0] _085_;
wire [16:0] _086_;
wire [15:0] _087_;
wire [15:0] _088_;
wire _089_;
wire [15:0] _090_;
wire [16:0] _091_;
wire [16:0] _092_;
wire [15:0] _093_;
wire [15:0] _094_;
wire _095_;
wire [15:0] _096_;
wire [16:0] _097_;
wire [16:0] _098_;
wire [15:0] _099_;
wire [15:0] _100_;
wire _101_;
wire [15:0] _102_;
wire [16:0] _103_;
wire [16:0] _104_;
wire [15:0] _105_;
wire [15:0] _106_;
wire _107_;
wire [15:0] _108_;
wire [16:0] _109_;
wire [16:0] _110_;
wire [15:0] _111_;
wire [15:0] _112_;
wire _113_;
wire [15:0] _114_;
wire [16:0] _115_;
wire [16:0] _116_;
wire [15:0] _117_;
wire [15:0] _118_;
wire _119_;
wire [15:0] _120_;
wire [16:0] _121_;
wire [16:0] _122_;
wire [15:0] _123_;
wire [15:0] _124_;
wire _125_;
wire [15:0] _126_;
wire [16:0] _127_;
wire [16:0] _128_;
wire [16:0] _129_;
wire [16:0] _130_;
wire _131_;
wire [16:0] _132_;
wire [17:0] _133_;
wire [17:0] _134_;
wire [16:0] _135_;
wire [16:0] _136_;
wire _137_;
wire [16:0] _138_;
wire [17:0] _139_;
wire [17:0] _140_;
wire [18:0] _141_;
wire [18:0] _142_;
wire _143_;
wire [18:0] _144_;
wire [19:0] _145_;
wire [19:0] _146_;
wire [19:0] _147_;
wire [19:0] _148_;
wire _149_;
wire [18:0] _150_;
wire [19:0] _151_;
wire [20:0] _152_;
wire [19:0] _153_;
wire [19:0] _154_;
wire _155_;
wire [19:0] _156_;
wire [20:0] _157_;
wire [20:0] _158_;
wire [26:0] _159_;
wire [26:0] _160_;
wire _161_;
wire [25:0] _162_;
wire [26:0] _163_;
wire [27:0] _164_;
wire _165_;
wire _166_;
wire _167_;
wire _168_;
wire _169_;
wire _170_;
wire _171_;
wire _172_;
wire _173_;
wire _174_;
wire _175_;
wire _176_;
wire _177_;
wire _178_;
wire _179_;
wire _180_;
wire _181_;
wire _182_;
wire _183_;
wire _184_;
wire _185_;
wire _186_;
wire _187_;
wire _188_;
wire _189_;
wire _190_;
wire _191_;
wire _192_;
wire _193_;
wire _194_;
wire _195_;
wire _196_;
wire _197_;
wire _198_;
wire _199_;
wire _200_;
wire _201_;
wire _202_;
wire _203_;
wire _204_;
wire _205_;
wire _206_;
wire _207_;
wire _208_;
wire _209_;
wire _210_;
wire [9:0] \add_10ns_10s_10_1_1_U5.din0 ;
wire [9:0] \add_10ns_10s_10_1_1_U5.din1 ;
wire [9:0] \add_10ns_10s_10_1_1_U5.dout ;
wire [9:0] \add_10ns_10s_10_1_1_U5.top_add_10ns_10s_10_1_1_Adder_4_U.a ;
wire [9:0] \add_10ns_10s_10_1_1_U5.top_add_10ns_10s_10_1_1_Adder_4_U.b ;
wire [9:0] \add_10ns_10s_10_1_1_U5.top_add_10ns_10s_10_1_1_Adder_4_U.s ;
wire [1:0] \add_2ns_2ns_2_1_1_U1.din0 ;
wire [1:0] \add_2ns_2ns_2_1_1_U1.din1 ;
wire [1:0] \add_2ns_2ns_2_1_1_U1.dout ;
wire [1:0] \add_2ns_2ns_2_1_1_U1.top_add_2ns_2ns_2_1_1_Adder_0_U.a ;
wire [1:0] \add_2ns_2ns_2_1_1_U1.top_add_2ns_2ns_2_1_1_Adder_0_U.b ;
wire [1:0] \add_2ns_2ns_2_1_1_U1.top_add_2ns_2ns_2_1_1_Adder_0_U.s ;
wire \add_32ns_32ns_32_2_1_U11.ce ;
wire \add_32ns_32ns_32_2_1_U11.clk ;
wire [31:0] \add_32ns_32ns_32_2_1_U11.din0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U11.din1 ;
wire [31:0] \add_32ns_32ns_32_2_1_U11.dout ;
wire \add_32ns_32ns_32_2_1_U11.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.a ;
wire [31:0] \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.b ;
wire [31:0] \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s0 ;
wire \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.ce ;
wire \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.clk ;
wire \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.facout_s1 ;
wire \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.facout_s2 ;
wire [15:0] \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s1 ;
wire [15:0] \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s2 ;
wire \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.b ;
wire \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cin ;
wire \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.b ;
wire \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cin ;
wire \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.s ;
wire \add_32ns_32ns_32_2_1_U13.ce ;
wire \add_32ns_32ns_32_2_1_U13.clk ;
wire [31:0] \add_32ns_32ns_32_2_1_U13.din0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U13.din1 ;
wire [31:0] \add_32ns_32ns_32_2_1_U13.dout ;
wire \add_32ns_32ns_32_2_1_U13.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_7_U.a ;
wire [31:0] \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_7_U.b ;
wire [31:0] \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s0 ;
wire \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_7_U.ce ;
wire \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_7_U.clk ;
wire \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_7_U.facout_s1 ;
wire \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_7_U.facout_s2 ;
wire [15:0] \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s1 ;
wire [15:0] \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s2 ;
wire \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_7_U.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_7_U.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.b ;
wire \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cin ;
wire \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.b ;
wire \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cin ;
wire \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.s ;
wire \add_32ns_32ns_32_2_1_U14.ce ;
wire \add_32ns_32ns_32_2_1_U14.clk ;
wire [31:0] \add_32ns_32ns_32_2_1_U14.din0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U14.din1 ;
wire [31:0] \add_32ns_32ns_32_2_1_U14.dout ;
wire \add_32ns_32ns_32_2_1_U14.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.a ;
wire [31:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.b ;
wire [31:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s0 ;
wire \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.ce ;
wire \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.clk ;
wire \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.facout_s1 ;
wire \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.facout_s2 ;
wire [15:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s1 ;
wire [15:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s2 ;
wire \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.b ;
wire \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cin ;
wire \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.b ;
wire \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cin ;
wire \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.s ;
wire \add_32ns_32ns_32_2_1_U16.ce ;
wire \add_32ns_32ns_32_2_1_U16.clk ;
wire [31:0] \add_32ns_32ns_32_2_1_U16.din0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U16.din1 ;
wire [31:0] \add_32ns_32ns_32_2_1_U16.dout ;
wire \add_32ns_32ns_32_2_1_U16.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.a ;
wire [31:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.b ;
wire [31:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s0 ;
wire \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.ce ;
wire \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.clk ;
wire \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.facout_s1 ;
wire \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.facout_s2 ;
wire [15:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s1 ;
wire [15:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s2 ;
wire \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.b ;
wire \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cin ;
wire \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.b ;
wire \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cin ;
wire \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.s ;
wire \add_32ns_32ns_32_2_1_U18.ce ;
wire \add_32ns_32ns_32_2_1_U18.clk ;
wire [31:0] \add_32ns_32ns_32_2_1_U18.din0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U18.din1 ;
wire [31:0] \add_32ns_32ns_32_2_1_U18.dout ;
wire \add_32ns_32ns_32_2_1_U18.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.a ;
wire [31:0] \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.b ;
wire [31:0] \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s0 ;
wire \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.ce ;
wire \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.clk ;
wire \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.facout_s1 ;
wire \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.facout_s2 ;
wire [15:0] \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s1 ;
wire [15:0] \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s2 ;
wire \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.b ;
wire \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cin ;
wire \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.b ;
wire \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cin ;
wire \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.s ;
wire \add_32ns_32ns_32_2_1_U9.ce ;
wire \add_32ns_32ns_32_2_1_U9.clk ;
wire [31:0] \add_32ns_32ns_32_2_1_U9.din0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U9.din1 ;
wire [31:0] \add_32ns_32ns_32_2_1_U9.dout ;
wire \add_32ns_32ns_32_2_1_U9.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.a ;
wire [31:0] \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.b ;
wire [31:0] \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s0 ;
wire \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.ce ;
wire \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.clk ;
wire \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.facout_s1 ;
wire \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.facout_s2 ;
wire [15:0] \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s1 ;
wire [15:0] \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s2 ;
wire \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.b ;
wire \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cin ;
wire \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.b ;
wire \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cin ;
wire \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.s ;
wire \add_32ns_32s_32_2_1_U20.ce ;
wire \add_32ns_32s_32_2_1_U20.clk ;
wire [31:0] \add_32ns_32s_32_2_1_U20.din0 ;
wire [31:0] \add_32ns_32s_32_2_1_U20.din1 ;
wire [31:0] \add_32ns_32s_32_2_1_U20.dout ;
wire \add_32ns_32s_32_2_1_U20.reset ;
wire [31:0] \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_12_U.a ;
wire [31:0] \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_12_U.ain_s0 ;
wire [31:0] \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_12_U.b ;
wire [31:0] \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_12_U.bin_s0 ;
wire \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_12_U.ce ;
wire \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_12_U.clk ;
wire \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_12_U.facout_s1 ;
wire \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_12_U.facout_s2 ;
wire [15:0] \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_12_U.fas_s1 ;
wire [15:0] \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_12_U.fas_s2 ;
wire \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_12_U.reset ;
wire [31:0] \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_12_U.s ;
wire [15:0] \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_12_U.u1.a ;
wire [15:0] \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_12_U.u1.b ;
wire \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_12_U.u1.cin ;
wire \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_12_U.u1.cout ;
wire [15:0] \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_12_U.u1.s ;
wire [15:0] \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_12_U.u2.a ;
wire [15:0] \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_12_U.u2.b ;
wire \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_12_U.u2.cin ;
wire \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_12_U.u2.cout ;
wire [15:0] \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_12_U.u2.s ;
wire \add_32ns_32s_32_2_1_U21.ce ;
wire \add_32ns_32s_32_2_1_U21.clk ;
wire [31:0] \add_32ns_32s_32_2_1_U21.din0 ;
wire [31:0] \add_32ns_32s_32_2_1_U21.din1 ;
wire [31:0] \add_32ns_32s_32_2_1_U21.dout ;
wire \add_32ns_32s_32_2_1_U21.reset ;
wire [31:0] \add_32ns_32s_32_2_1_U21.top_add_32ns_32s_32_2_1_Adder_12_U.a ;
wire [31:0] \add_32ns_32s_32_2_1_U21.top_add_32ns_32s_32_2_1_Adder_12_U.ain_s0 ;
wire [31:0] \add_32ns_32s_32_2_1_U21.top_add_32ns_32s_32_2_1_Adder_12_U.b ;
wire [31:0] \add_32ns_32s_32_2_1_U21.top_add_32ns_32s_32_2_1_Adder_12_U.bin_s0 ;
wire \add_32ns_32s_32_2_1_U21.top_add_32ns_32s_32_2_1_Adder_12_U.ce ;
wire \add_32ns_32s_32_2_1_U21.top_add_32ns_32s_32_2_1_Adder_12_U.clk ;
wire \add_32ns_32s_32_2_1_U21.top_add_32ns_32s_32_2_1_Adder_12_U.facout_s1 ;
wire \add_32ns_32s_32_2_1_U21.top_add_32ns_32s_32_2_1_Adder_12_U.facout_s2 ;
wire [15:0] \add_32ns_32s_32_2_1_U21.top_add_32ns_32s_32_2_1_Adder_12_U.fas_s1 ;
wire [15:0] \add_32ns_32s_32_2_1_U21.top_add_32ns_32s_32_2_1_Adder_12_U.fas_s2 ;
wire \add_32ns_32s_32_2_1_U21.top_add_32ns_32s_32_2_1_Adder_12_U.reset ;
wire [31:0] \add_32ns_32s_32_2_1_U21.top_add_32ns_32s_32_2_1_Adder_12_U.s ;
wire [15:0] \add_32ns_32s_32_2_1_U21.top_add_32ns_32s_32_2_1_Adder_12_U.u1.a ;
wire [15:0] \add_32ns_32s_32_2_1_U21.top_add_32ns_32s_32_2_1_Adder_12_U.u1.b ;
wire \add_32ns_32s_32_2_1_U21.top_add_32ns_32s_32_2_1_Adder_12_U.u1.cin ;
wire \add_32ns_32s_32_2_1_U21.top_add_32ns_32s_32_2_1_Adder_12_U.u1.cout ;
wire [15:0] \add_32ns_32s_32_2_1_U21.top_add_32ns_32s_32_2_1_Adder_12_U.u1.s ;
wire [15:0] \add_32ns_32s_32_2_1_U21.top_add_32ns_32s_32_2_1_Adder_12_U.u2.a ;
wire [15:0] \add_32ns_32s_32_2_1_U21.top_add_32ns_32s_32_2_1_Adder_12_U.u2.b ;
wire \add_32ns_32s_32_2_1_U21.top_add_32ns_32s_32_2_1_Adder_12_U.u2.cin ;
wire \add_32ns_32s_32_2_1_U21.top_add_32ns_32s_32_2_1_Adder_12_U.u2.cout ;
wire [15:0] \add_32ns_32s_32_2_1_U21.top_add_32ns_32s_32_2_1_Adder_12_U.u2.s ;
wire \add_32s_32ns_32_2_1_U7.ce ;
wire \add_32s_32ns_32_2_1_U7.clk ;
wire [31:0] \add_32s_32ns_32_2_1_U7.din0 ;
wire [31:0] \add_32s_32ns_32_2_1_U7.din1 ;
wire [31:0] \add_32s_32ns_32_2_1_U7.dout ;
wire \add_32s_32ns_32_2_1_U7.reset ;
wire [31:0] \add_32s_32ns_32_2_1_U7.top_add_32s_32ns_32_2_1_Adder_5_U.a ;
wire [31:0] \add_32s_32ns_32_2_1_U7.top_add_32s_32ns_32_2_1_Adder_5_U.ain_s0 ;
wire [31:0] \add_32s_32ns_32_2_1_U7.top_add_32s_32ns_32_2_1_Adder_5_U.b ;
wire [31:0] \add_32s_32ns_32_2_1_U7.top_add_32s_32ns_32_2_1_Adder_5_U.bin_s0 ;
wire \add_32s_32ns_32_2_1_U7.top_add_32s_32ns_32_2_1_Adder_5_U.ce ;
wire \add_32s_32ns_32_2_1_U7.top_add_32s_32ns_32_2_1_Adder_5_U.clk ;
wire \add_32s_32ns_32_2_1_U7.top_add_32s_32ns_32_2_1_Adder_5_U.facout_s1 ;
wire \add_32s_32ns_32_2_1_U7.top_add_32s_32ns_32_2_1_Adder_5_U.facout_s2 ;
wire [15:0] \add_32s_32ns_32_2_1_U7.top_add_32s_32ns_32_2_1_Adder_5_U.fas_s1 ;
wire [15:0] \add_32s_32ns_32_2_1_U7.top_add_32s_32ns_32_2_1_Adder_5_U.fas_s2 ;
wire \add_32s_32ns_32_2_1_U7.top_add_32s_32ns_32_2_1_Adder_5_U.reset ;
wire [31:0] \add_32s_32ns_32_2_1_U7.top_add_32s_32ns_32_2_1_Adder_5_U.s ;
wire [15:0] \add_32s_32ns_32_2_1_U7.top_add_32s_32ns_32_2_1_Adder_5_U.u1.a ;
wire [15:0] \add_32s_32ns_32_2_1_U7.top_add_32s_32ns_32_2_1_Adder_5_U.u1.b ;
wire \add_32s_32ns_32_2_1_U7.top_add_32s_32ns_32_2_1_Adder_5_U.u1.cin ;
wire \add_32s_32ns_32_2_1_U7.top_add_32s_32ns_32_2_1_Adder_5_U.u1.cout ;
wire [15:0] \add_32s_32ns_32_2_1_U7.top_add_32s_32ns_32_2_1_Adder_5_U.u1.s ;
wire [15:0] \add_32s_32ns_32_2_1_U7.top_add_32s_32ns_32_2_1_Adder_5_U.u2.a ;
wire [15:0] \add_32s_32ns_32_2_1_U7.top_add_32s_32ns_32_2_1_Adder_5_U.u2.b ;
wire \add_32s_32ns_32_2_1_U7.top_add_32s_32ns_32_2_1_Adder_5_U.u2.cin ;
wire \add_32s_32ns_32_2_1_U7.top_add_32s_32ns_32_2_1_Adder_5_U.u2.cout ;
wire [15:0] \add_32s_32ns_32_2_1_U7.top_add_32s_32ns_32_2_1_Adder_5_U.u2.s ;
wire \add_34ns_34s_34_2_1_U2.ce ;
wire \add_34ns_34s_34_2_1_U2.clk ;
wire [33:0] \add_34ns_34s_34_2_1_U2.din0 ;
wire [33:0] \add_34ns_34s_34_2_1_U2.din1 ;
wire [33:0] \add_34ns_34s_34_2_1_U2.dout ;
wire \add_34ns_34s_34_2_1_U2.reset ;
wire [33:0] \add_34ns_34s_34_2_1_U2.top_add_34ns_34s_34_2_1_Adder_1_U.a ;
wire [33:0] \add_34ns_34s_34_2_1_U2.top_add_34ns_34s_34_2_1_Adder_1_U.ain_s0 ;
wire [33:0] \add_34ns_34s_34_2_1_U2.top_add_34ns_34s_34_2_1_Adder_1_U.b ;
wire [33:0] \add_34ns_34s_34_2_1_U2.top_add_34ns_34s_34_2_1_Adder_1_U.bin_s0 ;
wire \add_34ns_34s_34_2_1_U2.top_add_34ns_34s_34_2_1_Adder_1_U.ce ;
wire \add_34ns_34s_34_2_1_U2.top_add_34ns_34s_34_2_1_Adder_1_U.clk ;
wire \add_34ns_34s_34_2_1_U2.top_add_34ns_34s_34_2_1_Adder_1_U.facout_s1 ;
wire \add_34ns_34s_34_2_1_U2.top_add_34ns_34s_34_2_1_Adder_1_U.facout_s2 ;
wire [16:0] \add_34ns_34s_34_2_1_U2.top_add_34ns_34s_34_2_1_Adder_1_U.fas_s1 ;
wire [16:0] \add_34ns_34s_34_2_1_U2.top_add_34ns_34s_34_2_1_Adder_1_U.fas_s2 ;
wire \add_34ns_34s_34_2_1_U2.top_add_34ns_34s_34_2_1_Adder_1_U.reset ;
wire [33:0] \add_34ns_34s_34_2_1_U2.top_add_34ns_34s_34_2_1_Adder_1_U.s ;
wire [16:0] \add_34ns_34s_34_2_1_U2.top_add_34ns_34s_34_2_1_Adder_1_U.u1.a ;
wire [16:0] \add_34ns_34s_34_2_1_U2.top_add_34ns_34s_34_2_1_Adder_1_U.u1.b ;
wire \add_34ns_34s_34_2_1_U2.top_add_34ns_34s_34_2_1_Adder_1_U.u1.cin ;
wire \add_34ns_34s_34_2_1_U2.top_add_34ns_34s_34_2_1_Adder_1_U.u1.cout ;
wire [16:0] \add_34ns_34s_34_2_1_U2.top_add_34ns_34s_34_2_1_Adder_1_U.u1.s ;
wire [16:0] \add_34ns_34s_34_2_1_U2.top_add_34ns_34s_34_2_1_Adder_1_U.u2.a ;
wire [16:0] \add_34ns_34s_34_2_1_U2.top_add_34ns_34s_34_2_1_Adder_1_U.u2.b ;
wire \add_34ns_34s_34_2_1_U2.top_add_34ns_34s_34_2_1_Adder_1_U.u2.cin ;
wire \add_34ns_34s_34_2_1_U2.top_add_34ns_34s_34_2_1_Adder_1_U.u2.cout ;
wire [16:0] \add_34ns_34s_34_2_1_U2.top_add_34ns_34s_34_2_1_Adder_1_U.u2.s ;
wire \add_34s_34s_34_2_1_U10.ce ;
wire \add_34s_34s_34_2_1_U10.clk ;
wire [33:0] \add_34s_34s_34_2_1_U10.din0 ;
wire [33:0] \add_34s_34s_34_2_1_U10.din1 ;
wire [33:0] \add_34s_34s_34_2_1_U10.dout ;
wire \add_34s_34s_34_2_1_U10.reset ;
wire [33:0] \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_8_U.a ;
wire [33:0] \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_8_U.ain_s0 ;
wire [33:0] \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_8_U.b ;
wire [33:0] \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_8_U.bin_s0 ;
wire \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_8_U.ce ;
wire \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_8_U.clk ;
wire \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_8_U.facout_s1 ;
wire \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_8_U.facout_s2 ;
wire [16:0] \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_8_U.fas_s1 ;
wire [16:0] \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_8_U.fas_s2 ;
wire \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_8_U.reset ;
wire [33:0] \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_8_U.s ;
wire [16:0] \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_8_U.u1.a ;
wire [16:0] \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_8_U.u1.b ;
wire \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_8_U.u1.cin ;
wire \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_8_U.u1.cout ;
wire [16:0] \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_8_U.u1.s ;
wire [16:0] \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_8_U.u2.a ;
wire [16:0] \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_8_U.u2.b ;
wire \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_8_U.u2.cin ;
wire \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_8_U.u2.cout ;
wire [16:0] \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_8_U.u2.s ;
wire \add_38s_38s_38_2_1_U15.ce ;
wire \add_38s_38s_38_2_1_U15.clk ;
wire [37:0] \add_38s_38s_38_2_1_U15.din0 ;
wire [37:0] \add_38s_38s_38_2_1_U15.din1 ;
wire [37:0] \add_38s_38s_38_2_1_U15.dout ;
wire \add_38s_38s_38_2_1_U15.reset ;
wire [37:0] \add_38s_38s_38_2_1_U15.top_add_38s_38s_38_2_1_Adder_10_U.a ;
wire [37:0] \add_38s_38s_38_2_1_U15.top_add_38s_38s_38_2_1_Adder_10_U.ain_s0 ;
wire [37:0] \add_38s_38s_38_2_1_U15.top_add_38s_38s_38_2_1_Adder_10_U.b ;
wire [37:0] \add_38s_38s_38_2_1_U15.top_add_38s_38s_38_2_1_Adder_10_U.bin_s0 ;
wire \add_38s_38s_38_2_1_U15.top_add_38s_38s_38_2_1_Adder_10_U.ce ;
wire \add_38s_38s_38_2_1_U15.top_add_38s_38s_38_2_1_Adder_10_U.clk ;
wire \add_38s_38s_38_2_1_U15.top_add_38s_38s_38_2_1_Adder_10_U.facout_s1 ;
wire \add_38s_38s_38_2_1_U15.top_add_38s_38s_38_2_1_Adder_10_U.facout_s2 ;
wire [18:0] \add_38s_38s_38_2_1_U15.top_add_38s_38s_38_2_1_Adder_10_U.fas_s1 ;
wire [18:0] \add_38s_38s_38_2_1_U15.top_add_38s_38s_38_2_1_Adder_10_U.fas_s2 ;
wire \add_38s_38s_38_2_1_U15.top_add_38s_38s_38_2_1_Adder_10_U.reset ;
wire [37:0] \add_38s_38s_38_2_1_U15.top_add_38s_38s_38_2_1_Adder_10_U.s ;
wire [18:0] \add_38s_38s_38_2_1_U15.top_add_38s_38s_38_2_1_Adder_10_U.u1.a ;
wire [18:0] \add_38s_38s_38_2_1_U15.top_add_38s_38s_38_2_1_Adder_10_U.u1.b ;
wire \add_38s_38s_38_2_1_U15.top_add_38s_38s_38_2_1_Adder_10_U.u1.cin ;
wire \add_38s_38s_38_2_1_U15.top_add_38s_38s_38_2_1_Adder_10_U.u1.cout ;
wire [18:0] \add_38s_38s_38_2_1_U15.top_add_38s_38s_38_2_1_Adder_10_U.u1.s ;
wire [18:0] \add_38s_38s_38_2_1_U15.top_add_38s_38s_38_2_1_Adder_10_U.u2.a ;
wire [18:0] \add_38s_38s_38_2_1_U15.top_add_38s_38s_38_2_1_Adder_10_U.u2.b ;
wire \add_38s_38s_38_2_1_U15.top_add_38s_38s_38_2_1_Adder_10_U.u2.cin ;
wire \add_38s_38s_38_2_1_U15.top_add_38s_38s_38_2_1_Adder_10_U.u2.cout ;
wire [18:0] \add_38s_38s_38_2_1_U15.top_add_38s_38s_38_2_1_Adder_10_U.u2.s ;
wire \add_39s_39s_39_2_1_U17.ce ;
wire \add_39s_39s_39_2_1_U17.clk ;
wire [38:0] \add_39s_39s_39_2_1_U17.din0 ;
wire [38:0] \add_39s_39s_39_2_1_U17.din1 ;
wire [38:0] \add_39s_39s_39_2_1_U17.dout ;
wire \add_39s_39s_39_2_1_U17.reset ;
wire [38:0] \add_39s_39s_39_2_1_U17.top_add_39s_39s_39_2_1_Adder_11_U.a ;
wire [38:0] \add_39s_39s_39_2_1_U17.top_add_39s_39s_39_2_1_Adder_11_U.ain_s0 ;
wire [38:0] \add_39s_39s_39_2_1_U17.top_add_39s_39s_39_2_1_Adder_11_U.b ;
wire [38:0] \add_39s_39s_39_2_1_U17.top_add_39s_39s_39_2_1_Adder_11_U.bin_s0 ;
wire \add_39s_39s_39_2_1_U17.top_add_39s_39s_39_2_1_Adder_11_U.ce ;
wire \add_39s_39s_39_2_1_U17.top_add_39s_39s_39_2_1_Adder_11_U.clk ;
wire \add_39s_39s_39_2_1_U17.top_add_39s_39s_39_2_1_Adder_11_U.facout_s1 ;
wire \add_39s_39s_39_2_1_U17.top_add_39s_39s_39_2_1_Adder_11_U.facout_s2 ;
wire [18:0] \add_39s_39s_39_2_1_U17.top_add_39s_39s_39_2_1_Adder_11_U.fas_s1 ;
wire [19:0] \add_39s_39s_39_2_1_U17.top_add_39s_39s_39_2_1_Adder_11_U.fas_s2 ;
wire \add_39s_39s_39_2_1_U17.top_add_39s_39s_39_2_1_Adder_11_U.reset ;
wire [38:0] \add_39s_39s_39_2_1_U17.top_add_39s_39s_39_2_1_Adder_11_U.s ;
wire [18:0] \add_39s_39s_39_2_1_U17.top_add_39s_39s_39_2_1_Adder_11_U.u1.a ;
wire [18:0] \add_39s_39s_39_2_1_U17.top_add_39s_39s_39_2_1_Adder_11_U.u1.b ;
wire \add_39s_39s_39_2_1_U17.top_add_39s_39s_39_2_1_Adder_11_U.u1.cin ;
wire \add_39s_39s_39_2_1_U17.top_add_39s_39s_39_2_1_Adder_11_U.u1.cout ;
wire [18:0] \add_39s_39s_39_2_1_U17.top_add_39s_39s_39_2_1_Adder_11_U.u1.s ;
wire [19:0] \add_39s_39s_39_2_1_U17.top_add_39s_39s_39_2_1_Adder_11_U.u2.a ;
wire [19:0] \add_39s_39s_39_2_1_U17.top_add_39s_39s_39_2_1_Adder_11_U.u2.b ;
wire \add_39s_39s_39_2_1_U17.top_add_39s_39s_39_2_1_Adder_11_U.u2.cin ;
wire \add_39s_39s_39_2_1_U17.top_add_39s_39s_39_2_1_Adder_11_U.u2.cout ;
wire [19:0] \add_39s_39s_39_2_1_U17.top_add_39s_39s_39_2_1_Adder_11_U.u2.s ;
wire \add_40s_40s_40_2_1_U8.ce ;
wire \add_40s_40s_40_2_1_U8.clk ;
wire [39:0] \add_40s_40s_40_2_1_U8.din0 ;
wire [39:0] \add_40s_40s_40_2_1_U8.din1 ;
wire [39:0] \add_40s_40s_40_2_1_U8.dout ;
wire \add_40s_40s_40_2_1_U8.reset ;
wire [39:0] \add_40s_40s_40_2_1_U8.top_add_40s_40s_40_2_1_Adder_6_U.a ;
wire [39:0] \add_40s_40s_40_2_1_U8.top_add_40s_40s_40_2_1_Adder_6_U.ain_s0 ;
wire [39:0] \add_40s_40s_40_2_1_U8.top_add_40s_40s_40_2_1_Adder_6_U.b ;
wire [39:0] \add_40s_40s_40_2_1_U8.top_add_40s_40s_40_2_1_Adder_6_U.bin_s0 ;
wire \add_40s_40s_40_2_1_U8.top_add_40s_40s_40_2_1_Adder_6_U.ce ;
wire \add_40s_40s_40_2_1_U8.top_add_40s_40s_40_2_1_Adder_6_U.clk ;
wire \add_40s_40s_40_2_1_U8.top_add_40s_40s_40_2_1_Adder_6_U.facout_s1 ;
wire \add_40s_40s_40_2_1_U8.top_add_40s_40s_40_2_1_Adder_6_U.facout_s2 ;
wire [19:0] \add_40s_40s_40_2_1_U8.top_add_40s_40s_40_2_1_Adder_6_U.fas_s1 ;
wire [19:0] \add_40s_40s_40_2_1_U8.top_add_40s_40s_40_2_1_Adder_6_U.fas_s2 ;
wire \add_40s_40s_40_2_1_U8.top_add_40s_40s_40_2_1_Adder_6_U.reset ;
wire [39:0] \add_40s_40s_40_2_1_U8.top_add_40s_40s_40_2_1_Adder_6_U.s ;
wire [19:0] \add_40s_40s_40_2_1_U8.top_add_40s_40s_40_2_1_Adder_6_U.u1.a ;
wire [19:0] \add_40s_40s_40_2_1_U8.top_add_40s_40s_40_2_1_Adder_6_U.u1.b ;
wire \add_40s_40s_40_2_1_U8.top_add_40s_40s_40_2_1_Adder_6_U.u1.cin ;
wire \add_40s_40s_40_2_1_U8.top_add_40s_40s_40_2_1_Adder_6_U.u1.cout ;
wire [19:0] \add_40s_40s_40_2_1_U8.top_add_40s_40s_40_2_1_Adder_6_U.u1.s ;
wire [19:0] \add_40s_40s_40_2_1_U8.top_add_40s_40s_40_2_1_Adder_6_U.u2.a ;
wire [19:0] \add_40s_40s_40_2_1_U8.top_add_40s_40s_40_2_1_Adder_6_U.u2.b ;
wire \add_40s_40s_40_2_1_U8.top_add_40s_40s_40_2_1_Adder_6_U.u2.cin ;
wire \add_40s_40s_40_2_1_U8.top_add_40s_40s_40_2_1_Adder_6_U.u2.cout ;
wire [19:0] \add_40s_40s_40_2_1_U8.top_add_40s_40s_40_2_1_Adder_6_U.u2.s ;
wire [3:0] \add_4ns_4ns_4_1_1_U19.din0 ;
wire [3:0] \add_4ns_4ns_4_1_1_U19.din1 ;
wire [3:0] \add_4ns_4ns_4_1_1_U19.dout ;
wire [3:0] \add_4ns_4ns_4_1_1_U19.top_add_4ns_4ns_4_1_1_Adder_3_U.a ;
wire [3:0] \add_4ns_4ns_4_1_1_U19.top_add_4ns_4ns_4_1_1_Adder_3_U.b ;
wire [3:0] \add_4ns_4ns_4_1_1_U19.top_add_4ns_4ns_4_1_1_Adder_3_U.s ;
wire [3:0] \add_4ns_4ns_4_1_1_U4.din0 ;
wire [3:0] \add_4ns_4ns_4_1_1_U4.din1 ;
wire [3:0] \add_4ns_4ns_4_1_1_U4.dout ;
wire [3:0] \add_4ns_4ns_4_1_1_U4.top_add_4ns_4ns_4_1_1_Adder_3_U.a ;
wire [3:0] \add_4ns_4ns_4_1_1_U4.top_add_4ns_4ns_4_1_1_Adder_3_U.b ;
wire [3:0] \add_4ns_4ns_4_1_1_U4.top_add_4ns_4ns_4_1_1_Adder_3_U.s ;
wire \add_53s_53s_53_2_1_U12.ce ;
wire \add_53s_53s_53_2_1_U12.clk ;
wire [52:0] \add_53s_53s_53_2_1_U12.din0 ;
wire [52:0] \add_53s_53s_53_2_1_U12.din1 ;
wire [52:0] \add_53s_53s_53_2_1_U12.dout ;
wire \add_53s_53s_53_2_1_U12.reset ;
wire [52:0] \add_53s_53s_53_2_1_U12.top_add_53s_53s_53_2_1_Adder_9_U.a ;
wire [52:0] \add_53s_53s_53_2_1_U12.top_add_53s_53s_53_2_1_Adder_9_U.ain_s0 ;
wire [52:0] \add_53s_53s_53_2_1_U12.top_add_53s_53s_53_2_1_Adder_9_U.b ;
wire [52:0] \add_53s_53s_53_2_1_U12.top_add_53s_53s_53_2_1_Adder_9_U.bin_s0 ;
wire \add_53s_53s_53_2_1_U12.top_add_53s_53s_53_2_1_Adder_9_U.ce ;
wire \add_53s_53s_53_2_1_U12.top_add_53s_53s_53_2_1_Adder_9_U.clk ;
wire \add_53s_53s_53_2_1_U12.top_add_53s_53s_53_2_1_Adder_9_U.facout_s1 ;
wire \add_53s_53s_53_2_1_U12.top_add_53s_53s_53_2_1_Adder_9_U.facout_s2 ;
wire [25:0] \add_53s_53s_53_2_1_U12.top_add_53s_53s_53_2_1_Adder_9_U.fas_s1 ;
wire [26:0] \add_53s_53s_53_2_1_U12.top_add_53s_53s_53_2_1_Adder_9_U.fas_s2 ;
wire \add_53s_53s_53_2_1_U12.top_add_53s_53s_53_2_1_Adder_9_U.reset ;
wire [52:0] \add_53s_53s_53_2_1_U12.top_add_53s_53s_53_2_1_Adder_9_U.s ;
wire [25:0] \add_53s_53s_53_2_1_U12.top_add_53s_53s_53_2_1_Adder_9_U.u1.a ;
wire [25:0] \add_53s_53s_53_2_1_U12.top_add_53s_53s_53_2_1_Adder_9_U.u1.b ;
wire \add_53s_53s_53_2_1_U12.top_add_53s_53s_53_2_1_Adder_9_U.u1.cin ;
wire \add_53s_53s_53_2_1_U12.top_add_53s_53s_53_2_1_Adder_9_U.u1.cout ;
wire [25:0] \add_53s_53s_53_2_1_U12.top_add_53s_53s_53_2_1_Adder_9_U.u1.s ;
wire [26:0] \add_53s_53s_53_2_1_U12.top_add_53s_53s_53_2_1_Adder_9_U.u2.a ;
wire [26:0] \add_53s_53s_53_2_1_U12.top_add_53s_53s_53_2_1_Adder_9_U.u2.b ;
wire \add_53s_53s_53_2_1_U12.top_add_53s_53s_53_2_1_Adder_9_U.u2.cin ;
wire \add_53s_53s_53_2_1_U12.top_add_53s_53s_53_2_1_Adder_9_U.u2.cout ;
wire [26:0] \add_53s_53s_53_2_1_U12.top_add_53s_53s_53_2_1_Adder_9_U.u2.s ;
wire [8:0] \add_9ns_9s_9_1_1_U3.din0 ;
wire [8:0] \add_9ns_9s_9_1_1_U3.din1 ;
wire [8:0] \add_9ns_9s_9_1_1_U3.dout ;
wire [8:0] \add_9ns_9s_9_1_1_U3.top_add_9ns_9s_9_1_1_Adder_2_U.a ;
wire [8:0] \add_9ns_9s_9_1_1_U3.top_add_9ns_9s_9_1_1_Adder_2_U.b ;
wire [8:0] \add_9ns_9s_9_1_1_U3.top_add_9ns_9s_9_1_1_Adder_2_U.s ;
wire [8:0] \add_9ns_9s_9_1_1_U6.din0 ;
wire [8:0] \add_9ns_9s_9_1_1_U6.din1 ;
wire [8:0] \add_9ns_9s_9_1_1_U6.dout ;
wire [8:0] \add_9ns_9s_9_1_1_U6.top_add_9ns_9s_9_1_1_Adder_2_U.a ;
wire [8:0] \add_9ns_9s_9_1_1_U6.top_add_9ns_9s_9_1_1_Adder_2_U.b ;
wire [8:0] \add_9ns_9s_9_1_1_U6.top_add_9ns_9s_9_1_1_Adder_2_U.s ;
wire [9:0] add_ln1346_1_fu_419_p1;
wire [9:0] add_ln1346_1_fu_419_p2;
wire [8:0] add_ln731_fu_424_p1;
wire [8:0] add_ln731_fu_424_p2;
wire and_ln340_1_fu_612_p2;
wire and_ln340_fu_576_p2;
wire and_ln785_1_fu_616_p2;
wire and_ln785_fu_599_p2;
wire and_ln786_1_fu_501_p2;
wire and_ln786_fu_396_p2;
wire ap_CS_fsm_state1;
wire ap_CS_fsm_state10;
wire ap_CS_fsm_state11;
wire ap_CS_fsm_state12;
wire ap_CS_fsm_state13;
wire ap_CS_fsm_state14;
wire ap_CS_fsm_state15;
wire ap_CS_fsm_state16;
wire ap_CS_fsm_state17;
wire ap_CS_fsm_state18;
wire ap_CS_fsm_state19;
wire ap_CS_fsm_state2;
wire ap_CS_fsm_state20;
wire ap_CS_fsm_state21;
wire ap_CS_fsm_state22;
wire ap_CS_fsm_state23;
wire ap_CS_fsm_state24;
wire ap_CS_fsm_state25;
wire ap_CS_fsm_state26;
wire ap_CS_fsm_state27;
wire ap_CS_fsm_state28;
wire ap_CS_fsm_state29;
wire ap_CS_fsm_state3;
wire ap_CS_fsm_state30;
wire ap_CS_fsm_state31;
wire ap_CS_fsm_state32;
wire ap_CS_fsm_state33;
wire ap_CS_fsm_state34;
wire ap_CS_fsm_state35;
wire ap_CS_fsm_state36;
wire ap_CS_fsm_state37;
wire ap_CS_fsm_state38;
wire ap_CS_fsm_state39;
wire ap_CS_fsm_state4;
wire ap_CS_fsm_state5;
wire ap_CS_fsm_state6;
wire ap_CS_fsm_state7;
wire ap_CS_fsm_state8;
wire ap_CS_fsm_state9;
wire [38:0] ap_NS_fsm;
wire ap_clk;
wire ap_done;
wire ap_idle;
wire ap_ready;
wire ap_rst;
wire ap_start;
wire [9:0] empty_fu_292_p1;
wire [31:0] grp_fu_1002_p1;
wire [31:0] grp_fu_1002_p2;
wire [31:0] grp_fu_1010_p1;
wire [31:0] grp_fu_1010_p2;
wire [33:0] grp_fu_316_p0;
wire [33:0] grp_fu_316_p1;
wire [33:0] grp_fu_316_p2;
wire [31:0] grp_fu_509_p0;
wire [31:0] grp_fu_509_p2;
wire [39:0] grp_fu_655_p0;
wire [39:0] grp_fu_655_p1;
wire [39:0] grp_fu_655_p2;
wire [31:0] grp_fu_676_p2;
wire [33:0] grp_fu_711_p0;
wire [33:0] grp_fu_711_p2;
wire [31:0] grp_fu_735_p2;
wire [52:0] grp_fu_760_p0;
wire [52:0] grp_fu_760_p1;
wire [52:0] grp_fu_760_p2;
wire [31:0] grp_fu_786_p2;
wire [31:0] grp_fu_822_p1;
wire [31:0] grp_fu_822_p2;
wire [37:0] grp_fu_842_p0;
wire [37:0] grp_fu_842_p1;
wire [37:0] grp_fu_842_p2;
wire [31:0] grp_fu_868_p2;
wire [38:0] grp_fu_907_p0;
wire [38:0] grp_fu_907_p1;
wire [38:0] grp_fu_907_p2;
wire [31:0] grp_fu_933_p2;
wire icmp_ln768_fu_437_p2;
wire icmp_ln786_fu_442_p2;
wire icmp_ln851_1_fu_245_p2;
wire icmp_ln851_2_fu_661_p2;
wire icmp_ln851_3_fu_770_p2;
wire icmp_ln851_4_fu_852_p2;
wire icmp_ln851_5_fu_917_p2;
wire icmp_ln851_fu_372_p2;
wire icmp_ln878_fu_299_p2;
wire [7:0] op_0;
wire op_1;
wire [2:0] op_10_V_fu_408_p3;
wire [15:0] op_11_V_fu_632_p3;
wire [31:0] op_13;
wire [4:0] op_14_V_fu_944_p3;
wire [7:0] op_16;
wire [7:0] op_17;
wire [3:0] op_18_V_fu_955_p0;
wire [3:0] op_18_V_fu_955_p2;
wire [3:0] op_2;
wire [31:0] op_29;
wire op_29_ap_vld;
wire [31:0] op_3;
wire [3:0] op_7;
wire [31:0] op_8;
wire or_ln340_fu_491_p2;
wire or_ln785_1_fu_466_p2;
wire or_ln785_2_fu_594_p2;
wire or_ln785_3_fu_620_p2;
wire or_ln785_fu_392_p2;
wire or_ln786_fu_486_p2;
wire overflow_fu_475_p2;
wire p_Result_10_fu_800_p3;
wire p_Result_11_fu_873_p3;
wire p_Result_12_fu_980_p3;
wire p_Result_16_fu_522_p3;
wire p_Result_1_fu_257_p3;
wire [15:0] p_Result_7_fu_561_p4;
wire p_Result_8_fu_681_p3;
wire p_Result_s_fu_447_p3;
wire [2:0] p_Val2_1_fu_385_p3;
wire [15:0] p_Val2_3_fu_515_p3;
wire [14:0] p_Val2_4_fu_555_p2;
wire [3:0] r_2_fu_938_p2;
wire [1:0] r_fu_794_p2;
wire [8:0] ret_V_16_fu_334_p0;
wire [8:0] ret_V_16_fu_334_p1;
wire [8:0] ret_V_16_fu_334_p2;
wire [3:0] ret_V_17_fu_459_p3;
wire [1:0] ret_V_18_fu_269_p3;
wire [31:0] ret_V_22_fu_812_p3;
wire [31:0] ret_V_25_fu_992_p3;
wire [3:0] ret_V_2_fu_377_p2;
wire [1:0] ret_V_5_fu_251_p0;
wire [1:0] ret_V_5_fu_251_p2;
wire [4:0] ret_V_7_fu_964_p2;
wire [38:0] rhs_3_fu_644_p3;
wire [32:0] rhs_4_fu_700_p3;
wire [51:0] rhs_5_fu_749_p3;
wire [36:0] rhs_7_fu_831_p3;
wire [37:0] rhs_8_fu_896_p3;
wire sel_tmp18_fu_626_p2;
wire select_ln1192_fu_326_p0;
wire [15:0] select_ln340_1_fu_581_p3;
wire [2:0] select_ln340_fu_400_p3;
wire [31:0] select_ln353_2_fu_885_p3;
wire [31:0] select_ln353_fu_693_p3;
wire [15:0] select_ln785_fu_604_p3;
wire [1:0] select_ln850_1_fu_264_p3;
wire [31:0] select_ln850_4_fu_807_p3;
wire [31:0] select_ln850_5_fu_688_p3;
wire [31:0] select_ln850_6_fu_987_p3;
wire [31:0] select_ln850_7_fu_740_p3;
wire [31:0] select_ln850_8_fu_880_p3;
wire [3:0] select_ln850_fu_454_p3;
wire [4:0] sext_ln1194_fu_961_p1;
wire [31:0] sext_ln703_2_fu_745_p0;
wire [7:0] sext_ln703_3_fu_827_p0;
wire [7:0] sext_ln703_4_fu_892_p0;
wire [31:0] sext_ln870_fu_296_p1;
wire tmp_7_fu_529_p3;
wire tmp_8_fu_536_p3;
wire [8:0] trunc_ln1346_fu_312_p1;
wire [1:0] trunc_ln851_1_fu_241_p1;
wire [6:0] trunc_ln851_2_fu_637_p1;
wire [31:0] trunc_ln851_3_fu_766_p0;
wire [19:0] trunc_ln851_3_fu_766_p1;
wire [7:0] trunc_ln851_4_fu_848_p0;
wire [4:0] trunc_ln851_4_fu_848_p1;
wire [7:0] trunc_ln851_5_fu_913_p0;
wire [5:0] trunc_ln851_5_fu_913_p1;
wire [4:0] trunc_ln851_fu_350_p1;
wire xor_ln340_fu_571_p2;
wire xor_ln365_1_fu_549_p2;
wire xor_ln365_fu_543_p2;
wire xor_ln785_1_fu_589_p2;
wire xor_ln785_fu_470_p2;
wire xor_ln786_1_fu_496_p2;
wire xor_ln786_fu_481_p2;
wire [1:0] zext_ln799_fu_791_p1;


assign _065_ = icmp_ln851_3_reg_1305 & ap_CS_fsm[21];
assign _066_ = icmp_ln851_4_reg_1357 & ap_CS_fsm[28];
assign _067_ = icmp_ln851_5_reg_1394 & ap_CS_fsm[33];
assign _068_ = ap_CS_fsm[11] & icmp_ln851_2_reg_1242;
assign _069_ = p_Result_9_reg_1274 & ap_CS_fsm[16];
assign _070_ = _072_ & ap_CS_fsm[0];
assign _071_ = ap_start & ap_CS_fsm[0];
assign and_ln340_1_fu_612_p2 = or_ln786_reg_1174 & or_ln340_reg_1180;
assign and_ln340_fu_576_p2 = xor_ln340_fu_571_p2 & or_ln786_reg_1174;
assign and_ln785_1_fu_616_p2 = xor_ln785_reg_1169 & and_ln786_1_reg_1186;
assign and_ln785_fu_599_p2 = or_ln785_2_fu_594_p2 & and_ln786_1_reg_1186;
assign and_ln786_1_fu_501_p2 = xor_ln786_1_fu_496_p2 & p_Result_15_reg_1141;
assign and_ln786_fu_396_p2 = tmp_3_reg_1052 & p_Result_13_reg_1046;
assign overflow_fu_475_p2 = xor_ln785_fu_470_p2 & or_ln785_1_fu_466_p2;
assign ret_V_7_fu_964_p2 = { op_10_V_reg_1124[2], op_10_V_reg_1124[2], op_10_V_reg_1124 } & { r_2_fu_938_p2, 1'h0 };
assign sel_tmp18_fu_626_p2 = xor_ln365_1_fu_549_p2 & or_ln785_3_fu_620_p2;
assign xor_ln340_fu_571_p2 = ~ or_ln340_reg_1180;
assign xor_ln785_1_fu_589_p2 = ~ or_ln785_1_reg_1164;
assign xor_ln786_1_fu_496_p2 = ~ icmp_ln786_reg_1153;
assign xor_ln785_fu_470_p2 = ~ p_Result_14_reg_1101;
assign xor_ln786_fu_481_p2 = ~ p_Result_15_reg_1141;
assign xor_ln365_1_fu_549_p2 = ~ xor_ln365_fu_543_p2;
assign p_Val2_4_fu_555_p2 = ~ { add_ln731_reg_1135[7:0], 7'h00 };
assign r_2_fu_938_p2 = ~ op_7;
assign _072_ = ~ ap_start;
assign _073_ = ! op_2[1:0];
assign _074_ = ! trunc_ln851_reg_1096;
assign \add_10ns_10s_10_1_1_U5.top_add_10ns_10s_10_1_1_Adder_4_U.s  = \add_10ns_10s_10_1_1_U5.top_add_10ns_10s_10_1_1_Adder_4_U.a  + \add_10ns_10s_10_1_1_U5.top_add_10ns_10s_10_1_1_Adder_4_U.b ;
assign \add_2ns_2ns_2_1_1_U1.top_add_2ns_2ns_2_1_1_Adder_0_U.s  = \add_2ns_2ns_2_1_1_U1.top_add_2ns_2ns_2_1_1_Adder_0_U.a  + \add_2ns_2ns_2_1_1_U1.top_add_2ns_2ns_2_1_1_Adder_0_U.b ;
always @(posedge \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.clk )
\add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s1  <= _076_;
always @(posedge \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.clk )
\add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s1  <= _075_;
always @(posedge \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.clk )
\add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.sum_s1  <= _078_;
always @(posedge \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.clk )
\add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.carry_s1  <= _077_;
assign _076_ = \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.ce  ? \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.b [31:16] : \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s1 ;
assign _075_ = \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.ce  ? \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.a [31:16] : \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s1 ;
assign _077_ = \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.ce  ? \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.facout_s1  : \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.carry_s1 ;
assign _078_ = \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.ce  ? \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s1  : \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.sum_s1 ;
assign _079_ = \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.a  + \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.b ;
assign { \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cout , \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.s  } = _079_ + \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cin ;
assign _080_ = \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.a  + \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.b ;
assign { \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cout , \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.s  } = _080_ + \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cin ;
always @(posedge \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_7_U.clk )
\add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s1  <= _082_;
always @(posedge \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_7_U.clk )
\add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s1  <= _081_;
always @(posedge \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_7_U.clk )
\add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_7_U.sum_s1  <= _084_;
always @(posedge \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_7_U.clk )
\add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_7_U.carry_s1  <= _083_;
assign _082_ = \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_7_U.ce  ? \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_7_U.b [31:16] : \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s1 ;
assign _081_ = \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_7_U.ce  ? \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_7_U.a [31:16] : \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s1 ;
assign _083_ = \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_7_U.ce  ? \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_7_U.facout_s1  : \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_7_U.carry_s1 ;
assign _084_ = \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_7_U.ce  ? \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s1  : \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_7_U.sum_s1 ;
assign _085_ = \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.a  + \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.b ;
assign { \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cout , \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.s  } = _085_ + \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cin ;
assign _086_ = \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.a  + \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.b ;
assign { \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cout , \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.s  } = _086_ + \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cin ;
always @(posedge \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.clk )
\add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s1  <= _088_;
always @(posedge \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.clk )
\add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s1  <= _087_;
always @(posedge \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.clk )
\add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.sum_s1  <= _090_;
always @(posedge \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.clk )
\add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.carry_s1  <= _089_;
assign _088_ = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.ce  ? \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.b [31:16] : \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s1 ;
assign _087_ = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.ce  ? \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.a [31:16] : \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s1 ;
assign _089_ = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.ce  ? \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.facout_s1  : \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.carry_s1 ;
assign _090_ = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.ce  ? \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s1  : \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.sum_s1 ;
assign _091_ = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.a  + \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.b ;
assign { \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cout , \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.s  } = _091_ + \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cin ;
assign _092_ = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.a  + \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.b ;
assign { \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cout , \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.s  } = _092_ + \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cin ;
always @(posedge \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.clk )
\add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s1  <= _094_;
always @(posedge \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.clk )
\add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s1  <= _093_;
always @(posedge \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.clk )
\add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.sum_s1  <= _096_;
always @(posedge \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.clk )
\add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.carry_s1  <= _095_;
assign _094_ = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.ce  ? \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.b [31:16] : \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s1 ;
assign _093_ = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.ce  ? \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.a [31:16] : \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s1 ;
assign _095_ = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.ce  ? \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.facout_s1  : \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.carry_s1 ;
assign _096_ = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.ce  ? \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s1  : \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.sum_s1 ;
assign _097_ = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.a  + \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.b ;
assign { \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cout , \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.s  } = _097_ + \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cin ;
assign _098_ = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.a  + \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.b ;
assign { \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cout , \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.s  } = _098_ + \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cin ;
always @(posedge \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.clk )
\add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s1  <= _100_;
always @(posedge \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.clk )
\add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s1  <= _099_;
always @(posedge \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.clk )
\add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.sum_s1  <= _102_;
always @(posedge \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.clk )
\add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.carry_s1  <= _101_;
assign _100_ = \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.ce  ? \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.b [31:16] : \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s1 ;
assign _099_ = \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.ce  ? \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.a [31:16] : \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s1 ;
assign _101_ = \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.ce  ? \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.facout_s1  : \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.carry_s1 ;
assign _102_ = \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.ce  ? \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s1  : \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.sum_s1 ;
assign _103_ = \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.a  + \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.b ;
assign { \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cout , \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.s  } = _103_ + \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cin ;
assign _104_ = \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.a  + \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.b ;
assign { \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cout , \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.s  } = _104_ + \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cin ;
always @(posedge \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.clk )
\add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s1  <= _106_;
always @(posedge \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.clk )
\add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s1  <= _105_;
always @(posedge \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.clk )
\add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.sum_s1  <= _108_;
always @(posedge \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.clk )
\add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.carry_s1  <= _107_;
assign _106_ = \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.ce  ? \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.b [31:16] : \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s1 ;
assign _105_ = \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.ce  ? \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.a [31:16] : \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s1 ;
assign _107_ = \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.ce  ? \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.facout_s1  : \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.carry_s1 ;
assign _108_ = \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.ce  ? \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s1  : \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.sum_s1 ;
assign _109_ = \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.a  + \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.b ;
assign { \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cout , \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.s  } = _109_ + \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cin ;
assign _110_ = \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.a  + \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.b ;
assign { \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cout , \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.s  } = _110_ + \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cin ;
always @(posedge \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_12_U.clk )
\add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_12_U.bin_s1  <= _112_;
always @(posedge \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_12_U.clk )
\add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_12_U.ain_s1  <= _111_;
always @(posedge \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_12_U.clk )
\add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_12_U.sum_s1  <= _114_;
always @(posedge \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_12_U.clk )
\add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_12_U.carry_s1  <= _113_;
assign _112_ = \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_12_U.ce  ? \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_12_U.b [31:16] : \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_12_U.bin_s1 ;
assign _111_ = \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_12_U.ce  ? \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_12_U.a [31:16] : \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_12_U.ain_s1 ;
assign _113_ = \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_12_U.ce  ? \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_12_U.facout_s1  : \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_12_U.carry_s1 ;
assign _114_ = \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_12_U.ce  ? \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_12_U.fas_s1  : \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_12_U.sum_s1 ;
assign _115_ = \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_12_U.u1.a  + \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_12_U.u1.b ;
assign { \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_12_U.u1.cout , \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_12_U.u1.s  } = _115_ + \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_12_U.u1.cin ;
assign _116_ = \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_12_U.u2.a  + \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_12_U.u2.b ;
assign { \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_12_U.u2.cout , \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_12_U.u2.s  } = _116_ + \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_12_U.u2.cin ;
always @(posedge \add_32ns_32s_32_2_1_U21.top_add_32ns_32s_32_2_1_Adder_12_U.clk )
\add_32ns_32s_32_2_1_U21.top_add_32ns_32s_32_2_1_Adder_12_U.bin_s1  <= _118_;
always @(posedge \add_32ns_32s_32_2_1_U21.top_add_32ns_32s_32_2_1_Adder_12_U.clk )
\add_32ns_32s_32_2_1_U21.top_add_32ns_32s_32_2_1_Adder_12_U.ain_s1  <= _117_;
always @(posedge \add_32ns_32s_32_2_1_U21.top_add_32ns_32s_32_2_1_Adder_12_U.clk )
\add_32ns_32s_32_2_1_U21.top_add_32ns_32s_32_2_1_Adder_12_U.sum_s1  <= _120_;
always @(posedge \add_32ns_32s_32_2_1_U21.top_add_32ns_32s_32_2_1_Adder_12_U.clk )
\add_32ns_32s_32_2_1_U21.top_add_32ns_32s_32_2_1_Adder_12_U.carry_s1  <= _119_;
assign _118_ = \add_32ns_32s_32_2_1_U21.top_add_32ns_32s_32_2_1_Adder_12_U.ce  ? \add_32ns_32s_32_2_1_U21.top_add_32ns_32s_32_2_1_Adder_12_U.b [31:16] : \add_32ns_32s_32_2_1_U21.top_add_32ns_32s_32_2_1_Adder_12_U.bin_s1 ;
assign _117_ = \add_32ns_32s_32_2_1_U21.top_add_32ns_32s_32_2_1_Adder_12_U.ce  ? \add_32ns_32s_32_2_1_U21.top_add_32ns_32s_32_2_1_Adder_12_U.a [31:16] : \add_32ns_32s_32_2_1_U21.top_add_32ns_32s_32_2_1_Adder_12_U.ain_s1 ;
assign _119_ = \add_32ns_32s_32_2_1_U21.top_add_32ns_32s_32_2_1_Adder_12_U.ce  ? \add_32ns_32s_32_2_1_U21.top_add_32ns_32s_32_2_1_Adder_12_U.facout_s1  : \add_32ns_32s_32_2_1_U21.top_add_32ns_32s_32_2_1_Adder_12_U.carry_s1 ;
assign _120_ = \add_32ns_32s_32_2_1_U21.top_add_32ns_32s_32_2_1_Adder_12_U.ce  ? \add_32ns_32s_32_2_1_U21.top_add_32ns_32s_32_2_1_Adder_12_U.fas_s1  : \add_32ns_32s_32_2_1_U21.top_add_32ns_32s_32_2_1_Adder_12_U.sum_s1 ;
assign _121_ = \add_32ns_32s_32_2_1_U21.top_add_32ns_32s_32_2_1_Adder_12_U.u1.a  + \add_32ns_32s_32_2_1_U21.top_add_32ns_32s_32_2_1_Adder_12_U.u1.b ;
assign { \add_32ns_32s_32_2_1_U21.top_add_32ns_32s_32_2_1_Adder_12_U.u1.cout , \add_32ns_32s_32_2_1_U21.top_add_32ns_32s_32_2_1_Adder_12_U.u1.s  } = _121_ + \add_32ns_32s_32_2_1_U21.top_add_32ns_32s_32_2_1_Adder_12_U.u1.cin ;
assign _122_ = \add_32ns_32s_32_2_1_U21.top_add_32ns_32s_32_2_1_Adder_12_U.u2.a  + \add_32ns_32s_32_2_1_U21.top_add_32ns_32s_32_2_1_Adder_12_U.u2.b ;
assign { \add_32ns_32s_32_2_1_U21.top_add_32ns_32s_32_2_1_Adder_12_U.u2.cout , \add_32ns_32s_32_2_1_U21.top_add_32ns_32s_32_2_1_Adder_12_U.u2.s  } = _122_ + \add_32ns_32s_32_2_1_U21.top_add_32ns_32s_32_2_1_Adder_12_U.u2.cin ;
always @(posedge \add_32s_32ns_32_2_1_U7.top_add_32s_32ns_32_2_1_Adder_5_U.clk )
\add_32s_32ns_32_2_1_U7.top_add_32s_32ns_32_2_1_Adder_5_U.bin_s1  <= _124_;
always @(posedge \add_32s_32ns_32_2_1_U7.top_add_32s_32ns_32_2_1_Adder_5_U.clk )
\add_32s_32ns_32_2_1_U7.top_add_32s_32ns_32_2_1_Adder_5_U.ain_s1  <= _123_;
always @(posedge \add_32s_32ns_32_2_1_U7.top_add_32s_32ns_32_2_1_Adder_5_U.clk )
\add_32s_32ns_32_2_1_U7.top_add_32s_32ns_32_2_1_Adder_5_U.sum_s1  <= _126_;
always @(posedge \add_32s_32ns_32_2_1_U7.top_add_32s_32ns_32_2_1_Adder_5_U.clk )
\add_32s_32ns_32_2_1_U7.top_add_32s_32ns_32_2_1_Adder_5_U.carry_s1  <= _125_;
assign _124_ = \add_32s_32ns_32_2_1_U7.top_add_32s_32ns_32_2_1_Adder_5_U.ce  ? \add_32s_32ns_32_2_1_U7.top_add_32s_32ns_32_2_1_Adder_5_U.b [31:16] : \add_32s_32ns_32_2_1_U7.top_add_32s_32ns_32_2_1_Adder_5_U.bin_s1 ;
assign _123_ = \add_32s_32ns_32_2_1_U7.top_add_32s_32ns_32_2_1_Adder_5_U.ce  ? \add_32s_32ns_32_2_1_U7.top_add_32s_32ns_32_2_1_Adder_5_U.a [31:16] : \add_32s_32ns_32_2_1_U7.top_add_32s_32ns_32_2_1_Adder_5_U.ain_s1 ;
assign _125_ = \add_32s_32ns_32_2_1_U7.top_add_32s_32ns_32_2_1_Adder_5_U.ce  ? \add_32s_32ns_32_2_1_U7.top_add_32s_32ns_32_2_1_Adder_5_U.facout_s1  : \add_32s_32ns_32_2_1_U7.top_add_32s_32ns_32_2_1_Adder_5_U.carry_s1 ;
assign _126_ = \add_32s_32ns_32_2_1_U7.top_add_32s_32ns_32_2_1_Adder_5_U.ce  ? \add_32s_32ns_32_2_1_U7.top_add_32s_32ns_32_2_1_Adder_5_U.fas_s1  : \add_32s_32ns_32_2_1_U7.top_add_32s_32ns_32_2_1_Adder_5_U.sum_s1 ;
assign _127_ = \add_32s_32ns_32_2_1_U7.top_add_32s_32ns_32_2_1_Adder_5_U.u1.a  + \add_32s_32ns_32_2_1_U7.top_add_32s_32ns_32_2_1_Adder_5_U.u1.b ;
assign { \add_32s_32ns_32_2_1_U7.top_add_32s_32ns_32_2_1_Adder_5_U.u1.cout , \add_32s_32ns_32_2_1_U7.top_add_32s_32ns_32_2_1_Adder_5_U.u1.s  } = _127_ + \add_32s_32ns_32_2_1_U7.top_add_32s_32ns_32_2_1_Adder_5_U.u1.cin ;
assign _128_ = \add_32s_32ns_32_2_1_U7.top_add_32s_32ns_32_2_1_Adder_5_U.u2.a  + \add_32s_32ns_32_2_1_U7.top_add_32s_32ns_32_2_1_Adder_5_U.u2.b ;
assign { \add_32s_32ns_32_2_1_U7.top_add_32s_32ns_32_2_1_Adder_5_U.u2.cout , \add_32s_32ns_32_2_1_U7.top_add_32s_32ns_32_2_1_Adder_5_U.u2.s  } = _128_ + \add_32s_32ns_32_2_1_U7.top_add_32s_32ns_32_2_1_Adder_5_U.u2.cin ;
always @(posedge \add_34ns_34s_34_2_1_U2.top_add_34ns_34s_34_2_1_Adder_1_U.clk )
\add_34ns_34s_34_2_1_U2.top_add_34ns_34s_34_2_1_Adder_1_U.bin_s1  <= _130_;
always @(posedge \add_34ns_34s_34_2_1_U2.top_add_34ns_34s_34_2_1_Adder_1_U.clk )
\add_34ns_34s_34_2_1_U2.top_add_34ns_34s_34_2_1_Adder_1_U.ain_s1  <= _129_;
always @(posedge \add_34ns_34s_34_2_1_U2.top_add_34ns_34s_34_2_1_Adder_1_U.clk )
\add_34ns_34s_34_2_1_U2.top_add_34ns_34s_34_2_1_Adder_1_U.sum_s1  <= _132_;
always @(posedge \add_34ns_34s_34_2_1_U2.top_add_34ns_34s_34_2_1_Adder_1_U.clk )
\add_34ns_34s_34_2_1_U2.top_add_34ns_34s_34_2_1_Adder_1_U.carry_s1  <= _131_;
assign _130_ = \add_34ns_34s_34_2_1_U2.top_add_34ns_34s_34_2_1_Adder_1_U.ce  ? \add_34ns_34s_34_2_1_U2.top_add_34ns_34s_34_2_1_Adder_1_U.b [33:17] : \add_34ns_34s_34_2_1_U2.top_add_34ns_34s_34_2_1_Adder_1_U.bin_s1 ;
assign _129_ = \add_34ns_34s_34_2_1_U2.top_add_34ns_34s_34_2_1_Adder_1_U.ce  ? \add_34ns_34s_34_2_1_U2.top_add_34ns_34s_34_2_1_Adder_1_U.a [33:17] : \add_34ns_34s_34_2_1_U2.top_add_34ns_34s_34_2_1_Adder_1_U.ain_s1 ;
assign _131_ = \add_34ns_34s_34_2_1_U2.top_add_34ns_34s_34_2_1_Adder_1_U.ce  ? \add_34ns_34s_34_2_1_U2.top_add_34ns_34s_34_2_1_Adder_1_U.facout_s1  : \add_34ns_34s_34_2_1_U2.top_add_34ns_34s_34_2_1_Adder_1_U.carry_s1 ;
assign _132_ = \add_34ns_34s_34_2_1_U2.top_add_34ns_34s_34_2_1_Adder_1_U.ce  ? \add_34ns_34s_34_2_1_U2.top_add_34ns_34s_34_2_1_Adder_1_U.fas_s1  : \add_34ns_34s_34_2_1_U2.top_add_34ns_34s_34_2_1_Adder_1_U.sum_s1 ;
assign _133_ = \add_34ns_34s_34_2_1_U2.top_add_34ns_34s_34_2_1_Adder_1_U.u1.a  + \add_34ns_34s_34_2_1_U2.top_add_34ns_34s_34_2_1_Adder_1_U.u1.b ;
assign { \add_34ns_34s_34_2_1_U2.top_add_34ns_34s_34_2_1_Adder_1_U.u1.cout , \add_34ns_34s_34_2_1_U2.top_add_34ns_34s_34_2_1_Adder_1_U.u1.s  } = _133_ + \add_34ns_34s_34_2_1_U2.top_add_34ns_34s_34_2_1_Adder_1_U.u1.cin ;
assign _134_ = \add_34ns_34s_34_2_1_U2.top_add_34ns_34s_34_2_1_Adder_1_U.u2.a  + \add_34ns_34s_34_2_1_U2.top_add_34ns_34s_34_2_1_Adder_1_U.u2.b ;
assign { \add_34ns_34s_34_2_1_U2.top_add_34ns_34s_34_2_1_Adder_1_U.u2.cout , \add_34ns_34s_34_2_1_U2.top_add_34ns_34s_34_2_1_Adder_1_U.u2.s  } = _134_ + \add_34ns_34s_34_2_1_U2.top_add_34ns_34s_34_2_1_Adder_1_U.u2.cin ;
always @(posedge \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_8_U.clk )
\add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_8_U.bin_s1  <= _136_;
always @(posedge \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_8_U.clk )
\add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_8_U.ain_s1  <= _135_;
always @(posedge \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_8_U.clk )
\add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_8_U.sum_s1  <= _138_;
always @(posedge \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_8_U.clk )
\add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_8_U.carry_s1  <= _137_;
assign _136_ = \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_8_U.ce  ? \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_8_U.b [33:17] : \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_8_U.bin_s1 ;
assign _135_ = \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_8_U.ce  ? \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_8_U.a [33:17] : \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_8_U.ain_s1 ;
assign _137_ = \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_8_U.ce  ? \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_8_U.facout_s1  : \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_8_U.carry_s1 ;
assign _138_ = \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_8_U.ce  ? \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_8_U.fas_s1  : \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_8_U.sum_s1 ;
assign _139_ = \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_8_U.u1.a  + \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_8_U.u1.b ;
assign { \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_8_U.u1.cout , \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_8_U.u1.s  } = _139_ + \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_8_U.u1.cin ;
assign _140_ = \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_8_U.u2.a  + \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_8_U.u2.b ;
assign { \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_8_U.u2.cout , \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_8_U.u2.s  } = _140_ + \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_8_U.u2.cin ;
always @(posedge \add_38s_38s_38_2_1_U15.top_add_38s_38s_38_2_1_Adder_10_U.clk )
\add_38s_38s_38_2_1_U15.top_add_38s_38s_38_2_1_Adder_10_U.bin_s1  <= _142_;
always @(posedge \add_38s_38s_38_2_1_U15.top_add_38s_38s_38_2_1_Adder_10_U.clk )
\add_38s_38s_38_2_1_U15.top_add_38s_38s_38_2_1_Adder_10_U.ain_s1  <= _141_;
always @(posedge \add_38s_38s_38_2_1_U15.top_add_38s_38s_38_2_1_Adder_10_U.clk )
\add_38s_38s_38_2_1_U15.top_add_38s_38s_38_2_1_Adder_10_U.sum_s1  <= _144_;
always @(posedge \add_38s_38s_38_2_1_U15.top_add_38s_38s_38_2_1_Adder_10_U.clk )
\add_38s_38s_38_2_1_U15.top_add_38s_38s_38_2_1_Adder_10_U.carry_s1  <= _143_;
assign _142_ = \add_38s_38s_38_2_1_U15.top_add_38s_38s_38_2_1_Adder_10_U.ce  ? \add_38s_38s_38_2_1_U15.top_add_38s_38s_38_2_1_Adder_10_U.b [37:19] : \add_38s_38s_38_2_1_U15.top_add_38s_38s_38_2_1_Adder_10_U.bin_s1 ;
assign _141_ = \add_38s_38s_38_2_1_U15.top_add_38s_38s_38_2_1_Adder_10_U.ce  ? \add_38s_38s_38_2_1_U15.top_add_38s_38s_38_2_1_Adder_10_U.a [37:19] : \add_38s_38s_38_2_1_U15.top_add_38s_38s_38_2_1_Adder_10_U.ain_s1 ;
assign _143_ = \add_38s_38s_38_2_1_U15.top_add_38s_38s_38_2_1_Adder_10_U.ce  ? \add_38s_38s_38_2_1_U15.top_add_38s_38s_38_2_1_Adder_10_U.facout_s1  : \add_38s_38s_38_2_1_U15.top_add_38s_38s_38_2_1_Adder_10_U.carry_s1 ;
assign _144_ = \add_38s_38s_38_2_1_U15.top_add_38s_38s_38_2_1_Adder_10_U.ce  ? \add_38s_38s_38_2_1_U15.top_add_38s_38s_38_2_1_Adder_10_U.fas_s1  : \add_38s_38s_38_2_1_U15.top_add_38s_38s_38_2_1_Adder_10_U.sum_s1 ;
assign _145_ = \add_38s_38s_38_2_1_U15.top_add_38s_38s_38_2_1_Adder_10_U.u1.a  + \add_38s_38s_38_2_1_U15.top_add_38s_38s_38_2_1_Adder_10_U.u1.b ;
assign { \add_38s_38s_38_2_1_U15.top_add_38s_38s_38_2_1_Adder_10_U.u1.cout , \add_38s_38s_38_2_1_U15.top_add_38s_38s_38_2_1_Adder_10_U.u1.s  } = _145_ + \add_38s_38s_38_2_1_U15.top_add_38s_38s_38_2_1_Adder_10_U.u1.cin ;
assign _146_ = \add_38s_38s_38_2_1_U15.top_add_38s_38s_38_2_1_Adder_10_U.u2.a  + \add_38s_38s_38_2_1_U15.top_add_38s_38s_38_2_1_Adder_10_U.u2.b ;
assign { \add_38s_38s_38_2_1_U15.top_add_38s_38s_38_2_1_Adder_10_U.u2.cout , \add_38s_38s_38_2_1_U15.top_add_38s_38s_38_2_1_Adder_10_U.u2.s  } = _146_ + \add_38s_38s_38_2_1_U15.top_add_38s_38s_38_2_1_Adder_10_U.u2.cin ;
always @(posedge \add_39s_39s_39_2_1_U17.top_add_39s_39s_39_2_1_Adder_11_U.clk )
\add_39s_39s_39_2_1_U17.top_add_39s_39s_39_2_1_Adder_11_U.bin_s1  <= _148_;
always @(posedge \add_39s_39s_39_2_1_U17.top_add_39s_39s_39_2_1_Adder_11_U.clk )
\add_39s_39s_39_2_1_U17.top_add_39s_39s_39_2_1_Adder_11_U.ain_s1  <= _147_;
always @(posedge \add_39s_39s_39_2_1_U17.top_add_39s_39s_39_2_1_Adder_11_U.clk )
\add_39s_39s_39_2_1_U17.top_add_39s_39s_39_2_1_Adder_11_U.sum_s1  <= _150_;
always @(posedge \add_39s_39s_39_2_1_U17.top_add_39s_39s_39_2_1_Adder_11_U.clk )
\add_39s_39s_39_2_1_U17.top_add_39s_39s_39_2_1_Adder_11_U.carry_s1  <= _149_;
assign _148_ = \add_39s_39s_39_2_1_U17.top_add_39s_39s_39_2_1_Adder_11_U.ce  ? \add_39s_39s_39_2_1_U17.top_add_39s_39s_39_2_1_Adder_11_U.b [38:19] : \add_39s_39s_39_2_1_U17.top_add_39s_39s_39_2_1_Adder_11_U.bin_s1 ;
assign _147_ = \add_39s_39s_39_2_1_U17.top_add_39s_39s_39_2_1_Adder_11_U.ce  ? \add_39s_39s_39_2_1_U17.top_add_39s_39s_39_2_1_Adder_11_U.a [38:19] : \add_39s_39s_39_2_1_U17.top_add_39s_39s_39_2_1_Adder_11_U.ain_s1 ;
assign _149_ = \add_39s_39s_39_2_1_U17.top_add_39s_39s_39_2_1_Adder_11_U.ce  ? \add_39s_39s_39_2_1_U17.top_add_39s_39s_39_2_1_Adder_11_U.facout_s1  : \add_39s_39s_39_2_1_U17.top_add_39s_39s_39_2_1_Adder_11_U.carry_s1 ;
assign _150_ = \add_39s_39s_39_2_1_U17.top_add_39s_39s_39_2_1_Adder_11_U.ce  ? \add_39s_39s_39_2_1_U17.top_add_39s_39s_39_2_1_Adder_11_U.fas_s1  : \add_39s_39s_39_2_1_U17.top_add_39s_39s_39_2_1_Adder_11_U.sum_s1 ;
assign _151_ = \add_39s_39s_39_2_1_U17.top_add_39s_39s_39_2_1_Adder_11_U.u1.a  + \add_39s_39s_39_2_1_U17.top_add_39s_39s_39_2_1_Adder_11_U.u1.b ;
assign { \add_39s_39s_39_2_1_U17.top_add_39s_39s_39_2_1_Adder_11_U.u1.cout , \add_39s_39s_39_2_1_U17.top_add_39s_39s_39_2_1_Adder_11_U.u1.s  } = _151_ + \add_39s_39s_39_2_1_U17.top_add_39s_39s_39_2_1_Adder_11_U.u1.cin ;
assign _152_ = \add_39s_39s_39_2_1_U17.top_add_39s_39s_39_2_1_Adder_11_U.u2.a  + \add_39s_39s_39_2_1_U17.top_add_39s_39s_39_2_1_Adder_11_U.u2.b ;
assign { \add_39s_39s_39_2_1_U17.top_add_39s_39s_39_2_1_Adder_11_U.u2.cout , \add_39s_39s_39_2_1_U17.top_add_39s_39s_39_2_1_Adder_11_U.u2.s  } = _152_ + \add_39s_39s_39_2_1_U17.top_add_39s_39s_39_2_1_Adder_11_U.u2.cin ;
always @(posedge \add_40s_40s_40_2_1_U8.top_add_40s_40s_40_2_1_Adder_6_U.clk )
\add_40s_40s_40_2_1_U8.top_add_40s_40s_40_2_1_Adder_6_U.bin_s1  <= _154_;
always @(posedge \add_40s_40s_40_2_1_U8.top_add_40s_40s_40_2_1_Adder_6_U.clk )
\add_40s_40s_40_2_1_U8.top_add_40s_40s_40_2_1_Adder_6_U.ain_s1  <= _153_;
always @(posedge \add_40s_40s_40_2_1_U8.top_add_40s_40s_40_2_1_Adder_6_U.clk )
\add_40s_40s_40_2_1_U8.top_add_40s_40s_40_2_1_Adder_6_U.sum_s1  <= _156_;
always @(posedge \add_40s_40s_40_2_1_U8.top_add_40s_40s_40_2_1_Adder_6_U.clk )
\add_40s_40s_40_2_1_U8.top_add_40s_40s_40_2_1_Adder_6_U.carry_s1  <= _155_;
assign _154_ = \add_40s_40s_40_2_1_U8.top_add_40s_40s_40_2_1_Adder_6_U.ce  ? \add_40s_40s_40_2_1_U8.top_add_40s_40s_40_2_1_Adder_6_U.b [39:20] : \add_40s_40s_40_2_1_U8.top_add_40s_40s_40_2_1_Adder_6_U.bin_s1 ;
assign _153_ = \add_40s_40s_40_2_1_U8.top_add_40s_40s_40_2_1_Adder_6_U.ce  ? \add_40s_40s_40_2_1_U8.top_add_40s_40s_40_2_1_Adder_6_U.a [39:20] : \add_40s_40s_40_2_1_U8.top_add_40s_40s_40_2_1_Adder_6_U.ain_s1 ;
assign _155_ = \add_40s_40s_40_2_1_U8.top_add_40s_40s_40_2_1_Adder_6_U.ce  ? \add_40s_40s_40_2_1_U8.top_add_40s_40s_40_2_1_Adder_6_U.facout_s1  : \add_40s_40s_40_2_1_U8.top_add_40s_40s_40_2_1_Adder_6_U.carry_s1 ;
assign _156_ = \add_40s_40s_40_2_1_U8.top_add_40s_40s_40_2_1_Adder_6_U.ce  ? \add_40s_40s_40_2_1_U8.top_add_40s_40s_40_2_1_Adder_6_U.fas_s1  : \add_40s_40s_40_2_1_U8.top_add_40s_40s_40_2_1_Adder_6_U.sum_s1 ;
assign _157_ = \add_40s_40s_40_2_1_U8.top_add_40s_40s_40_2_1_Adder_6_U.u1.a  + \add_40s_40s_40_2_1_U8.top_add_40s_40s_40_2_1_Adder_6_U.u1.b ;
assign { \add_40s_40s_40_2_1_U8.top_add_40s_40s_40_2_1_Adder_6_U.u1.cout , \add_40s_40s_40_2_1_U8.top_add_40s_40s_40_2_1_Adder_6_U.u1.s  } = _157_ + \add_40s_40s_40_2_1_U8.top_add_40s_40s_40_2_1_Adder_6_U.u1.cin ;
assign _158_ = \add_40s_40s_40_2_1_U8.top_add_40s_40s_40_2_1_Adder_6_U.u2.a  + \add_40s_40s_40_2_1_U8.top_add_40s_40s_40_2_1_Adder_6_U.u2.b ;
assign { \add_40s_40s_40_2_1_U8.top_add_40s_40s_40_2_1_Adder_6_U.u2.cout , \add_40s_40s_40_2_1_U8.top_add_40s_40s_40_2_1_Adder_6_U.u2.s  } = _158_ + \add_40s_40s_40_2_1_U8.top_add_40s_40s_40_2_1_Adder_6_U.u2.cin ;
assign \add_4ns_4ns_4_1_1_U19.top_add_4ns_4ns_4_1_1_Adder_3_U.s  = \add_4ns_4ns_4_1_1_U19.top_add_4ns_4ns_4_1_1_Adder_3_U.a  + \add_4ns_4ns_4_1_1_U19.top_add_4ns_4ns_4_1_1_Adder_3_U.b ;
assign \add_4ns_4ns_4_1_1_U4.top_add_4ns_4ns_4_1_1_Adder_3_U.s  = \add_4ns_4ns_4_1_1_U4.top_add_4ns_4ns_4_1_1_Adder_3_U.a  + \add_4ns_4ns_4_1_1_U4.top_add_4ns_4ns_4_1_1_Adder_3_U.b ;
always @(posedge \add_53s_53s_53_2_1_U12.top_add_53s_53s_53_2_1_Adder_9_U.clk )
\add_53s_53s_53_2_1_U12.top_add_53s_53s_53_2_1_Adder_9_U.bin_s1  <= _160_;
always @(posedge \add_53s_53s_53_2_1_U12.top_add_53s_53s_53_2_1_Adder_9_U.clk )
\add_53s_53s_53_2_1_U12.top_add_53s_53s_53_2_1_Adder_9_U.ain_s1  <= _159_;
always @(posedge \add_53s_53s_53_2_1_U12.top_add_53s_53s_53_2_1_Adder_9_U.clk )
\add_53s_53s_53_2_1_U12.top_add_53s_53s_53_2_1_Adder_9_U.sum_s1  <= _162_;
always @(posedge \add_53s_53s_53_2_1_U12.top_add_53s_53s_53_2_1_Adder_9_U.clk )
\add_53s_53s_53_2_1_U12.top_add_53s_53s_53_2_1_Adder_9_U.carry_s1  <= _161_;
assign _160_ = \add_53s_53s_53_2_1_U12.top_add_53s_53s_53_2_1_Adder_9_U.ce  ? \add_53s_53s_53_2_1_U12.top_add_53s_53s_53_2_1_Adder_9_U.b [52:26] : \add_53s_53s_53_2_1_U12.top_add_53s_53s_53_2_1_Adder_9_U.bin_s1 ;
assign _159_ = \add_53s_53s_53_2_1_U12.top_add_53s_53s_53_2_1_Adder_9_U.ce  ? \add_53s_53s_53_2_1_U12.top_add_53s_53s_53_2_1_Adder_9_U.a [52:26] : \add_53s_53s_53_2_1_U12.top_add_53s_53s_53_2_1_Adder_9_U.ain_s1 ;
assign _161_ = \add_53s_53s_53_2_1_U12.top_add_53s_53s_53_2_1_Adder_9_U.ce  ? \add_53s_53s_53_2_1_U12.top_add_53s_53s_53_2_1_Adder_9_U.facout_s1  : \add_53s_53s_53_2_1_U12.top_add_53s_53s_53_2_1_Adder_9_U.carry_s1 ;
assign _162_ = \add_53s_53s_53_2_1_U12.top_add_53s_53s_53_2_1_Adder_9_U.ce  ? \add_53s_53s_53_2_1_U12.top_add_53s_53s_53_2_1_Adder_9_U.fas_s1  : \add_53s_53s_53_2_1_U12.top_add_53s_53s_53_2_1_Adder_9_U.sum_s1 ;
assign _163_ = \add_53s_53s_53_2_1_U12.top_add_53s_53s_53_2_1_Adder_9_U.u1.a  + \add_53s_53s_53_2_1_U12.top_add_53s_53s_53_2_1_Adder_9_U.u1.b ;
assign { \add_53s_53s_53_2_1_U12.top_add_53s_53s_53_2_1_Adder_9_U.u1.cout , \add_53s_53s_53_2_1_U12.top_add_53s_53s_53_2_1_Adder_9_U.u1.s  } = _163_ + \add_53s_53s_53_2_1_U12.top_add_53s_53s_53_2_1_Adder_9_U.u1.cin ;
assign _164_ = \add_53s_53s_53_2_1_U12.top_add_53s_53s_53_2_1_Adder_9_U.u2.a  + \add_53s_53s_53_2_1_U12.top_add_53s_53s_53_2_1_Adder_9_U.u2.b ;
assign { \add_53s_53s_53_2_1_U12.top_add_53s_53s_53_2_1_Adder_9_U.u2.cout , \add_53s_53s_53_2_1_U12.top_add_53s_53s_53_2_1_Adder_9_U.u2.s  } = _164_ + \add_53s_53s_53_2_1_U12.top_add_53s_53s_53_2_1_Adder_9_U.u2.cin ;
assign \add_9ns_9s_9_1_1_U3.top_add_9ns_9s_9_1_1_Adder_2_U.s  = \add_9ns_9s_9_1_1_U3.top_add_9ns_9s_9_1_1_Adder_2_U.a  + \add_9ns_9s_9_1_1_U3.top_add_9ns_9s_9_1_1_Adder_2_U.b ;
assign \add_9ns_9s_9_1_1_U6.top_add_9ns_9s_9_1_1_Adder_2_U.s  = \add_9ns_9s_9_1_1_U6.top_add_9ns_9s_9_1_1_Adder_2_U.a  + \add_9ns_9s_9_1_1_U6.top_add_9ns_9s_9_1_1_Adder_2_U.b ;
assign _165_ = { ret_V_18_reg_1037[1], ret_V_18_reg_1037[1], ret_V_18_reg_1037[1], ret_V_18_reg_1037[1], ret_V_18_reg_1037[1], ret_V_18_reg_1037[1], ret_V_18_reg_1037[1], ret_V_18_reg_1037[1], ret_V_18_reg_1037[1], ret_V_18_reg_1037[1], ret_V_18_reg_1037[1], ret_V_18_reg_1037[1], ret_V_18_reg_1037[1], ret_V_18_reg_1037[1], ret_V_18_reg_1037[1], ret_V_18_reg_1037[1], ret_V_18_reg_1037[1], ret_V_18_reg_1037[1], ret_V_18_reg_1037[1], ret_V_18_reg_1037[1], ret_V_18_reg_1037[1], ret_V_18_reg_1037[1], ret_V_18_reg_1037[1], ret_V_18_reg_1037[1], ret_V_18_reg_1037[1], ret_V_18_reg_1037[1], ret_V_18_reg_1037[1], ret_V_18_reg_1037[1], ret_V_18_reg_1037[1], ret_V_18_reg_1037[1], ret_V_18_reg_1037 } > op_3;
assign _166_ = | p_Result_s_20_reg_1108;
assign _167_ = p_Result_s_20_reg_1108 != 25'h1ffffff;
assign _168_ = | trunc_ln851_2_reg_1227;
assign _169_ = | op_13[19:0];
assign _170_ = | op_16[4:0];
assign _171_ = | op_17[5:0];
assign or_ln340_fu_491_p2 = p_Result_14_reg_1101 | overflow_fu_475_p2;
assign or_ln785_1_fu_466_p2 = p_Result_15_reg_1141 | icmp_ln768_reg_1148;
assign or_ln785_2_fu_594_p2 = xor_ln785_1_fu_589_p2 | p_Result_14_reg_1101;
assign or_ln785_3_fu_620_p2 = and_ln785_1_fu_616_p2 | and_ln340_1_fu_612_p2;
assign or_ln785_fu_392_p2 = tmp_3_reg_1052 | p_Result_13_reg_1046;
assign or_ln786_fu_486_p2 = xor_ln786_fu_481_p2 | icmp_ln786_reg_1153;
always @(posedge ap_clk)
op_10_V_reg_1124[0] <= 1'h0;
always @(posedge ap_clk)
p_Val2_3_reg_1202[6:0] <= 7'h00;
always @(posedge ap_clk)
select_ln850_7_reg_1290 <= _056_;
always @(posedge ap_clk)
select_ln353_reg_1264 <= _054_;
always @(posedge ap_clk)
select_ln353_2_reg_1379 <= _053_;
always @(posedge ap_clk)
ret_V_24_reg_1399 <= _044_;
always @(posedge ap_clk)
ret_V_26_cast_reg_1404 <= _046_;
always @(posedge ap_clk)
ret_V_23_reg_1362 <= _042_;
always @(posedge ap_clk)
ret_V_24_cast_reg_1367 <= _043_;
always @(posedge ap_clk)
ret_V_21_reg_1310 <= _039_;
always @(posedge ap_clk)
ret_V_22_cast_reg_1315 <= _040_;
always @(posedge ap_clk)
ret_V_19_reg_1247 <= _038_;
always @(posedge ap_clk)
ret_V_8_cast_reg_1252 <= _050_;
always @(posedge ap_clk)
r_reg_1327 <= _034_;
always @(posedge ap_clk)
ret_V_22_reg_1332 <= _041_;
always @(posedge ap_clk)
p_Val2_3_reg_1202[15:7] <= _033_;
always @(posedge ap_clk)
select_ln785_reg_1207 <= _055_;
always @(posedge ap_clk)
sel_tmp18_reg_1212 <= _052_;
always @(posedge ap_clk)
p_Result_9_reg_1274 <= _031_;
always @(posedge ap_clk)
tmp_2_reg_1279 <= _057_;
always @(posedge ap_clk)
ret_V_16_reg_1084 <= _035_;
always @(posedge ap_clk)
ret_V_reg_1089 <= _051_;
always @(posedge ap_clk)
trunc_ln851_reg_1096 <= _062_;
always @(posedge ap_clk)
p_Result_14_reg_1101 <= _029_;
always @(posedge ap_clk)
p_Result_s_20_reg_1108 <= _032_;
always @(posedge ap_clk)
ret_V_18_reg_1037 <= _037_;
always @(posedge ap_clk)
p_Result_13_reg_1046 <= _028_;
always @(posedge ap_clk)
tmp_3_reg_1052 <= _058_;
always @(posedge ap_clk)
op_28_V_reg_1436 <= _024_;
always @(posedge ap_clk)
op_25_V_reg_1342 <= _023_;
always @(posedge ap_clk)
op_18_V_reg_1416 <= _021_;
always @(posedge ap_clk)
trunc_ln2_reg_1421 <= _060_;
always @(posedge ap_clk)
ret_V_25_reg_1426 <= _045_;
always @(posedge ap_clk)
op_21_V_reg_1217 <= _022_;
always @(posedge ap_clk)
op_11_V_reg_1222 <= _020_;
always @(posedge ap_clk)
trunc_ln851_2_reg_1227 <= _061_;
always @(posedge ap_clk)
icmp_ln851_5_reg_1394 <= _016_;
always @(posedge ap_clk)
icmp_ln851_4_reg_1357 <= _015_;
always @(posedge ap_clk)
icmp_ln851_3_reg_1305 <= _014_;
always @(posedge ap_clk)
icmp_ln851_2_reg_1242 <= _013_;
always @(posedge ap_clk)
ret_V_3_reg_1021 <= _048_;
always @(posedge ap_clk)
icmp_ln851_1_reg_1027 <= _012_;
always @(posedge ap_clk)
ret_V_5_reg_1032 <= _049_;
always @(posedge ap_clk)
empty_reg_1058 <= _009_;
always @(posedge ap_clk)
icmp_ln878_reg_1063 <= _018_;
always @(posedge ap_clk)
trunc_ln1346_reg_1079 <= _059_;
always @(posedge ap_clk)
ret_V_17_reg_1159 <= _036_;
always @(posedge ap_clk)
or_ln785_1_reg_1164 <= _026_;
always @(posedge ap_clk)
xor_ln785_reg_1169 <= _063_;
always @(posedge ap_clk)
or_ln786_reg_1174 <= _027_;
always @(posedge ap_clk)
or_ln340_reg_1180 <= _025_;
always @(posedge ap_clk)
and_ln786_1_reg_1186 <= _007_;
always @(posedge ap_clk)
add_ln850_reg_1285 <= _006_;
always @(posedge ap_clk)
add_ln691_reg_1259 <= _004_;
always @(posedge ap_clk)
add_ln691_4_reg_1411 <= _003_;
always @(posedge ap_clk)
add_ln691_3_reg_1374 <= _002_;
always @(posedge ap_clk)
add_ln691_2_reg_1322 <= _001_;
always @(posedge ap_clk)
icmp_ln851_reg_1114 <= _017_;
always @(posedge ap_clk)
ret_V_2_reg_1119 <= _047_;
always @(posedge ap_clk)
op_10_V_reg_1124[2:1] <= _019_;
always @(posedge ap_clk)
add_ln1346_1_reg_1129 <= _000_;
always @(posedge ap_clk)
add_ln731_reg_1135 <= _005_;
always @(posedge ap_clk)
p_Result_15_reg_1141 <= _030_;
always @(posedge ap_clk)
icmp_ln768_reg_1148 <= _010_;
always @(posedge ap_clk)
icmp_ln786_reg_1153 <= _011_;
always @(posedge ap_clk)
ap_CS_fsm <= _008_;
assign _064_ = _071_ ? 2'h2 : 2'h1;
assign _172_ = ap_CS_fsm == 1'h1;
function [38:0] _505_;
input [38:0] a;
input [1520:0] b;
input [38:0] s;
case (s)
39'b000000000000000000000000000000000000001:
_505_ = b[38:0];
39'b000000000000000000000000000000000000010:
_505_ = b[77:39];
39'b000000000000000000000000000000000000100:
_505_ = b[116:78];
39'b000000000000000000000000000000000001000:
_505_ = b[155:117];
39'b000000000000000000000000000000000010000:
_505_ = b[194:156];
39'b000000000000000000000000000000000100000:
_505_ = b[233:195];
39'b000000000000000000000000000000001000000:
_505_ = b[272:234];
39'b000000000000000000000000000000010000000:
_505_ = b[311:273];
39'b000000000000000000000000000000100000000:
_505_ = b[350:312];
39'b000000000000000000000000000001000000000:
_505_ = b[389:351];
39'b000000000000000000000000000010000000000:
_505_ = b[428:390];
39'b000000000000000000000000000100000000000:
_505_ = b[467:429];
39'b000000000000000000000000001000000000000:
_505_ = b[506:468];
39'b000000000000000000000000010000000000000:
_505_ = b[545:507];
39'b000000000000000000000000100000000000000:
_505_ = b[584:546];
39'b000000000000000000000001000000000000000:
_505_ = b[623:585];
39'b000000000000000000000010000000000000000:
_505_ = b[662:624];
39'b000000000000000000000100000000000000000:
_505_ = b[701:663];
39'b000000000000000000001000000000000000000:
_505_ = b[740:702];
39'b000000000000000000010000000000000000000:
_505_ = b[779:741];
39'b000000000000000000100000000000000000000:
_505_ = b[818:780];
39'b000000000000000001000000000000000000000:
_505_ = b[857:819];
39'b000000000000000010000000000000000000000:
_505_ = b[896:858];
39'b000000000000000100000000000000000000000:
_505_ = b[935:897];
39'b000000000000001000000000000000000000000:
_505_ = b[974:936];
39'b000000000000010000000000000000000000000:
_505_ = b[1013:975];
39'b000000000000100000000000000000000000000:
_505_ = b[1052:1014];
39'b000000000001000000000000000000000000000:
_505_ = b[1091:1053];
39'b000000000010000000000000000000000000000:
_505_ = b[1130:1092];
39'b000000000100000000000000000000000000000:
_505_ = b[1169:1131];
39'b000000001000000000000000000000000000000:
_505_ = b[1208:1170];
39'b000000010000000000000000000000000000000:
_505_ = b[1247:1209];
39'b000000100000000000000000000000000000000:
_505_ = b[1286:1248];
39'b000001000000000000000000000000000000000:
_505_ = b[1325:1287];
39'b000010000000000000000000000000000000000:
_505_ = b[1364:1326];
39'b000100000000000000000000000000000000000:
_505_ = b[1403:1365];
39'b001000000000000000000000000000000000000:
_505_ = b[1442:1404];
39'b010000000000000000000000000000000000000:
_505_ = b[1481:1443];
39'b100000000000000000000000000000000000000:
_505_ = b[1520:1482];
39'b000000000000000000000000000000000000000:
_505_ = a;
default:
_505_ = 39'bx;
endcase
endfunction
assign ap_NS_fsm = _505_(39'hxxxxxxxxxx, { 37'h0000000000, _064_, 1482'h00000000020000000008000000002000000000800000000200000000080000000020000000008000000002000000000800000000200000000080000000020000000008000000002000000000800000000200000000080000000020000000008000000002000000000800000000200000000080000000020000000008000000002000000000800000000200000000080000000020000000008000000002000000000800000000200000000080000000020000000000000000001 }, { _172_, _210_, _209_, _208_, _207_, _206_, _205_, _204_, _203_, _202_, _201_, _200_, _199_, _198_, _197_, _196_, _195_, _194_, _193_, _192_, _191_, _190_, _189_, _188_, _187_, _186_, _185_, _184_, _183_, _182_, _181_, _180_, _179_, _178_, _177_, _176_, _175_, _174_, _173_ });
assign _173_ = ap_CS_fsm == 39'h4000000000;
assign _174_ = ap_CS_fsm == 38'h2000000000;
assign _175_ = ap_CS_fsm == 37'h1000000000;
assign _176_ = ap_CS_fsm == 36'h800000000;
assign _177_ = ap_CS_fsm == 35'h400000000;
assign _178_ = ap_CS_fsm == 34'h200000000;
assign _179_ = ap_CS_fsm == 33'h100000000;
assign _180_ = ap_CS_fsm == 32'd2147483648;
assign _181_ = ap_CS_fsm == 31'h40000000;
assign _182_ = ap_CS_fsm == 30'h20000000;
assign _183_ = ap_CS_fsm == 29'h10000000;
assign _184_ = ap_CS_fsm == 28'h8000000;
assign _185_ = ap_CS_fsm == 27'h4000000;
assign _186_ = ap_CS_fsm == 26'h2000000;
assign _187_ = ap_CS_fsm == 25'h1000000;
assign _188_ = ap_CS_fsm == 24'h800000;
assign _189_ = ap_CS_fsm == 23'h400000;
assign _190_ = ap_CS_fsm == 22'h200000;
assign _191_ = ap_CS_fsm == 21'h100000;
assign _192_ = ap_CS_fsm == 20'h80000;
assign _193_ = ap_CS_fsm == 19'h40000;
assign _194_ = ap_CS_fsm == 18'h20000;
assign _195_ = ap_CS_fsm == 17'h10000;
assign _196_ = ap_CS_fsm == 16'h8000;
assign _197_ = ap_CS_fsm == 15'h4000;
assign _198_ = ap_CS_fsm == 14'h2000;
assign _199_ = ap_CS_fsm == 13'h1000;
assign _200_ = ap_CS_fsm == 12'h800;
assign _201_ = ap_CS_fsm == 11'h400;
assign _202_ = ap_CS_fsm == 10'h200;
assign _203_ = ap_CS_fsm == 9'h100;
assign _204_ = ap_CS_fsm == 8'h80;
assign _205_ = ap_CS_fsm == 7'h40;
assign _206_ = ap_CS_fsm == 6'h20;
assign _207_ = ap_CS_fsm == 5'h10;
assign _208_ = ap_CS_fsm == 4'h8;
assign _209_ = ap_CS_fsm == 3'h4;
assign _210_ = ap_CS_fsm == 2'h2;
assign op_29_ap_vld = ap_CS_fsm[38] ? 1'h1 : 1'h0;
assign ap_idle = _070_ ? 1'h1 : 1'h0;
assign _056_ = ap_CS_fsm[17] ? select_ln850_7_fu_740_p3 : select_ln850_7_reg_1290;
assign _054_ = ap_CS_fsm[12] ? select_ln353_fu_693_p3 : select_ln353_reg_1264;
assign _053_ = ap_CS_fsm[29] ? select_ln353_2_fu_885_p3 : select_ln353_2_reg_1379;
assign _046_ = ap_CS_fsm[31] ? grp_fu_907_p2[37:6] : ret_V_26_cast_reg_1404;
assign _044_ = ap_CS_fsm[31] ? grp_fu_907_p2 : ret_V_24_reg_1399;
assign _043_ = ap_CS_fsm[26] ? grp_fu_842_p2[36:5] : ret_V_24_cast_reg_1367;
assign _042_ = ap_CS_fsm[26] ? grp_fu_842_p2 : ret_V_23_reg_1362;
assign _040_ = ap_CS_fsm[19] ? grp_fu_760_p2[51:20] : ret_V_22_cast_reg_1315;
assign _039_ = ap_CS_fsm[19] ? grp_fu_760_p2 : ret_V_21_reg_1310;
assign _050_ = ap_CS_fsm[9] ? grp_fu_655_p2[38:7] : ret_V_8_cast_reg_1252;
assign _038_ = ap_CS_fsm[9] ? grp_fu_655_p2 : ret_V_19_reg_1247;
assign _041_ = ap_CS_fsm[22] ? ret_V_22_fu_812_p3 : ret_V_22_reg_1332;
assign _034_ = ap_CS_fsm[22] ? r_fu_794_p2 : r_reg_1327;
assign _052_ = ap_CS_fsm[6] ? sel_tmp18_fu_626_p2 : sel_tmp18_reg_1212;
assign _055_ = ap_CS_fsm[6] ? select_ln785_fu_604_p3 : select_ln785_reg_1207;
assign _033_ = ap_CS_fsm[6] ? add_ln731_reg_1135 : p_Val2_3_reg_1202[15:7];
assign _057_ = ap_CS_fsm[14] ? grp_fu_711_p2[32:1] : tmp_2_reg_1279;
assign _031_ = ap_CS_fsm[14] ? grp_fu_711_p2[33] : p_Result_9_reg_1274;
assign _032_ = ap_CS_fsm[3] ? grp_fu_316_p2[33:9] : p_Result_s_20_reg_1108;
assign _029_ = ap_CS_fsm[3] ? grp_fu_316_p2[33] : p_Result_14_reg_1101;
assign _062_ = ap_CS_fsm[3] ? ret_V_16_fu_334_p2[4:0] : trunc_ln851_reg_1096;
assign _051_ = ap_CS_fsm[3] ? ret_V_16_fu_334_p2[8:5] : ret_V_reg_1089;
assign _035_ = ap_CS_fsm[3] ? ret_V_16_fu_334_p2 : ret_V_16_reg_1084;
assign _058_ = ap_CS_fsm[1] ? ret_V_18_fu_269_p3[1] : tmp_3_reg_1052;
assign _028_ = ap_CS_fsm[1] ? ret_V_18_fu_269_p3[1] : p_Result_13_reg_1046;
assign _037_ = ap_CS_fsm[1] ? ret_V_18_fu_269_p3 : ret_V_18_reg_1037;
assign _024_ = ap_CS_fsm[36] ? grp_fu_1002_p2 : op_28_V_reg_1436;
assign _023_ = ap_CS_fsm[24] ? grp_fu_822_p2 : op_25_V_reg_1342;
assign _045_ = ap_CS_fsm[34] ? ret_V_25_fu_992_p3 : ret_V_25_reg_1426;
assign _060_ = ap_CS_fsm[34] ? ret_V_7_fu_964_p2[4:1] : trunc_ln2_reg_1421;
assign _021_ = ap_CS_fsm[34] ? op_18_V_fu_955_p2 : op_18_V_reg_1416;
assign _061_ = ap_CS_fsm[7] ? op_11_V_fu_632_p3[6:0] : trunc_ln851_2_reg_1227;
assign _020_ = ap_CS_fsm[7] ? op_11_V_fu_632_p3 : op_11_V_reg_1222;
assign _022_ = ap_CS_fsm[7] ? grp_fu_509_p2 : op_21_V_reg_1217;
assign _016_ = ap_CS_fsm[30] ? icmp_ln851_5_fu_917_p2 : icmp_ln851_5_reg_1394;
assign _015_ = ap_CS_fsm[25] ? icmp_ln851_4_fu_852_p2 : icmp_ln851_4_reg_1357;
assign _014_ = ap_CS_fsm[18] ? icmp_ln851_3_fu_770_p2 : icmp_ln851_3_reg_1305;
assign _013_ = ap_CS_fsm[8] ? icmp_ln851_2_fu_661_p2 : icmp_ln851_2_reg_1242;
assign _049_ = ap_CS_fsm[0] ? ret_V_5_fu_251_p2 : ret_V_5_reg_1032;
assign _012_ = ap_CS_fsm[0] ? icmp_ln851_1_fu_245_p2 : icmp_ln851_1_reg_1027;
assign _048_ = ap_CS_fsm[0] ? op_2[3:2] : ret_V_3_reg_1021;
assign _059_ = ap_CS_fsm[2] ? op_3[8:0] : trunc_ln1346_reg_1079;
assign _018_ = ap_CS_fsm[2] ? icmp_ln878_fu_299_p2 : icmp_ln878_reg_1063;
assign _009_ = ap_CS_fsm[2] ? op_3[9:0] : empty_reg_1058;
assign _007_ = ap_CS_fsm[5] ? and_ln786_1_fu_501_p2 : and_ln786_1_reg_1186;
assign _025_ = ap_CS_fsm[5] ? or_ln340_fu_491_p2 : or_ln340_reg_1180;
assign _027_ = ap_CS_fsm[5] ? or_ln786_fu_486_p2 : or_ln786_reg_1174;
assign _063_ = ap_CS_fsm[5] ? xor_ln785_fu_470_p2 : xor_ln785_reg_1169;
assign _026_ = ap_CS_fsm[5] ? or_ln785_1_fu_466_p2 : or_ln785_1_reg_1164;
assign _036_ = ap_CS_fsm[5] ? ret_V_17_fu_459_p3 : ret_V_17_reg_1159;
assign _006_ = _069_ ? grp_fu_735_p2 : add_ln850_reg_1285;
assign _004_ = _068_ ? grp_fu_676_p2 : add_ln691_reg_1259;
assign _003_ = _067_ ? grp_fu_933_p2 : add_ln691_4_reg_1411;
assign _002_ = _066_ ? grp_fu_868_p2 : add_ln691_3_reg_1374;
assign _001_ = _065_ ? grp_fu_786_p2 : add_ln691_2_reg_1322;
assign _011_ = ap_CS_fsm[4] ? icmp_ln786_fu_442_p2 : icmp_ln786_reg_1153;
assign _010_ = ap_CS_fsm[4] ? icmp_ln768_fu_437_p2 : icmp_ln768_reg_1148;
assign _030_ = ap_CS_fsm[4] ? add_ln731_fu_424_p2[8] : p_Result_15_reg_1141;
assign _005_ = ap_CS_fsm[4] ? add_ln731_fu_424_p2 : add_ln731_reg_1135;
assign _000_ = ap_CS_fsm[4] ? add_ln1346_1_fu_419_p2 : add_ln1346_1_reg_1129;
assign _019_ = ap_CS_fsm[4] ? op_10_V_fu_408_p3[2:1] : op_10_V_reg_1124[2:1];
assign _047_ = ap_CS_fsm[4] ? ret_V_2_fu_377_p2 : ret_V_2_reg_1119;
assign _017_ = ap_CS_fsm[4] ? icmp_ln851_fu_372_p2 : icmp_ln851_reg_1114;
assign _008_ = ap_rst ? 39'h0000000001 : ap_NS_fsm;
assign r_fu_794_p2 = icmp_ln878_reg_1063 >> icmp_ln878_reg_1063;
assign icmp_ln768_fu_437_p2 = _166_ ? 1'h1 : 1'h0;
assign icmp_ln786_fu_442_p2 = _167_ ? 1'h1 : 1'h0;
assign icmp_ln851_1_fu_245_p2 = _073_ ? 1'h1 : 1'h0;
assign icmp_ln851_2_fu_661_p2 = _168_ ? 1'h1 : 1'h0;
assign icmp_ln851_3_fu_770_p2 = _169_ ? 1'h1 : 1'h0;
assign icmp_ln851_4_fu_852_p2 = _170_ ? 1'h1 : 1'h0;
assign icmp_ln851_5_fu_917_p2 = _171_ ? 1'h1 : 1'h0;
assign icmp_ln851_fu_372_p2 = _074_ ? 1'h1 : 1'h0;
assign icmp_ln878_fu_299_p2 = _165_ ? 1'h1 : 1'h0;
assign op_10_V_fu_408_p3 = and_ln786_fu_396_p2 ? { ret_V_18_reg_1037, 1'h0 } : select_ln340_fu_400_p3;
assign op_11_V_fu_632_p3 = sel_tmp18_reg_1212 ? p_Val2_3_reg_1202 : select_ln785_reg_1207;
assign ret_V_16_fu_334_p0 = op_1 ? 9'h1e0 : 9'h000;
assign ret_V_17_fu_459_p3 = ret_V_16_reg_1084[8] ? select_ln850_fu_454_p3 : ret_V_reg_1089;
assign ret_V_18_fu_269_p3 = op_2[3] ? select_ln850_1_fu_264_p3 : ret_V_3_reg_1021;
assign ret_V_22_fu_812_p3 = ret_V_21_reg_1310[52] ? select_ln850_4_fu_807_p3 : ret_V_22_cast_reg_1315;
assign ret_V_25_fu_992_p3 = ret_V_24_reg_1399[38] ? select_ln850_6_fu_987_p3 : ret_V_26_cast_reg_1404;
assign select_ln340_1_fu_581_p3 = and_ln340_fu_576_p2 ? { add_ln731_reg_1135, 7'h00 } : { add_ln1346_1_reg_1129[9], p_Val2_4_fu_555_p2 };
assign select_ln340_fu_400_p3 = or_ln785_fu_392_p2 ? 3'h0 : { ret_V_18_reg_1037, 1'h0 };
assign select_ln353_2_fu_885_p3 = ret_V_23_reg_1362[37] ? select_ln850_8_fu_880_p3 : ret_V_24_cast_reg_1367;
assign select_ln353_fu_693_p3 = ret_V_19_reg_1247[39] ? select_ln850_5_fu_688_p3 : ret_V_8_cast_reg_1252;
assign select_ln785_fu_604_p3 = and_ln785_fu_599_p2 ? { add_ln731_reg_1135, 7'h00 } : select_ln340_1_fu_581_p3;
assign select_ln850_1_fu_264_p3 = icmp_ln851_1_reg_1027 ? ret_V_3_reg_1021 : ret_V_5_reg_1032;
assign select_ln850_4_fu_807_p3 = icmp_ln851_3_reg_1305 ? add_ln691_2_reg_1322 : ret_V_22_cast_reg_1315;
assign select_ln850_5_fu_688_p3 = icmp_ln851_2_reg_1242 ? add_ln691_reg_1259 : ret_V_8_cast_reg_1252;
assign select_ln850_6_fu_987_p3 = icmp_ln851_5_reg_1394 ? add_ln691_4_reg_1411 : ret_V_26_cast_reg_1404;
assign select_ln850_7_fu_740_p3 = p_Result_9_reg_1274 ? add_ln850_reg_1285 : tmp_2_reg_1279;
assign select_ln850_8_fu_880_p3 = icmp_ln851_4_reg_1357 ? add_ln691_3_reg_1374 : ret_V_24_cast_reg_1367;
assign select_ln850_fu_454_p3 = icmp_ln851_reg_1114 ? ret_V_reg_1089 : ret_V_2_reg_1119;
assign xor_ln365_fu_543_p2 = add_ln731_reg_1135[8] ^ add_ln1346_1_reg_1129[9];
assign add_ln1346_1_fu_419_p1 = { ret_V_18_reg_1037[1], ret_V_18_reg_1037[1], ret_V_18_reg_1037[1], ret_V_18_reg_1037[1], ret_V_18_reg_1037[1], ret_V_18_reg_1037[1], ret_V_18_reg_1037[1], ret_V_18_reg_1037[1], ret_V_18_reg_1037 };
assign add_ln731_fu_424_p1 = { ret_V_18_reg_1037[1], ret_V_18_reg_1037[1], ret_V_18_reg_1037[1], ret_V_18_reg_1037[1], ret_V_18_reg_1037[1], ret_V_18_reg_1037[1], ret_V_18_reg_1037[1], ret_V_18_reg_1037 };
assign ap_CS_fsm_state1 = ap_CS_fsm[0];
assign ap_CS_fsm_state10 = ap_CS_fsm[9];
assign ap_CS_fsm_state11 = ap_CS_fsm[10];
assign ap_CS_fsm_state12 = ap_CS_fsm[11];
assign ap_CS_fsm_state13 = ap_CS_fsm[12];
assign ap_CS_fsm_state14 = ap_CS_fsm[13];
assign ap_CS_fsm_state15 = ap_CS_fsm[14];
assign ap_CS_fsm_state16 = ap_CS_fsm[15];
assign ap_CS_fsm_state17 = ap_CS_fsm[16];
assign ap_CS_fsm_state18 = ap_CS_fsm[17];
assign ap_CS_fsm_state19 = ap_CS_fsm[18];
assign ap_CS_fsm_state2 = ap_CS_fsm[1];
assign ap_CS_fsm_state20 = ap_CS_fsm[19];
assign ap_CS_fsm_state21 = ap_CS_fsm[20];
assign ap_CS_fsm_state22 = ap_CS_fsm[21];
assign ap_CS_fsm_state23 = ap_CS_fsm[22];
assign ap_CS_fsm_state24 = ap_CS_fsm[23];
assign ap_CS_fsm_state25 = ap_CS_fsm[24];
assign ap_CS_fsm_state26 = ap_CS_fsm[25];
assign ap_CS_fsm_state27 = ap_CS_fsm[26];
assign ap_CS_fsm_state28 = ap_CS_fsm[27];
assign ap_CS_fsm_state29 = ap_CS_fsm[28];
assign ap_CS_fsm_state3 = ap_CS_fsm[2];
assign ap_CS_fsm_state30 = ap_CS_fsm[29];
assign ap_CS_fsm_state31 = ap_CS_fsm[30];
assign ap_CS_fsm_state32 = ap_CS_fsm[31];
assign ap_CS_fsm_state33 = ap_CS_fsm[32];
assign ap_CS_fsm_state34 = ap_CS_fsm[33];
assign ap_CS_fsm_state35 = ap_CS_fsm[34];
assign ap_CS_fsm_state36 = ap_CS_fsm[35];
assign ap_CS_fsm_state37 = ap_CS_fsm[36];
assign ap_CS_fsm_state38 = ap_CS_fsm[37];
assign ap_CS_fsm_state39 = ap_CS_fsm[38];
assign ap_CS_fsm_state4 = ap_CS_fsm[3];
assign ap_CS_fsm_state5 = ap_CS_fsm[4];
assign ap_CS_fsm_state6 = ap_CS_fsm[5];
assign ap_CS_fsm_state7 = ap_CS_fsm[6];
assign ap_CS_fsm_state8 = ap_CS_fsm[7];
assign ap_CS_fsm_state9 = ap_CS_fsm[8];
assign ap_done = op_29_ap_vld;
assign ap_ready = op_29_ap_vld;
assign empty_fu_292_p1 = op_3[9:0];
assign grp_fu_1002_p1 = { op_18_V_reg_1416[3], op_18_V_reg_1416[3], op_18_V_reg_1416[3], op_18_V_reg_1416[3], op_18_V_reg_1416[3], op_18_V_reg_1416[3], op_18_V_reg_1416[3], op_18_V_reg_1416[3], op_18_V_reg_1416[3], op_18_V_reg_1416[3], op_18_V_reg_1416[3], op_18_V_reg_1416[3], op_18_V_reg_1416[3], op_18_V_reg_1416[3], op_18_V_reg_1416[3], op_18_V_reg_1416[3], op_18_V_reg_1416[3], op_18_V_reg_1416[3], op_18_V_reg_1416[3], op_18_V_reg_1416[3], op_18_V_reg_1416[3], op_18_V_reg_1416[3], op_18_V_reg_1416[3], op_18_V_reg_1416[3], op_18_V_reg_1416[3], op_18_V_reg_1416[3], op_18_V_reg_1416[3], op_18_V_reg_1416[3], op_18_V_reg_1416 };
assign grp_fu_1010_p1 = { trunc_ln2_reg_1421[3], trunc_ln2_reg_1421[3], trunc_ln2_reg_1421[3], trunc_ln2_reg_1421[3], trunc_ln2_reg_1421[3], trunc_ln2_reg_1421[3], trunc_ln2_reg_1421[3], trunc_ln2_reg_1421[3], trunc_ln2_reg_1421[3], trunc_ln2_reg_1421[3], trunc_ln2_reg_1421[3], trunc_ln2_reg_1421[3], trunc_ln2_reg_1421[3], trunc_ln2_reg_1421[3], trunc_ln2_reg_1421[3], trunc_ln2_reg_1421[3], trunc_ln2_reg_1421[3], trunc_ln2_reg_1421[3], trunc_ln2_reg_1421[3], trunc_ln2_reg_1421[3], trunc_ln2_reg_1421[3], trunc_ln2_reg_1421[3], trunc_ln2_reg_1421[3], trunc_ln2_reg_1421[3], trunc_ln2_reg_1421[3], trunc_ln2_reg_1421[3], trunc_ln2_reg_1421[3], trunc_ln2_reg_1421[3], trunc_ln2_reg_1421 };
assign grp_fu_316_p0 = { 2'h0, op_3 };
assign grp_fu_316_p1 = { ret_V_18_reg_1037[1], ret_V_18_reg_1037[1], ret_V_18_reg_1037[1], ret_V_18_reg_1037[1], ret_V_18_reg_1037[1], ret_V_18_reg_1037[1], ret_V_18_reg_1037[1], ret_V_18_reg_1037[1], ret_V_18_reg_1037[1], ret_V_18_reg_1037[1], ret_V_18_reg_1037[1], ret_V_18_reg_1037[1], ret_V_18_reg_1037[1], ret_V_18_reg_1037[1], ret_V_18_reg_1037[1], ret_V_18_reg_1037[1], ret_V_18_reg_1037[1], ret_V_18_reg_1037[1], ret_V_18_reg_1037[1], ret_V_18_reg_1037[1], ret_V_18_reg_1037[1], ret_V_18_reg_1037[1], ret_V_18_reg_1037[1], ret_V_18_reg_1037[1], ret_V_18_reg_1037[1], ret_V_18_reg_1037[1], ret_V_18_reg_1037[1], ret_V_18_reg_1037[1], ret_V_18_reg_1037[1], ret_V_18_reg_1037[1], ret_V_18_reg_1037[1], ret_V_18_reg_1037[1], ret_V_18_reg_1037 };
assign grp_fu_509_p0 = { ret_V_17_reg_1159[3], ret_V_17_reg_1159[3], ret_V_17_reg_1159[3], ret_V_17_reg_1159[3], ret_V_17_reg_1159[3], ret_V_17_reg_1159[3], ret_V_17_reg_1159[3], ret_V_17_reg_1159[3], ret_V_17_reg_1159[3], ret_V_17_reg_1159[3], ret_V_17_reg_1159[3], ret_V_17_reg_1159[3], ret_V_17_reg_1159[3], ret_V_17_reg_1159[3], ret_V_17_reg_1159[3], ret_V_17_reg_1159[3], ret_V_17_reg_1159[3], ret_V_17_reg_1159[3], ret_V_17_reg_1159[3], ret_V_17_reg_1159[3], ret_V_17_reg_1159[3], ret_V_17_reg_1159[3], ret_V_17_reg_1159[3], ret_V_17_reg_1159[3], ret_V_17_reg_1159[3], ret_V_17_reg_1159[3], ret_V_17_reg_1159[3], ret_V_17_reg_1159[3], ret_V_17_reg_1159 };
assign grp_fu_655_p0 = { op_21_V_reg_1217[31], op_21_V_reg_1217, 7'h00 };
assign grp_fu_655_p1 = { op_11_V_reg_1222[15], op_11_V_reg_1222[15], op_11_V_reg_1222[15], op_11_V_reg_1222[15], op_11_V_reg_1222[15], op_11_V_reg_1222[15], op_11_V_reg_1222[15], op_11_V_reg_1222[15], op_11_V_reg_1222[15], op_11_V_reg_1222[15], op_11_V_reg_1222[15], op_11_V_reg_1222[15], op_11_V_reg_1222[15], op_11_V_reg_1222[15], op_11_V_reg_1222[15], op_11_V_reg_1222[15], op_11_V_reg_1222[15], op_11_V_reg_1222[15], op_11_V_reg_1222[15], op_11_V_reg_1222[15], op_11_V_reg_1222[15], op_11_V_reg_1222[15], op_11_V_reg_1222[15], op_11_V_reg_1222[15], op_11_V_reg_1222 };
assign grp_fu_711_p0 = { select_ln353_reg_1264[31], select_ln353_reg_1264, 1'h0 };
assign grp_fu_760_p0 = { select_ln850_7_reg_1290[31], select_ln850_7_reg_1290, 20'h00000 };
assign grp_fu_760_p1 = { op_13[31], op_13[31], op_13[31], op_13[31], op_13[31], op_13[31], op_13[31], op_13[31], op_13[31], op_13[31], op_13[31], op_13[31], op_13[31], op_13[31], op_13[31], op_13[31], op_13[31], op_13[31], op_13[31], op_13[31], op_13[31], op_13 };
assign grp_fu_822_p1 = { 30'h00000000, r_reg_1327 };
assign grp_fu_842_p0 = { op_25_V_reg_1342[31], op_25_V_reg_1342, 5'h00 };
assign grp_fu_842_p1 = { op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16 };
assign grp_fu_907_p0 = { select_ln353_2_reg_1379[31], select_ln353_2_reg_1379, 6'h00 };
assign grp_fu_907_p1 = { op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17 };
assign op_14_V_fu_944_p3 = { r_2_fu_938_p2, 1'h0 };
assign op_18_V_fu_955_p0 = { 3'h0, icmp_ln878_reg_1063 };
assign op_29 = grp_fu_1010_p2;
assign p_Result_10_fu_800_p3 = ret_V_21_reg_1310[52];
assign p_Result_11_fu_873_p3 = ret_V_23_reg_1362[37];
assign p_Result_12_fu_980_p3 = ret_V_24_reg_1399[38];
assign p_Result_16_fu_522_p3 = add_ln1346_1_reg_1129[9];
assign p_Result_1_fu_257_p3 = op_2[3];
assign p_Result_7_fu_561_p4 = { add_ln1346_1_reg_1129[9], p_Val2_4_fu_555_p2 };
assign p_Result_8_fu_681_p3 = ret_V_19_reg_1247[39];
assign p_Result_s_fu_447_p3 = ret_V_16_reg_1084[8];
assign p_Val2_1_fu_385_p3 = { ret_V_18_reg_1037, 1'h0 };
assign p_Val2_3_fu_515_p3 = { add_ln731_reg_1135, 7'h00 };
assign ret_V_16_fu_334_p1 = { op_0[7], op_0 };
assign ret_V_5_fu_251_p0 = op_2[3:2];
assign rhs_3_fu_644_p3 = { op_21_V_reg_1217, 7'h00 };
assign rhs_4_fu_700_p3 = { select_ln353_reg_1264, 1'h0 };
assign rhs_5_fu_749_p3 = { select_ln850_7_reg_1290, 20'h00000 };
assign rhs_7_fu_831_p3 = { op_25_V_reg_1342, 5'h00 };
assign rhs_8_fu_896_p3 = { select_ln353_2_reg_1379, 6'h00 };
assign select_ln1192_fu_326_p0 = op_1;
assign sext_ln1194_fu_961_p1 = { op_10_V_reg_1124[2], op_10_V_reg_1124[2], op_10_V_reg_1124 };
assign sext_ln703_2_fu_745_p0 = op_13;
assign sext_ln703_3_fu_827_p0 = op_16;
assign sext_ln703_4_fu_892_p0 = op_17;
assign sext_ln870_fu_296_p1 = { ret_V_18_reg_1037[1], ret_V_18_reg_1037[1], ret_V_18_reg_1037[1], ret_V_18_reg_1037[1], ret_V_18_reg_1037[1], ret_V_18_reg_1037[1], ret_V_18_reg_1037[1], ret_V_18_reg_1037[1], ret_V_18_reg_1037[1], ret_V_18_reg_1037[1], ret_V_18_reg_1037[1], ret_V_18_reg_1037[1], ret_V_18_reg_1037[1], ret_V_18_reg_1037[1], ret_V_18_reg_1037[1], ret_V_18_reg_1037[1], ret_V_18_reg_1037[1], ret_V_18_reg_1037[1], ret_V_18_reg_1037[1], ret_V_18_reg_1037[1], ret_V_18_reg_1037[1], ret_V_18_reg_1037[1], ret_V_18_reg_1037[1], ret_V_18_reg_1037[1], ret_V_18_reg_1037[1], ret_V_18_reg_1037[1], ret_V_18_reg_1037[1], ret_V_18_reg_1037[1], ret_V_18_reg_1037[1], ret_V_18_reg_1037[1], ret_V_18_reg_1037 };
assign tmp_7_fu_529_p3 = add_ln1346_1_reg_1129[9];
assign tmp_8_fu_536_p3 = add_ln731_reg_1135[8];
assign trunc_ln1346_fu_312_p1 = op_3[8:0];
assign trunc_ln851_1_fu_241_p1 = op_2[1:0];
assign trunc_ln851_2_fu_637_p1 = op_11_V_fu_632_p3[6:0];
assign trunc_ln851_3_fu_766_p0 = op_13;
assign trunc_ln851_3_fu_766_p1 = op_13[19:0];
assign trunc_ln851_4_fu_848_p0 = op_16;
assign trunc_ln851_4_fu_848_p1 = op_16[4:0];
assign trunc_ln851_5_fu_913_p0 = op_17;
assign trunc_ln851_5_fu_913_p1 = op_17[5:0];
assign trunc_ln851_fu_350_p1 = ret_V_16_fu_334_p2[4:0];
assign zext_ln799_fu_791_p1 = { 1'h0, icmp_ln878_reg_1063 };
assign \add_9ns_9s_9_1_1_U6.top_add_9ns_9s_9_1_1_Adder_2_U.a  = \add_9ns_9s_9_1_1_U6.din0 ;
assign \add_9ns_9s_9_1_1_U6.top_add_9ns_9s_9_1_1_Adder_2_U.b  = \add_9ns_9s_9_1_1_U6.din1 ;
assign \add_9ns_9s_9_1_1_U6.dout  = \add_9ns_9s_9_1_1_U6.top_add_9ns_9s_9_1_1_Adder_2_U.s ;
assign \add_9ns_9s_9_1_1_U6.din0  = trunc_ln1346_reg_1079;
assign \add_9ns_9s_9_1_1_U6.din1  = { ret_V_18_reg_1037[1], ret_V_18_reg_1037[1], ret_V_18_reg_1037[1], ret_V_18_reg_1037[1], ret_V_18_reg_1037[1], ret_V_18_reg_1037[1], ret_V_18_reg_1037[1], ret_V_18_reg_1037 };
assign add_ln731_fu_424_p2 = \add_9ns_9s_9_1_1_U6.dout ;
assign \add_9ns_9s_9_1_1_U3.top_add_9ns_9s_9_1_1_Adder_2_U.a  = \add_9ns_9s_9_1_1_U3.din0 ;
assign \add_9ns_9s_9_1_1_U3.top_add_9ns_9s_9_1_1_Adder_2_U.b  = \add_9ns_9s_9_1_1_U3.din1 ;
assign \add_9ns_9s_9_1_1_U3.dout  = \add_9ns_9s_9_1_1_U3.top_add_9ns_9s_9_1_1_Adder_2_U.s ;
assign \add_9ns_9s_9_1_1_U3.din0  = ret_V_16_fu_334_p0;
assign \add_9ns_9s_9_1_1_U3.din1  = { op_0[7], op_0 };
assign ret_V_16_fu_334_p2 = \add_9ns_9s_9_1_1_U3.dout ;
assign \add_53s_53s_53_2_1_U12.top_add_53s_53s_53_2_1_Adder_9_U.ain_s0  = \add_53s_53s_53_2_1_U12.top_add_53s_53s_53_2_1_Adder_9_U.a ;
assign \add_53s_53s_53_2_1_U12.top_add_53s_53s_53_2_1_Adder_9_U.bin_s0  = \add_53s_53s_53_2_1_U12.top_add_53s_53s_53_2_1_Adder_9_U.b ;
assign \add_53s_53s_53_2_1_U12.top_add_53s_53s_53_2_1_Adder_9_U.s  = { \add_53s_53s_53_2_1_U12.top_add_53s_53s_53_2_1_Adder_9_U.fas_s2 , \add_53s_53s_53_2_1_U12.top_add_53s_53s_53_2_1_Adder_9_U.sum_s1  };
assign \add_53s_53s_53_2_1_U12.top_add_53s_53s_53_2_1_Adder_9_U.u2.a  = \add_53s_53s_53_2_1_U12.top_add_53s_53s_53_2_1_Adder_9_U.ain_s1 ;
assign \add_53s_53s_53_2_1_U12.top_add_53s_53s_53_2_1_Adder_9_U.u2.b  = \add_53s_53s_53_2_1_U12.top_add_53s_53s_53_2_1_Adder_9_U.bin_s1 ;
assign \add_53s_53s_53_2_1_U12.top_add_53s_53s_53_2_1_Adder_9_U.u2.cin  = \add_53s_53s_53_2_1_U12.top_add_53s_53s_53_2_1_Adder_9_U.carry_s1 ;
assign \add_53s_53s_53_2_1_U12.top_add_53s_53s_53_2_1_Adder_9_U.facout_s2  = \add_53s_53s_53_2_1_U12.top_add_53s_53s_53_2_1_Adder_9_U.u2.cout ;
assign \add_53s_53s_53_2_1_U12.top_add_53s_53s_53_2_1_Adder_9_U.fas_s2  = \add_53s_53s_53_2_1_U12.top_add_53s_53s_53_2_1_Adder_9_U.u2.s ;
assign \add_53s_53s_53_2_1_U12.top_add_53s_53s_53_2_1_Adder_9_U.u1.a  = \add_53s_53s_53_2_1_U12.top_add_53s_53s_53_2_1_Adder_9_U.a [25:0];
assign \add_53s_53s_53_2_1_U12.top_add_53s_53s_53_2_1_Adder_9_U.u1.b  = \add_53s_53s_53_2_1_U12.top_add_53s_53s_53_2_1_Adder_9_U.b [25:0];
assign \add_53s_53s_53_2_1_U12.top_add_53s_53s_53_2_1_Adder_9_U.u1.cin  = 1'h0;
assign \add_53s_53s_53_2_1_U12.top_add_53s_53s_53_2_1_Adder_9_U.facout_s1  = \add_53s_53s_53_2_1_U12.top_add_53s_53s_53_2_1_Adder_9_U.u1.cout ;
assign \add_53s_53s_53_2_1_U12.top_add_53s_53s_53_2_1_Adder_9_U.fas_s1  = \add_53s_53s_53_2_1_U12.top_add_53s_53s_53_2_1_Adder_9_U.u1.s ;
assign \add_53s_53s_53_2_1_U12.top_add_53s_53s_53_2_1_Adder_9_U.a  = \add_53s_53s_53_2_1_U12.din0 ;
assign \add_53s_53s_53_2_1_U12.top_add_53s_53s_53_2_1_Adder_9_U.b  = \add_53s_53s_53_2_1_U12.din1 ;
assign \add_53s_53s_53_2_1_U12.top_add_53s_53s_53_2_1_Adder_9_U.ce  = \add_53s_53s_53_2_1_U12.ce ;
assign \add_53s_53s_53_2_1_U12.top_add_53s_53s_53_2_1_Adder_9_U.clk  = \add_53s_53s_53_2_1_U12.clk ;
assign \add_53s_53s_53_2_1_U12.top_add_53s_53s_53_2_1_Adder_9_U.reset  = \add_53s_53s_53_2_1_U12.reset ;
assign \add_53s_53s_53_2_1_U12.dout  = \add_53s_53s_53_2_1_U12.top_add_53s_53s_53_2_1_Adder_9_U.s ;
assign \add_53s_53s_53_2_1_U12.ce  = 1'h1;
assign \add_53s_53s_53_2_1_U12.clk  = ap_clk;
assign \add_53s_53s_53_2_1_U12.din0  = { select_ln850_7_reg_1290[31], select_ln850_7_reg_1290, 20'h00000 };
assign \add_53s_53s_53_2_1_U12.din1  = { op_13[31], op_13[31], op_13[31], op_13[31], op_13[31], op_13[31], op_13[31], op_13[31], op_13[31], op_13[31], op_13[31], op_13[31], op_13[31], op_13[31], op_13[31], op_13[31], op_13[31], op_13[31], op_13[31], op_13[31], op_13[31], op_13 };
assign grp_fu_760_p2 = \add_53s_53s_53_2_1_U12.dout ;
assign \add_53s_53s_53_2_1_U12.reset  = ap_rst;
assign \add_4ns_4ns_4_1_1_U4.top_add_4ns_4ns_4_1_1_Adder_3_U.a  = \add_4ns_4ns_4_1_1_U4.din0 ;
assign \add_4ns_4ns_4_1_1_U4.top_add_4ns_4ns_4_1_1_Adder_3_U.b  = \add_4ns_4ns_4_1_1_U4.din1 ;
assign \add_4ns_4ns_4_1_1_U4.dout  = \add_4ns_4ns_4_1_1_U4.top_add_4ns_4ns_4_1_1_Adder_3_U.s ;
assign \add_4ns_4ns_4_1_1_U4.din0  = ret_V_reg_1089;
assign \add_4ns_4ns_4_1_1_U4.din1  = 4'h1;
assign ret_V_2_fu_377_p2 = \add_4ns_4ns_4_1_1_U4.dout ;
assign \add_4ns_4ns_4_1_1_U19.top_add_4ns_4ns_4_1_1_Adder_3_U.a  = \add_4ns_4ns_4_1_1_U19.din0 ;
assign \add_4ns_4ns_4_1_1_U19.top_add_4ns_4ns_4_1_1_Adder_3_U.b  = \add_4ns_4ns_4_1_1_U19.din1 ;
assign \add_4ns_4ns_4_1_1_U19.dout  = \add_4ns_4ns_4_1_1_U19.top_add_4ns_4ns_4_1_1_Adder_3_U.s ;
assign \add_4ns_4ns_4_1_1_U19.din0  = { 3'h0, icmp_ln878_reg_1063 };
assign \add_4ns_4ns_4_1_1_U19.din1  = op_7;
assign op_18_V_fu_955_p2 = \add_4ns_4ns_4_1_1_U19.dout ;
assign \add_40s_40s_40_2_1_U8.top_add_40s_40s_40_2_1_Adder_6_U.ain_s0  = \add_40s_40s_40_2_1_U8.top_add_40s_40s_40_2_1_Adder_6_U.a ;
assign \add_40s_40s_40_2_1_U8.top_add_40s_40s_40_2_1_Adder_6_U.bin_s0  = \add_40s_40s_40_2_1_U8.top_add_40s_40s_40_2_1_Adder_6_U.b ;
assign \add_40s_40s_40_2_1_U8.top_add_40s_40s_40_2_1_Adder_6_U.s  = { \add_40s_40s_40_2_1_U8.top_add_40s_40s_40_2_1_Adder_6_U.fas_s2 , \add_40s_40s_40_2_1_U8.top_add_40s_40s_40_2_1_Adder_6_U.sum_s1  };
assign \add_40s_40s_40_2_1_U8.top_add_40s_40s_40_2_1_Adder_6_U.u2.a  = \add_40s_40s_40_2_1_U8.top_add_40s_40s_40_2_1_Adder_6_U.ain_s1 ;
assign \add_40s_40s_40_2_1_U8.top_add_40s_40s_40_2_1_Adder_6_U.u2.b  = \add_40s_40s_40_2_1_U8.top_add_40s_40s_40_2_1_Adder_6_U.bin_s1 ;
assign \add_40s_40s_40_2_1_U8.top_add_40s_40s_40_2_1_Adder_6_U.u2.cin  = \add_40s_40s_40_2_1_U8.top_add_40s_40s_40_2_1_Adder_6_U.carry_s1 ;
assign \add_40s_40s_40_2_1_U8.top_add_40s_40s_40_2_1_Adder_6_U.facout_s2  = \add_40s_40s_40_2_1_U8.top_add_40s_40s_40_2_1_Adder_6_U.u2.cout ;
assign \add_40s_40s_40_2_1_U8.top_add_40s_40s_40_2_1_Adder_6_U.fas_s2  = \add_40s_40s_40_2_1_U8.top_add_40s_40s_40_2_1_Adder_6_U.u2.s ;
assign \add_40s_40s_40_2_1_U8.top_add_40s_40s_40_2_1_Adder_6_U.u1.a  = \add_40s_40s_40_2_1_U8.top_add_40s_40s_40_2_1_Adder_6_U.a [19:0];
assign \add_40s_40s_40_2_1_U8.top_add_40s_40s_40_2_1_Adder_6_U.u1.b  = \add_40s_40s_40_2_1_U8.top_add_40s_40s_40_2_1_Adder_6_U.b [19:0];
assign \add_40s_40s_40_2_1_U8.top_add_40s_40s_40_2_1_Adder_6_U.u1.cin  = 1'h0;
assign \add_40s_40s_40_2_1_U8.top_add_40s_40s_40_2_1_Adder_6_U.facout_s1  = \add_40s_40s_40_2_1_U8.top_add_40s_40s_40_2_1_Adder_6_U.u1.cout ;
assign \add_40s_40s_40_2_1_U8.top_add_40s_40s_40_2_1_Adder_6_U.fas_s1  = \add_40s_40s_40_2_1_U8.top_add_40s_40s_40_2_1_Adder_6_U.u1.s ;
assign \add_40s_40s_40_2_1_U8.top_add_40s_40s_40_2_1_Adder_6_U.a  = \add_40s_40s_40_2_1_U8.din0 ;
assign \add_40s_40s_40_2_1_U8.top_add_40s_40s_40_2_1_Adder_6_U.b  = \add_40s_40s_40_2_1_U8.din1 ;
assign \add_40s_40s_40_2_1_U8.top_add_40s_40s_40_2_1_Adder_6_U.ce  = \add_40s_40s_40_2_1_U8.ce ;
assign \add_40s_40s_40_2_1_U8.top_add_40s_40s_40_2_1_Adder_6_U.clk  = \add_40s_40s_40_2_1_U8.clk ;
assign \add_40s_40s_40_2_1_U8.top_add_40s_40s_40_2_1_Adder_6_U.reset  = \add_40s_40s_40_2_1_U8.reset ;
assign \add_40s_40s_40_2_1_U8.dout  = \add_40s_40s_40_2_1_U8.top_add_40s_40s_40_2_1_Adder_6_U.s ;
assign \add_40s_40s_40_2_1_U8.ce  = 1'h1;
assign \add_40s_40s_40_2_1_U8.clk  = ap_clk;
assign \add_40s_40s_40_2_1_U8.din0  = { op_21_V_reg_1217[31], op_21_V_reg_1217, 7'h00 };
assign \add_40s_40s_40_2_1_U8.din1  = { op_11_V_reg_1222[15], op_11_V_reg_1222[15], op_11_V_reg_1222[15], op_11_V_reg_1222[15], op_11_V_reg_1222[15], op_11_V_reg_1222[15], op_11_V_reg_1222[15], op_11_V_reg_1222[15], op_11_V_reg_1222[15], op_11_V_reg_1222[15], op_11_V_reg_1222[15], op_11_V_reg_1222[15], op_11_V_reg_1222[15], op_11_V_reg_1222[15], op_11_V_reg_1222[15], op_11_V_reg_1222[15], op_11_V_reg_1222[15], op_11_V_reg_1222[15], op_11_V_reg_1222[15], op_11_V_reg_1222[15], op_11_V_reg_1222[15], op_11_V_reg_1222[15], op_11_V_reg_1222[15], op_11_V_reg_1222[15], op_11_V_reg_1222 };
assign grp_fu_655_p2 = \add_40s_40s_40_2_1_U8.dout ;
assign \add_40s_40s_40_2_1_U8.reset  = ap_rst;
assign \add_39s_39s_39_2_1_U17.top_add_39s_39s_39_2_1_Adder_11_U.ain_s0  = \add_39s_39s_39_2_1_U17.top_add_39s_39s_39_2_1_Adder_11_U.a ;
assign \add_39s_39s_39_2_1_U17.top_add_39s_39s_39_2_1_Adder_11_U.bin_s0  = \add_39s_39s_39_2_1_U17.top_add_39s_39s_39_2_1_Adder_11_U.b ;
assign \add_39s_39s_39_2_1_U17.top_add_39s_39s_39_2_1_Adder_11_U.s  = { \add_39s_39s_39_2_1_U17.top_add_39s_39s_39_2_1_Adder_11_U.fas_s2 , \add_39s_39s_39_2_1_U17.top_add_39s_39s_39_2_1_Adder_11_U.sum_s1  };
assign \add_39s_39s_39_2_1_U17.top_add_39s_39s_39_2_1_Adder_11_U.u2.a  = \add_39s_39s_39_2_1_U17.top_add_39s_39s_39_2_1_Adder_11_U.ain_s1 ;
assign \add_39s_39s_39_2_1_U17.top_add_39s_39s_39_2_1_Adder_11_U.u2.b  = \add_39s_39s_39_2_1_U17.top_add_39s_39s_39_2_1_Adder_11_U.bin_s1 ;
assign \add_39s_39s_39_2_1_U17.top_add_39s_39s_39_2_1_Adder_11_U.u2.cin  = \add_39s_39s_39_2_1_U17.top_add_39s_39s_39_2_1_Adder_11_U.carry_s1 ;
assign \add_39s_39s_39_2_1_U17.top_add_39s_39s_39_2_1_Adder_11_U.facout_s2  = \add_39s_39s_39_2_1_U17.top_add_39s_39s_39_2_1_Adder_11_U.u2.cout ;
assign \add_39s_39s_39_2_1_U17.top_add_39s_39s_39_2_1_Adder_11_U.fas_s2  = \add_39s_39s_39_2_1_U17.top_add_39s_39s_39_2_1_Adder_11_U.u2.s ;
assign \add_39s_39s_39_2_1_U17.top_add_39s_39s_39_2_1_Adder_11_U.u1.a  = \add_39s_39s_39_2_1_U17.top_add_39s_39s_39_2_1_Adder_11_U.a [18:0];
assign \add_39s_39s_39_2_1_U17.top_add_39s_39s_39_2_1_Adder_11_U.u1.b  = \add_39s_39s_39_2_1_U17.top_add_39s_39s_39_2_1_Adder_11_U.b [18:0];
assign \add_39s_39s_39_2_1_U17.top_add_39s_39s_39_2_1_Adder_11_U.u1.cin  = 1'h0;
assign \add_39s_39s_39_2_1_U17.top_add_39s_39s_39_2_1_Adder_11_U.facout_s1  = \add_39s_39s_39_2_1_U17.top_add_39s_39s_39_2_1_Adder_11_U.u1.cout ;
assign \add_39s_39s_39_2_1_U17.top_add_39s_39s_39_2_1_Adder_11_U.fas_s1  = \add_39s_39s_39_2_1_U17.top_add_39s_39s_39_2_1_Adder_11_U.u1.s ;
assign \add_39s_39s_39_2_1_U17.top_add_39s_39s_39_2_1_Adder_11_U.a  = \add_39s_39s_39_2_1_U17.din0 ;
assign \add_39s_39s_39_2_1_U17.top_add_39s_39s_39_2_1_Adder_11_U.b  = \add_39s_39s_39_2_1_U17.din1 ;
assign \add_39s_39s_39_2_1_U17.top_add_39s_39s_39_2_1_Adder_11_U.ce  = \add_39s_39s_39_2_1_U17.ce ;
assign \add_39s_39s_39_2_1_U17.top_add_39s_39s_39_2_1_Adder_11_U.clk  = \add_39s_39s_39_2_1_U17.clk ;
assign \add_39s_39s_39_2_1_U17.top_add_39s_39s_39_2_1_Adder_11_U.reset  = \add_39s_39s_39_2_1_U17.reset ;
assign \add_39s_39s_39_2_1_U17.dout  = \add_39s_39s_39_2_1_U17.top_add_39s_39s_39_2_1_Adder_11_U.s ;
assign \add_39s_39s_39_2_1_U17.ce  = 1'h1;
assign \add_39s_39s_39_2_1_U17.clk  = ap_clk;
assign \add_39s_39s_39_2_1_U17.din0  = { select_ln353_2_reg_1379[31], select_ln353_2_reg_1379, 6'h00 };
assign \add_39s_39s_39_2_1_U17.din1  = { op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17[7], op_17 };
assign grp_fu_907_p2 = \add_39s_39s_39_2_1_U17.dout ;
assign \add_39s_39s_39_2_1_U17.reset  = ap_rst;
assign \add_38s_38s_38_2_1_U15.top_add_38s_38s_38_2_1_Adder_10_U.ain_s0  = \add_38s_38s_38_2_1_U15.top_add_38s_38s_38_2_1_Adder_10_U.a ;
assign \add_38s_38s_38_2_1_U15.top_add_38s_38s_38_2_1_Adder_10_U.bin_s0  = \add_38s_38s_38_2_1_U15.top_add_38s_38s_38_2_1_Adder_10_U.b ;
assign \add_38s_38s_38_2_1_U15.top_add_38s_38s_38_2_1_Adder_10_U.s  = { \add_38s_38s_38_2_1_U15.top_add_38s_38s_38_2_1_Adder_10_U.fas_s2 , \add_38s_38s_38_2_1_U15.top_add_38s_38s_38_2_1_Adder_10_U.sum_s1  };
assign \add_38s_38s_38_2_1_U15.top_add_38s_38s_38_2_1_Adder_10_U.u2.a  = \add_38s_38s_38_2_1_U15.top_add_38s_38s_38_2_1_Adder_10_U.ain_s1 ;
assign \add_38s_38s_38_2_1_U15.top_add_38s_38s_38_2_1_Adder_10_U.u2.b  = \add_38s_38s_38_2_1_U15.top_add_38s_38s_38_2_1_Adder_10_U.bin_s1 ;
assign \add_38s_38s_38_2_1_U15.top_add_38s_38s_38_2_1_Adder_10_U.u2.cin  = \add_38s_38s_38_2_1_U15.top_add_38s_38s_38_2_1_Adder_10_U.carry_s1 ;
assign \add_38s_38s_38_2_1_U15.top_add_38s_38s_38_2_1_Adder_10_U.facout_s2  = \add_38s_38s_38_2_1_U15.top_add_38s_38s_38_2_1_Adder_10_U.u2.cout ;
assign \add_38s_38s_38_2_1_U15.top_add_38s_38s_38_2_1_Adder_10_U.fas_s2  = \add_38s_38s_38_2_1_U15.top_add_38s_38s_38_2_1_Adder_10_U.u2.s ;
assign \add_38s_38s_38_2_1_U15.top_add_38s_38s_38_2_1_Adder_10_U.u1.a  = \add_38s_38s_38_2_1_U15.top_add_38s_38s_38_2_1_Adder_10_U.a [18:0];
assign \add_38s_38s_38_2_1_U15.top_add_38s_38s_38_2_1_Adder_10_U.u1.b  = \add_38s_38s_38_2_1_U15.top_add_38s_38s_38_2_1_Adder_10_U.b [18:0];
assign \add_38s_38s_38_2_1_U15.top_add_38s_38s_38_2_1_Adder_10_U.u1.cin  = 1'h0;
assign \add_38s_38s_38_2_1_U15.top_add_38s_38s_38_2_1_Adder_10_U.facout_s1  = \add_38s_38s_38_2_1_U15.top_add_38s_38s_38_2_1_Adder_10_U.u1.cout ;
assign \add_38s_38s_38_2_1_U15.top_add_38s_38s_38_2_1_Adder_10_U.fas_s1  = \add_38s_38s_38_2_1_U15.top_add_38s_38s_38_2_1_Adder_10_U.u1.s ;
assign \add_38s_38s_38_2_1_U15.top_add_38s_38s_38_2_1_Adder_10_U.a  = \add_38s_38s_38_2_1_U15.din0 ;
assign \add_38s_38s_38_2_1_U15.top_add_38s_38s_38_2_1_Adder_10_U.b  = \add_38s_38s_38_2_1_U15.din1 ;
assign \add_38s_38s_38_2_1_U15.top_add_38s_38s_38_2_1_Adder_10_U.ce  = \add_38s_38s_38_2_1_U15.ce ;
assign \add_38s_38s_38_2_1_U15.top_add_38s_38s_38_2_1_Adder_10_U.clk  = \add_38s_38s_38_2_1_U15.clk ;
assign \add_38s_38s_38_2_1_U15.top_add_38s_38s_38_2_1_Adder_10_U.reset  = \add_38s_38s_38_2_1_U15.reset ;
assign \add_38s_38s_38_2_1_U15.dout  = \add_38s_38s_38_2_1_U15.top_add_38s_38s_38_2_1_Adder_10_U.s ;
assign \add_38s_38s_38_2_1_U15.ce  = 1'h1;
assign \add_38s_38s_38_2_1_U15.clk  = ap_clk;
assign \add_38s_38s_38_2_1_U15.din0  = { op_25_V_reg_1342[31], op_25_V_reg_1342, 5'h00 };
assign \add_38s_38s_38_2_1_U15.din1  = { op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16[7], op_16 };
assign grp_fu_842_p2 = \add_38s_38s_38_2_1_U15.dout ;
assign \add_38s_38s_38_2_1_U15.reset  = ap_rst;
assign \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_8_U.ain_s0  = \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_8_U.a ;
assign \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_8_U.bin_s0  = \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_8_U.b ;
assign \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_8_U.s  = { \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_8_U.fas_s2 , \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_8_U.sum_s1  };
assign \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_8_U.u2.a  = \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_8_U.ain_s1 ;
assign \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_8_U.u2.b  = \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_8_U.bin_s1 ;
assign \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_8_U.u2.cin  = \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_8_U.carry_s1 ;
assign \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_8_U.facout_s2  = \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_8_U.u2.cout ;
assign \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_8_U.fas_s2  = \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_8_U.u2.s ;
assign \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_8_U.u1.a  = \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_8_U.a [16:0];
assign \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_8_U.u1.b  = \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_8_U.b [16:0];
assign \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_8_U.u1.cin  = 1'h0;
assign \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_8_U.facout_s1  = \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_8_U.u1.cout ;
assign \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_8_U.fas_s1  = \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_8_U.u1.s ;
assign \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_8_U.a  = \add_34s_34s_34_2_1_U10.din0 ;
assign \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_8_U.b  = \add_34s_34s_34_2_1_U10.din1 ;
assign \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_8_U.ce  = \add_34s_34s_34_2_1_U10.ce ;
assign \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_8_U.clk  = \add_34s_34s_34_2_1_U10.clk ;
assign \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_8_U.reset  = \add_34s_34s_34_2_1_U10.reset ;
assign \add_34s_34s_34_2_1_U10.dout  = \add_34s_34s_34_2_1_U10.top_add_34s_34s_34_2_1_Adder_8_U.s ;
assign \add_34s_34s_34_2_1_U10.ce  = 1'h1;
assign \add_34s_34s_34_2_1_U10.clk  = ap_clk;
assign \add_34s_34s_34_2_1_U10.din0  = { select_ln353_reg_1264[31], select_ln353_reg_1264, 1'h0 };
assign \add_34s_34s_34_2_1_U10.din1  = 34'h3ffffffff;
assign grp_fu_711_p2 = \add_34s_34s_34_2_1_U10.dout ;
assign \add_34s_34s_34_2_1_U10.reset  = ap_rst;
assign \add_34ns_34s_34_2_1_U2.top_add_34ns_34s_34_2_1_Adder_1_U.ain_s0  = \add_34ns_34s_34_2_1_U2.top_add_34ns_34s_34_2_1_Adder_1_U.a ;
assign \add_34ns_34s_34_2_1_U2.top_add_34ns_34s_34_2_1_Adder_1_U.bin_s0  = \add_34ns_34s_34_2_1_U2.top_add_34ns_34s_34_2_1_Adder_1_U.b ;
assign \add_34ns_34s_34_2_1_U2.top_add_34ns_34s_34_2_1_Adder_1_U.s  = { \add_34ns_34s_34_2_1_U2.top_add_34ns_34s_34_2_1_Adder_1_U.fas_s2 , \add_34ns_34s_34_2_1_U2.top_add_34ns_34s_34_2_1_Adder_1_U.sum_s1  };
assign \add_34ns_34s_34_2_1_U2.top_add_34ns_34s_34_2_1_Adder_1_U.u2.a  = \add_34ns_34s_34_2_1_U2.top_add_34ns_34s_34_2_1_Adder_1_U.ain_s1 ;
assign \add_34ns_34s_34_2_1_U2.top_add_34ns_34s_34_2_1_Adder_1_U.u2.b  = \add_34ns_34s_34_2_1_U2.top_add_34ns_34s_34_2_1_Adder_1_U.bin_s1 ;
assign \add_34ns_34s_34_2_1_U2.top_add_34ns_34s_34_2_1_Adder_1_U.u2.cin  = \add_34ns_34s_34_2_1_U2.top_add_34ns_34s_34_2_1_Adder_1_U.carry_s1 ;
assign \add_34ns_34s_34_2_1_U2.top_add_34ns_34s_34_2_1_Adder_1_U.facout_s2  = \add_34ns_34s_34_2_1_U2.top_add_34ns_34s_34_2_1_Adder_1_U.u2.cout ;
assign \add_34ns_34s_34_2_1_U2.top_add_34ns_34s_34_2_1_Adder_1_U.fas_s2  = \add_34ns_34s_34_2_1_U2.top_add_34ns_34s_34_2_1_Adder_1_U.u2.s ;
assign \add_34ns_34s_34_2_1_U2.top_add_34ns_34s_34_2_1_Adder_1_U.u1.a  = \add_34ns_34s_34_2_1_U2.top_add_34ns_34s_34_2_1_Adder_1_U.a [16:0];
assign \add_34ns_34s_34_2_1_U2.top_add_34ns_34s_34_2_1_Adder_1_U.u1.b  = \add_34ns_34s_34_2_1_U2.top_add_34ns_34s_34_2_1_Adder_1_U.b [16:0];
assign \add_34ns_34s_34_2_1_U2.top_add_34ns_34s_34_2_1_Adder_1_U.u1.cin  = 1'h0;
assign \add_34ns_34s_34_2_1_U2.top_add_34ns_34s_34_2_1_Adder_1_U.facout_s1  = \add_34ns_34s_34_2_1_U2.top_add_34ns_34s_34_2_1_Adder_1_U.u1.cout ;
assign \add_34ns_34s_34_2_1_U2.top_add_34ns_34s_34_2_1_Adder_1_U.fas_s1  = \add_34ns_34s_34_2_1_U2.top_add_34ns_34s_34_2_1_Adder_1_U.u1.s ;
assign \add_34ns_34s_34_2_1_U2.top_add_34ns_34s_34_2_1_Adder_1_U.a  = \add_34ns_34s_34_2_1_U2.din0 ;
assign \add_34ns_34s_34_2_1_U2.top_add_34ns_34s_34_2_1_Adder_1_U.b  = \add_34ns_34s_34_2_1_U2.din1 ;
assign \add_34ns_34s_34_2_1_U2.top_add_34ns_34s_34_2_1_Adder_1_U.ce  = \add_34ns_34s_34_2_1_U2.ce ;
assign \add_34ns_34s_34_2_1_U2.top_add_34ns_34s_34_2_1_Adder_1_U.clk  = \add_34ns_34s_34_2_1_U2.clk ;
assign \add_34ns_34s_34_2_1_U2.top_add_34ns_34s_34_2_1_Adder_1_U.reset  = \add_34ns_34s_34_2_1_U2.reset ;
assign \add_34ns_34s_34_2_1_U2.dout  = \add_34ns_34s_34_2_1_U2.top_add_34ns_34s_34_2_1_Adder_1_U.s ;
assign \add_34ns_34s_34_2_1_U2.ce  = 1'h1;
assign \add_34ns_34s_34_2_1_U2.clk  = ap_clk;
assign \add_34ns_34s_34_2_1_U2.din0  = { 2'h0, op_3 };
assign \add_34ns_34s_34_2_1_U2.din1  = { ret_V_18_reg_1037[1], ret_V_18_reg_1037[1], ret_V_18_reg_1037[1], ret_V_18_reg_1037[1], ret_V_18_reg_1037[1], ret_V_18_reg_1037[1], ret_V_18_reg_1037[1], ret_V_18_reg_1037[1], ret_V_18_reg_1037[1], ret_V_18_reg_1037[1], ret_V_18_reg_1037[1], ret_V_18_reg_1037[1], ret_V_18_reg_1037[1], ret_V_18_reg_1037[1], ret_V_18_reg_1037[1], ret_V_18_reg_1037[1], ret_V_18_reg_1037[1], ret_V_18_reg_1037[1], ret_V_18_reg_1037[1], ret_V_18_reg_1037[1], ret_V_18_reg_1037[1], ret_V_18_reg_1037[1], ret_V_18_reg_1037[1], ret_V_18_reg_1037[1], ret_V_18_reg_1037[1], ret_V_18_reg_1037[1], ret_V_18_reg_1037[1], ret_V_18_reg_1037[1], ret_V_18_reg_1037[1], ret_V_18_reg_1037[1], ret_V_18_reg_1037[1], ret_V_18_reg_1037[1], ret_V_18_reg_1037 };
assign grp_fu_316_p2 = \add_34ns_34s_34_2_1_U2.dout ;
assign \add_34ns_34s_34_2_1_U2.reset  = ap_rst;
assign \add_32s_32ns_32_2_1_U7.top_add_32s_32ns_32_2_1_Adder_5_U.ain_s0  = \add_32s_32ns_32_2_1_U7.top_add_32s_32ns_32_2_1_Adder_5_U.a ;
assign \add_32s_32ns_32_2_1_U7.top_add_32s_32ns_32_2_1_Adder_5_U.bin_s0  = \add_32s_32ns_32_2_1_U7.top_add_32s_32ns_32_2_1_Adder_5_U.b ;
assign \add_32s_32ns_32_2_1_U7.top_add_32s_32ns_32_2_1_Adder_5_U.s  = { \add_32s_32ns_32_2_1_U7.top_add_32s_32ns_32_2_1_Adder_5_U.fas_s2 , \add_32s_32ns_32_2_1_U7.top_add_32s_32ns_32_2_1_Adder_5_U.sum_s1  };
assign \add_32s_32ns_32_2_1_U7.top_add_32s_32ns_32_2_1_Adder_5_U.u2.a  = \add_32s_32ns_32_2_1_U7.top_add_32s_32ns_32_2_1_Adder_5_U.ain_s1 ;
assign \add_32s_32ns_32_2_1_U7.top_add_32s_32ns_32_2_1_Adder_5_U.u2.b  = \add_32s_32ns_32_2_1_U7.top_add_32s_32ns_32_2_1_Adder_5_U.bin_s1 ;
assign \add_32s_32ns_32_2_1_U7.top_add_32s_32ns_32_2_1_Adder_5_U.u2.cin  = \add_32s_32ns_32_2_1_U7.top_add_32s_32ns_32_2_1_Adder_5_U.carry_s1 ;
assign \add_32s_32ns_32_2_1_U7.top_add_32s_32ns_32_2_1_Adder_5_U.facout_s2  = \add_32s_32ns_32_2_1_U7.top_add_32s_32ns_32_2_1_Adder_5_U.u2.cout ;
assign \add_32s_32ns_32_2_1_U7.top_add_32s_32ns_32_2_1_Adder_5_U.fas_s2  = \add_32s_32ns_32_2_1_U7.top_add_32s_32ns_32_2_1_Adder_5_U.u2.s ;
assign \add_32s_32ns_32_2_1_U7.top_add_32s_32ns_32_2_1_Adder_5_U.u1.a  = \add_32s_32ns_32_2_1_U7.top_add_32s_32ns_32_2_1_Adder_5_U.a [15:0];
assign \add_32s_32ns_32_2_1_U7.top_add_32s_32ns_32_2_1_Adder_5_U.u1.b  = \add_32s_32ns_32_2_1_U7.top_add_32s_32ns_32_2_1_Adder_5_U.b [15:0];
assign \add_32s_32ns_32_2_1_U7.top_add_32s_32ns_32_2_1_Adder_5_U.u1.cin  = 1'h0;
assign \add_32s_32ns_32_2_1_U7.top_add_32s_32ns_32_2_1_Adder_5_U.facout_s1  = \add_32s_32ns_32_2_1_U7.top_add_32s_32ns_32_2_1_Adder_5_U.u1.cout ;
assign \add_32s_32ns_32_2_1_U7.top_add_32s_32ns_32_2_1_Adder_5_U.fas_s1  = \add_32s_32ns_32_2_1_U7.top_add_32s_32ns_32_2_1_Adder_5_U.u1.s ;
assign \add_32s_32ns_32_2_1_U7.top_add_32s_32ns_32_2_1_Adder_5_U.a  = \add_32s_32ns_32_2_1_U7.din0 ;
assign \add_32s_32ns_32_2_1_U7.top_add_32s_32ns_32_2_1_Adder_5_U.b  = \add_32s_32ns_32_2_1_U7.din1 ;
assign \add_32s_32ns_32_2_1_U7.top_add_32s_32ns_32_2_1_Adder_5_U.ce  = \add_32s_32ns_32_2_1_U7.ce ;
assign \add_32s_32ns_32_2_1_U7.top_add_32s_32ns_32_2_1_Adder_5_U.clk  = \add_32s_32ns_32_2_1_U7.clk ;
assign \add_32s_32ns_32_2_1_U7.top_add_32s_32ns_32_2_1_Adder_5_U.reset  = \add_32s_32ns_32_2_1_U7.reset ;
assign \add_32s_32ns_32_2_1_U7.dout  = \add_32s_32ns_32_2_1_U7.top_add_32s_32ns_32_2_1_Adder_5_U.s ;
assign \add_32s_32ns_32_2_1_U7.ce  = 1'h1;
assign \add_32s_32ns_32_2_1_U7.clk  = ap_clk;
assign \add_32s_32ns_32_2_1_U7.din0  = { ret_V_17_reg_1159[3], ret_V_17_reg_1159[3], ret_V_17_reg_1159[3], ret_V_17_reg_1159[3], ret_V_17_reg_1159[3], ret_V_17_reg_1159[3], ret_V_17_reg_1159[3], ret_V_17_reg_1159[3], ret_V_17_reg_1159[3], ret_V_17_reg_1159[3], ret_V_17_reg_1159[3], ret_V_17_reg_1159[3], ret_V_17_reg_1159[3], ret_V_17_reg_1159[3], ret_V_17_reg_1159[3], ret_V_17_reg_1159[3], ret_V_17_reg_1159[3], ret_V_17_reg_1159[3], ret_V_17_reg_1159[3], ret_V_17_reg_1159[3], ret_V_17_reg_1159[3], ret_V_17_reg_1159[3], ret_V_17_reg_1159[3], ret_V_17_reg_1159[3], ret_V_17_reg_1159[3], ret_V_17_reg_1159[3], ret_V_17_reg_1159[3], ret_V_17_reg_1159[3], ret_V_17_reg_1159 };
assign \add_32s_32ns_32_2_1_U7.din1  = op_8;
assign grp_fu_509_p2 = \add_32s_32ns_32_2_1_U7.dout ;
assign \add_32s_32ns_32_2_1_U7.reset  = ap_rst;
assign \add_32ns_32s_32_2_1_U21.top_add_32ns_32s_32_2_1_Adder_12_U.ain_s0  = \add_32ns_32s_32_2_1_U21.top_add_32ns_32s_32_2_1_Adder_12_U.a ;
assign \add_32ns_32s_32_2_1_U21.top_add_32ns_32s_32_2_1_Adder_12_U.bin_s0  = \add_32ns_32s_32_2_1_U21.top_add_32ns_32s_32_2_1_Adder_12_U.b ;
assign \add_32ns_32s_32_2_1_U21.top_add_32ns_32s_32_2_1_Adder_12_U.s  = { \add_32ns_32s_32_2_1_U21.top_add_32ns_32s_32_2_1_Adder_12_U.fas_s2 , \add_32ns_32s_32_2_1_U21.top_add_32ns_32s_32_2_1_Adder_12_U.sum_s1  };
assign \add_32ns_32s_32_2_1_U21.top_add_32ns_32s_32_2_1_Adder_12_U.u2.a  = \add_32ns_32s_32_2_1_U21.top_add_32ns_32s_32_2_1_Adder_12_U.ain_s1 ;
assign \add_32ns_32s_32_2_1_U21.top_add_32ns_32s_32_2_1_Adder_12_U.u2.b  = \add_32ns_32s_32_2_1_U21.top_add_32ns_32s_32_2_1_Adder_12_U.bin_s1 ;
assign \add_32ns_32s_32_2_1_U21.top_add_32ns_32s_32_2_1_Adder_12_U.u2.cin  = \add_32ns_32s_32_2_1_U21.top_add_32ns_32s_32_2_1_Adder_12_U.carry_s1 ;
assign \add_32ns_32s_32_2_1_U21.top_add_32ns_32s_32_2_1_Adder_12_U.facout_s2  = \add_32ns_32s_32_2_1_U21.top_add_32ns_32s_32_2_1_Adder_12_U.u2.cout ;
assign \add_32ns_32s_32_2_1_U21.top_add_32ns_32s_32_2_1_Adder_12_U.fas_s2  = \add_32ns_32s_32_2_1_U21.top_add_32ns_32s_32_2_1_Adder_12_U.u2.s ;
assign \add_32ns_32s_32_2_1_U21.top_add_32ns_32s_32_2_1_Adder_12_U.u1.a  = \add_32ns_32s_32_2_1_U21.top_add_32ns_32s_32_2_1_Adder_12_U.a [15:0];
assign \add_32ns_32s_32_2_1_U21.top_add_32ns_32s_32_2_1_Adder_12_U.u1.b  = \add_32ns_32s_32_2_1_U21.top_add_32ns_32s_32_2_1_Adder_12_U.b [15:0];
assign \add_32ns_32s_32_2_1_U21.top_add_32ns_32s_32_2_1_Adder_12_U.u1.cin  = 1'h0;
assign \add_32ns_32s_32_2_1_U21.top_add_32ns_32s_32_2_1_Adder_12_U.facout_s1  = \add_32ns_32s_32_2_1_U21.top_add_32ns_32s_32_2_1_Adder_12_U.u1.cout ;
assign \add_32ns_32s_32_2_1_U21.top_add_32ns_32s_32_2_1_Adder_12_U.fas_s1  = \add_32ns_32s_32_2_1_U21.top_add_32ns_32s_32_2_1_Adder_12_U.u1.s ;
assign \add_32ns_32s_32_2_1_U21.top_add_32ns_32s_32_2_1_Adder_12_U.a  = \add_32ns_32s_32_2_1_U21.din0 ;
assign \add_32ns_32s_32_2_1_U21.top_add_32ns_32s_32_2_1_Adder_12_U.b  = \add_32ns_32s_32_2_1_U21.din1 ;
assign \add_32ns_32s_32_2_1_U21.top_add_32ns_32s_32_2_1_Adder_12_U.ce  = \add_32ns_32s_32_2_1_U21.ce ;
assign \add_32ns_32s_32_2_1_U21.top_add_32ns_32s_32_2_1_Adder_12_U.clk  = \add_32ns_32s_32_2_1_U21.clk ;
assign \add_32ns_32s_32_2_1_U21.top_add_32ns_32s_32_2_1_Adder_12_U.reset  = \add_32ns_32s_32_2_1_U21.reset ;
assign \add_32ns_32s_32_2_1_U21.dout  = \add_32ns_32s_32_2_1_U21.top_add_32ns_32s_32_2_1_Adder_12_U.s ;
assign \add_32ns_32s_32_2_1_U21.ce  = 1'h1;
assign \add_32ns_32s_32_2_1_U21.clk  = ap_clk;
assign \add_32ns_32s_32_2_1_U21.din0  = op_28_V_reg_1436;
assign \add_32ns_32s_32_2_1_U21.din1  = { trunc_ln2_reg_1421[3], trunc_ln2_reg_1421[3], trunc_ln2_reg_1421[3], trunc_ln2_reg_1421[3], trunc_ln2_reg_1421[3], trunc_ln2_reg_1421[3], trunc_ln2_reg_1421[3], trunc_ln2_reg_1421[3], trunc_ln2_reg_1421[3], trunc_ln2_reg_1421[3], trunc_ln2_reg_1421[3], trunc_ln2_reg_1421[3], trunc_ln2_reg_1421[3], trunc_ln2_reg_1421[3], trunc_ln2_reg_1421[3], trunc_ln2_reg_1421[3], trunc_ln2_reg_1421[3], trunc_ln2_reg_1421[3], trunc_ln2_reg_1421[3], trunc_ln2_reg_1421[3], trunc_ln2_reg_1421[3], trunc_ln2_reg_1421[3], trunc_ln2_reg_1421[3], trunc_ln2_reg_1421[3], trunc_ln2_reg_1421[3], trunc_ln2_reg_1421[3], trunc_ln2_reg_1421[3], trunc_ln2_reg_1421[3], trunc_ln2_reg_1421 };
assign grp_fu_1010_p2 = \add_32ns_32s_32_2_1_U21.dout ;
assign \add_32ns_32s_32_2_1_U21.reset  = ap_rst;
assign \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_12_U.ain_s0  = \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_12_U.a ;
assign \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_12_U.bin_s0  = \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_12_U.b ;
assign \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_12_U.s  = { \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_12_U.fas_s2 , \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_12_U.sum_s1  };
assign \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_12_U.u2.a  = \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_12_U.ain_s1 ;
assign \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_12_U.u2.b  = \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_12_U.bin_s1 ;
assign \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_12_U.u2.cin  = \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_12_U.carry_s1 ;
assign \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_12_U.facout_s2  = \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_12_U.u2.cout ;
assign \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_12_U.fas_s2  = \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_12_U.u2.s ;
assign \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_12_U.u1.a  = \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_12_U.a [15:0];
assign \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_12_U.u1.b  = \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_12_U.b [15:0];
assign \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_12_U.u1.cin  = 1'h0;
assign \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_12_U.facout_s1  = \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_12_U.u1.cout ;
assign \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_12_U.fas_s1  = \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_12_U.u1.s ;
assign \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_12_U.a  = \add_32ns_32s_32_2_1_U20.din0 ;
assign \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_12_U.b  = \add_32ns_32s_32_2_1_U20.din1 ;
assign \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_12_U.ce  = \add_32ns_32s_32_2_1_U20.ce ;
assign \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_12_U.clk  = \add_32ns_32s_32_2_1_U20.clk ;
assign \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_12_U.reset  = \add_32ns_32s_32_2_1_U20.reset ;
assign \add_32ns_32s_32_2_1_U20.dout  = \add_32ns_32s_32_2_1_U20.top_add_32ns_32s_32_2_1_Adder_12_U.s ;
assign \add_32ns_32s_32_2_1_U20.ce  = 1'h1;
assign \add_32ns_32s_32_2_1_U20.clk  = ap_clk;
assign \add_32ns_32s_32_2_1_U20.din0  = ret_V_25_reg_1426;
assign \add_32ns_32s_32_2_1_U20.din1  = { op_18_V_reg_1416[3], op_18_V_reg_1416[3], op_18_V_reg_1416[3], op_18_V_reg_1416[3], op_18_V_reg_1416[3], op_18_V_reg_1416[3], op_18_V_reg_1416[3], op_18_V_reg_1416[3], op_18_V_reg_1416[3], op_18_V_reg_1416[3], op_18_V_reg_1416[3], op_18_V_reg_1416[3], op_18_V_reg_1416[3], op_18_V_reg_1416[3], op_18_V_reg_1416[3], op_18_V_reg_1416[3], op_18_V_reg_1416[3], op_18_V_reg_1416[3], op_18_V_reg_1416[3], op_18_V_reg_1416[3], op_18_V_reg_1416[3], op_18_V_reg_1416[3], op_18_V_reg_1416[3], op_18_V_reg_1416[3], op_18_V_reg_1416[3], op_18_V_reg_1416[3], op_18_V_reg_1416[3], op_18_V_reg_1416[3], op_18_V_reg_1416 };
assign grp_fu_1002_p2 = \add_32ns_32s_32_2_1_U20.dout ;
assign \add_32ns_32s_32_2_1_U20.reset  = ap_rst;
assign \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s0  = \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.a ;
assign \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s0  = \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.b ;
assign \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.s  = { \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s2 , \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.sum_s1  };
assign \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.a  = \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s1 ;
assign \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.b  = \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s1 ;
assign \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cin  = \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.carry_s1 ;
assign \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.facout_s2  = \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cout ;
assign \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s2  = \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.s ;
assign \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.a  = \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.a [15:0];
assign \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.b  = \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.b [15:0];
assign \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cin  = 1'h0;
assign \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.facout_s1  = \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cout ;
assign \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s1  = \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.s ;
assign \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.a  = \add_32ns_32ns_32_2_1_U9.din0 ;
assign \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.b  = \add_32ns_32ns_32_2_1_U9.din1 ;
assign \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.ce  = \add_32ns_32ns_32_2_1_U9.ce ;
assign \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.clk  = \add_32ns_32ns_32_2_1_U9.clk ;
assign \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.reset  = \add_32ns_32ns_32_2_1_U9.reset ;
assign \add_32ns_32ns_32_2_1_U9.dout  = \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.s ;
assign \add_32ns_32ns_32_2_1_U9.ce  = 1'h1;
assign \add_32ns_32ns_32_2_1_U9.clk  = ap_clk;
assign \add_32ns_32ns_32_2_1_U9.din0  = ret_V_8_cast_reg_1252;
assign \add_32ns_32ns_32_2_1_U9.din1  = 32'd1;
assign grp_fu_676_p2 = \add_32ns_32ns_32_2_1_U9.dout ;
assign \add_32ns_32ns_32_2_1_U9.reset  = ap_rst;
assign \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s0  = \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.a ;
assign \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s0  = \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.b ;
assign \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.s  = { \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s2 , \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.sum_s1  };
assign \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.a  = \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s1 ;
assign \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.b  = \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s1 ;
assign \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cin  = \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.carry_s1 ;
assign \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.facout_s2  = \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cout ;
assign \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s2  = \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.s ;
assign \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.a  = \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.a [15:0];
assign \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.b  = \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.b [15:0];
assign \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cin  = 1'h0;
assign \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.facout_s1  = \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cout ;
assign \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s1  = \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.s ;
assign \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.a  = \add_32ns_32ns_32_2_1_U18.din0 ;
assign \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.b  = \add_32ns_32ns_32_2_1_U18.din1 ;
assign \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.ce  = \add_32ns_32ns_32_2_1_U18.ce ;
assign \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.clk  = \add_32ns_32ns_32_2_1_U18.clk ;
assign \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.reset  = \add_32ns_32ns_32_2_1_U18.reset ;
assign \add_32ns_32ns_32_2_1_U18.dout  = \add_32ns_32ns_32_2_1_U18.top_add_32ns_32ns_32_2_1_Adder_7_U.s ;
assign \add_32ns_32ns_32_2_1_U18.ce  = 1'h1;
assign \add_32ns_32ns_32_2_1_U18.clk  = ap_clk;
assign \add_32ns_32ns_32_2_1_U18.din0  = ret_V_26_cast_reg_1404;
assign \add_32ns_32ns_32_2_1_U18.din1  = 32'd1;
assign grp_fu_933_p2 = \add_32ns_32ns_32_2_1_U18.dout ;
assign \add_32ns_32ns_32_2_1_U18.reset  = ap_rst;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s0  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.a ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s0  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.b ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.s  = { \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s2 , \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.sum_s1  };
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.a  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s1 ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.b  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s1 ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cin  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.carry_s1 ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.facout_s2  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cout ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s2  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.s ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.a  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.a [15:0];
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.b  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.b [15:0];
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cin  = 1'h0;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.facout_s1  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cout ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s1  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.s ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.a  = \add_32ns_32ns_32_2_1_U16.din0 ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.b  = \add_32ns_32ns_32_2_1_U16.din1 ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.ce  = \add_32ns_32ns_32_2_1_U16.ce ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.clk  = \add_32ns_32ns_32_2_1_U16.clk ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.reset  = \add_32ns_32ns_32_2_1_U16.reset ;
assign \add_32ns_32ns_32_2_1_U16.dout  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.s ;
assign \add_32ns_32ns_32_2_1_U16.ce  = 1'h1;
assign \add_32ns_32ns_32_2_1_U16.clk  = ap_clk;
assign \add_32ns_32ns_32_2_1_U16.din0  = ret_V_24_cast_reg_1367;
assign \add_32ns_32ns_32_2_1_U16.din1  = 32'd1;
assign grp_fu_868_p2 = \add_32ns_32ns_32_2_1_U16.dout ;
assign \add_32ns_32ns_32_2_1_U16.reset  = ap_rst;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s0  = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.a ;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s0  = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.b ;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.s  = { \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s2 , \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.sum_s1  };
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.a  = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s1 ;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.b  = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s1 ;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cin  = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.carry_s1 ;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.facout_s2  = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cout ;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s2  = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.s ;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.a  = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.a [15:0];
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.b  = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.b [15:0];
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cin  = 1'h0;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.facout_s1  = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cout ;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s1  = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.s ;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.a  = \add_32ns_32ns_32_2_1_U14.din0 ;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.b  = \add_32ns_32ns_32_2_1_U14.din1 ;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.ce  = \add_32ns_32ns_32_2_1_U14.ce ;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.clk  = \add_32ns_32ns_32_2_1_U14.clk ;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.reset  = \add_32ns_32ns_32_2_1_U14.reset ;
assign \add_32ns_32ns_32_2_1_U14.dout  = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.s ;
assign \add_32ns_32ns_32_2_1_U14.ce  = 1'h1;
assign \add_32ns_32ns_32_2_1_U14.clk  = ap_clk;
assign \add_32ns_32ns_32_2_1_U14.din0  = ret_V_22_reg_1332;
assign \add_32ns_32ns_32_2_1_U14.din1  = { 30'h00000000, r_reg_1327 };
assign grp_fu_822_p2 = \add_32ns_32ns_32_2_1_U14.dout ;
assign \add_32ns_32ns_32_2_1_U14.reset  = ap_rst;
assign \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s0  = \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_7_U.a ;
assign \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s0  = \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_7_U.b ;
assign \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_7_U.s  = { \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s2 , \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_7_U.sum_s1  };
assign \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.a  = \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s1 ;
assign \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.b  = \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s1 ;
assign \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cin  = \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_7_U.carry_s1 ;
assign \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_7_U.facout_s2  = \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cout ;
assign \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s2  = \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.s ;
assign \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.a  = \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_7_U.a [15:0];
assign \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.b  = \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_7_U.b [15:0];
assign \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cin  = 1'h0;
assign \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_7_U.facout_s1  = \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cout ;
assign \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s1  = \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.s ;
assign \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_7_U.a  = \add_32ns_32ns_32_2_1_U13.din0 ;
assign \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_7_U.b  = \add_32ns_32ns_32_2_1_U13.din1 ;
assign \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_7_U.ce  = \add_32ns_32ns_32_2_1_U13.ce ;
assign \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_7_U.clk  = \add_32ns_32ns_32_2_1_U13.clk ;
assign \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_7_U.reset  = \add_32ns_32ns_32_2_1_U13.reset ;
assign \add_32ns_32ns_32_2_1_U13.dout  = \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_7_U.s ;
assign \add_32ns_32ns_32_2_1_U13.ce  = 1'h1;
assign \add_32ns_32ns_32_2_1_U13.clk  = ap_clk;
assign \add_32ns_32ns_32_2_1_U13.din0  = ret_V_22_cast_reg_1315;
assign \add_32ns_32ns_32_2_1_U13.din1  = 32'd1;
assign grp_fu_786_p2 = \add_32ns_32ns_32_2_1_U13.dout ;
assign \add_32ns_32ns_32_2_1_U13.reset  = ap_rst;
assign \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s0  = \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.a ;
assign \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s0  = \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.b ;
assign \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.s  = { \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s2 , \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.sum_s1  };
assign \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.a  = \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s1 ;
assign \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.b  = \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s1 ;
assign \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cin  = \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.carry_s1 ;
assign \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.facout_s2  = \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cout ;
assign \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s2  = \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.s ;
assign \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.a  = \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.a [15:0];
assign \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.b  = \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.b [15:0];
assign \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cin  = 1'h0;
assign \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.facout_s1  = \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cout ;
assign \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s1  = \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.s ;
assign \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.a  = \add_32ns_32ns_32_2_1_U11.din0 ;
assign \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.b  = \add_32ns_32ns_32_2_1_U11.din1 ;
assign \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.ce  = \add_32ns_32ns_32_2_1_U11.ce ;
assign \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.clk  = \add_32ns_32ns_32_2_1_U11.clk ;
assign \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.reset  = \add_32ns_32ns_32_2_1_U11.reset ;
assign \add_32ns_32ns_32_2_1_U11.dout  = \add_32ns_32ns_32_2_1_U11.top_add_32ns_32ns_32_2_1_Adder_7_U.s ;
assign \add_32ns_32ns_32_2_1_U11.ce  = 1'h1;
assign \add_32ns_32ns_32_2_1_U11.clk  = ap_clk;
assign \add_32ns_32ns_32_2_1_U11.din0  = tmp_2_reg_1279;
assign \add_32ns_32ns_32_2_1_U11.din1  = 32'd1;
assign grp_fu_735_p2 = \add_32ns_32ns_32_2_1_U11.dout ;
assign \add_32ns_32ns_32_2_1_U11.reset  = ap_rst;
assign \add_2ns_2ns_2_1_1_U1.top_add_2ns_2ns_2_1_1_Adder_0_U.a  = \add_2ns_2ns_2_1_1_U1.din0 ;
assign \add_2ns_2ns_2_1_1_U1.top_add_2ns_2ns_2_1_1_Adder_0_U.b  = \add_2ns_2ns_2_1_1_U1.din1 ;
assign \add_2ns_2ns_2_1_1_U1.dout  = \add_2ns_2ns_2_1_1_U1.top_add_2ns_2ns_2_1_1_Adder_0_U.s ;
assign \add_2ns_2ns_2_1_1_U1.din0  = op_2[3:2];
assign \add_2ns_2ns_2_1_1_U1.din1  = 2'h1;
assign ret_V_5_fu_251_p2 = \add_2ns_2ns_2_1_1_U1.dout ;
assign \add_10ns_10s_10_1_1_U5.top_add_10ns_10s_10_1_1_Adder_4_U.a  = \add_10ns_10s_10_1_1_U5.din0 ;
assign \add_10ns_10s_10_1_1_U5.top_add_10ns_10s_10_1_1_Adder_4_U.b  = \add_10ns_10s_10_1_1_U5.din1 ;
assign \add_10ns_10s_10_1_1_U5.dout  = \add_10ns_10s_10_1_1_U5.top_add_10ns_10s_10_1_1_Adder_4_U.s ;
assign \add_10ns_10s_10_1_1_U5.din0  = empty_reg_1058;
assign \add_10ns_10s_10_1_1_U5.din1  = { ret_V_18_reg_1037[1], ret_V_18_reg_1037[1], ret_V_18_reg_1037[1], ret_V_18_reg_1037[1], ret_V_18_reg_1037[1], ret_V_18_reg_1037[1], ret_V_18_reg_1037[1], ret_V_18_reg_1037[1], ret_V_18_reg_1037 };
assign add_ln1346_1_fu_419_p2 = \add_10ns_10s_10_1_1_U5.dout ;
endmodule


// Product machine:
module top_A_times_top_B (ap_start, op_0, op_1, op_13, op_16, op_17, op_2, op_3, op_7, op_8, ap_clk, unsafe_signal);
input ap_start;
input [7:0] op_0;
input op_1;
input [31:0] op_13;
input [7:0] op_16;
input [7:0] op_17;
input [3:0] op_2;
input [31:0] op_3;
input [3:0] op_7;
input [31:0] op_8;
input ap_clk;
output unsafe_signal;
reg _setup;
initial _setup = 1'b0;
always @ (posedge ap_clk) _setup <= 1'b1;
reg ap_start_internal;
always @ (posedge ap_clk) if (!_setup) ap_start_internal <= ap_start;
reg [7:0] op_0_internal;
always @ (posedge ap_clk) if (!_setup) op_0_internal <= op_0;
reg op_1_internal;
always @ (posedge ap_clk) if (!_setup) op_1_internal <= op_1;
reg [31:0] op_13_internal;
always @ (posedge ap_clk) if (!_setup) op_13_internal <= op_13;
reg [7:0] op_16_internal;
always @ (posedge ap_clk) if (!_setup) op_16_internal <= op_16;
reg [7:0] op_17_internal;
always @ (posedge ap_clk) if (!_setup) op_17_internal <= op_17;
reg [3:0] op_2_internal;
always @ (posedge ap_clk) if (!_setup) op_2_internal <= op_2;
reg [31:0] op_3_internal;
always @ (posedge ap_clk) if (!_setup) op_3_internal <= op_3;
reg [3:0] op_7_internal;
always @ (posedge ap_clk) if (!_setup) op_7_internal <= op_7;
reg [31:0] op_8_internal;
always @ (posedge ap_clk) if (!_setup) op_8_internal <= op_8;
wire ap_done_A;
wire ap_done_B;
wire ap_done_eq;
assign ap_done_eq = ap_done_A == ap_done_B;
wire ap_idle_A;
wire ap_idle_B;
wire ap_idle_eq;
assign ap_idle_eq = ap_idle_A == ap_idle_B;
wire ap_ready_A;
wire ap_ready_B;
wire ap_ready_eq;
assign ap_ready_eq = ap_ready_A == ap_ready_B;
wire [31:0] op_29_A;
wire [31:0] op_29_B;
wire op_29_eq;
assign op_29_eq = op_29_A == op_29_B;
wire op_29_ap_vld_A;
wire op_29_ap_vld_B;
wire clk_enable_A;
wire clk_enable_B;
assign clk_enable_A = _setup & (~op_29_ap_vld_A | op_29_ap_vld_B);
assign clk_enable_B = _setup;
wire divergent;
assign divergent = ~(ap_done_eq & ap_idle_eq & ap_ready_eq & op_29_eq);
assign unsafe_signal = op_29_ap_vld_A & op_29_ap_vld_B & divergent;
top_A instance_A (
    .ap_clk(ap_clk),
    .clk_enable(clk_enable_A),
    .ap_start(ap_start_internal),
    .op_0(op_0_internal),
    .op_1(op_1_internal),
    .op_13(op_13_internal),
    .op_16(op_16_internal),
    .op_17(op_17_internal),
    .op_2(op_2_internal),
    .op_3(op_3_internal),
    .op_7(op_7_internal),
    .op_8(op_8_internal),
    .ap_done(ap_done_A),
    .ap_idle(ap_idle_A),
    .ap_ready(ap_ready_A),
    .op_29(op_29_A),
    .op_29_ap_vld(op_29_ap_vld_A)
);
top_B instance_B (
    .ap_clk(ap_clk),
    .clk_enable(clk_enable_B),
    .ap_start(ap_start_internal),
    .op_0(op_0_internal),
    .op_1(op_1_internal),
    .op_13(op_13_internal),
    .op_16(op_16_internal),
    .op_17(op_17_internal),
    .op_2(op_2_internal),
    .op_3(op_3_internal),
    .op_7(op_7_internal),
    .op_8(op_8_internal),
    .ap_done(ap_done_B),
    .ap_idle(ap_idle_B),
    .ap_ready(ap_ready_B),
    .op_29(op_29_B),
    .op_29_ap_vld(op_29_ap_vld_B)
);
endmodule
