// Processed by function `construct_kairos` in `verilog_tricks.py`.
// Machine A:
// Processed by function `add_clk_enable_signal` in `verilog_tricks.py`.
// Processed by function `remove_reset_signal` in `verilog_tricks.py`.
module top_A (
  ap_clk,
  ap_start,
  ap_done,
  ap_idle,
  ap_ready,
  op_0,
  op_3,
  op_4,
  op_5,
  op_9,
  op_10,
  op_11,
  op_13,
  op_15,
  op_16,
  op_17,
  op_19,
  op_29,
  op_29_ap_vld,
clk_enable
);
input clk_enable;


input ap_clk;
wire ap_rst;
assign ap_rst = op_29_ap_vld;
input ap_start;
input op_0;
input [1:0] op_10;
input [15:0] op_11;
input [1:0] op_13;
input [3:0] op_15;
input [31:0] op_16;
input [3:0] op_17;
input [3:0] op_19;
input [3:0] op_3;
input [3:0] op_4;
input [3:0] op_5;
input [7:0] op_9;
output ap_done;
output ap_idle;
output ap_ready;
output [31:0] op_29;
output op_29_ap_vld;


reg [8:0] \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.ain_s1 ;
reg [8:0] \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.bin_s1 ;
reg \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.carry_s1 ;
reg [7:0] \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.sum_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s1 ;
reg \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.carry_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.sum_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s1 ;
reg \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.carry_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.sum_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s1 ;
reg \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.carry_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.sum_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s1 ;
reg \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.carry_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.sum_s1 ;
reg [15:0] \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.ain_s1 ;
reg [15:0] \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.bin_s1 ;
reg \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.carry_s1 ;
reg [15:0] \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.sum_s1 ;
reg [15:0] \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.ain_s1 ;
reg [15:0] \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.bin_s1 ;
reg \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.carry_s1 ;
reg [15:0] \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.sum_s1 ;
reg [16:0] \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.ain_s1 ;
reg [16:0] \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.bin_s1 ;
reg \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.carry_s1 ;
reg [16:0] \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.sum_s1 ;
reg [17:0] \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.ain_s1 ;
reg [17:0] \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.bin_s1 ;
reg \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.carry_s1 ;
reg [16:0] \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.sum_s1 ;
reg [17:0] \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.ain_s1 ;
reg [17:0] \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.bin_s1 ;
reg \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.carry_s1 ;
reg [16:0] \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.sum_s1 ;
reg [1:0] \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.ain_s1 ;
reg [1:0] \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.bin_s1 ;
reg \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.carry_s1 ;
reg \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.sum_s1 ;
reg [1:0] \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.ain_s1 ;
reg [1:0] \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.bin_s1 ;
reg \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.carry_s1 ;
reg [1:0] \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.sum_s1 ;
reg [2:0] \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.ain_s1 ;
reg [2:0] \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.bin_s1 ;
reg \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.carry_s1 ;
reg [1:0] \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.sum_s1 ;
reg [2:0] \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.ain_s1 ;
reg [2:0] \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.bin_s1 ;
reg \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.carry_s1 ;
reg [1:0] \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.sum_s1 ;
reg [2:0] \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.ain_s1 ;
reg [2:0] \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.bin_s1 ;
reg \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.carry_s1 ;
reg [1:0] \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.sum_s1 ;
reg [2:0] \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.ain_s1 ;
reg [2:0] \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.bin_s1 ;
reg \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.carry_s1 ;
reg [2:0] \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.sum_s1 ;
reg [4:0] \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.ain_s1 ;
reg [4:0] \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.bin_s1 ;
reg \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.carry_s1 ;
reg [3:0] \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.sum_s1 ;
reg [31:0] add_ln691_1_reg_1073;
reg [31:0] add_ln691_2_reg_1160;
reg [31:0] add_ln691_reg_953;
reg [31:0] add_ln69_2_reg_1098;
reg [8:0] add_ln69_reg_978;
reg [26:0] ap_CS_fsm = 27'h0000001;
reg icmp_ln785_reg_846;
reg icmp_ln786_1_reg_858;
reg icmp_ln786_reg_852;
reg icmp_ln851_1_reg_921;
reg icmp_ln851_2_reg_1143;
reg icmp_ln851_reg_906;
reg [3:0] op_14_V_reg_1083;
reg [31:0] op_24_V_reg_1008;
reg [31:0] op_27_V_reg_1113;
reg [1:0] p_Result_s_16_reg_840;
reg [4:0] ret_V_13_reg_1108;
reg [4:0] ret_V_21_reg_1055;
reg [5:0] ret_V_24_reg_941;
reg [4:0] ret_V_25_reg_995;
reg [2:0] ret_V_27_reg_901;
reg [16:0] ret_V_28_reg_931;
reg [31:0] ret_V_29_reg_973;
reg [33:0] ret_V_30_reg_1033;
reg [31:0] ret_V_31_reg_1093;
reg [34:0] ret_V_32_reg_1148;
reg [31:0] ret_V_33_cast_reg_1038;
reg [31:0] ret_V_36_cast_reg_1153;
reg [5:0] ret_V_3_reg_889;
reg [5:0] ret_V_5_reg_926;
reg [3:0] ret_V_8_cast_reg_1001;
reg [3:0] ret_V_8_reg_1028;
reg [1:0] ret_V_9_reg_869;
reg [4:0] select_ln1192_reg_968;
reg [1:0] select_ln340_reg_864;
reg [3:0] select_ln353_reg_1045;
reg [4:0] select_ln703_reg_1088;
reg [4:0] sext_ln703_reg_983;
reg [31:0] sext_ln831_reg_946;
reg tmp_2_reg_822;
reg tmp_3_reg_834;
reg [31:0] tmp_5_reg_1128;
reg [11:0] tmp_8_reg_936;
reg tmp_reg_1061;
reg [1:0] trunc_ln731_reg_828;
reg [1:0] trunc_ln851_1_reg_896;
reg [5:0] _428_;
wire [31:0] _000_;
wire [31:0] _001_;
wire [31:0] _002_;
wire [31:0] _003_;
wire [8:0] _004_;
wire [26:0] _005_;
wire _006_;
wire _007_;
wire _008_;
wire _009_;
wire _010_;
wire _011_;
wire [3:0] _012_;
wire [31:0] _013_;
wire [31:0] _014_;
wire [1:0] _015_;
wire [4:0] _016_;
wire [4:0] _017_;
wire [5:0] _018_;
wire [5:0] _019_;
wire [4:0] _020_;
wire [2:0] _021_;
wire [16:0] _022_;
wire [31:0] _023_;
wire [33:0] _024_;
wire [31:0] _025_;
wire [34:0] _026_;
wire [31:0] _027_;
wire [31:0] _028_;
wire [5:0] _029_;
wire [5:0] _030_;
wire [3:0] _031_;
wire [3:0] _032_;
wire [1:0] _033_;
wire [3:0] _034_;
wire [1:0] _035_;
wire [3:0] _036_;
wire [4:0] _037_;
wire [4:0] _038_;
wire [31:0] _039_;
wire _040_;
wire _041_;
wire [31:0] _042_;
wire [11:0] _043_;
wire _044_;
wire [1:0] _045_;
wire [1:0] _046_;
wire _047_;
wire _048_;
wire _049_;
wire _050_;
wire _051_;
wire _052_;
wire _053_;
wire [8:0] _054_;
wire [8:0] _055_;
wire _056_;
wire [7:0] _057_;
wire [8:0] _058_;
wire [9:0] _059_;
wire [15:0] _060_;
wire [15:0] _061_;
wire _062_;
wire [15:0] _063_;
wire [16:0] _064_;
wire [16:0] _065_;
wire [15:0] _066_;
wire [15:0] _067_;
wire _068_;
wire [15:0] _069_;
wire [16:0] _070_;
wire [16:0] _071_;
wire [15:0] _072_;
wire [15:0] _073_;
wire _074_;
wire [15:0] _075_;
wire [16:0] _076_;
wire [16:0] _077_;
wire [15:0] _078_;
wire [15:0] _079_;
wire _080_;
wire [15:0] _081_;
wire [16:0] _082_;
wire [16:0] _083_;
wire [15:0] _084_;
wire [15:0] _085_;
wire _086_;
wire [15:0] _087_;
wire [16:0] _088_;
wire [16:0] _089_;
wire [15:0] _090_;
wire [15:0] _091_;
wire _092_;
wire [15:0] _093_;
wire [16:0] _094_;
wire [16:0] _095_;
wire [16:0] _096_;
wire [16:0] _097_;
wire _098_;
wire [16:0] _099_;
wire [17:0] _100_;
wire [17:0] _101_;
wire [17:0] _102_;
wire [17:0] _103_;
wire _104_;
wire [16:0] _105_;
wire [17:0] _106_;
wire [18:0] _107_;
wire [17:0] _108_;
wire [17:0] _109_;
wire _110_;
wire [16:0] _111_;
wire [17:0] _112_;
wire [18:0] _113_;
wire [1:0] _114_;
wire [1:0] _115_;
wire _116_;
wire _117_;
wire [1:0] _118_;
wire [2:0] _119_;
wire [1:0] _120_;
wire [1:0] _121_;
wire _122_;
wire [1:0] _123_;
wire [2:0] _124_;
wire [2:0] _125_;
wire [2:0] _126_;
wire [2:0] _127_;
wire _128_;
wire [1:0] _129_;
wire [2:0] _130_;
wire [3:0] _131_;
wire [2:0] _132_;
wire [2:0] _133_;
wire _134_;
wire [1:0] _135_;
wire [2:0] _136_;
wire [3:0] _137_;
wire [2:0] _138_;
wire [2:0] _139_;
wire _140_;
wire [1:0] _141_;
wire [2:0] _142_;
wire [3:0] _143_;
wire [2:0] _144_;
wire [2:0] _145_;
wire _146_;
wire [2:0] _147_;
wire [3:0] _148_;
wire [3:0] _149_;
wire [4:0] _150_;
wire [4:0] _151_;
wire _152_;
wire [3:0] _153_;
wire [4:0] _154_;
wire [5:0] _155_;
wire _156_;
wire _157_;
wire _158_;
wire _159_;
wire _160_;
wire _161_;
wire _162_;
wire _163_;
wire _164_;
wire _165_;
wire _166_;
wire _167_;
wire _168_;
wire _169_;
wire _170_;
wire _171_;
wire _172_;
wire _173_;
wire _174_;
wire _175_;
wire _176_;
wire _177_;
wire _178_;
wire _179_;
wire _180_;
wire _181_;
wire _182_;
wire _183_;
wire _184_;
wire _185_;
wire _186_;
wire \add_17s_17s_17_2_1_U3.ce ;
wire \add_17s_17s_17_2_1_U3.clk ;
wire [16:0] \add_17s_17s_17_2_1_U3.din0 ;
wire [16:0] \add_17s_17s_17_2_1_U3.din1 ;
wire [16:0] \add_17s_17s_17_2_1_U3.dout ;
wire \add_17s_17s_17_2_1_U3.reset ;
wire [16:0] \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.a ;
wire [16:0] \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.ain_s0 ;
wire [16:0] \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.b ;
wire [16:0] \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.bin_s0 ;
wire \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.ce ;
wire \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.clk ;
wire \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.facout_s1 ;
wire \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.facout_s2 ;
wire [7:0] \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.fas_s1 ;
wire [8:0] \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.fas_s2 ;
wire \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.reset ;
wire [16:0] \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.s ;
wire [7:0] \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.u1.a ;
wire [7:0] \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.u1.b ;
wire \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.u1.cin ;
wire \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.u1.cout ;
wire [7:0] \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.u1.s ;
wire [8:0] \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.u2.a ;
wire [8:0] \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.u2.b ;
wire \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.u2.cin ;
wire \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.u2.cout ;
wire [8:0] \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.u2.s ;
wire \add_32ns_32ns_32_2_1_U10.ce ;
wire \add_32ns_32ns_32_2_1_U10.clk ;
wire [31:0] \add_32ns_32ns_32_2_1_U10.din0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U10.din1 ;
wire [31:0] \add_32ns_32ns_32_2_1_U10.dout ;
wire \add_32ns_32ns_32_2_1_U10.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.a ;
wire [31:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.b ;
wire [31:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s0 ;
wire \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.ce ;
wire \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.clk ;
wire \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s1 ;
wire \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s2 ;
wire [15:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s1 ;
wire [15:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s2 ;
wire \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.b ;
wire \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cin ;
wire \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.b ;
wire \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cin ;
wire \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.s ;
wire \add_32ns_32ns_32_2_1_U14.ce ;
wire \add_32ns_32ns_32_2_1_U14.clk ;
wire [31:0] \add_32ns_32ns_32_2_1_U14.din0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U14.din1 ;
wire [31:0] \add_32ns_32ns_32_2_1_U14.dout ;
wire \add_32ns_32ns_32_2_1_U14.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.a ;
wire [31:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.b ;
wire [31:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s0 ;
wire \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.ce ;
wire \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.clk ;
wire \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s1 ;
wire \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s2 ;
wire [15:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s1 ;
wire [15:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s2 ;
wire \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.b ;
wire \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cin ;
wire \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.b ;
wire \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cin ;
wire \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.s ;
wire \add_32ns_32ns_32_2_1_U17.ce ;
wire \add_32ns_32ns_32_2_1_U17.clk ;
wire [31:0] \add_32ns_32ns_32_2_1_U17.din0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U17.din1 ;
wire [31:0] \add_32ns_32ns_32_2_1_U17.dout ;
wire \add_32ns_32ns_32_2_1_U17.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.a ;
wire [31:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.b ;
wire [31:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s0 ;
wire \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.ce ;
wire \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.clk ;
wire \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s1 ;
wire \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s2 ;
wire [15:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s1 ;
wire [15:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s2 ;
wire \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.b ;
wire \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cin ;
wire \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.b ;
wire \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cin ;
wire \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.s ;
wire \add_32ns_32ns_32_2_1_U7.ce ;
wire \add_32ns_32ns_32_2_1_U7.clk ;
wire [31:0] \add_32ns_32ns_32_2_1_U7.din0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U7.din1 ;
wire [31:0] \add_32ns_32ns_32_2_1_U7.dout ;
wire \add_32ns_32ns_32_2_1_U7.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.a ;
wire [31:0] \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.b ;
wire [31:0] \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s0 ;
wire \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.ce ;
wire \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.clk ;
wire \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s1 ;
wire \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s2 ;
wire [15:0] \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s1 ;
wire [15:0] \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s2 ;
wire \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.b ;
wire \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cin ;
wire \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.b ;
wire \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cin ;
wire \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.s ;
wire \add_32s_32ns_32_2_1_U12.ce ;
wire \add_32s_32ns_32_2_1_U12.clk ;
wire [31:0] \add_32s_32ns_32_2_1_U12.din0 ;
wire [31:0] \add_32s_32ns_32_2_1_U12.din1 ;
wire [31:0] \add_32s_32ns_32_2_1_U12.dout ;
wire \add_32s_32ns_32_2_1_U12.reset ;
wire [31:0] \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.a ;
wire [31:0] \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.ain_s0 ;
wire [31:0] \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.b ;
wire [31:0] \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.bin_s0 ;
wire \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.ce ;
wire \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.clk ;
wire \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.facout_s1 ;
wire \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.facout_s2 ;
wire [15:0] \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.fas_s1 ;
wire [15:0] \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.fas_s2 ;
wire \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.reset ;
wire [31:0] \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.s ;
wire [15:0] \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.u1.a ;
wire [15:0] \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.u1.b ;
wire \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.u1.cin ;
wire \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.u1.cout ;
wire [15:0] \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.u1.s ;
wire [15:0] \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.u2.a ;
wire [15:0] \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.u2.b ;
wire \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.u2.cin ;
wire \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.u2.cout ;
wire [15:0] \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.u2.s ;
wire \add_32s_32ns_32_2_1_U4.ce ;
wire \add_32s_32ns_32_2_1_U4.clk ;
wire [31:0] \add_32s_32ns_32_2_1_U4.din0 ;
wire [31:0] \add_32s_32ns_32_2_1_U4.din1 ;
wire [31:0] \add_32s_32ns_32_2_1_U4.dout ;
wire \add_32s_32ns_32_2_1_U4.reset ;
wire [31:0] \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.a ;
wire [31:0] \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.ain_s0 ;
wire [31:0] \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.b ;
wire [31:0] \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.bin_s0 ;
wire \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.ce ;
wire \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.clk ;
wire \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.facout_s1 ;
wire \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.facout_s2 ;
wire [15:0] \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.fas_s1 ;
wire [15:0] \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.fas_s2 ;
wire \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.reset ;
wire [31:0] \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.s ;
wire [15:0] \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.u1.a ;
wire [15:0] \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.u1.b ;
wire \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.u1.cin ;
wire \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.u1.cout ;
wire [15:0] \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.u1.s ;
wire [15:0] \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.u2.a ;
wire [15:0] \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.u2.b ;
wire \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.u2.cin ;
wire \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.u2.cout ;
wire [15:0] \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.u2.s ;
wire \add_34s_34s_34_2_1_U9.ce ;
wire \add_34s_34s_34_2_1_U9.clk ;
wire [33:0] \add_34s_34s_34_2_1_U9.din0 ;
wire [33:0] \add_34s_34s_34_2_1_U9.din1 ;
wire [33:0] \add_34s_34s_34_2_1_U9.dout ;
wire \add_34s_34s_34_2_1_U9.reset ;
wire [33:0] \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.a ;
wire [33:0] \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.ain_s0 ;
wire [33:0] \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.b ;
wire [33:0] \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.bin_s0 ;
wire \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.ce ;
wire \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.clk ;
wire \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.facout_s1 ;
wire \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.facout_s2 ;
wire [16:0] \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.fas_s1 ;
wire [16:0] \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.fas_s2 ;
wire \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.reset ;
wire [33:0] \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.s ;
wire [16:0] \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.u1.a ;
wire [16:0] \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.u1.b ;
wire \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.u1.cin ;
wire \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.u1.cout ;
wire [16:0] \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.u1.s ;
wire [16:0] \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.u2.a ;
wire [16:0] \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.u2.b ;
wire \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.u2.cin ;
wire \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.u2.cout ;
wire [16:0] \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.u2.s ;
wire \add_35ns_35s_35_2_1_U15.ce ;
wire \add_35ns_35s_35_2_1_U15.clk ;
wire [34:0] \add_35ns_35s_35_2_1_U15.din0 ;
wire [34:0] \add_35ns_35s_35_2_1_U15.din1 ;
wire [34:0] \add_35ns_35s_35_2_1_U15.dout ;
wire \add_35ns_35s_35_2_1_U15.reset ;
wire [34:0] \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.a ;
wire [34:0] \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.ain_s0 ;
wire [34:0] \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.b ;
wire [34:0] \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.bin_s0 ;
wire \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.ce ;
wire \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.clk ;
wire \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.facout_s1 ;
wire \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.facout_s2 ;
wire [16:0] \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.fas_s1 ;
wire [17:0] \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.fas_s2 ;
wire \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.reset ;
wire [34:0] \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.s ;
wire [16:0] \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.u1.a ;
wire [16:0] \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.u1.b ;
wire \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.u1.cin ;
wire \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.u1.cout ;
wire [16:0] \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.u1.s ;
wire [17:0] \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.u2.a ;
wire [17:0] \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.u2.b ;
wire \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.u2.cin ;
wire \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.u2.cout ;
wire [17:0] \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.u2.s ;
wire \add_35s_35s_35_2_1_U16.ce ;
wire \add_35s_35s_35_2_1_U16.clk ;
wire [34:0] \add_35s_35s_35_2_1_U16.din0 ;
wire [34:0] \add_35s_35s_35_2_1_U16.din1 ;
wire [34:0] \add_35s_35s_35_2_1_U16.dout ;
wire \add_35s_35s_35_2_1_U16.reset ;
wire [34:0] \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.a ;
wire [34:0] \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.ain_s0 ;
wire [34:0] \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.b ;
wire [34:0] \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.bin_s0 ;
wire \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.ce ;
wire \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.clk ;
wire \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.facout_s1 ;
wire \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.facout_s2 ;
wire [16:0] \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.fas_s1 ;
wire [17:0] \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.fas_s2 ;
wire \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.reset ;
wire [34:0] \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.s ;
wire [16:0] \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.u1.a ;
wire [16:0] \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.u1.b ;
wire \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.u1.cin ;
wire \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.u1.cout ;
wire [16:0] \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.u1.s ;
wire [17:0] \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.u2.a ;
wire [17:0] \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.u2.b ;
wire \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.u2.cin ;
wire \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.u2.cout ;
wire [17:0] \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.u2.s ;
wire \add_3s_3s_3_2_1_U1.ce ;
wire \add_3s_3s_3_2_1_U1.clk ;
wire [2:0] \add_3s_3s_3_2_1_U1.din0 ;
wire [2:0] \add_3s_3s_3_2_1_U1.din1 ;
wire [2:0] \add_3s_3s_3_2_1_U1.dout ;
wire \add_3s_3s_3_2_1_U1.reset ;
wire [2:0] \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.a ;
wire [2:0] \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.ain_s0 ;
wire [2:0] \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.b ;
wire [2:0] \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.bin_s0 ;
wire \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.ce ;
wire \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.clk ;
wire \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.facout_s1 ;
wire \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.facout_s2 ;
wire \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.fas_s1 ;
wire [1:0] \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.fas_s2 ;
wire \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.reset ;
wire [2:0] \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.s ;
wire \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.u1.a ;
wire \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.u1.b ;
wire \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.u1.cin ;
wire \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.u1.cout ;
wire \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.u1.s ;
wire [1:0] \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.u2.a ;
wire [1:0] \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.u2.b ;
wire \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.u2.cin ;
wire \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.u2.cout ;
wire [1:0] \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.u2.s ;
wire \add_4ns_4ns_4_2_1_U8.ce ;
wire \add_4ns_4ns_4_2_1_U8.clk ;
wire [3:0] \add_4ns_4ns_4_2_1_U8.din0 ;
wire [3:0] \add_4ns_4ns_4_2_1_U8.din1 ;
wire [3:0] \add_4ns_4ns_4_2_1_U8.dout ;
wire \add_4ns_4ns_4_2_1_U8.reset ;
wire [3:0] \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.a ;
wire [3:0] \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.ain_s0 ;
wire [3:0] \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.b ;
wire [3:0] \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.bin_s0 ;
wire \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.ce ;
wire \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.clk ;
wire \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.facout_s1 ;
wire \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.facout_s2 ;
wire [1:0] \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.fas_s1 ;
wire [1:0] \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.fas_s2 ;
wire \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.reset ;
wire [3:0] \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.s ;
wire [1:0] \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.u1.a ;
wire [1:0] \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.u1.b ;
wire \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.u1.cin ;
wire \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.u1.cout ;
wire [1:0] \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.u1.s ;
wire [1:0] \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.u2.a ;
wire [1:0] \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.u2.b ;
wire \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.u2.cin ;
wire \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.u2.cout ;
wire [1:0] \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.u2.s ;
wire \add_5ns_5s_5_2_1_U11.ce ;
wire \add_5ns_5s_5_2_1_U11.clk ;
wire [4:0] \add_5ns_5s_5_2_1_U11.din0 ;
wire [4:0] \add_5ns_5s_5_2_1_U11.din1 ;
wire [4:0] \add_5ns_5s_5_2_1_U11.dout ;
wire \add_5ns_5s_5_2_1_U11.reset ;
wire [4:0] \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.a ;
wire [4:0] \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.ain_s0 ;
wire [4:0] \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.b ;
wire [4:0] \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.bin_s0 ;
wire \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.ce ;
wire \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.clk ;
wire \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.facout_s1 ;
wire \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.facout_s2 ;
wire [1:0] \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.fas_s1 ;
wire [2:0] \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.fas_s2 ;
wire \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.reset ;
wire [4:0] \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.s ;
wire [1:0] \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.u1.a ;
wire [1:0] \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.u1.b ;
wire \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.u1.cin ;
wire \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.u1.cout ;
wire [1:0] \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.u1.s ;
wire [2:0] \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.u2.a ;
wire [2:0] \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.u2.b ;
wire \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.u2.cin ;
wire \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.u2.cout ;
wire [2:0] \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.u2.s ;
wire \add_5ns_5s_5_2_1_U6.ce ;
wire \add_5ns_5s_5_2_1_U6.clk ;
wire [4:0] \add_5ns_5s_5_2_1_U6.din0 ;
wire [4:0] \add_5ns_5s_5_2_1_U6.din1 ;
wire [4:0] \add_5ns_5s_5_2_1_U6.dout ;
wire \add_5ns_5s_5_2_1_U6.reset ;
wire [4:0] \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.a ;
wire [4:0] \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.ain_s0 ;
wire [4:0] \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.b ;
wire [4:0] \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.bin_s0 ;
wire \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.ce ;
wire \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.clk ;
wire \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.facout_s1 ;
wire \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.facout_s2 ;
wire [1:0] \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.fas_s1 ;
wire [2:0] \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.fas_s2 ;
wire \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.reset ;
wire [4:0] \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.s ;
wire [1:0] \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.u1.a ;
wire [1:0] \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.u1.b ;
wire \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.u1.cin ;
wire \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.u1.cout ;
wire [1:0] \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.u1.s ;
wire [2:0] \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.u2.a ;
wire [2:0] \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.u2.b ;
wire \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.u2.cin ;
wire \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.u2.cout ;
wire [2:0] \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.u2.s ;
wire \add_5s_5ns_5_2_1_U13.ce ;
wire \add_5s_5ns_5_2_1_U13.clk ;
wire [4:0] \add_5s_5ns_5_2_1_U13.din0 ;
wire [4:0] \add_5s_5ns_5_2_1_U13.din1 ;
wire [4:0] \add_5s_5ns_5_2_1_U13.dout ;
wire \add_5s_5ns_5_2_1_U13.reset ;
wire [4:0] \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.a ;
wire [4:0] \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.ain_s0 ;
wire [4:0] \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.b ;
wire [4:0] \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.bin_s0 ;
wire \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.ce ;
wire \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.clk ;
wire \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.facout_s1 ;
wire \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.facout_s2 ;
wire [1:0] \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.fas_s1 ;
wire [2:0] \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.fas_s2 ;
wire \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.reset ;
wire [4:0] \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.s ;
wire [1:0] \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.u1.a ;
wire [1:0] \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.u1.b ;
wire \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.u1.cin ;
wire \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.u1.cout ;
wire [1:0] \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.u1.s ;
wire [2:0] \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.u2.a ;
wire [2:0] \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.u2.b ;
wire \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.u2.cin ;
wire \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.u2.cout ;
wire [2:0] \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.u2.s ;
wire \add_6ns_6ns_6_2_1_U2.ce ;
wire \add_6ns_6ns_6_2_1_U2.clk ;
wire [5:0] \add_6ns_6ns_6_2_1_U2.din0 ;
wire [5:0] \add_6ns_6ns_6_2_1_U2.din1 ;
wire [5:0] \add_6ns_6ns_6_2_1_U2.dout ;
wire \add_6ns_6ns_6_2_1_U2.reset ;
wire [5:0] \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.a ;
wire [5:0] \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.ain_s0 ;
wire [5:0] \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.b ;
wire [5:0] \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.bin_s0 ;
wire \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.ce ;
wire \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.clk ;
wire \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.facout_s1 ;
wire \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.facout_s2 ;
wire [2:0] \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.fas_s1 ;
wire [2:0] \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.fas_s2 ;
wire \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.reset ;
wire [5:0] \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.s ;
wire [2:0] \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.u1.a ;
wire [2:0] \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.u1.b ;
wire \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.u1.cin ;
wire \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.u1.cout ;
wire [2:0] \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.u1.s ;
wire [2:0] \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.u2.a ;
wire [2:0] \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.u2.b ;
wire \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.u2.cin ;
wire \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.u2.cout ;
wire [2:0] \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.u2.s ;
wire \add_9ns_9ns_9_2_1_U5.ce ;
wire \add_9ns_9ns_9_2_1_U5.clk ;
wire [8:0] \add_9ns_9ns_9_2_1_U5.din0 ;
wire [8:0] \add_9ns_9ns_9_2_1_U5.din1 ;
wire [8:0] \add_9ns_9ns_9_2_1_U5.dout ;
wire \add_9ns_9ns_9_2_1_U5.reset ;
wire [8:0] \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.a ;
wire [8:0] \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.ain_s0 ;
wire [8:0] \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.b ;
wire [8:0] \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.bin_s0 ;
wire \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.ce ;
wire \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.clk ;
wire \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.facout_s1 ;
wire \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.facout_s2 ;
wire [3:0] \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.fas_s1 ;
wire [4:0] \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.fas_s2 ;
wire \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.reset ;
wire [8:0] \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.s ;
wire [3:0] \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.u1.a ;
wire [3:0] \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.u1.b ;
wire \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.u1.cin ;
wire \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.u1.cout ;
wire [3:0] \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.u1.s ;
wire [4:0] \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.u2.a ;
wire [4:0] \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.u2.b ;
wire \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.u2.cin ;
wire \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.u2.cout ;
wire [4:0] \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.u2.s ;
wire and_ln340_1_fu_296_p2;
wire and_ln340_fu_301_p2;
wire and_ln785_fu_318_p2;
wire [3:0] and_ln_fu_255_p3;
wire ap_CS_fsm_state1;
wire ap_CS_fsm_state10;
wire ap_CS_fsm_state11;
wire ap_CS_fsm_state12;
wire ap_CS_fsm_state13;
wire ap_CS_fsm_state14;
wire ap_CS_fsm_state15;
wire ap_CS_fsm_state16;
wire ap_CS_fsm_state17;
wire ap_CS_fsm_state18;
wire ap_CS_fsm_state19;
wire ap_CS_fsm_state2;
wire ap_CS_fsm_state20;
wire ap_CS_fsm_state21;
wire ap_CS_fsm_state22;
wire ap_CS_fsm_state23;
wire ap_CS_fsm_state24;
wire ap_CS_fsm_state25;
wire ap_CS_fsm_state26;
wire ap_CS_fsm_state27;
wire ap_CS_fsm_state3;
wire ap_CS_fsm_state4;
wire ap_CS_fsm_state5;
wire ap_CS_fsm_state6;
wire ap_CS_fsm_state7;
wire ap_CS_fsm_state8;
wire ap_CS_fsm_state9;
wire [26:0] ap_NS_fsm;
wire ap_clk;
wire ap_done;
wire ap_idle;
wire ap_ready;
wire ap_rst;
wire ap_start;
wire [2:0] grp_fu_341_p0;
wire [2:0] grp_fu_341_p1;
wire [2:0] grp_fu_341_p2;
wire [5:0] grp_fu_384_p2;
wire [16:0] grp_fu_404_p0;
wire [16:0] grp_fu_404_p1;
wire [16:0] grp_fu_404_p2;
wire [31:0] grp_fu_452_p0;
wire [31:0] grp_fu_452_p2;
wire [8:0] grp_fu_469_p0;
wire [8:0] grp_fu_469_p1;
wire [8:0] grp_fu_469_p2;
wire [4:0] grp_fu_506_p1;
wire [4:0] grp_fu_506_p2;
wire [31:0] grp_fu_514_p0;
wire [31:0] grp_fu_514_p2;
wire [3:0] grp_fu_529_p2;
wire [33:0] grp_fu_549_p0;
wire [33:0] grp_fu_549_p1;
wire [33:0] grp_fu_549_p2;
wire [31:0] grp_fu_588_p2;
wire [4:0] grp_fu_620_p0;
wire [4:0] grp_fu_620_p2;
wire [31:0] grp_fu_629_p0;
wire [31:0] grp_fu_629_p2;
wire [4:0] grp_fu_708_p0;
wire [4:0] grp_fu_708_p2;
wire [31:0] grp_fu_713_p2;
wire [34:0] grp_fu_735_p0;
wire [34:0] grp_fu_735_p1;
wire [34:0] grp_fu_735_p2;
wire [34:0] grp_fu_766_p0;
wire [34:0] grp_fu_766_p1;
wire [34:0] grp_fu_766_p2;
wire [31:0] grp_fu_792_p2;
wire icmp_ln785_fu_270_p2;
wire icmp_ln786_1_fu_282_p2;
wire icmp_ln786_fu_276_p2;
wire icmp_ln851_1_fu_414_p2;
wire icmp_ln851_2_fu_776_p2;
wire icmp_ln851_fu_379_p2;
wire [5:0] lhs_fu_347_p3;
wire op_0;
wire [1:0] op_10;
wire [15:0] op_11;
wire [1:0] op_13;
wire [3:0] op_15;
wire [31:0] op_16;
wire [3:0] op_17;
wire [7:0] op_18_V_fu_717_p3;
wire [3:0] op_19;
wire [31:0] op_29;
wire op_29_ap_vld;
wire [3:0] op_3;
wire [3:0] op_4;
wire [3:0] op_5;
wire [7:0] op_9;
wire or_ln785_fu_322_p2;
wire or_ln786_1_fu_314_p2;
wire or_ln786_fu_287_p2;
wire [3:0] or_ln_fu_262_p4;
wire p_Result_1_fu_430_p3;
wire p_Result_2_fu_565_p3;
wire p_Result_3_fu_483_p3;
wire p_Result_4_fu_682_p3;
wire p_Result_5_fu_797_p3;
wire p_Result_s_fu_635_p3;
wire [3:0] r_fu_219_p2;
wire [4:0] ret_V_21_fu_600_p2;
wire ret_V_22_fu_657_p3;
wire [7:0] ret_V_23_fu_359_p2;
wire [7:0] ret_V_23_reg_884;
wire [5:0] ret_V_24_fu_442_p3;
wire [31:0] ret_V_29_fu_495_p3;
wire [31:0] ret_V_31_fu_698_p3;
wire [1:0] ret_V_9_fu_328_p3;
wire ret_V_fu_645_p2;
wire [32:0] rhs_5_fu_538_p3;
wire [33:0] rhs_8_fu_755_p3;
wire [4:0] rhs_fu_593_p3;
wire [4:0] select_ln1192_fu_475_p3;
wire [1:0] select_ln340_fu_307_p3;
wire [3:0] select_ln353_fu_581_p3;
wire [4:0] select_ln703_fu_674_p3;
wire [5:0] select_ln850_1_fu_437_p3;
wire [3:0] select_ln850_3_fu_575_p3;
wire [31:0] select_ln850_4_fu_490_p3;
wire [31:0] select_ln850_5_fu_692_p3;
wire [31:0] select_ln850_6_fu_804_p3;
wire select_ln850_fu_650_p3;
wire [15:0] sext_ln1192_1_fu_389_p0;
wire [7:0] sext_ln1194_fu_355_p1;
wire [7:0] sext_ln69_1_fu_458_p1;
wire [3:0] sext_ln703_2_fu_534_p0;
wire [3:0] sext_ln703_3_fu_751_p0;
wire [4:0] sext_ln703_fu_502_p1;
wire [31:0] sext_ln831_fu_449_p1;
wire [7:0] tmp_4_fu_393_p3;
wire [1:0] trunc_ln731_fu_233_p1;
wire [1:0] trunc_ln851_1_fu_375_p1;
wire trunc_ln851_2_fu_572_p1;
wire [15:0] trunc_ln851_3_fu_410_p0;
wire [4:0] trunc_ln851_3_fu_410_p1;
wire [3:0] trunc_ln851_4_fu_689_p0;
wire trunc_ln851_4_fu_689_p1;
wire [3:0] trunc_ln851_5_fu_772_p0;
wire [1:0] trunc_ln851_5_fu_772_p1;
wire trunc_ln851_fu_642_p1;
wire xor_ln340_1_fu_291_p2;


assign _047_ = icmp_ln851_2_reg_1143 & ap_CS_fsm[25];
assign _048_ = ap_CS_fsm[9] & icmp_ln851_1_reg_921;
assign _049_ = _051_ & ap_CS_fsm[0];
assign _050_ = ap_start & ap_CS_fsm[0];
assign and_ln340_1_fu_296_p2 = xor_ln340_1_fu_291_p2 & tmp_2_reg_822;
assign and_ln340_fu_301_p2 = or_ln786_1_fu_314_p2 & and_ln340_1_fu_296_p2;
assign and_ln785_fu_318_p2 = tmp_2_reg_822 & icmp_ln785_reg_846;
assign ret_V_23_fu_359_p2 = { op_5[3], op_5[3], op_5, 2'h0 } & op_9;
assign xor_ln340_1_fu_291_p2 = ~ icmp_ln785_reg_846;
assign ret_V_fu_645_p2 = ~ tmp_reg_1061;
assign r_fu_219_p2 = ~ op_4;
assign _051_ = ~ ap_start;
assign _052_ = ! { tmp_3_reg_834, 3'h0 };
assign _053_ = ! trunc_ln851_1_reg_896;
always @(posedge \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.clk )
\add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.bin_s1  <= _055_;
always @(posedge \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.clk )
\add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.ain_s1  <= _054_;
always @(posedge \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.clk )
\add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.sum_s1  <= _057_;
always @(posedge \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.clk )
\add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.carry_s1  <= _056_;
assign _055_ = \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.ce  ? \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.b [16:8] : \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.bin_s1 ;
assign _054_ = \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.ce  ? \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.a [16:8] : \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.ain_s1 ;
assign _056_ = \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.ce  ? \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.facout_s1  : \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.carry_s1 ;
assign _057_ = \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.ce  ? \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.fas_s1  : \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.sum_s1 ;
assign _058_ = \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.u1.a  + \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.u1.b ;
assign { \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.u1.cout , \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.u1.s  } = _058_ + \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.u1.cin ;
assign _059_ = \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.u2.a  + \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.u2.b ;
assign { \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.u2.cout , \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.u2.s  } = _059_ + \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.u2.cin ;
always @(posedge \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.clk )
\add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s1  <= _061_;
always @(posedge \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.clk )
\add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s1  <= _060_;
always @(posedge \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.clk )
\add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.sum_s1  <= _063_;
always @(posedge \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.clk )
\add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.carry_s1  <= _062_;
assign _061_ = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  ? \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.b [31:16] : \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s1 ;
assign _060_ = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  ? \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.a [31:16] : \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s1 ;
assign _062_ = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  ? \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s1  : \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.carry_s1 ;
assign _063_ = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  ? \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s1  : \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.sum_s1 ;
assign _064_ = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.a  + \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.b ;
assign { \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cout , \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.s  } = _064_ + \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cin ;
assign _065_ = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.a  + \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.b ;
assign { \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cout , \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.s  } = _065_ + \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cin ;
always @(posedge \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.clk )
\add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s1  <= _067_;
always @(posedge \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.clk )
\add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s1  <= _066_;
always @(posedge \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.clk )
\add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.sum_s1  <= _069_;
always @(posedge \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.clk )
\add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.carry_s1  <= _068_;
assign _067_ = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  ? \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.b [31:16] : \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s1 ;
assign _066_ = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  ? \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.a [31:16] : \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s1 ;
assign _068_ = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  ? \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s1  : \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.carry_s1 ;
assign _069_ = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  ? \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s1  : \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.sum_s1 ;
assign _070_ = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.a  + \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.b ;
assign { \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cout , \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.s  } = _070_ + \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cin ;
assign _071_ = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.a  + \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.b ;
assign { \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cout , \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.s  } = _071_ + \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cin ;
always @(posedge \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.clk )
\add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s1  <= _073_;
always @(posedge \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.clk )
\add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s1  <= _072_;
always @(posedge \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.clk )
\add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.sum_s1  <= _075_;
always @(posedge \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.clk )
\add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.carry_s1  <= _074_;
assign _073_ = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  ? \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.b [31:16] : \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s1 ;
assign _072_ = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  ? \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.a [31:16] : \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s1 ;
assign _074_ = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  ? \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s1  : \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.carry_s1 ;
assign _075_ = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  ? \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s1  : \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.sum_s1 ;
assign _076_ = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.a  + \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.b ;
assign { \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cout , \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.s  } = _076_ + \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cin ;
assign _077_ = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.a  + \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.b ;
assign { \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cout , \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.s  } = _077_ + \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cin ;
always @(posedge \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.clk )
\add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s1  <= _079_;
always @(posedge \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.clk )
\add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s1  <= _078_;
always @(posedge \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.clk )
\add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.sum_s1  <= _081_;
always @(posedge \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.clk )
\add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.carry_s1  <= _080_;
assign _079_ = \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  ? \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.b [31:16] : \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s1 ;
assign _078_ = \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  ? \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.a [31:16] : \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s1 ;
assign _080_ = \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  ? \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s1  : \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.carry_s1 ;
assign _081_ = \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  ? \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s1  : \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.sum_s1 ;
assign _082_ = \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.a  + \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.b ;
assign { \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cout , \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.s  } = _082_ + \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cin ;
assign _083_ = \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.a  + \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.b ;
assign { \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cout , \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.s  } = _083_ + \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cin ;
always @(posedge \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.clk )
\add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.bin_s1  <= _085_;
always @(posedge \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.clk )
\add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.ain_s1  <= _084_;
always @(posedge \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.clk )
\add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.sum_s1  <= _087_;
always @(posedge \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.clk )
\add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.carry_s1  <= _086_;
assign _085_ = \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.ce  ? \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.b [31:16] : \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.bin_s1 ;
assign _084_ = \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.ce  ? \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.a [31:16] : \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.ain_s1 ;
assign _086_ = \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.ce  ? \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.facout_s1  : \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.carry_s1 ;
assign _087_ = \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.ce  ? \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.fas_s1  : \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.sum_s1 ;
assign _088_ = \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.u1.a  + \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.u1.b ;
assign { \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.u1.cout , \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.u1.s  } = _088_ + \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.u1.cin ;
assign _089_ = \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.u2.a  + \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.u2.b ;
assign { \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.u2.cout , \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.u2.s  } = _089_ + \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.u2.cin ;
always @(posedge \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.clk )
\add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.bin_s1  <= _091_;
always @(posedge \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.clk )
\add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.ain_s1  <= _090_;
always @(posedge \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.clk )
\add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.sum_s1  <= _093_;
always @(posedge \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.clk )
\add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.carry_s1  <= _092_;
assign _091_ = \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.ce  ? \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.b [31:16] : \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.bin_s1 ;
assign _090_ = \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.ce  ? \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.a [31:16] : \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.ain_s1 ;
assign _092_ = \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.ce  ? \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.facout_s1  : \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.carry_s1 ;
assign _093_ = \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.ce  ? \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.fas_s1  : \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.sum_s1 ;
assign _094_ = \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.u1.a  + \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.u1.b ;
assign { \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.u1.cout , \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.u1.s  } = _094_ + \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.u1.cin ;
assign _095_ = \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.u2.a  + \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.u2.b ;
assign { \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.u2.cout , \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.u2.s  } = _095_ + \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.u2.cin ;
always @(posedge \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.clk )
\add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.bin_s1  <= _097_;
always @(posedge \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.clk )
\add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.ain_s1  <= _096_;
always @(posedge \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.clk )
\add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.sum_s1  <= _099_;
always @(posedge \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.clk )
\add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.carry_s1  <= _098_;
assign _097_ = \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.ce  ? \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.b [33:17] : \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.bin_s1 ;
assign _096_ = \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.ce  ? \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.a [33:17] : \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.ain_s1 ;
assign _098_ = \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.ce  ? \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.facout_s1  : \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.carry_s1 ;
assign _099_ = \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.ce  ? \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.fas_s1  : \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.sum_s1 ;
assign _100_ = \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.u1.a  + \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.u1.b ;
assign { \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.u1.cout , \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.u1.s  } = _100_ + \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.u1.cin ;
assign _101_ = \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.u2.a  + \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.u2.b ;
assign { \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.u2.cout , \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.u2.s  } = _101_ + \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.u2.cin ;
always @(posedge \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.clk )
\add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.bin_s1  <= _103_;
always @(posedge \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.clk )
\add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.ain_s1  <= _102_;
always @(posedge \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.clk )
\add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.sum_s1  <= _105_;
always @(posedge \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.clk )
\add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.carry_s1  <= _104_;
assign _103_ = \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.ce  ? \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.b [34:17] : \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.bin_s1 ;
assign _102_ = \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.ce  ? \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.a [34:17] : \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.ain_s1 ;
assign _104_ = \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.ce  ? \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.facout_s1  : \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.carry_s1 ;
assign _105_ = \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.ce  ? \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.fas_s1  : \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.sum_s1 ;
assign _106_ = \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.u1.a  + \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.u1.b ;
assign { \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.u1.cout , \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.u1.s  } = _106_ + \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.u1.cin ;
assign _107_ = \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.u2.a  + \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.u2.b ;
assign { \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.u2.cout , \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.u2.s  } = _107_ + \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.u2.cin ;
always @(posedge \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.clk )
\add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.bin_s1  <= _109_;
always @(posedge \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.clk )
\add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.ain_s1  <= _108_;
always @(posedge \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.clk )
\add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.sum_s1  <= _111_;
always @(posedge \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.clk )
\add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.carry_s1  <= _110_;
assign _109_ = \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.ce  ? \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.b [34:17] : \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.bin_s1 ;
assign _108_ = \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.ce  ? \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.a [34:17] : \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.ain_s1 ;
assign _110_ = \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.ce  ? \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.facout_s1  : \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.carry_s1 ;
assign _111_ = \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.ce  ? \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.fas_s1  : \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.sum_s1 ;
assign _112_ = \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.u1.a  + \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.u1.b ;
assign { \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.u1.cout , \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.u1.s  } = _112_ + \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.u1.cin ;
assign _113_ = \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.u2.a  + \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.u2.b ;
assign { \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.u2.cout , \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.u2.s  } = _113_ + \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.u2.cin ;
always @(posedge \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.clk )
\add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.bin_s1  <= _115_;
always @(posedge \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.clk )
\add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.ain_s1  <= _114_;
always @(posedge \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.clk )
\add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.sum_s1  <= _117_;
always @(posedge \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.clk )
\add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.carry_s1  <= _116_;
assign _115_ = \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.ce  ? \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.b [2:1] : \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.bin_s1 ;
assign _114_ = \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.ce  ? \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.a [2:1] : \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.ain_s1 ;
assign _116_ = \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.ce  ? \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.facout_s1  : \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.carry_s1 ;
assign _117_ = \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.ce  ? \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.fas_s1  : \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.sum_s1 ;
assign _118_ = \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.u1.a  + \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.u1.b ;
assign { \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.u1.cout , \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.u1.s  } = _118_ + \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.u1.cin ;
assign _119_ = \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.u2.a  + \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.u2.b ;
assign { \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.u2.cout , \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.u2.s  } = _119_ + \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.u2.cin ;
always @(posedge \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.clk )
\add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.bin_s1  <= _121_;
always @(posedge \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.clk )
\add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.ain_s1  <= _120_;
always @(posedge \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.clk )
\add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.sum_s1  <= _123_;
always @(posedge \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.clk )
\add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.carry_s1  <= _122_;
assign _121_ = \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.ce  ? \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.b [3:2] : \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.bin_s1 ;
assign _120_ = \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.ce  ? \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.a [3:2] : \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.ain_s1 ;
assign _122_ = \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.ce  ? \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.facout_s1  : \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.carry_s1 ;
assign _123_ = \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.ce  ? \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.fas_s1  : \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.sum_s1 ;
assign _124_ = \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.u1.a  + \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.u1.b ;
assign { \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.u1.cout , \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.u1.s  } = _124_ + \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.u1.cin ;
assign _125_ = \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.u2.a  + \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.u2.b ;
assign { \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.u2.cout , \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.u2.s  } = _125_ + \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.u2.cin ;
always @(posedge \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.clk )
\add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.bin_s1  <= _127_;
always @(posedge \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.clk )
\add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.ain_s1  <= _126_;
always @(posedge \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.clk )
\add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.sum_s1  <= _129_;
always @(posedge \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.clk )
\add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.carry_s1  <= _128_;
assign _127_ = \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.ce  ? \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.b [4:2] : \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.bin_s1 ;
assign _126_ = \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.ce  ? \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.a [4:2] : \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.ain_s1 ;
assign _128_ = \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.ce  ? \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.facout_s1  : \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.carry_s1 ;
assign _129_ = \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.ce  ? \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.fas_s1  : \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.sum_s1 ;
assign _130_ = \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.u1.a  + \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.u1.b ;
assign { \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.u1.cout , \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.u1.s  } = _130_ + \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.u1.cin ;
assign _131_ = \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.u2.a  + \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.u2.b ;
assign { \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.u2.cout , \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.u2.s  } = _131_ + \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.u2.cin ;
always @(posedge \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.clk )
\add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.bin_s1  <= _133_;
always @(posedge \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.clk )
\add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.ain_s1  <= _132_;
always @(posedge \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.clk )
\add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.sum_s1  <= _135_;
always @(posedge \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.clk )
\add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.carry_s1  <= _134_;
assign _133_ = \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.ce  ? \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.b [4:2] : \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.bin_s1 ;
assign _132_ = \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.ce  ? \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.a [4:2] : \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.ain_s1 ;
assign _134_ = \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.ce  ? \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.facout_s1  : \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.carry_s1 ;
assign _135_ = \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.ce  ? \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.fas_s1  : \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.sum_s1 ;
assign _136_ = \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.u1.a  + \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.u1.b ;
assign { \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.u1.cout , \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.u1.s  } = _136_ + \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.u1.cin ;
assign _137_ = \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.u2.a  + \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.u2.b ;
assign { \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.u2.cout , \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.u2.s  } = _137_ + \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.u2.cin ;
always @(posedge \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.clk )
\add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.bin_s1  <= _139_;
always @(posedge \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.clk )
\add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.ain_s1  <= _138_;
always @(posedge \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.clk )
\add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.sum_s1  <= _141_;
always @(posedge \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.clk )
\add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.carry_s1  <= _140_;
assign _139_ = \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.ce  ? \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.b [4:2] : \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.bin_s1 ;
assign _138_ = \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.ce  ? \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.a [4:2] : \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.ain_s1 ;
assign _140_ = \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.ce  ? \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.facout_s1  : \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.carry_s1 ;
assign _141_ = \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.ce  ? \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.fas_s1  : \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.sum_s1 ;
assign _142_ = \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.u1.a  + \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.u1.b ;
assign { \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.u1.cout , \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.u1.s  } = _142_ + \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.u1.cin ;
assign _143_ = \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.u2.a  + \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.u2.b ;
assign { \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.u2.cout , \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.u2.s  } = _143_ + \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.u2.cin ;
always @(posedge \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.clk )
\add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.bin_s1  <= _145_;
always @(posedge \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.clk )
\add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.ain_s1  <= _144_;
always @(posedge \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.clk )
\add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.sum_s1  <= _147_;
always @(posedge \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.clk )
\add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.carry_s1  <= _146_;
assign _145_ = \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.ce  ? \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.b [5:3] : \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.bin_s1 ;
assign _144_ = \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.ce  ? \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.a [5:3] : \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.ain_s1 ;
assign _146_ = \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.ce  ? \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.facout_s1  : \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.carry_s1 ;
assign _147_ = \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.ce  ? \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.fas_s1  : \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.sum_s1 ;
assign _148_ = \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.u1.a  + \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.u1.b ;
assign { \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.u1.cout , \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.u1.s  } = _148_ + \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.u1.cin ;
assign _149_ = \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.u2.a  + \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.u2.b ;
assign { \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.u2.cout , \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.u2.s  } = _149_ + \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.u2.cin ;
always @(posedge \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.clk )
\add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.bin_s1  <= _151_;
always @(posedge \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.clk )
\add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.ain_s1  <= _150_;
always @(posedge \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.clk )
\add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.sum_s1  <= _153_;
always @(posedge \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.clk )
\add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.carry_s1  <= _152_;
assign _151_ = \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.ce  ? \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.b [8:4] : \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.bin_s1 ;
assign _150_ = \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.ce  ? \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.a [8:4] : \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.ain_s1 ;
assign _152_ = \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.ce  ? \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.facout_s1  : \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.carry_s1 ;
assign _153_ = \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.ce  ? \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.fas_s1  : \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.sum_s1 ;
assign _154_ = \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.u1.a  + \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.u1.b ;
assign { \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.u1.cout , \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.u1.s  } = _154_ + \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.u1.cin ;
assign _155_ = \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.u2.a  + \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.u2.b ;
assign { \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.u2.cout , \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.u2.s  } = _155_ + \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.u2.cin ;
assign _156_ = | { tmp_3_reg_834, 1'h0, p_Result_s_16_reg_840 };
assign _157_ = p_Result_s_16_reg_840 != 2'h3;
assign _158_ = | op_11[4:0];
assign _159_ = | op_19[1:0];
assign or_ln785_fu_322_p2 = or_ln786_1_fu_314_p2 | and_ln785_fu_318_p2;
assign or_ln786_1_fu_314_p2 = icmp_ln786_reg_852 | icmp_ln786_1_reg_858;
always @(posedge ap_clk)
trunc_ln851_1_reg_896 <= 2'h0;
always @(posedge ap_clk)
select_ln1192_reg_968[0] <= 1'h0;
always @(posedge ap_clk)
tmp_5_reg_1128 <= _042_;
always @(posedge ap_clk)
sext_ln703_reg_983 <= _038_;
always @(posedge ap_clk)
select_ln353_reg_1045 <= _036_;
always @(posedge ap_clk)
select_ln340_reg_864 <= _035_;
always @(posedge ap_clk)
ret_V_9_reg_869 <= _033_;
always @(posedge ap_clk)
ret_V_32_reg_1148 <= _026_;
always @(posedge ap_clk)
ret_V_36_cast_reg_1153 <= _028_;
always @(posedge ap_clk)
ret_V_8_reg_1028 <= _032_;
always @(posedge ap_clk)
ret_V_30_reg_1033 <= _024_;
always @(posedge ap_clk)
ret_V_33_cast_reg_1038 <= _027_;
always @(posedge ap_clk)
ret_V_5_reg_926 <= _030_;
always @(posedge ap_clk)
ret_V_28_reg_931 <= _022_;
always @(posedge ap_clk)
tmp_8_reg_936 <= _043_;
always @(posedge ap_clk)
ret_V_24_reg_941 <= _019_;
always @(posedge ap_clk)
sext_ln831_reg_946 <= _039_;
always @(posedge ap_clk)
_428_ <= _018_;
assign ret_V_23_reg_884[7:2] = _428_;
always @(posedge ap_clk)
ret_V_3_reg_889 <= _029_;
always @(posedge ap_clk)
ret_V_27_reg_901 <= _021_;
always @(posedge ap_clk)
tmp_2_reg_822 <= _040_;
always @(posedge ap_clk)
trunc_ln731_reg_828 <= _045_;
always @(posedge ap_clk)
tmp_3_reg_834 <= _041_;
always @(posedge ap_clk)
p_Result_s_16_reg_840 <= _015_;
always @(posedge ap_clk)
ret_V_13_reg_1108 <= _016_;
always @(posedge ap_clk)
op_27_V_reg_1113 <= _014_;
always @(posedge ap_clk)
ret_V_25_reg_995 <= _020_;
always @(posedge ap_clk)
ret_V_8_cast_reg_1001 <= _031_;
always @(posedge ap_clk)
op_24_V_reg_1008 <= _013_;
always @(posedge ap_clk)
icmp_ln851_2_reg_1143 <= _010_;
always @(posedge ap_clk)
icmp_ln851_reg_906 <= _011_;
always @(posedge ap_clk)
icmp_ln851_1_reg_921 <= _009_;
always @(posedge ap_clk)
icmp_ln785_reg_846 <= _006_;
always @(posedge ap_clk)
icmp_ln786_reg_852 <= _008_;
always @(posedge ap_clk)
icmp_ln786_1_reg_858 <= _007_;
always @(posedge ap_clk)
select_ln1192_reg_968[4:1] <= _034_;
always @(posedge ap_clk)
ret_V_29_reg_973 <= _023_;
always @(posedge ap_clk)
add_ln69_reg_978 <= _004_;
always @(posedge ap_clk)
op_14_V_reg_1083 <= _012_;
always @(posedge ap_clk)
select_ln703_reg_1088 <= _037_;
always @(posedge ap_clk)
ret_V_31_reg_1093 <= _025_;
always @(posedge ap_clk)
add_ln69_2_reg_1098 <= _003_;
always @(posedge ap_clk)
add_ln691_reg_953 <= _002_;
always @(posedge ap_clk)
add_ln691_2_reg_1160 <= _001_;
always @(posedge ap_clk)
ret_V_21_reg_1055 <= _017_;
always @(posedge ap_clk)
tmp_reg_1061 <= _044_;
always @(posedge ap_clk)
add_ln691_1_reg_1073 <= _000_;
always @(posedge ap_clk)
ap_CS_fsm <= _005_;
assign _046_ = _050_ ? 2'h2 : 2'h1;
assign _160_ = ap_CS_fsm == 1'h1;
function [26:0] _461_;
input [26:0] a;
input [728:0] b;
input [26:0] s;
case (s)
27'b000000000000000000000000001:
_461_ = b[26:0];
27'b000000000000000000000000010:
_461_ = b[53:27];
27'b000000000000000000000000100:
_461_ = b[80:54];
27'b000000000000000000000001000:
_461_ = b[107:81];
27'b000000000000000000000010000:
_461_ = b[134:108];
27'b000000000000000000000100000:
_461_ = b[161:135];
27'b000000000000000000001000000:
_461_ = b[188:162];
27'b000000000000000000010000000:
_461_ = b[215:189];
27'b000000000000000000100000000:
_461_ = b[242:216];
27'b000000000000000001000000000:
_461_ = b[269:243];
27'b000000000000000010000000000:
_461_ = b[296:270];
27'b000000000000000100000000000:
_461_ = b[323:297];
27'b000000000000001000000000000:
_461_ = b[350:324];
27'b000000000000010000000000000:
_461_ = b[377:351];
27'b000000000000100000000000000:
_461_ = b[404:378];
27'b000000000001000000000000000:
_461_ = b[431:405];
27'b000000000010000000000000000:
_461_ = b[458:432];
27'b000000000100000000000000000:
_461_ = b[485:459];
27'b000000001000000000000000000:
_461_ = b[512:486];
27'b000000010000000000000000000:
_461_ = b[539:513];
27'b000000100000000000000000000:
_461_ = b[566:540];
27'b000001000000000000000000000:
_461_ = b[593:567];
27'b000010000000000000000000000:
_461_ = b[620:594];
27'b000100000000000000000000000:
_461_ = b[647:621];
27'b001000000000000000000000000:
_461_ = b[674:648];
27'b010000000000000000000000000:
_461_ = b[701:675];
27'b100000000000000000000000000:
_461_ = b[728:702];
27'b000000000000000000000000000:
_461_ = a;
default:
_461_ = 27'bx;
endcase
endfunction
assign ap_NS_fsm = _461_(27'hxxxxxxx, { 25'h0000000, _046_, 702'h00000020000008000002000000800000200000080000020000008000002000000800000200000080000020000008000002000000800000200000080000020000008000002000000800000200000080000020000000000001 }, { _160_, _186_, _185_, _184_, _183_, _182_, _181_, _180_, _179_, _178_, _177_, _176_, _175_, _174_, _173_, _172_, _171_, _170_, _169_, _168_, _167_, _166_, _165_, _164_, _163_, _162_, _161_ });
assign _161_ = ap_CS_fsm == 27'h4000000;
assign _162_ = ap_CS_fsm == 26'h2000000;
assign _163_ = ap_CS_fsm == 25'h1000000;
assign _164_ = ap_CS_fsm == 24'h800000;
assign _165_ = ap_CS_fsm == 23'h400000;
assign _166_ = ap_CS_fsm == 22'h200000;
assign _167_ = ap_CS_fsm == 21'h100000;
assign _168_ = ap_CS_fsm == 20'h80000;
assign _169_ = ap_CS_fsm == 19'h40000;
assign _170_ = ap_CS_fsm == 18'h20000;
assign _171_ = ap_CS_fsm == 17'h10000;
assign _172_ = ap_CS_fsm == 16'h8000;
assign _173_ = ap_CS_fsm == 15'h4000;
assign _174_ = ap_CS_fsm == 14'h2000;
assign _175_ = ap_CS_fsm == 13'h1000;
assign _176_ = ap_CS_fsm == 12'h800;
assign _177_ = ap_CS_fsm == 11'h400;
assign _178_ = ap_CS_fsm == 10'h200;
assign _179_ = ap_CS_fsm == 9'h100;
assign _180_ = ap_CS_fsm == 8'h80;
assign _181_ = ap_CS_fsm == 7'h40;
assign _182_ = ap_CS_fsm == 6'h20;
assign _183_ = ap_CS_fsm == 5'h10;
assign _184_ = ap_CS_fsm == 4'h8;
assign _185_ = ap_CS_fsm == 3'h4;
assign _186_ = ap_CS_fsm == 2'h2;
assign op_29_ap_vld = ap_CS_fsm[26] ? 1'h1 : 1'h0;
assign ap_idle = _049_ ? 1'h1 : 1'h0;
assign _042_ = ap_CS_fsm[21] ? grp_fu_735_p2[34:3] : tmp_5_reg_1128;
assign _038_ = ap_CS_fsm[11] ? { op_3[3], op_3 } : sext_ln703_reg_983;
assign _036_ = ap_CS_fsm[15] ? select_ln353_fu_581_p3 : select_ln353_reg_1045;
assign _035_ = ap_CS_fsm[2] ? select_ln340_fu_307_p3 : select_ln340_reg_864;
assign _033_ = ap_CS_fsm[3] ? ret_V_9_fu_328_p3 : ret_V_9_reg_869;
assign _028_ = ap_CS_fsm[23] ? grp_fu_766_p2[33:2] : ret_V_36_cast_reg_1153;
assign _026_ = ap_CS_fsm[23] ? grp_fu_766_p2 : ret_V_32_reg_1148;
assign _027_ = ap_CS_fsm[14] ? grp_fu_549_p2[32:1] : ret_V_33_cast_reg_1038;
assign _024_ = ap_CS_fsm[14] ? grp_fu_549_p2 : ret_V_30_reg_1033;
assign _032_ = ap_CS_fsm[14] ? grp_fu_529_p2 : ret_V_8_reg_1028;
assign _043_ = ap_CS_fsm[7] ? grp_fu_404_p2[16:5] : tmp_8_reg_936;
assign _022_ = ap_CS_fsm[7] ? grp_fu_404_p2 : ret_V_28_reg_931;
assign _030_ = ap_CS_fsm[7] ? grp_fu_384_p2 : ret_V_5_reg_926;
assign _039_ = ap_CS_fsm[8] ? { tmp_8_reg_936[11], tmp_8_reg_936[11], tmp_8_reg_936[11], tmp_8_reg_936[11], tmp_8_reg_936[11], tmp_8_reg_936[11], tmp_8_reg_936[11], tmp_8_reg_936[11], tmp_8_reg_936[11], tmp_8_reg_936[11], tmp_8_reg_936[11], tmp_8_reg_936[11], tmp_8_reg_936[11], tmp_8_reg_936[11], tmp_8_reg_936[11], tmp_8_reg_936[11], tmp_8_reg_936[11], tmp_8_reg_936[11], tmp_8_reg_936[11], tmp_8_reg_936[11], tmp_8_reg_936 } : sext_ln831_reg_946;
assign _019_ = ap_CS_fsm[8] ? ret_V_24_fu_442_p3 : ret_V_24_reg_941;
assign _021_ = ap_CS_fsm[5] ? grp_fu_341_p2 : ret_V_27_reg_901;
assign _029_ = ap_CS_fsm[5] ? ret_V_23_fu_359_p2[7:2] : ret_V_3_reg_889;
assign _018_ = ap_CS_fsm[5] ? ret_V_23_fu_359_p2[7:2] : ret_V_23_reg_884[7:2];
assign _015_ = ap_CS_fsm[0] ? r_fu_219_p2[3:2] : p_Result_s_16_reg_840;
assign _041_ = ap_CS_fsm[0] ? r_fu_219_p2[1] : tmp_3_reg_834;
assign _045_ = ap_CS_fsm[0] ? r_fu_219_p2[1:0] : trunc_ln731_reg_828;
assign _040_ = ap_CS_fsm[0] ? op_4[3] : tmp_2_reg_822;
assign _014_ = ap_CS_fsm[19] ? grp_fu_713_p2 : op_27_V_reg_1113;
assign _016_ = ap_CS_fsm[19] ? grp_fu_708_p2 : ret_V_13_reg_1108;
assign _013_ = ap_CS_fsm[12] ? grp_fu_514_p2 : op_24_V_reg_1008;
assign _031_ = ap_CS_fsm[12] ? grp_fu_506_p2[4:1] : ret_V_8_cast_reg_1001;
assign _020_ = ap_CS_fsm[12] ? grp_fu_506_p2 : ret_V_25_reg_995;
assign _010_ = ap_CS_fsm[22] ? icmp_ln851_2_fu_776_p2 : icmp_ln851_2_reg_1143;
assign _009_ = ap_CS_fsm[6] ? icmp_ln851_1_fu_414_p2 : icmp_ln851_1_reg_921;
assign _011_ = ap_CS_fsm[6] ? icmp_ln851_fu_379_p2 : icmp_ln851_reg_906;
assign _007_ = ap_CS_fsm[1] ? icmp_ln786_1_fu_282_p2 : icmp_ln786_1_reg_858;
assign _008_ = ap_CS_fsm[1] ? icmp_ln786_fu_276_p2 : icmp_ln786_reg_852;
assign _006_ = ap_CS_fsm[1] ? icmp_ln785_fu_270_p2 : icmp_ln785_reg_846;
assign _004_ = ap_CS_fsm[10] ? grp_fu_469_p2 : add_ln69_reg_978;
assign _023_ = ap_CS_fsm[10] ? ret_V_29_fu_495_p3 : ret_V_29_reg_973;
assign _034_ = ap_CS_fsm[10] ? select_ln1192_fu_475_p3[4:1] : select_ln1192_reg_968[4:1];
assign _003_ = ap_CS_fsm[17] ? grp_fu_629_p2 : add_ln69_2_reg_1098;
assign _025_ = ap_CS_fsm[17] ? ret_V_31_fu_698_p3 : ret_V_31_reg_1093;
assign _037_ = ap_CS_fsm[17] ? select_ln703_fu_674_p3 : select_ln703_reg_1088;
assign _012_ = ap_CS_fsm[17] ? grp_fu_620_p2[4:1] : op_14_V_reg_1083;
assign _002_ = _048_ ? grp_fu_452_p2 : add_ln691_reg_953;
assign _001_ = _047_ ? grp_fu_792_p2 : add_ln691_2_reg_1160;
assign _000_ = ap_CS_fsm[16] ? grp_fu_588_p2 : add_ln691_1_reg_1073;
assign _044_ = ap_CS_fsm[16] ? ret_V_21_fu_600_p2[1] : tmp_reg_1061;
assign _017_ = ap_CS_fsm[16] ? ret_V_21_fu_600_p2 : ret_V_21_reg_1055;
assign _005_ = ap_rst ? 27'h0000001 : ap_NS_fsm;
assign icmp_ln785_fu_270_p2 = _156_ ? 1'h1 : 1'h0;
assign icmp_ln786_1_fu_282_p2 = _157_ ? 1'h1 : 1'h0;
assign icmp_ln786_fu_276_p2 = _052_ ? 1'h1 : 1'h0;
assign icmp_ln851_1_fu_414_p2 = _158_ ? 1'h1 : 1'h0;
assign icmp_ln851_2_fu_776_p2 = _159_ ? 1'h1 : 1'h0;
assign icmp_ln851_fu_379_p2 = _053_ ? 1'h1 : 1'h0;
assign op_29 = ret_V_32_reg_1148[34] ? select_ln850_6_fu_804_p3 : ret_V_36_cast_reg_1153;
assign ret_V_22_fu_657_p3 = ret_V_21_reg_1055[4] ? select_ln850_fu_650_p3 : tmp_reg_1061;
assign ret_V_24_fu_442_p3 = ret_V_23_reg_884[7] ? select_ln850_1_fu_437_p3 : ret_V_3_reg_889;
assign ret_V_29_fu_495_p3 = ret_V_28_reg_931[16] ? select_ln850_4_fu_490_p3 : sext_ln831_reg_946;
assign ret_V_31_fu_698_p3 = ret_V_30_reg_1033[33] ? select_ln850_5_fu_692_p3 : ret_V_33_cast_reg_1038;
assign ret_V_9_fu_328_p3 = or_ln785_fu_322_p2 ? select_ln340_reg_864 : trunc_ln731_reg_828;
assign select_ln1192_fu_475_p3 = op_0 ? 5'h00 : 5'h1e;
assign select_ln340_fu_307_p3 = and_ln340_fu_301_p2 ? trunc_ln731_reg_828 : 2'h0;
assign select_ln353_fu_581_p3 = ret_V_25_reg_995[4] ? select_ln850_3_fu_575_p3 : ret_V_8_cast_reg_1001;
assign select_ln703_fu_674_p3 = ret_V_22_fu_657_p3 ? 5'h1f : 5'h00;
assign select_ln850_1_fu_437_p3 = icmp_ln851_reg_906 ? ret_V_3_reg_889 : ret_V_5_reg_926;
assign select_ln850_3_fu_575_p3 = ret_V_25_reg_995[0] ? ret_V_8_reg_1028 : ret_V_8_cast_reg_1001;
assign select_ln850_4_fu_490_p3 = icmp_ln851_1_reg_921 ? add_ln691_reg_953 : sext_ln831_reg_946;
assign select_ln850_5_fu_692_p3 = op_15[0] ? add_ln691_1_reg_1073 : ret_V_33_cast_reg_1038;
assign select_ln850_6_fu_804_p3 = icmp_ln851_2_reg_1143 ? add_ln691_2_reg_1160 : ret_V_36_cast_reg_1153;
assign select_ln850_fu_650_p3 = ret_V_21_reg_1055[0] ? ret_V_fu_645_p2 : tmp_reg_1061;
assign ret_V_21_fu_600_p2 = sext_ln703_reg_983 ^ { op_4, 1'h0 };
assign and_ln_fu_255_p3 = { tmp_3_reg_834, 3'h0 };
assign ap_CS_fsm_state1 = ap_CS_fsm[0];
assign ap_CS_fsm_state10 = ap_CS_fsm[9];
assign ap_CS_fsm_state11 = ap_CS_fsm[10];
assign ap_CS_fsm_state12 = ap_CS_fsm[11];
assign ap_CS_fsm_state13 = ap_CS_fsm[12];
assign ap_CS_fsm_state14 = ap_CS_fsm[13];
assign ap_CS_fsm_state15 = ap_CS_fsm[14];
assign ap_CS_fsm_state16 = ap_CS_fsm[15];
assign ap_CS_fsm_state17 = ap_CS_fsm[16];
assign ap_CS_fsm_state18 = ap_CS_fsm[17];
assign ap_CS_fsm_state19 = ap_CS_fsm[18];
assign ap_CS_fsm_state2 = ap_CS_fsm[1];
assign ap_CS_fsm_state20 = ap_CS_fsm[19];
assign ap_CS_fsm_state21 = ap_CS_fsm[20];
assign ap_CS_fsm_state22 = ap_CS_fsm[21];
assign ap_CS_fsm_state23 = ap_CS_fsm[22];
assign ap_CS_fsm_state24 = ap_CS_fsm[23];
assign ap_CS_fsm_state25 = ap_CS_fsm[24];
assign ap_CS_fsm_state26 = ap_CS_fsm[25];
assign ap_CS_fsm_state27 = ap_CS_fsm[26];
assign ap_CS_fsm_state3 = ap_CS_fsm[2];
assign ap_CS_fsm_state4 = ap_CS_fsm[3];
assign ap_CS_fsm_state5 = ap_CS_fsm[4];
assign ap_CS_fsm_state6 = ap_CS_fsm[5];
assign ap_CS_fsm_state7 = ap_CS_fsm[6];
assign ap_CS_fsm_state8 = ap_CS_fsm[7];
assign ap_CS_fsm_state9 = ap_CS_fsm[8];
assign ap_done = op_29_ap_vld;
assign ap_ready = op_29_ap_vld;
assign grp_fu_341_p0 = { ret_V_9_reg_869[1], ret_V_9_reg_869 };
assign grp_fu_341_p1 = { op_10[1], op_10 };
assign grp_fu_404_p0 = { ret_V_27_reg_901[2], ret_V_27_reg_901[2], ret_V_27_reg_901[2], ret_V_27_reg_901[2], ret_V_27_reg_901[2], ret_V_27_reg_901[2], ret_V_27_reg_901[2], ret_V_27_reg_901[2], ret_V_27_reg_901[2], ret_V_27_reg_901, 5'h00 };
assign grp_fu_404_p1 = { op_11[15], op_11 };
assign grp_fu_452_p0 = { tmp_8_reg_936[11], tmp_8_reg_936[11], tmp_8_reg_936[11], tmp_8_reg_936[11], tmp_8_reg_936[11], tmp_8_reg_936[11], tmp_8_reg_936[11], tmp_8_reg_936[11], tmp_8_reg_936[11], tmp_8_reg_936[11], tmp_8_reg_936[11], tmp_8_reg_936[11], tmp_8_reg_936[11], tmp_8_reg_936[11], tmp_8_reg_936[11], tmp_8_reg_936[11], tmp_8_reg_936[11], tmp_8_reg_936[11], tmp_8_reg_936[11], tmp_8_reg_936[11], tmp_8_reg_936 };
assign grp_fu_469_p0 = { 1'h0, ret_V_24_reg_941[5], ret_V_24_reg_941[5], ret_V_24_reg_941 };
assign grp_fu_469_p1 = { 7'h00, op_13 };
assign grp_fu_506_p1 = { op_3[3], op_3 };
assign grp_fu_514_p0 = { 23'h000000, add_ln69_reg_978 };
assign grp_fu_549_p0 = { op_24_V_reg_1008[31], op_24_V_reg_1008, 1'h0 };
assign grp_fu_549_p1 = { op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15 };
assign grp_fu_620_p0 = { select_ln353_reg_1045, 1'h0 };
assign grp_fu_629_p0 = { op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17 };
assign grp_fu_708_p0 = { op_14_V_reg_1083[3], op_14_V_reg_1083 };
assign grp_fu_735_p0 = { op_27_V_reg_1113, 3'h0 };
assign grp_fu_735_p1 = { ret_V_13_reg_1108[4], ret_V_13_reg_1108[4], ret_V_13_reg_1108[4], ret_V_13_reg_1108[4], ret_V_13_reg_1108[4], ret_V_13_reg_1108[4], ret_V_13_reg_1108[4], ret_V_13_reg_1108[4], ret_V_13_reg_1108[4], ret_V_13_reg_1108[4], ret_V_13_reg_1108[4], ret_V_13_reg_1108[4], ret_V_13_reg_1108[4], ret_V_13_reg_1108[4], ret_V_13_reg_1108[4], ret_V_13_reg_1108[4], ret_V_13_reg_1108[4], ret_V_13_reg_1108[4], ret_V_13_reg_1108[4], ret_V_13_reg_1108[4], ret_V_13_reg_1108[4], ret_V_13_reg_1108[4], ret_V_13_reg_1108[4], ret_V_13_reg_1108[4], ret_V_13_reg_1108[4], ret_V_13_reg_1108[4], ret_V_13_reg_1108[4], ret_V_13_reg_1108, 3'h0 };
assign grp_fu_766_p0 = { tmp_5_reg_1128[31], tmp_5_reg_1128, 2'h0 };
assign grp_fu_766_p1 = { op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19 };
assign lhs_fu_347_p3 = { op_5, 2'h0 };
assign op_18_V_fu_717_p3 = { ret_V_13_reg_1108, 3'h0 };
assign or_ln786_fu_287_p2 = or_ln786_1_fu_314_p2;
assign or_ln_fu_262_p4 = { tmp_3_reg_834, 1'h0, p_Result_s_16_reg_840 };
assign p_Result_1_fu_430_p3 = ret_V_23_reg_884[7];
assign p_Result_2_fu_565_p3 = ret_V_25_reg_995[4];
assign p_Result_3_fu_483_p3 = ret_V_28_reg_931[16];
assign p_Result_4_fu_682_p3 = ret_V_30_reg_1033[33];
assign p_Result_5_fu_797_p3 = ret_V_32_reg_1148[34];
assign p_Result_s_fu_635_p3 = ret_V_21_reg_1055[4];
assign rhs_5_fu_538_p3 = { op_24_V_reg_1008, 1'h0 };
assign rhs_8_fu_755_p3 = { tmp_5_reg_1128, 2'h0 };
assign rhs_fu_593_p3 = { op_4, 1'h0 };
assign sext_ln1192_1_fu_389_p0 = op_11;
assign sext_ln1194_fu_355_p1 = { op_5[3], op_5[3], op_5, 2'h0 };
assign sext_ln69_1_fu_458_p1 = { ret_V_24_reg_941[5], ret_V_24_reg_941[5], ret_V_24_reg_941 };
assign sext_ln703_2_fu_534_p0 = op_15;
assign sext_ln703_3_fu_751_p0 = op_19;
assign sext_ln703_fu_502_p1 = { op_3[3], op_3 };
assign sext_ln831_fu_449_p1 = { tmp_8_reg_936[11], tmp_8_reg_936[11], tmp_8_reg_936[11], tmp_8_reg_936[11], tmp_8_reg_936[11], tmp_8_reg_936[11], tmp_8_reg_936[11], tmp_8_reg_936[11], tmp_8_reg_936[11], tmp_8_reg_936[11], tmp_8_reg_936[11], tmp_8_reg_936[11], tmp_8_reg_936[11], tmp_8_reg_936[11], tmp_8_reg_936[11], tmp_8_reg_936[11], tmp_8_reg_936[11], tmp_8_reg_936[11], tmp_8_reg_936[11], tmp_8_reg_936[11], tmp_8_reg_936 };
assign tmp_4_fu_393_p3 = { ret_V_27_reg_901, 5'h00 };
assign trunc_ln731_fu_233_p1 = r_fu_219_p2[1:0];
assign trunc_ln851_1_fu_375_p1 = ret_V_23_fu_359_p2[1:0];
assign trunc_ln851_2_fu_572_p1 = ret_V_25_reg_995[0];
assign trunc_ln851_3_fu_410_p0 = op_11;
assign trunc_ln851_3_fu_410_p1 = op_11[4:0];
assign trunc_ln851_4_fu_689_p0 = op_15;
assign trunc_ln851_4_fu_689_p1 = op_15[0];
assign trunc_ln851_5_fu_772_p0 = op_19;
assign trunc_ln851_5_fu_772_p1 = op_19[1:0];
assign trunc_ln851_fu_642_p1 = ret_V_21_reg_1055[0];
assign \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.ain_s0  = \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.a ;
assign \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.bin_s0  = \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.b ;
assign \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.s  = { \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.fas_s2 , \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.sum_s1  };
assign \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.u2.a  = \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.ain_s1 ;
assign \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.u2.b  = \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.bin_s1 ;
assign \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.u2.cin  = \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.carry_s1 ;
assign \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.facout_s2  = \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.u2.cout ;
assign \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.fas_s2  = \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.u2.s ;
assign \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.u1.a  = \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.a [3:0];
assign \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.u1.b  = \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.b [3:0];
assign \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.u1.cin  = 1'h0;
assign \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.facout_s1  = \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.u1.cout ;
assign \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.fas_s1  = \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.u1.s ;
assign \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.a  = \add_9ns_9ns_9_2_1_U5.din0 ;
assign \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.b  = \add_9ns_9ns_9_2_1_U5.din1 ;
assign \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.ce  = \add_9ns_9ns_9_2_1_U5.ce ;
assign \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.clk  = \add_9ns_9ns_9_2_1_U5.clk ;
assign \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.reset  = \add_9ns_9ns_9_2_1_U5.reset ;
assign \add_9ns_9ns_9_2_1_U5.dout  = \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.s ;
assign \add_9ns_9ns_9_2_1_U5.ce  = 1'h1;
assign \add_9ns_9ns_9_2_1_U5.clk  = ap_clk;
assign \add_9ns_9ns_9_2_1_U5.din0  = { 1'h0, ret_V_24_reg_941[5], ret_V_24_reg_941[5], ret_V_24_reg_941 };
assign \add_9ns_9ns_9_2_1_U5.din1  = { 7'h00, op_13 };
assign grp_fu_469_p2 = \add_9ns_9ns_9_2_1_U5.dout ;
assign \add_9ns_9ns_9_2_1_U5.reset  = ap_rst;
assign \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.ain_s0  = \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.a ;
assign \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.bin_s0  = \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.b ;
assign \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.s  = { \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.fas_s2 , \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.sum_s1  };
assign \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.u2.a  = \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.ain_s1 ;
assign \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.u2.b  = \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.bin_s1 ;
assign \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.u2.cin  = \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.carry_s1 ;
assign \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.facout_s2  = \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.u2.cout ;
assign \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.fas_s2  = \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.u2.s ;
assign \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.u1.a  = \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.a [2:0];
assign \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.u1.b  = \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.b [2:0];
assign \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.u1.cin  = 1'h0;
assign \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.facout_s1  = \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.u1.cout ;
assign \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.fas_s1  = \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.u1.s ;
assign \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.a  = \add_6ns_6ns_6_2_1_U2.din0 ;
assign \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.b  = \add_6ns_6ns_6_2_1_U2.din1 ;
assign \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.ce  = \add_6ns_6ns_6_2_1_U2.ce ;
assign \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.clk  = \add_6ns_6ns_6_2_1_U2.clk ;
assign \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.reset  = \add_6ns_6ns_6_2_1_U2.reset ;
assign \add_6ns_6ns_6_2_1_U2.dout  = \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.s ;
assign \add_6ns_6ns_6_2_1_U2.ce  = 1'h1;
assign \add_6ns_6ns_6_2_1_U2.clk  = ap_clk;
assign \add_6ns_6ns_6_2_1_U2.din0  = ret_V_3_reg_889;
assign \add_6ns_6ns_6_2_1_U2.din1  = 6'h01;
assign grp_fu_384_p2 = \add_6ns_6ns_6_2_1_U2.dout ;
assign \add_6ns_6ns_6_2_1_U2.reset  = ap_rst;
assign \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.ain_s0  = \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.a ;
assign \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.bin_s0  = \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.b ;
assign \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.s  = { \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.fas_s2 , \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.sum_s1  };
assign \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.u2.a  = \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.ain_s1 ;
assign \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.u2.b  = \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.bin_s1 ;
assign \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.u2.cin  = \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.carry_s1 ;
assign \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.facout_s2  = \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.u2.cout ;
assign \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.fas_s2  = \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.u2.s ;
assign \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.u1.a  = \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.a [1:0];
assign \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.u1.b  = \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.b [1:0];
assign \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.u1.cin  = 1'h0;
assign \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.facout_s1  = \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.u1.cout ;
assign \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.fas_s1  = \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.u1.s ;
assign \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.a  = \add_5s_5ns_5_2_1_U13.din0 ;
assign \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.b  = \add_5s_5ns_5_2_1_U13.din1 ;
assign \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.ce  = \add_5s_5ns_5_2_1_U13.ce ;
assign \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.clk  = \add_5s_5ns_5_2_1_U13.clk ;
assign \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.reset  = \add_5s_5ns_5_2_1_U13.reset ;
assign \add_5s_5ns_5_2_1_U13.dout  = \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.s ;
assign \add_5s_5ns_5_2_1_U13.ce  = 1'h1;
assign \add_5s_5ns_5_2_1_U13.clk  = ap_clk;
assign \add_5s_5ns_5_2_1_U13.din0  = { op_14_V_reg_1083[3], op_14_V_reg_1083 };
assign \add_5s_5ns_5_2_1_U13.din1  = select_ln703_reg_1088;
assign grp_fu_708_p2 = \add_5s_5ns_5_2_1_U13.dout ;
assign \add_5s_5ns_5_2_1_U13.reset  = ap_rst;
assign \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.ain_s0  = \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.a ;
assign \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.bin_s0  = \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.b ;
assign \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.s  = { \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.fas_s2 , \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.sum_s1  };
assign \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.u2.a  = \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.ain_s1 ;
assign \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.u2.b  = \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.bin_s1 ;
assign \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.u2.cin  = \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.carry_s1 ;
assign \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.facout_s2  = \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.u2.cout ;
assign \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.fas_s2  = \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.u2.s ;
assign \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.u1.a  = \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.a [1:0];
assign \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.u1.b  = \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.b [1:0];
assign \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.u1.cin  = 1'h0;
assign \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.facout_s1  = \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.u1.cout ;
assign \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.fas_s1  = \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.u1.s ;
assign \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.a  = \add_5ns_5s_5_2_1_U6.din0 ;
assign \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.b  = \add_5ns_5s_5_2_1_U6.din1 ;
assign \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.ce  = \add_5ns_5s_5_2_1_U6.ce ;
assign \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.clk  = \add_5ns_5s_5_2_1_U6.clk ;
assign \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.reset  = \add_5ns_5s_5_2_1_U6.reset ;
assign \add_5ns_5s_5_2_1_U6.dout  = \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.s ;
assign \add_5ns_5s_5_2_1_U6.ce  = 1'h1;
assign \add_5ns_5s_5_2_1_U6.clk  = ap_clk;
assign \add_5ns_5s_5_2_1_U6.din0  = select_ln1192_reg_968;
assign \add_5ns_5s_5_2_1_U6.din1  = { op_3[3], op_3 };
assign grp_fu_506_p2 = \add_5ns_5s_5_2_1_U6.dout ;
assign \add_5ns_5s_5_2_1_U6.reset  = ap_rst;
assign \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.ain_s0  = \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.a ;
assign \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.bin_s0  = \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.b ;
assign \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.s  = { \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.fas_s2 , \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.sum_s1  };
assign \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.u2.a  = \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.ain_s1 ;
assign \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.u2.b  = \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.bin_s1 ;
assign \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.u2.cin  = \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.carry_s1 ;
assign \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.facout_s2  = \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.u2.cout ;
assign \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.fas_s2  = \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.u2.s ;
assign \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.u1.a  = \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.a [1:0];
assign \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.u1.b  = \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.b [1:0];
assign \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.u1.cin  = 1'h0;
assign \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.facout_s1  = \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.u1.cout ;
assign \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.fas_s1  = \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.u1.s ;
assign \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.a  = \add_5ns_5s_5_2_1_U11.din0 ;
assign \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.b  = \add_5ns_5s_5_2_1_U11.din1 ;
assign \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.ce  = \add_5ns_5s_5_2_1_U11.ce ;
assign \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.clk  = \add_5ns_5s_5_2_1_U11.clk ;
assign \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.reset  = \add_5ns_5s_5_2_1_U11.reset ;
assign \add_5ns_5s_5_2_1_U11.dout  = \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.s ;
assign \add_5ns_5s_5_2_1_U11.ce  = 1'h1;
assign \add_5ns_5s_5_2_1_U11.clk  = ap_clk;
assign \add_5ns_5s_5_2_1_U11.din0  = { select_ln353_reg_1045, 1'h0 };
assign \add_5ns_5s_5_2_1_U11.din1  = sext_ln703_reg_983;
assign grp_fu_620_p2 = \add_5ns_5s_5_2_1_U11.dout ;
assign \add_5ns_5s_5_2_1_U11.reset  = ap_rst;
assign \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.ain_s0  = \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.a ;
assign \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.bin_s0  = \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.b ;
assign \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.s  = { \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.fas_s2 , \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.sum_s1  };
assign \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.u2.a  = \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.ain_s1 ;
assign \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.u2.b  = \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.bin_s1 ;
assign \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.u2.cin  = \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.carry_s1 ;
assign \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.facout_s2  = \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.u2.cout ;
assign \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.fas_s2  = \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.u2.s ;
assign \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.u1.a  = \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.a [1:0];
assign \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.u1.b  = \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.b [1:0];
assign \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.u1.cin  = 1'h0;
assign \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.facout_s1  = \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.u1.cout ;
assign \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.fas_s1  = \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.u1.s ;
assign \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.a  = \add_4ns_4ns_4_2_1_U8.din0 ;
assign \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.b  = \add_4ns_4ns_4_2_1_U8.din1 ;
assign \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.ce  = \add_4ns_4ns_4_2_1_U8.ce ;
assign \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.clk  = \add_4ns_4ns_4_2_1_U8.clk ;
assign \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.reset  = \add_4ns_4ns_4_2_1_U8.reset ;
assign \add_4ns_4ns_4_2_1_U8.dout  = \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.s ;
assign \add_4ns_4ns_4_2_1_U8.ce  = 1'h1;
assign \add_4ns_4ns_4_2_1_U8.clk  = ap_clk;
assign \add_4ns_4ns_4_2_1_U8.din0  = ret_V_8_cast_reg_1001;
assign \add_4ns_4ns_4_2_1_U8.din1  = 4'h1;
assign grp_fu_529_p2 = \add_4ns_4ns_4_2_1_U8.dout ;
assign \add_4ns_4ns_4_2_1_U8.reset  = ap_rst;
assign \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.ain_s0  = \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.a ;
assign \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.bin_s0  = \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.b ;
assign \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.s  = { \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.fas_s2 , \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.sum_s1  };
assign \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.u2.a  = \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.ain_s1 ;
assign \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.u2.b  = \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.bin_s1 ;
assign \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.u2.cin  = \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.carry_s1 ;
assign \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.facout_s2  = \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.u2.cout ;
assign \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.fas_s2  = \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.u2.s ;
assign \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.u1.a  = \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.a [0];
assign \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.u1.b  = \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.b [0];
assign \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.u1.cin  = 1'h0;
assign \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.facout_s1  = \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.u1.cout ;
assign \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.fas_s1  = \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.u1.s ;
assign \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.a  = \add_3s_3s_3_2_1_U1.din0 ;
assign \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.b  = \add_3s_3s_3_2_1_U1.din1 ;
assign \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.ce  = \add_3s_3s_3_2_1_U1.ce ;
assign \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.clk  = \add_3s_3s_3_2_1_U1.clk ;
assign \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.reset  = \add_3s_3s_3_2_1_U1.reset ;
assign \add_3s_3s_3_2_1_U1.dout  = \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.s ;
assign \add_3s_3s_3_2_1_U1.ce  = 1'h1;
assign \add_3s_3s_3_2_1_U1.clk  = ap_clk;
assign \add_3s_3s_3_2_1_U1.din0  = { ret_V_9_reg_869[1], ret_V_9_reg_869 };
assign \add_3s_3s_3_2_1_U1.din1  = { op_10[1], op_10 };
assign grp_fu_341_p2 = \add_3s_3s_3_2_1_U1.dout ;
assign \add_3s_3s_3_2_1_U1.reset  = ap_rst;
assign \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.ain_s0  = \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.a ;
assign \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.bin_s0  = \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.b ;
assign \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.s  = { \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.fas_s2 , \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.sum_s1  };
assign \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.u2.a  = \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.ain_s1 ;
assign \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.u2.b  = \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.bin_s1 ;
assign \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.u2.cin  = \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.carry_s1 ;
assign \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.facout_s2  = \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.u2.cout ;
assign \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.fas_s2  = \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.u2.s ;
assign \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.u1.a  = \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.a [16:0];
assign \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.u1.b  = \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.b [16:0];
assign \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.u1.cin  = 1'h0;
assign \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.facout_s1  = \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.u1.cout ;
assign \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.fas_s1  = \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.u1.s ;
assign \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.a  = \add_35s_35s_35_2_1_U16.din0 ;
assign \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.b  = \add_35s_35s_35_2_1_U16.din1 ;
assign \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.ce  = \add_35s_35s_35_2_1_U16.ce ;
assign \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.clk  = \add_35s_35s_35_2_1_U16.clk ;
assign \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.reset  = \add_35s_35s_35_2_1_U16.reset ;
assign \add_35s_35s_35_2_1_U16.dout  = \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.s ;
assign \add_35s_35s_35_2_1_U16.ce  = 1'h1;
assign \add_35s_35s_35_2_1_U16.clk  = ap_clk;
assign \add_35s_35s_35_2_1_U16.din0  = { tmp_5_reg_1128[31], tmp_5_reg_1128, 2'h0 };
assign \add_35s_35s_35_2_1_U16.din1  = { op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19 };
assign grp_fu_766_p2 = \add_35s_35s_35_2_1_U16.dout ;
assign \add_35s_35s_35_2_1_U16.reset  = ap_rst;
assign \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.ain_s0  = \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.a ;
assign \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.bin_s0  = \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.b ;
assign \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.s  = { \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.fas_s2 , \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.sum_s1  };
assign \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.u2.a  = \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.ain_s1 ;
assign \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.u2.b  = \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.bin_s1 ;
assign \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.u2.cin  = \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.carry_s1 ;
assign \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.facout_s2  = \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.u2.cout ;
assign \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.fas_s2  = \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.u2.s ;
assign \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.u1.a  = \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.a [16:0];
assign \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.u1.b  = \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.b [16:0];
assign \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.u1.cin  = 1'h0;
assign \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.facout_s1  = \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.u1.cout ;
assign \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.fas_s1  = \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.u1.s ;
assign \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.a  = \add_35ns_35s_35_2_1_U15.din0 ;
assign \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.b  = \add_35ns_35s_35_2_1_U15.din1 ;
assign \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.ce  = \add_35ns_35s_35_2_1_U15.ce ;
assign \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.clk  = \add_35ns_35s_35_2_1_U15.clk ;
assign \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.reset  = \add_35ns_35s_35_2_1_U15.reset ;
assign \add_35ns_35s_35_2_1_U15.dout  = \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.s ;
assign \add_35ns_35s_35_2_1_U15.ce  = 1'h1;
assign \add_35ns_35s_35_2_1_U15.clk  = ap_clk;
assign \add_35ns_35s_35_2_1_U15.din0  = { op_27_V_reg_1113, 3'h0 };
assign \add_35ns_35s_35_2_1_U15.din1  = { ret_V_13_reg_1108[4], ret_V_13_reg_1108[4], ret_V_13_reg_1108[4], ret_V_13_reg_1108[4], ret_V_13_reg_1108[4], ret_V_13_reg_1108[4], ret_V_13_reg_1108[4], ret_V_13_reg_1108[4], ret_V_13_reg_1108[4], ret_V_13_reg_1108[4], ret_V_13_reg_1108[4], ret_V_13_reg_1108[4], ret_V_13_reg_1108[4], ret_V_13_reg_1108[4], ret_V_13_reg_1108[4], ret_V_13_reg_1108[4], ret_V_13_reg_1108[4], ret_V_13_reg_1108[4], ret_V_13_reg_1108[4], ret_V_13_reg_1108[4], ret_V_13_reg_1108[4], ret_V_13_reg_1108[4], ret_V_13_reg_1108[4], ret_V_13_reg_1108[4], ret_V_13_reg_1108[4], ret_V_13_reg_1108[4], ret_V_13_reg_1108[4], ret_V_13_reg_1108, 3'h0 };
assign grp_fu_735_p2 = \add_35ns_35s_35_2_1_U15.dout ;
assign \add_35ns_35s_35_2_1_U15.reset  = ap_rst;
assign \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.ain_s0  = \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.a ;
assign \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.bin_s0  = \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.b ;
assign \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.s  = { \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.fas_s2 , \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.sum_s1  };
assign \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.u2.a  = \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.ain_s1 ;
assign \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.u2.b  = \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.bin_s1 ;
assign \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.u2.cin  = \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.carry_s1 ;
assign \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.facout_s2  = \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.u2.cout ;
assign \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.fas_s2  = \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.u2.s ;
assign \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.u1.a  = \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.a [16:0];
assign \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.u1.b  = \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.b [16:0];
assign \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.u1.cin  = 1'h0;
assign \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.facout_s1  = \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.u1.cout ;
assign \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.fas_s1  = \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.u1.s ;
assign \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.a  = \add_34s_34s_34_2_1_U9.din0 ;
assign \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.b  = \add_34s_34s_34_2_1_U9.din1 ;
assign \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.ce  = \add_34s_34s_34_2_1_U9.ce ;
assign \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.clk  = \add_34s_34s_34_2_1_U9.clk ;
assign \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.reset  = \add_34s_34s_34_2_1_U9.reset ;
assign \add_34s_34s_34_2_1_U9.dout  = \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.s ;
assign \add_34s_34s_34_2_1_U9.ce  = 1'h1;
assign \add_34s_34s_34_2_1_U9.clk  = ap_clk;
assign \add_34s_34s_34_2_1_U9.din0  = { op_24_V_reg_1008[31], op_24_V_reg_1008, 1'h0 };
assign \add_34s_34s_34_2_1_U9.din1  = { op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15 };
assign grp_fu_549_p2 = \add_34s_34s_34_2_1_U9.dout ;
assign \add_34s_34s_34_2_1_U9.reset  = ap_rst;
assign \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.ain_s0  = \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.a ;
assign \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.bin_s0  = \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.b ;
assign \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.s  = { \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.fas_s2 , \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.sum_s1  };
assign \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.u2.a  = \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.ain_s1 ;
assign \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.u2.b  = \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.bin_s1 ;
assign \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.u2.cin  = \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.carry_s1 ;
assign \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.facout_s2  = \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.u2.cout ;
assign \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.fas_s2  = \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.u2.s ;
assign \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.u1.a  = \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.a [15:0];
assign \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.u1.b  = \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.b [15:0];
assign \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.u1.cin  = 1'h0;
assign \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.facout_s1  = \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.u1.cout ;
assign \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.fas_s1  = \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.u1.s ;
assign \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.a  = \add_32s_32ns_32_2_1_U4.din0 ;
assign \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.b  = \add_32s_32ns_32_2_1_U4.din1 ;
assign \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.ce  = \add_32s_32ns_32_2_1_U4.ce ;
assign \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.clk  = \add_32s_32ns_32_2_1_U4.clk ;
assign \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.reset  = \add_32s_32ns_32_2_1_U4.reset ;
assign \add_32s_32ns_32_2_1_U4.dout  = \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.s ;
assign \add_32s_32ns_32_2_1_U4.ce  = 1'h1;
assign \add_32s_32ns_32_2_1_U4.clk  = ap_clk;
assign \add_32s_32ns_32_2_1_U4.din0  = { tmp_8_reg_936[11], tmp_8_reg_936[11], tmp_8_reg_936[11], tmp_8_reg_936[11], tmp_8_reg_936[11], tmp_8_reg_936[11], tmp_8_reg_936[11], tmp_8_reg_936[11], tmp_8_reg_936[11], tmp_8_reg_936[11], tmp_8_reg_936[11], tmp_8_reg_936[11], tmp_8_reg_936[11], tmp_8_reg_936[11], tmp_8_reg_936[11], tmp_8_reg_936[11], tmp_8_reg_936[11], tmp_8_reg_936[11], tmp_8_reg_936[11], tmp_8_reg_936[11], tmp_8_reg_936 };
assign \add_32s_32ns_32_2_1_U4.din1  = 32'd1;
assign grp_fu_452_p2 = \add_32s_32ns_32_2_1_U4.dout ;
assign \add_32s_32ns_32_2_1_U4.reset  = ap_rst;
assign \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.ain_s0  = \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.a ;
assign \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.bin_s0  = \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.b ;
assign \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.s  = { \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.fas_s2 , \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.sum_s1  };
assign \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.u2.a  = \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.ain_s1 ;
assign \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.u2.b  = \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.bin_s1 ;
assign \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.u2.cin  = \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.carry_s1 ;
assign \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.facout_s2  = \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.u2.cout ;
assign \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.fas_s2  = \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.u2.s ;
assign \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.u1.a  = \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.a [15:0];
assign \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.u1.b  = \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.b [15:0];
assign \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.u1.cin  = 1'h0;
assign \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.facout_s1  = \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.u1.cout ;
assign \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.fas_s1  = \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.u1.s ;
assign \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.a  = \add_32s_32ns_32_2_1_U12.din0 ;
assign \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.b  = \add_32s_32ns_32_2_1_U12.din1 ;
assign \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.ce  = \add_32s_32ns_32_2_1_U12.ce ;
assign \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.clk  = \add_32s_32ns_32_2_1_U12.clk ;
assign \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.reset  = \add_32s_32ns_32_2_1_U12.reset ;
assign \add_32s_32ns_32_2_1_U12.dout  = \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.s ;
assign \add_32s_32ns_32_2_1_U12.ce  = 1'h1;
assign \add_32s_32ns_32_2_1_U12.clk  = ap_clk;
assign \add_32s_32ns_32_2_1_U12.din0  = { op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17 };
assign \add_32s_32ns_32_2_1_U12.din1  = op_16;
assign grp_fu_629_p2 = \add_32s_32ns_32_2_1_U12.dout ;
assign \add_32s_32ns_32_2_1_U12.reset  = ap_rst;
assign \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s0  = \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.a ;
assign \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s0  = \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.b ;
assign \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.s  = { \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s2 , \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.sum_s1  };
assign \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.a  = \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s1 ;
assign \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.b  = \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s1 ;
assign \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cin  = \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.carry_s1 ;
assign \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s2  = \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cout ;
assign \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s2  = \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.s ;
assign \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.a  = \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.a [15:0];
assign \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.b  = \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.b [15:0];
assign \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cin  = 1'h0;
assign \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s1  = \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cout ;
assign \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s1  = \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.s ;
assign \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.a  = \add_32ns_32ns_32_2_1_U7.din0 ;
assign \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.b  = \add_32ns_32ns_32_2_1_U7.din1 ;
assign \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  = \add_32ns_32ns_32_2_1_U7.ce ;
assign \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.clk  = \add_32ns_32ns_32_2_1_U7.clk ;
assign \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.reset  = \add_32ns_32ns_32_2_1_U7.reset ;
assign \add_32ns_32ns_32_2_1_U7.dout  = \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.s ;
assign \add_32ns_32ns_32_2_1_U7.ce  = 1'h1;
assign \add_32ns_32ns_32_2_1_U7.clk  = ap_clk;
assign \add_32ns_32ns_32_2_1_U7.din0  = { 23'h000000, add_ln69_reg_978 };
assign \add_32ns_32ns_32_2_1_U7.din1  = ret_V_29_reg_973;
assign grp_fu_514_p2 = \add_32ns_32ns_32_2_1_U7.dout ;
assign \add_32ns_32ns_32_2_1_U7.reset  = ap_rst;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s0  = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.a ;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s0  = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.b ;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.s  = { \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s2 , \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.sum_s1  };
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.a  = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s1 ;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.b  = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s1 ;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cin  = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.carry_s1 ;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s2  = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cout ;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s2  = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.s ;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.a  = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.a [15:0];
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.b  = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.b [15:0];
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cin  = 1'h0;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s1  = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cout ;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s1  = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.s ;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.a  = \add_32ns_32ns_32_2_1_U17.din0 ;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.b  = \add_32ns_32ns_32_2_1_U17.din1 ;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  = \add_32ns_32ns_32_2_1_U17.ce ;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.clk  = \add_32ns_32ns_32_2_1_U17.clk ;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.reset  = \add_32ns_32ns_32_2_1_U17.reset ;
assign \add_32ns_32ns_32_2_1_U17.dout  = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.s ;
assign \add_32ns_32ns_32_2_1_U17.ce  = 1'h1;
assign \add_32ns_32ns_32_2_1_U17.clk  = ap_clk;
assign \add_32ns_32ns_32_2_1_U17.din0  = ret_V_36_cast_reg_1153;
assign \add_32ns_32ns_32_2_1_U17.din1  = 32'd1;
assign grp_fu_792_p2 = \add_32ns_32ns_32_2_1_U17.dout ;
assign \add_32ns_32ns_32_2_1_U17.reset  = ap_rst;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s0  = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.a ;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s0  = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.b ;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.s  = { \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s2 , \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.sum_s1  };
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.a  = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s1 ;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.b  = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s1 ;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cin  = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.carry_s1 ;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s2  = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cout ;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s2  = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.s ;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.a  = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.a [15:0];
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.b  = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.b [15:0];
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cin  = 1'h0;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s1  = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cout ;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s1  = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.s ;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.a  = \add_32ns_32ns_32_2_1_U14.din0 ;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.b  = \add_32ns_32ns_32_2_1_U14.din1 ;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  = \add_32ns_32ns_32_2_1_U14.ce ;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.clk  = \add_32ns_32ns_32_2_1_U14.clk ;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.reset  = \add_32ns_32ns_32_2_1_U14.reset ;
assign \add_32ns_32ns_32_2_1_U14.dout  = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.s ;
assign \add_32ns_32ns_32_2_1_U14.ce  = 1'h1;
assign \add_32ns_32ns_32_2_1_U14.clk  = ap_clk;
assign \add_32ns_32ns_32_2_1_U14.din0  = add_ln69_2_reg_1098;
assign \add_32ns_32ns_32_2_1_U14.din1  = ret_V_31_reg_1093;
assign grp_fu_713_p2 = \add_32ns_32ns_32_2_1_U14.dout ;
assign \add_32ns_32ns_32_2_1_U14.reset  = ap_rst;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s0  = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.a ;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s0  = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.b ;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.s  = { \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s2 , \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.sum_s1  };
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.a  = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s1 ;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.b  = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s1 ;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cin  = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.carry_s1 ;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s2  = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cout ;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s2  = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.s ;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.a  = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.a [15:0];
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.b  = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.b [15:0];
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cin  = 1'h0;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s1  = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cout ;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s1  = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.s ;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.a  = \add_32ns_32ns_32_2_1_U10.din0 ;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.b  = \add_32ns_32ns_32_2_1_U10.din1 ;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  = \add_32ns_32ns_32_2_1_U10.ce ;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.clk  = \add_32ns_32ns_32_2_1_U10.clk ;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.reset  = \add_32ns_32ns_32_2_1_U10.reset ;
assign \add_32ns_32ns_32_2_1_U10.dout  = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.s ;
assign \add_32ns_32ns_32_2_1_U10.ce  = 1'h1;
assign \add_32ns_32ns_32_2_1_U10.clk  = ap_clk;
assign \add_32ns_32ns_32_2_1_U10.din0  = ret_V_33_cast_reg_1038;
assign \add_32ns_32ns_32_2_1_U10.din1  = 32'd1;
assign grp_fu_588_p2 = \add_32ns_32ns_32_2_1_U10.dout ;
assign \add_32ns_32ns_32_2_1_U10.reset  = ap_rst;
assign \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.ain_s0  = \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.a ;
assign \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.bin_s0  = \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.b ;
assign \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.s  = { \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.fas_s2 , \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.sum_s1  };
assign \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.u2.a  = \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.ain_s1 ;
assign \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.u2.b  = \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.bin_s1 ;
assign \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.u2.cin  = \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.carry_s1 ;
assign \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.facout_s2  = \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.u2.cout ;
assign \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.fas_s2  = \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.u2.s ;
assign \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.u1.a  = \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.a [7:0];
assign \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.u1.b  = \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.b [7:0];
assign \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.u1.cin  = 1'h0;
assign \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.facout_s1  = \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.u1.cout ;
assign \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.fas_s1  = \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.u1.s ;
assign \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.a  = \add_17s_17s_17_2_1_U3.din0 ;
assign \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.b  = \add_17s_17s_17_2_1_U3.din1 ;
assign \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.ce  = \add_17s_17s_17_2_1_U3.ce ;
assign \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.clk  = \add_17s_17s_17_2_1_U3.clk ;
assign \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.reset  = \add_17s_17s_17_2_1_U3.reset ;
assign \add_17s_17s_17_2_1_U3.dout  = \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.s ;
assign \add_17s_17s_17_2_1_U3.ce  = 1'h1;
assign \add_17s_17s_17_2_1_U3.clk  = ap_clk;
assign \add_17s_17s_17_2_1_U3.din0  = { ret_V_27_reg_901[2], ret_V_27_reg_901[2], ret_V_27_reg_901[2], ret_V_27_reg_901[2], ret_V_27_reg_901[2], ret_V_27_reg_901[2], ret_V_27_reg_901[2], ret_V_27_reg_901[2], ret_V_27_reg_901[2], ret_V_27_reg_901, 5'h00 };
assign \add_17s_17s_17_2_1_U3.din1  = { op_11[15], op_11 };
assign grp_fu_404_p2 = \add_17s_17s_17_2_1_U3.dout ;
assign \add_17s_17s_17_2_1_U3.reset  = ap_rst;
endmodule


// Machine B:
// Processed by function `add_clk_enable_signal` in `verilog_tricks.py`.
// Processed by function `remove_reset_signal` in `verilog_tricks.py`.
module top_B (
  ap_clk,
  ap_start,
  ap_done,
  ap_idle,
  ap_ready,
  op_0,
  op_3,
  op_4,
  op_5,
  op_9,
  op_10,
  op_11,
  op_13,
  op_15,
  op_16,
  op_17,
  op_19,
  op_29,
  op_29_ap_vld,
clk_enable
);
input clk_enable;


input ap_clk;
wire ap_rst;
assign ap_rst = op_29_ap_vld;
input ap_start;
input op_0;
input [1:0] op_10;
input [15:0] op_11;
input [1:0] op_13;
input [3:0] op_15;
input [31:0] op_16;
input [3:0] op_17;
input [3:0] op_19;
input [3:0] op_3;
input [3:0] op_4;
input [3:0] op_5;
input [7:0] op_9;
output ap_done;
output ap_idle;
output ap_ready;
output [31:0] op_29;
output op_29_ap_vld;


reg [8:0] \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.ain_s1 ;
reg [8:0] \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.bin_s1 ;
reg \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.carry_s1 ;
reg [7:0] \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.sum_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s1 ;
reg \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.carry_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.sum_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s1 ;
reg \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.carry_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.sum_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s1 ;
reg \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.carry_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.sum_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s1 ;
reg \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.carry_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.sum_s1 ;
reg [15:0] \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.ain_s1 ;
reg [15:0] \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.bin_s1 ;
reg \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.carry_s1 ;
reg [15:0] \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.sum_s1 ;
reg [15:0] \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.ain_s1 ;
reg [15:0] \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.bin_s1 ;
reg \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.carry_s1 ;
reg [15:0] \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.sum_s1 ;
reg [16:0] \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.ain_s1 ;
reg [16:0] \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.bin_s1 ;
reg \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.carry_s1 ;
reg [16:0] \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.sum_s1 ;
reg [17:0] \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.ain_s1 ;
reg [17:0] \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.bin_s1 ;
reg \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.carry_s1 ;
reg [16:0] \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.sum_s1 ;
reg [17:0] \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.ain_s1 ;
reg [17:0] \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.bin_s1 ;
reg \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.carry_s1 ;
reg [16:0] \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.sum_s1 ;
reg [1:0] \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.ain_s1 ;
reg [1:0] \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.bin_s1 ;
reg \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.carry_s1 ;
reg \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.sum_s1 ;
reg [1:0] \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.ain_s1 ;
reg [1:0] \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.bin_s1 ;
reg \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.carry_s1 ;
reg [1:0] \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.sum_s1 ;
reg [2:0] \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.ain_s1 ;
reg [2:0] \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.bin_s1 ;
reg \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.carry_s1 ;
reg [1:0] \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.sum_s1 ;
reg [2:0] \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.ain_s1 ;
reg [2:0] \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.bin_s1 ;
reg \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.carry_s1 ;
reg [1:0] \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.sum_s1 ;
reg [2:0] \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.ain_s1 ;
reg [2:0] \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.bin_s1 ;
reg \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.carry_s1 ;
reg [1:0] \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.sum_s1 ;
reg [2:0] \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.ain_s1 ;
reg [2:0] \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.bin_s1 ;
reg \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.carry_s1 ;
reg [2:0] \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.sum_s1 ;
reg [4:0] \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.ain_s1 ;
reg [4:0] \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.bin_s1 ;
reg \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.carry_s1 ;
reg [3:0] \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.sum_s1 ;
reg [31:0] add_ln691_1_reg_1073;
reg [31:0] add_ln691_2_reg_1160;
reg [31:0] add_ln691_reg_953;
reg [31:0] add_ln69_2_reg_1098;
reg [8:0] add_ln69_reg_978;
reg [26:0] ap_CS_fsm = 27'h0000001;
reg icmp_ln785_reg_846;
reg icmp_ln786_1_reg_858;
reg icmp_ln786_reg_852;
reg icmp_ln851_1_reg_921;
reg icmp_ln851_2_reg_1143;
reg icmp_ln851_reg_906;
reg [3:0] op_14_V_reg_1083;
reg [31:0] op_24_V_reg_1008;
reg [31:0] op_27_V_reg_1113;
reg [1:0] p_Result_s_16_reg_840;
reg [4:0] ret_V_13_reg_1108;
reg [4:0] ret_V_21_reg_1055;
reg [5:0] ret_V_24_reg_941;
reg [4:0] ret_V_25_reg_995;
reg [2:0] ret_V_27_reg_901;
reg [16:0] ret_V_28_reg_931;
reg [31:0] ret_V_29_reg_973;
reg [33:0] ret_V_30_reg_1033;
reg [31:0] ret_V_31_reg_1093;
reg [34:0] ret_V_32_reg_1148;
reg [31:0] ret_V_33_cast_reg_1038;
reg [31:0] ret_V_36_cast_reg_1153;
reg [5:0] ret_V_3_reg_889;
reg [5:0] ret_V_5_reg_926;
reg [3:0] ret_V_8_cast_reg_1001;
reg [3:0] ret_V_8_reg_1028;
reg [1:0] ret_V_9_reg_869;
reg [4:0] select_ln1192_reg_968;
reg [1:0] select_ln340_reg_864;
reg [3:0] select_ln353_reg_1045;
reg [4:0] select_ln703_reg_1088;
reg [4:0] sext_ln703_reg_983;
reg [31:0] sext_ln831_reg_946;
reg tmp_2_reg_822;
reg tmp_3_reg_834;
reg [31:0] tmp_5_reg_1128;
reg [11:0] tmp_8_reg_936;
reg tmp_reg_1061;
reg [1:0] trunc_ln731_reg_828;
reg [1:0] trunc_ln851_1_reg_896;
reg [5:0] _428_;
wire [31:0] _000_;
wire [31:0] _001_;
wire [31:0] _002_;
wire [31:0] _003_;
wire [8:0] _004_;
wire [26:0] _005_;
wire _006_;
wire _007_;
wire _008_;
wire _009_;
wire _010_;
wire _011_;
wire [3:0] _012_;
wire [31:0] _013_;
wire [31:0] _014_;
wire [1:0] _015_;
wire [4:0] _016_;
wire [4:0] _017_;
wire [5:0] _018_;
wire [5:0] _019_;
wire [4:0] _020_;
wire [2:0] _021_;
wire [16:0] _022_;
wire [31:0] _023_;
wire [33:0] _024_;
wire [31:0] _025_;
wire [34:0] _026_;
wire [31:0] _027_;
wire [31:0] _028_;
wire [5:0] _029_;
wire [5:0] _030_;
wire [3:0] _031_;
wire [3:0] _032_;
wire [1:0] _033_;
wire [3:0] _034_;
wire [1:0] _035_;
wire [3:0] _036_;
wire [4:0] _037_;
wire [4:0] _038_;
wire [31:0] _039_;
wire _040_;
wire _041_;
wire [31:0] _042_;
wire [11:0] _043_;
wire _044_;
wire [1:0] _045_;
wire [1:0] _046_;
wire _047_;
wire _048_;
wire _049_;
wire _050_;
wire _051_;
wire _052_;
wire _053_;
wire [8:0] _054_;
wire [8:0] _055_;
wire _056_;
wire [7:0] _057_;
wire [8:0] _058_;
wire [9:0] _059_;
wire [15:0] _060_;
wire [15:0] _061_;
wire _062_;
wire [15:0] _063_;
wire [16:0] _064_;
wire [16:0] _065_;
wire [15:0] _066_;
wire [15:0] _067_;
wire _068_;
wire [15:0] _069_;
wire [16:0] _070_;
wire [16:0] _071_;
wire [15:0] _072_;
wire [15:0] _073_;
wire _074_;
wire [15:0] _075_;
wire [16:0] _076_;
wire [16:0] _077_;
wire [15:0] _078_;
wire [15:0] _079_;
wire _080_;
wire [15:0] _081_;
wire [16:0] _082_;
wire [16:0] _083_;
wire [15:0] _084_;
wire [15:0] _085_;
wire _086_;
wire [15:0] _087_;
wire [16:0] _088_;
wire [16:0] _089_;
wire [15:0] _090_;
wire [15:0] _091_;
wire _092_;
wire [15:0] _093_;
wire [16:0] _094_;
wire [16:0] _095_;
wire [16:0] _096_;
wire [16:0] _097_;
wire _098_;
wire [16:0] _099_;
wire [17:0] _100_;
wire [17:0] _101_;
wire [17:0] _102_;
wire [17:0] _103_;
wire _104_;
wire [16:0] _105_;
wire [17:0] _106_;
wire [18:0] _107_;
wire [17:0] _108_;
wire [17:0] _109_;
wire _110_;
wire [16:0] _111_;
wire [17:0] _112_;
wire [18:0] _113_;
wire [1:0] _114_;
wire [1:0] _115_;
wire _116_;
wire _117_;
wire [1:0] _118_;
wire [2:0] _119_;
wire [1:0] _120_;
wire [1:0] _121_;
wire _122_;
wire [1:0] _123_;
wire [2:0] _124_;
wire [2:0] _125_;
wire [2:0] _126_;
wire [2:0] _127_;
wire _128_;
wire [1:0] _129_;
wire [2:0] _130_;
wire [3:0] _131_;
wire [2:0] _132_;
wire [2:0] _133_;
wire _134_;
wire [1:0] _135_;
wire [2:0] _136_;
wire [3:0] _137_;
wire [2:0] _138_;
wire [2:0] _139_;
wire _140_;
wire [1:0] _141_;
wire [2:0] _142_;
wire [3:0] _143_;
wire [2:0] _144_;
wire [2:0] _145_;
wire _146_;
wire [2:0] _147_;
wire [3:0] _148_;
wire [3:0] _149_;
wire [4:0] _150_;
wire [4:0] _151_;
wire _152_;
wire [3:0] _153_;
wire [4:0] _154_;
wire [5:0] _155_;
wire _156_;
wire _157_;
wire _158_;
wire _159_;
wire _160_;
wire _161_;
wire _162_;
wire _163_;
wire _164_;
wire _165_;
wire _166_;
wire _167_;
wire _168_;
wire _169_;
wire _170_;
wire _171_;
wire _172_;
wire _173_;
wire _174_;
wire _175_;
wire _176_;
wire _177_;
wire _178_;
wire _179_;
wire _180_;
wire _181_;
wire _182_;
wire _183_;
wire _184_;
wire _185_;
wire _186_;
wire \add_17s_17s_17_2_1_U3.ce ;
wire \add_17s_17s_17_2_1_U3.clk ;
wire [16:0] \add_17s_17s_17_2_1_U3.din0 ;
wire [16:0] \add_17s_17s_17_2_1_U3.din1 ;
wire [16:0] \add_17s_17s_17_2_1_U3.dout ;
wire \add_17s_17s_17_2_1_U3.reset ;
wire [16:0] \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.a ;
wire [16:0] \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.ain_s0 ;
wire [16:0] \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.b ;
wire [16:0] \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.bin_s0 ;
wire \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.ce ;
wire \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.clk ;
wire \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.facout_s1 ;
wire \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.facout_s2 ;
wire [7:0] \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.fas_s1 ;
wire [8:0] \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.fas_s2 ;
wire \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.reset ;
wire [16:0] \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.s ;
wire [7:0] \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.u1.a ;
wire [7:0] \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.u1.b ;
wire \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.u1.cin ;
wire \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.u1.cout ;
wire [7:0] \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.u1.s ;
wire [8:0] \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.u2.a ;
wire [8:0] \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.u2.b ;
wire \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.u2.cin ;
wire \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.u2.cout ;
wire [8:0] \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.u2.s ;
wire \add_32ns_32ns_32_2_1_U10.ce ;
wire \add_32ns_32ns_32_2_1_U10.clk ;
wire [31:0] \add_32ns_32ns_32_2_1_U10.din0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U10.din1 ;
wire [31:0] \add_32ns_32ns_32_2_1_U10.dout ;
wire \add_32ns_32ns_32_2_1_U10.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.a ;
wire [31:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.b ;
wire [31:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s0 ;
wire \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.ce ;
wire \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.clk ;
wire \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s1 ;
wire \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s2 ;
wire [15:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s1 ;
wire [15:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s2 ;
wire \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.b ;
wire \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cin ;
wire \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.b ;
wire \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cin ;
wire \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.s ;
wire \add_32ns_32ns_32_2_1_U14.ce ;
wire \add_32ns_32ns_32_2_1_U14.clk ;
wire [31:0] \add_32ns_32ns_32_2_1_U14.din0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U14.din1 ;
wire [31:0] \add_32ns_32ns_32_2_1_U14.dout ;
wire \add_32ns_32ns_32_2_1_U14.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.a ;
wire [31:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.b ;
wire [31:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s0 ;
wire \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.ce ;
wire \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.clk ;
wire \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s1 ;
wire \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s2 ;
wire [15:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s1 ;
wire [15:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s2 ;
wire \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.b ;
wire \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cin ;
wire \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.b ;
wire \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cin ;
wire \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.s ;
wire \add_32ns_32ns_32_2_1_U17.ce ;
wire \add_32ns_32ns_32_2_1_U17.clk ;
wire [31:0] \add_32ns_32ns_32_2_1_U17.din0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U17.din1 ;
wire [31:0] \add_32ns_32ns_32_2_1_U17.dout ;
wire \add_32ns_32ns_32_2_1_U17.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.a ;
wire [31:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.b ;
wire [31:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s0 ;
wire \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.ce ;
wire \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.clk ;
wire \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s1 ;
wire \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s2 ;
wire [15:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s1 ;
wire [15:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s2 ;
wire \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.b ;
wire \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cin ;
wire \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.b ;
wire \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cin ;
wire \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.s ;
wire \add_32ns_32ns_32_2_1_U7.ce ;
wire \add_32ns_32ns_32_2_1_U7.clk ;
wire [31:0] \add_32ns_32ns_32_2_1_U7.din0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U7.din1 ;
wire [31:0] \add_32ns_32ns_32_2_1_U7.dout ;
wire \add_32ns_32ns_32_2_1_U7.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.a ;
wire [31:0] \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.b ;
wire [31:0] \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s0 ;
wire \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.ce ;
wire \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.clk ;
wire \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s1 ;
wire \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s2 ;
wire [15:0] \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s1 ;
wire [15:0] \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s2 ;
wire \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.b ;
wire \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cin ;
wire \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.b ;
wire \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cin ;
wire \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.s ;
wire \add_32s_32ns_32_2_1_U12.ce ;
wire \add_32s_32ns_32_2_1_U12.clk ;
wire [31:0] \add_32s_32ns_32_2_1_U12.din0 ;
wire [31:0] \add_32s_32ns_32_2_1_U12.din1 ;
wire [31:0] \add_32s_32ns_32_2_1_U12.dout ;
wire \add_32s_32ns_32_2_1_U12.reset ;
wire [31:0] \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.a ;
wire [31:0] \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.ain_s0 ;
wire [31:0] \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.b ;
wire [31:0] \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.bin_s0 ;
wire \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.ce ;
wire \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.clk ;
wire \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.facout_s1 ;
wire \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.facout_s2 ;
wire [15:0] \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.fas_s1 ;
wire [15:0] \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.fas_s2 ;
wire \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.reset ;
wire [31:0] \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.s ;
wire [15:0] \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.u1.a ;
wire [15:0] \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.u1.b ;
wire \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.u1.cin ;
wire \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.u1.cout ;
wire [15:0] \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.u1.s ;
wire [15:0] \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.u2.a ;
wire [15:0] \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.u2.b ;
wire \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.u2.cin ;
wire \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.u2.cout ;
wire [15:0] \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.u2.s ;
wire \add_32s_32ns_32_2_1_U4.ce ;
wire \add_32s_32ns_32_2_1_U4.clk ;
wire [31:0] \add_32s_32ns_32_2_1_U4.din0 ;
wire [31:0] \add_32s_32ns_32_2_1_U4.din1 ;
wire [31:0] \add_32s_32ns_32_2_1_U4.dout ;
wire \add_32s_32ns_32_2_1_U4.reset ;
wire [31:0] \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.a ;
wire [31:0] \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.ain_s0 ;
wire [31:0] \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.b ;
wire [31:0] \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.bin_s0 ;
wire \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.ce ;
wire \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.clk ;
wire \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.facout_s1 ;
wire \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.facout_s2 ;
wire [15:0] \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.fas_s1 ;
wire [15:0] \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.fas_s2 ;
wire \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.reset ;
wire [31:0] \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.s ;
wire [15:0] \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.u1.a ;
wire [15:0] \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.u1.b ;
wire \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.u1.cin ;
wire \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.u1.cout ;
wire [15:0] \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.u1.s ;
wire [15:0] \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.u2.a ;
wire [15:0] \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.u2.b ;
wire \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.u2.cin ;
wire \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.u2.cout ;
wire [15:0] \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.u2.s ;
wire \add_34s_34s_34_2_1_U9.ce ;
wire \add_34s_34s_34_2_1_U9.clk ;
wire [33:0] \add_34s_34s_34_2_1_U9.din0 ;
wire [33:0] \add_34s_34s_34_2_1_U9.din1 ;
wire [33:0] \add_34s_34s_34_2_1_U9.dout ;
wire \add_34s_34s_34_2_1_U9.reset ;
wire [33:0] \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.a ;
wire [33:0] \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.ain_s0 ;
wire [33:0] \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.b ;
wire [33:0] \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.bin_s0 ;
wire \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.ce ;
wire \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.clk ;
wire \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.facout_s1 ;
wire \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.facout_s2 ;
wire [16:0] \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.fas_s1 ;
wire [16:0] \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.fas_s2 ;
wire \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.reset ;
wire [33:0] \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.s ;
wire [16:0] \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.u1.a ;
wire [16:0] \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.u1.b ;
wire \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.u1.cin ;
wire \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.u1.cout ;
wire [16:0] \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.u1.s ;
wire [16:0] \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.u2.a ;
wire [16:0] \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.u2.b ;
wire \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.u2.cin ;
wire \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.u2.cout ;
wire [16:0] \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.u2.s ;
wire \add_35ns_35s_35_2_1_U15.ce ;
wire \add_35ns_35s_35_2_1_U15.clk ;
wire [34:0] \add_35ns_35s_35_2_1_U15.din0 ;
wire [34:0] \add_35ns_35s_35_2_1_U15.din1 ;
wire [34:0] \add_35ns_35s_35_2_1_U15.dout ;
wire \add_35ns_35s_35_2_1_U15.reset ;
wire [34:0] \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.a ;
wire [34:0] \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.ain_s0 ;
wire [34:0] \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.b ;
wire [34:0] \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.bin_s0 ;
wire \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.ce ;
wire \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.clk ;
wire \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.facout_s1 ;
wire \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.facout_s2 ;
wire [16:0] \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.fas_s1 ;
wire [17:0] \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.fas_s2 ;
wire \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.reset ;
wire [34:0] \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.s ;
wire [16:0] \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.u1.a ;
wire [16:0] \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.u1.b ;
wire \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.u1.cin ;
wire \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.u1.cout ;
wire [16:0] \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.u1.s ;
wire [17:0] \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.u2.a ;
wire [17:0] \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.u2.b ;
wire \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.u2.cin ;
wire \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.u2.cout ;
wire [17:0] \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.u2.s ;
wire \add_35s_35s_35_2_1_U16.ce ;
wire \add_35s_35s_35_2_1_U16.clk ;
wire [34:0] \add_35s_35s_35_2_1_U16.din0 ;
wire [34:0] \add_35s_35s_35_2_1_U16.din1 ;
wire [34:0] \add_35s_35s_35_2_1_U16.dout ;
wire \add_35s_35s_35_2_1_U16.reset ;
wire [34:0] \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.a ;
wire [34:0] \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.ain_s0 ;
wire [34:0] \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.b ;
wire [34:0] \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.bin_s0 ;
wire \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.ce ;
wire \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.clk ;
wire \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.facout_s1 ;
wire \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.facout_s2 ;
wire [16:0] \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.fas_s1 ;
wire [17:0] \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.fas_s2 ;
wire \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.reset ;
wire [34:0] \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.s ;
wire [16:0] \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.u1.a ;
wire [16:0] \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.u1.b ;
wire \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.u1.cin ;
wire \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.u1.cout ;
wire [16:0] \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.u1.s ;
wire [17:0] \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.u2.a ;
wire [17:0] \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.u2.b ;
wire \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.u2.cin ;
wire \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.u2.cout ;
wire [17:0] \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.u2.s ;
wire \add_3s_3s_3_2_1_U1.ce ;
wire \add_3s_3s_3_2_1_U1.clk ;
wire [2:0] \add_3s_3s_3_2_1_U1.din0 ;
wire [2:0] \add_3s_3s_3_2_1_U1.din1 ;
wire [2:0] \add_3s_3s_3_2_1_U1.dout ;
wire \add_3s_3s_3_2_1_U1.reset ;
wire [2:0] \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.a ;
wire [2:0] \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.ain_s0 ;
wire [2:0] \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.b ;
wire [2:0] \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.bin_s0 ;
wire \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.ce ;
wire \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.clk ;
wire \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.facout_s1 ;
wire \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.facout_s2 ;
wire \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.fas_s1 ;
wire [1:0] \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.fas_s2 ;
wire \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.reset ;
wire [2:0] \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.s ;
wire \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.u1.a ;
wire \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.u1.b ;
wire \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.u1.cin ;
wire \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.u1.cout ;
wire \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.u1.s ;
wire [1:0] \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.u2.a ;
wire [1:0] \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.u2.b ;
wire \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.u2.cin ;
wire \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.u2.cout ;
wire [1:0] \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.u2.s ;
wire \add_4ns_4ns_4_2_1_U8.ce ;
wire \add_4ns_4ns_4_2_1_U8.clk ;
wire [3:0] \add_4ns_4ns_4_2_1_U8.din0 ;
wire [3:0] \add_4ns_4ns_4_2_1_U8.din1 ;
wire [3:0] \add_4ns_4ns_4_2_1_U8.dout ;
wire \add_4ns_4ns_4_2_1_U8.reset ;
wire [3:0] \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.a ;
wire [3:0] \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.ain_s0 ;
wire [3:0] \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.b ;
wire [3:0] \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.bin_s0 ;
wire \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.ce ;
wire \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.clk ;
wire \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.facout_s1 ;
wire \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.facout_s2 ;
wire [1:0] \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.fas_s1 ;
wire [1:0] \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.fas_s2 ;
wire \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.reset ;
wire [3:0] \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.s ;
wire [1:0] \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.u1.a ;
wire [1:0] \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.u1.b ;
wire \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.u1.cin ;
wire \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.u1.cout ;
wire [1:0] \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.u1.s ;
wire [1:0] \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.u2.a ;
wire [1:0] \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.u2.b ;
wire \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.u2.cin ;
wire \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.u2.cout ;
wire [1:0] \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.u2.s ;
wire \add_5ns_5s_5_2_1_U11.ce ;
wire \add_5ns_5s_5_2_1_U11.clk ;
wire [4:0] \add_5ns_5s_5_2_1_U11.din0 ;
wire [4:0] \add_5ns_5s_5_2_1_U11.din1 ;
wire [4:0] \add_5ns_5s_5_2_1_U11.dout ;
wire \add_5ns_5s_5_2_1_U11.reset ;
wire [4:0] \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.a ;
wire [4:0] \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.ain_s0 ;
wire [4:0] \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.b ;
wire [4:0] \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.bin_s0 ;
wire \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.ce ;
wire \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.clk ;
wire \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.facout_s1 ;
wire \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.facout_s2 ;
wire [1:0] \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.fas_s1 ;
wire [2:0] \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.fas_s2 ;
wire \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.reset ;
wire [4:0] \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.s ;
wire [1:0] \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.u1.a ;
wire [1:0] \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.u1.b ;
wire \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.u1.cin ;
wire \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.u1.cout ;
wire [1:0] \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.u1.s ;
wire [2:0] \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.u2.a ;
wire [2:0] \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.u2.b ;
wire \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.u2.cin ;
wire \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.u2.cout ;
wire [2:0] \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.u2.s ;
wire \add_5ns_5s_5_2_1_U6.ce ;
wire \add_5ns_5s_5_2_1_U6.clk ;
wire [4:0] \add_5ns_5s_5_2_1_U6.din0 ;
wire [4:0] \add_5ns_5s_5_2_1_U6.din1 ;
wire [4:0] \add_5ns_5s_5_2_1_U6.dout ;
wire \add_5ns_5s_5_2_1_U6.reset ;
wire [4:0] \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.a ;
wire [4:0] \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.ain_s0 ;
wire [4:0] \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.b ;
wire [4:0] \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.bin_s0 ;
wire \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.ce ;
wire \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.clk ;
wire \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.facout_s1 ;
wire \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.facout_s2 ;
wire [1:0] \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.fas_s1 ;
wire [2:0] \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.fas_s2 ;
wire \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.reset ;
wire [4:0] \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.s ;
wire [1:0] \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.u1.a ;
wire [1:0] \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.u1.b ;
wire \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.u1.cin ;
wire \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.u1.cout ;
wire [1:0] \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.u1.s ;
wire [2:0] \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.u2.a ;
wire [2:0] \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.u2.b ;
wire \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.u2.cin ;
wire \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.u2.cout ;
wire [2:0] \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.u2.s ;
wire \add_5s_5ns_5_2_1_U13.ce ;
wire \add_5s_5ns_5_2_1_U13.clk ;
wire [4:0] \add_5s_5ns_5_2_1_U13.din0 ;
wire [4:0] \add_5s_5ns_5_2_1_U13.din1 ;
wire [4:0] \add_5s_5ns_5_2_1_U13.dout ;
wire \add_5s_5ns_5_2_1_U13.reset ;
wire [4:0] \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.a ;
wire [4:0] \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.ain_s0 ;
wire [4:0] \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.b ;
wire [4:0] \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.bin_s0 ;
wire \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.ce ;
wire \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.clk ;
wire \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.facout_s1 ;
wire \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.facout_s2 ;
wire [1:0] \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.fas_s1 ;
wire [2:0] \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.fas_s2 ;
wire \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.reset ;
wire [4:0] \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.s ;
wire [1:0] \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.u1.a ;
wire [1:0] \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.u1.b ;
wire \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.u1.cin ;
wire \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.u1.cout ;
wire [1:0] \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.u1.s ;
wire [2:0] \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.u2.a ;
wire [2:0] \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.u2.b ;
wire \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.u2.cin ;
wire \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.u2.cout ;
wire [2:0] \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.u2.s ;
wire \add_6ns_6ns_6_2_1_U2.ce ;
wire \add_6ns_6ns_6_2_1_U2.clk ;
wire [5:0] \add_6ns_6ns_6_2_1_U2.din0 ;
wire [5:0] \add_6ns_6ns_6_2_1_U2.din1 ;
wire [5:0] \add_6ns_6ns_6_2_1_U2.dout ;
wire \add_6ns_6ns_6_2_1_U2.reset ;
wire [5:0] \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.a ;
wire [5:0] \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.ain_s0 ;
wire [5:0] \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.b ;
wire [5:0] \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.bin_s0 ;
wire \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.ce ;
wire \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.clk ;
wire \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.facout_s1 ;
wire \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.facout_s2 ;
wire [2:0] \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.fas_s1 ;
wire [2:0] \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.fas_s2 ;
wire \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.reset ;
wire [5:0] \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.s ;
wire [2:0] \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.u1.a ;
wire [2:0] \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.u1.b ;
wire \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.u1.cin ;
wire \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.u1.cout ;
wire [2:0] \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.u1.s ;
wire [2:0] \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.u2.a ;
wire [2:0] \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.u2.b ;
wire \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.u2.cin ;
wire \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.u2.cout ;
wire [2:0] \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.u2.s ;
wire \add_9ns_9ns_9_2_1_U5.ce ;
wire \add_9ns_9ns_9_2_1_U5.clk ;
wire [8:0] \add_9ns_9ns_9_2_1_U5.din0 ;
wire [8:0] \add_9ns_9ns_9_2_1_U5.din1 ;
wire [8:0] \add_9ns_9ns_9_2_1_U5.dout ;
wire \add_9ns_9ns_9_2_1_U5.reset ;
wire [8:0] \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.a ;
wire [8:0] \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.ain_s0 ;
wire [8:0] \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.b ;
wire [8:0] \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.bin_s0 ;
wire \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.ce ;
wire \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.clk ;
wire \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.facout_s1 ;
wire \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.facout_s2 ;
wire [3:0] \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.fas_s1 ;
wire [4:0] \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.fas_s2 ;
wire \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.reset ;
wire [8:0] \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.s ;
wire [3:0] \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.u1.a ;
wire [3:0] \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.u1.b ;
wire \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.u1.cin ;
wire \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.u1.cout ;
wire [3:0] \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.u1.s ;
wire [4:0] \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.u2.a ;
wire [4:0] \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.u2.b ;
wire \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.u2.cin ;
wire \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.u2.cout ;
wire [4:0] \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.u2.s ;
wire and_ln340_1_fu_296_p2;
wire and_ln340_fu_301_p2;
wire and_ln785_fu_318_p2;
wire [3:0] and_ln_fu_255_p3;
wire ap_CS_fsm_state1;
wire ap_CS_fsm_state10;
wire ap_CS_fsm_state11;
wire ap_CS_fsm_state12;
wire ap_CS_fsm_state13;
wire ap_CS_fsm_state14;
wire ap_CS_fsm_state15;
wire ap_CS_fsm_state16;
wire ap_CS_fsm_state17;
wire ap_CS_fsm_state18;
wire ap_CS_fsm_state19;
wire ap_CS_fsm_state2;
wire ap_CS_fsm_state20;
wire ap_CS_fsm_state21;
wire ap_CS_fsm_state22;
wire ap_CS_fsm_state23;
wire ap_CS_fsm_state24;
wire ap_CS_fsm_state25;
wire ap_CS_fsm_state26;
wire ap_CS_fsm_state27;
wire ap_CS_fsm_state3;
wire ap_CS_fsm_state4;
wire ap_CS_fsm_state5;
wire ap_CS_fsm_state6;
wire ap_CS_fsm_state7;
wire ap_CS_fsm_state8;
wire ap_CS_fsm_state9;
wire [26:0] ap_NS_fsm;
wire ap_clk;
wire ap_done;
wire ap_idle;
wire ap_ready;
wire ap_rst;
wire ap_start;
wire [2:0] grp_fu_341_p0;
wire [2:0] grp_fu_341_p1;
wire [2:0] grp_fu_341_p2;
wire [5:0] grp_fu_384_p2;
wire [16:0] grp_fu_404_p0;
wire [16:0] grp_fu_404_p1;
wire [16:0] grp_fu_404_p2;
wire [31:0] grp_fu_452_p0;
wire [31:0] grp_fu_452_p2;
wire [8:0] grp_fu_469_p0;
wire [8:0] grp_fu_469_p1;
wire [8:0] grp_fu_469_p2;
wire [4:0] grp_fu_506_p1;
wire [4:0] grp_fu_506_p2;
wire [31:0] grp_fu_514_p0;
wire [31:0] grp_fu_514_p2;
wire [3:0] grp_fu_529_p2;
wire [33:0] grp_fu_549_p0;
wire [33:0] grp_fu_549_p1;
wire [33:0] grp_fu_549_p2;
wire [31:0] grp_fu_588_p2;
wire [4:0] grp_fu_620_p0;
wire [4:0] grp_fu_620_p2;
wire [31:0] grp_fu_629_p0;
wire [31:0] grp_fu_629_p2;
wire [4:0] grp_fu_708_p0;
wire [4:0] grp_fu_708_p2;
wire [31:0] grp_fu_713_p2;
wire [34:0] grp_fu_735_p0;
wire [34:0] grp_fu_735_p1;
wire [34:0] grp_fu_735_p2;
wire [34:0] grp_fu_766_p0;
wire [34:0] grp_fu_766_p1;
wire [34:0] grp_fu_766_p2;
wire [31:0] grp_fu_792_p2;
wire icmp_ln785_fu_270_p2;
wire icmp_ln786_1_fu_282_p2;
wire icmp_ln786_fu_276_p2;
wire icmp_ln851_1_fu_414_p2;
wire icmp_ln851_2_fu_776_p2;
wire icmp_ln851_fu_379_p2;
wire [5:0] lhs_fu_347_p3;
wire op_0;
wire [1:0] op_10;
wire [15:0] op_11;
wire [1:0] op_13;
wire [3:0] op_15;
wire [31:0] op_16;
wire [3:0] op_17;
wire [7:0] op_18_V_fu_717_p3;
wire [3:0] op_19;
wire [31:0] op_29;
wire op_29_ap_vld;
wire [3:0] op_3;
wire [3:0] op_4;
wire [3:0] op_5;
wire [7:0] op_9;
wire or_ln785_fu_322_p2;
wire or_ln786_1_fu_314_p2;
wire or_ln786_fu_287_p2;
wire [3:0] or_ln_fu_262_p4;
wire p_Result_1_fu_430_p3;
wire p_Result_2_fu_565_p3;
wire p_Result_3_fu_483_p3;
wire p_Result_4_fu_682_p3;
wire p_Result_5_fu_797_p3;
wire p_Result_s_fu_635_p3;
wire [3:0] r_fu_219_p2;
wire [4:0] ret_V_21_fu_600_p2;
wire ret_V_22_fu_657_p3;
wire [7:0] ret_V_23_fu_359_p2;
wire [7:0] ret_V_23_reg_884;
wire [5:0] ret_V_24_fu_442_p3;
wire [31:0] ret_V_29_fu_495_p3;
wire [31:0] ret_V_31_fu_698_p3;
wire [1:0] ret_V_9_fu_328_p3;
wire ret_V_fu_645_p2;
wire [32:0] rhs_5_fu_538_p3;
wire [33:0] rhs_8_fu_755_p3;
wire [4:0] rhs_fu_593_p3;
wire [4:0] select_ln1192_fu_475_p3;
wire [1:0] select_ln340_fu_307_p3;
wire [3:0] select_ln353_fu_581_p3;
wire [4:0] select_ln703_fu_674_p3;
wire [5:0] select_ln850_1_fu_437_p3;
wire [3:0] select_ln850_3_fu_575_p3;
wire [31:0] select_ln850_4_fu_490_p3;
wire [31:0] select_ln850_5_fu_692_p3;
wire [31:0] select_ln850_6_fu_804_p3;
wire select_ln850_fu_650_p3;
wire [15:0] sext_ln1192_1_fu_389_p0;
wire [7:0] sext_ln1194_fu_355_p1;
wire [7:0] sext_ln69_1_fu_458_p1;
wire [3:0] sext_ln703_2_fu_534_p0;
wire [3:0] sext_ln703_3_fu_751_p0;
wire [4:0] sext_ln703_fu_502_p1;
wire [31:0] sext_ln831_fu_449_p1;
wire [7:0] tmp_4_fu_393_p3;
wire [1:0] trunc_ln731_fu_233_p1;
wire [1:0] trunc_ln851_1_fu_375_p1;
wire trunc_ln851_2_fu_572_p1;
wire [15:0] trunc_ln851_3_fu_410_p0;
wire [4:0] trunc_ln851_3_fu_410_p1;
wire [3:0] trunc_ln851_4_fu_689_p0;
wire trunc_ln851_4_fu_689_p1;
wire [3:0] trunc_ln851_5_fu_772_p0;
wire [1:0] trunc_ln851_5_fu_772_p1;
wire trunc_ln851_fu_642_p1;
wire xor_ln340_1_fu_291_p2;


assign _047_ = icmp_ln851_2_reg_1143 & ap_CS_fsm[25];
assign _048_ = ap_CS_fsm[9] & icmp_ln851_1_reg_921;
assign _049_ = _051_ & ap_CS_fsm[0];
assign _050_ = ap_start & ap_CS_fsm[0];
assign and_ln340_1_fu_296_p2 = xor_ln340_1_fu_291_p2 & tmp_2_reg_822;
assign and_ln340_fu_301_p2 = or_ln786_1_fu_314_p2 & and_ln340_1_fu_296_p2;
assign and_ln785_fu_318_p2 = tmp_2_reg_822 & icmp_ln785_reg_846;
assign ret_V_23_fu_359_p2 = { op_5[3], op_5[3], op_5, 2'h0 } & op_9;
assign xor_ln340_1_fu_291_p2 = ~ icmp_ln785_reg_846;
assign ret_V_fu_645_p2 = ~ tmp_reg_1061;
assign r_fu_219_p2 = ~ op_4;
assign _051_ = ~ ap_start;
assign _052_ = ! { tmp_3_reg_834, 3'h0 };
assign _053_ = ! trunc_ln851_1_reg_896;
always @(posedge \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.clk )
\add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.bin_s1  <= _055_;
always @(posedge \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.clk )
\add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.ain_s1  <= _054_;
always @(posedge \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.clk )
\add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.sum_s1  <= _057_;
always @(posedge \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.clk )
\add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.carry_s1  <= _056_;
assign _055_ = \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.ce  ? \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.b [16:8] : \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.bin_s1 ;
assign _054_ = \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.ce  ? \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.a [16:8] : \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.ain_s1 ;
assign _056_ = \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.ce  ? \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.facout_s1  : \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.carry_s1 ;
assign _057_ = \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.ce  ? \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.fas_s1  : \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.sum_s1 ;
assign _058_ = \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.u1.a  + \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.u1.b ;
assign { \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.u1.cout , \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.u1.s  } = _058_ + \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.u1.cin ;
assign _059_ = \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.u2.a  + \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.u2.b ;
assign { \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.u2.cout , \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.u2.s  } = _059_ + \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.u2.cin ;
always @(posedge \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.clk )
\add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s1  <= _061_;
always @(posedge \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.clk )
\add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s1  <= _060_;
always @(posedge \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.clk )
\add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.sum_s1  <= _063_;
always @(posedge \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.clk )
\add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.carry_s1  <= _062_;
assign _061_ = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  ? \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.b [31:16] : \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s1 ;
assign _060_ = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  ? \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.a [31:16] : \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s1 ;
assign _062_ = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  ? \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s1  : \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.carry_s1 ;
assign _063_ = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  ? \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s1  : \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.sum_s1 ;
assign _064_ = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.a  + \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.b ;
assign { \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cout , \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.s  } = _064_ + \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cin ;
assign _065_ = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.a  + \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.b ;
assign { \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cout , \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.s  } = _065_ + \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cin ;
always @(posedge \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.clk )
\add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s1  <= _067_;
always @(posedge \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.clk )
\add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s1  <= _066_;
always @(posedge \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.clk )
\add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.sum_s1  <= _069_;
always @(posedge \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.clk )
\add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.carry_s1  <= _068_;
assign _067_ = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  ? \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.b [31:16] : \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s1 ;
assign _066_ = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  ? \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.a [31:16] : \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s1 ;
assign _068_ = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  ? \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s1  : \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.carry_s1 ;
assign _069_ = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  ? \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s1  : \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.sum_s1 ;
assign _070_ = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.a  + \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.b ;
assign { \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cout , \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.s  } = _070_ + \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cin ;
assign _071_ = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.a  + \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.b ;
assign { \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cout , \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.s  } = _071_ + \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cin ;
always @(posedge \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.clk )
\add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s1  <= _073_;
always @(posedge \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.clk )
\add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s1  <= _072_;
always @(posedge \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.clk )
\add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.sum_s1  <= _075_;
always @(posedge \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.clk )
\add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.carry_s1  <= _074_;
assign _073_ = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  ? \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.b [31:16] : \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s1 ;
assign _072_ = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  ? \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.a [31:16] : \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s1 ;
assign _074_ = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  ? \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s1  : \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.carry_s1 ;
assign _075_ = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  ? \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s1  : \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.sum_s1 ;
assign _076_ = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.a  + \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.b ;
assign { \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cout , \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.s  } = _076_ + \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cin ;
assign _077_ = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.a  + \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.b ;
assign { \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cout , \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.s  } = _077_ + \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cin ;
always @(posedge \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.clk )
\add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s1  <= _079_;
always @(posedge \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.clk )
\add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s1  <= _078_;
always @(posedge \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.clk )
\add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.sum_s1  <= _081_;
always @(posedge \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.clk )
\add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.carry_s1  <= _080_;
assign _079_ = \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  ? \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.b [31:16] : \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s1 ;
assign _078_ = \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  ? \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.a [31:16] : \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s1 ;
assign _080_ = \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  ? \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s1  : \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.carry_s1 ;
assign _081_ = \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  ? \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s1  : \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.sum_s1 ;
assign _082_ = \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.a  + \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.b ;
assign { \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cout , \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.s  } = _082_ + \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cin ;
assign _083_ = \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.a  + \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.b ;
assign { \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cout , \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.s  } = _083_ + \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cin ;
always @(posedge \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.clk )
\add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.bin_s1  <= _085_;
always @(posedge \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.clk )
\add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.ain_s1  <= _084_;
always @(posedge \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.clk )
\add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.sum_s1  <= _087_;
always @(posedge \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.clk )
\add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.carry_s1  <= _086_;
assign _085_ = \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.ce  ? \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.b [31:16] : \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.bin_s1 ;
assign _084_ = \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.ce  ? \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.a [31:16] : \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.ain_s1 ;
assign _086_ = \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.ce  ? \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.facout_s1  : \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.carry_s1 ;
assign _087_ = \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.ce  ? \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.fas_s1  : \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.sum_s1 ;
assign _088_ = \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.u1.a  + \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.u1.b ;
assign { \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.u1.cout , \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.u1.s  } = _088_ + \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.u1.cin ;
assign _089_ = \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.u2.a  + \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.u2.b ;
assign { \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.u2.cout , \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.u2.s  } = _089_ + \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.u2.cin ;
always @(posedge \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.clk )
\add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.bin_s1  <= _091_;
always @(posedge \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.clk )
\add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.ain_s1  <= _090_;
always @(posedge \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.clk )
\add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.sum_s1  <= _093_;
always @(posedge \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.clk )
\add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.carry_s1  <= _092_;
assign _091_ = \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.ce  ? \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.b [31:16] : \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.bin_s1 ;
assign _090_ = \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.ce  ? \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.a [31:16] : \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.ain_s1 ;
assign _092_ = \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.ce  ? \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.facout_s1  : \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.carry_s1 ;
assign _093_ = \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.ce  ? \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.fas_s1  : \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.sum_s1 ;
assign _094_ = \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.u1.a  + \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.u1.b ;
assign { \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.u1.cout , \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.u1.s  } = _094_ + \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.u1.cin ;
assign _095_ = \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.u2.a  + \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.u2.b ;
assign { \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.u2.cout , \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.u2.s  } = _095_ + \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.u2.cin ;
always @(posedge \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.clk )
\add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.bin_s1  <= _097_;
always @(posedge \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.clk )
\add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.ain_s1  <= _096_;
always @(posedge \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.clk )
\add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.sum_s1  <= _099_;
always @(posedge \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.clk )
\add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.carry_s1  <= _098_;
assign _097_ = \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.ce  ? \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.b [33:17] : \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.bin_s1 ;
assign _096_ = \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.ce  ? \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.a [33:17] : \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.ain_s1 ;
assign _098_ = \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.ce  ? \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.facout_s1  : \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.carry_s1 ;
assign _099_ = \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.ce  ? \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.fas_s1  : \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.sum_s1 ;
assign _100_ = \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.u1.a  + \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.u1.b ;
assign { \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.u1.cout , \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.u1.s  } = _100_ + \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.u1.cin ;
assign _101_ = \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.u2.a  + \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.u2.b ;
assign { \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.u2.cout , \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.u2.s  } = _101_ + \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.u2.cin ;
always @(posedge \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.clk )
\add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.bin_s1  <= _103_;
always @(posedge \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.clk )
\add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.ain_s1  <= _102_;
always @(posedge \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.clk )
\add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.sum_s1  <= _105_;
always @(posedge \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.clk )
\add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.carry_s1  <= _104_;
assign _103_ = \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.ce  ? \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.b [34:17] : \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.bin_s1 ;
assign _102_ = \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.ce  ? \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.a [34:17] : \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.ain_s1 ;
assign _104_ = \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.ce  ? \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.facout_s1  : \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.carry_s1 ;
assign _105_ = \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.ce  ? \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.fas_s1  : \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.sum_s1 ;
assign _106_ = \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.u1.a  + \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.u1.b ;
assign { \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.u1.cout , \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.u1.s  } = _106_ + \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.u1.cin ;
assign _107_ = \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.u2.a  + \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.u2.b ;
assign { \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.u2.cout , \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.u2.s  } = _107_ + \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.u2.cin ;
always @(posedge \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.clk )
\add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.bin_s1  <= _109_;
always @(posedge \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.clk )
\add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.ain_s1  <= _108_;
always @(posedge \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.clk )
\add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.sum_s1  <= _111_;
always @(posedge \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.clk )
\add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.carry_s1  <= _110_;
assign _109_ = \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.ce  ? \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.b [34:17] : \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.bin_s1 ;
assign _108_ = \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.ce  ? \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.a [34:17] : \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.ain_s1 ;
assign _110_ = \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.ce  ? \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.facout_s1  : \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.carry_s1 ;
assign _111_ = \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.ce  ? \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.fas_s1  : \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.sum_s1 ;
assign _112_ = \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.u1.a  + \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.u1.b ;
assign { \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.u1.cout , \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.u1.s  } = _112_ + \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.u1.cin ;
assign _113_ = \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.u2.a  + \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.u2.b ;
assign { \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.u2.cout , \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.u2.s  } = _113_ + \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.u2.cin ;
always @(posedge \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.clk )
\add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.bin_s1  <= _115_;
always @(posedge \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.clk )
\add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.ain_s1  <= _114_;
always @(posedge \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.clk )
\add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.sum_s1  <= _117_;
always @(posedge \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.clk )
\add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.carry_s1  <= _116_;
assign _115_ = \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.ce  ? \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.b [2:1] : \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.bin_s1 ;
assign _114_ = \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.ce  ? \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.a [2:1] : \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.ain_s1 ;
assign _116_ = \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.ce  ? \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.facout_s1  : \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.carry_s1 ;
assign _117_ = \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.ce  ? \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.fas_s1  : \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.sum_s1 ;
assign _118_ = \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.u1.a  + \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.u1.b ;
assign { \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.u1.cout , \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.u1.s  } = _118_ + \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.u1.cin ;
assign _119_ = \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.u2.a  + \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.u2.b ;
assign { \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.u2.cout , \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.u2.s  } = _119_ + \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.u2.cin ;
always @(posedge \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.clk )
\add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.bin_s1  <= _121_;
always @(posedge \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.clk )
\add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.ain_s1  <= _120_;
always @(posedge \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.clk )
\add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.sum_s1  <= _123_;
always @(posedge \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.clk )
\add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.carry_s1  <= _122_;
assign _121_ = \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.ce  ? \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.b [3:2] : \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.bin_s1 ;
assign _120_ = \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.ce  ? \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.a [3:2] : \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.ain_s1 ;
assign _122_ = \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.ce  ? \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.facout_s1  : \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.carry_s1 ;
assign _123_ = \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.ce  ? \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.fas_s1  : \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.sum_s1 ;
assign _124_ = \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.u1.a  + \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.u1.b ;
assign { \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.u1.cout , \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.u1.s  } = _124_ + \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.u1.cin ;
assign _125_ = \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.u2.a  + \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.u2.b ;
assign { \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.u2.cout , \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.u2.s  } = _125_ + \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.u2.cin ;
always @(posedge \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.clk )
\add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.bin_s1  <= _127_;
always @(posedge \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.clk )
\add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.ain_s1  <= _126_;
always @(posedge \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.clk )
\add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.sum_s1  <= _129_;
always @(posedge \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.clk )
\add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.carry_s1  <= _128_;
assign _127_ = \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.ce  ? \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.b [4:2] : \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.bin_s1 ;
assign _126_ = \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.ce  ? \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.a [4:2] : \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.ain_s1 ;
assign _128_ = \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.ce  ? \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.facout_s1  : \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.carry_s1 ;
assign _129_ = \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.ce  ? \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.fas_s1  : \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.sum_s1 ;
assign _130_ = \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.u1.a  + \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.u1.b ;
assign { \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.u1.cout , \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.u1.s  } = _130_ + \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.u1.cin ;
assign _131_ = \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.u2.a  + \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.u2.b ;
assign { \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.u2.cout , \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.u2.s  } = _131_ + \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.u2.cin ;
always @(posedge \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.clk )
\add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.bin_s1  <= _133_;
always @(posedge \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.clk )
\add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.ain_s1  <= _132_;
always @(posedge \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.clk )
\add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.sum_s1  <= _135_;
always @(posedge \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.clk )
\add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.carry_s1  <= _134_;
assign _133_ = \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.ce  ? \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.b [4:2] : \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.bin_s1 ;
assign _132_ = \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.ce  ? \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.a [4:2] : \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.ain_s1 ;
assign _134_ = \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.ce  ? \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.facout_s1  : \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.carry_s1 ;
assign _135_ = \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.ce  ? \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.fas_s1  : \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.sum_s1 ;
assign _136_ = \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.u1.a  + \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.u1.b ;
assign { \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.u1.cout , \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.u1.s  } = _136_ + \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.u1.cin ;
assign _137_ = \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.u2.a  + \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.u2.b ;
assign { \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.u2.cout , \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.u2.s  } = _137_ + \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.u2.cin ;
always @(posedge \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.clk )
\add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.bin_s1  <= _139_;
always @(posedge \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.clk )
\add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.ain_s1  <= _138_;
always @(posedge \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.clk )
\add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.sum_s1  <= _141_;
always @(posedge \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.clk )
\add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.carry_s1  <= _140_;
assign _139_ = \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.ce  ? \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.b [4:2] : \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.bin_s1 ;
assign _138_ = \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.ce  ? \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.a [4:2] : \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.ain_s1 ;
assign _140_ = \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.ce  ? \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.facout_s1  : \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.carry_s1 ;
assign _141_ = \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.ce  ? \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.fas_s1  : \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.sum_s1 ;
assign _142_ = \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.u1.a  + \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.u1.b ;
assign { \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.u1.cout , \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.u1.s  } = _142_ + \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.u1.cin ;
assign _143_ = \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.u2.a  + \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.u2.b ;
assign { \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.u2.cout , \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.u2.s  } = _143_ + \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.u2.cin ;
always @(posedge \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.clk )
\add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.bin_s1  <= _145_;
always @(posedge \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.clk )
\add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.ain_s1  <= _144_;
always @(posedge \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.clk )
\add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.sum_s1  <= _147_;
always @(posedge \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.clk )
\add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.carry_s1  <= _146_;
assign _145_ = \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.ce  ? \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.b [5:3] : \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.bin_s1 ;
assign _144_ = \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.ce  ? \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.a [5:3] : \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.ain_s1 ;
assign _146_ = \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.ce  ? \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.facout_s1  : \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.carry_s1 ;
assign _147_ = \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.ce  ? \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.fas_s1  : \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.sum_s1 ;
assign _148_ = \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.u1.a  + \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.u1.b ;
assign { \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.u1.cout , \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.u1.s  } = _148_ + \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.u1.cin ;
assign _149_ = \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.u2.a  + \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.u2.b ;
assign { \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.u2.cout , \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.u2.s  } = _149_ + \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.u2.cin ;
always @(posedge \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.clk )
\add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.bin_s1  <= _151_;
always @(posedge \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.clk )
\add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.ain_s1  <= _150_;
always @(posedge \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.clk )
\add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.sum_s1  <= _153_;
always @(posedge \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.clk )
\add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.carry_s1  <= _152_;
assign _151_ = \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.ce  ? \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.b [8:4] : \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.bin_s1 ;
assign _150_ = \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.ce  ? \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.a [8:4] : \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.ain_s1 ;
assign _152_ = \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.ce  ? \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.facout_s1  : \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.carry_s1 ;
assign _153_ = \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.ce  ? \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.fas_s1  : \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.sum_s1 ;
assign _154_ = \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.u1.a  + \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.u1.b ;
assign { \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.u1.cout , \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.u1.s  } = _154_ + \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.u1.cin ;
assign _155_ = \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.u2.a  + \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.u2.b ;
assign { \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.u2.cout , \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.u2.s  } = _155_ + \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.u2.cin ;
assign _156_ = | { tmp_3_reg_834, 1'h0, p_Result_s_16_reg_840 };
assign _157_ = p_Result_s_16_reg_840 != 2'h3;
assign _158_ = | op_11[4:0];
assign _159_ = | op_19[1:0];
assign or_ln785_fu_322_p2 = or_ln786_1_fu_314_p2 | and_ln785_fu_318_p2;
assign or_ln786_1_fu_314_p2 = icmp_ln786_reg_852 | icmp_ln786_1_reg_858;
always @(posedge ap_clk)
trunc_ln851_1_reg_896 <= 2'h0;
always @(posedge ap_clk)
select_ln1192_reg_968[0] <= 1'h0;
always @(posedge ap_clk)
tmp_5_reg_1128 <= _042_;
always @(posedge ap_clk)
sext_ln703_reg_983 <= _038_;
always @(posedge ap_clk)
select_ln353_reg_1045 <= _036_;
always @(posedge ap_clk)
select_ln340_reg_864 <= _035_;
always @(posedge ap_clk)
ret_V_9_reg_869 <= _033_;
always @(posedge ap_clk)
ret_V_32_reg_1148 <= _026_;
always @(posedge ap_clk)
ret_V_36_cast_reg_1153 <= _028_;
always @(posedge ap_clk)
ret_V_8_reg_1028 <= _032_;
always @(posedge ap_clk)
ret_V_30_reg_1033 <= _024_;
always @(posedge ap_clk)
ret_V_33_cast_reg_1038 <= _027_;
always @(posedge ap_clk)
ret_V_5_reg_926 <= _030_;
always @(posedge ap_clk)
ret_V_28_reg_931 <= _022_;
always @(posedge ap_clk)
tmp_8_reg_936 <= _043_;
always @(posedge ap_clk)
ret_V_24_reg_941 <= _019_;
always @(posedge ap_clk)
sext_ln831_reg_946 <= _039_;
always @(posedge ap_clk)
_428_ <= _018_;
assign ret_V_23_reg_884[7:2] = _428_;
always @(posedge ap_clk)
ret_V_3_reg_889 <= _029_;
always @(posedge ap_clk)
ret_V_27_reg_901 <= _021_;
always @(posedge ap_clk)
tmp_2_reg_822 <= _040_;
always @(posedge ap_clk)
trunc_ln731_reg_828 <= _045_;
always @(posedge ap_clk)
tmp_3_reg_834 <= _041_;
always @(posedge ap_clk)
p_Result_s_16_reg_840 <= _015_;
always @(posedge ap_clk)
ret_V_13_reg_1108 <= _016_;
always @(posedge ap_clk)
op_27_V_reg_1113 <= _014_;
always @(posedge ap_clk)
ret_V_25_reg_995 <= _020_;
always @(posedge ap_clk)
ret_V_8_cast_reg_1001 <= _031_;
always @(posedge ap_clk)
op_24_V_reg_1008 <= _013_;
always @(posedge ap_clk)
icmp_ln851_2_reg_1143 <= _010_;
always @(posedge ap_clk)
icmp_ln851_reg_906 <= _011_;
always @(posedge ap_clk)
icmp_ln851_1_reg_921 <= _009_;
always @(posedge ap_clk)
icmp_ln785_reg_846 <= _006_;
always @(posedge ap_clk)
icmp_ln786_reg_852 <= _008_;
always @(posedge ap_clk)
icmp_ln786_1_reg_858 <= _007_;
always @(posedge ap_clk)
select_ln1192_reg_968[4:1] <= _034_;
always @(posedge ap_clk)
ret_V_29_reg_973 <= _023_;
always @(posedge ap_clk)
add_ln69_reg_978 <= _004_;
always @(posedge ap_clk)
op_14_V_reg_1083 <= _012_;
always @(posedge ap_clk)
select_ln703_reg_1088 <= _037_;
always @(posedge ap_clk)
ret_V_31_reg_1093 <= _025_;
always @(posedge ap_clk)
add_ln69_2_reg_1098 <= _003_;
always @(posedge ap_clk)
add_ln691_reg_953 <= _002_;
always @(posedge ap_clk)
add_ln691_2_reg_1160 <= _001_;
always @(posedge ap_clk)
ret_V_21_reg_1055 <= _017_;
always @(posedge ap_clk)
tmp_reg_1061 <= _044_;
always @(posedge ap_clk)
add_ln691_1_reg_1073 <= _000_;
always @(posedge ap_clk)
ap_CS_fsm <= _005_;
assign _046_ = _050_ ? 2'h2 : 2'h1;
assign _160_ = ap_CS_fsm == 1'h1;
function [26:0] _461_;
input [26:0] a;
input [728:0] b;
input [26:0] s;
case (s)
27'b000000000000000000000000001:
_461_ = b[26:0];
27'b000000000000000000000000010:
_461_ = b[53:27];
27'b000000000000000000000000100:
_461_ = b[80:54];
27'b000000000000000000000001000:
_461_ = b[107:81];
27'b000000000000000000000010000:
_461_ = b[134:108];
27'b000000000000000000000100000:
_461_ = b[161:135];
27'b000000000000000000001000000:
_461_ = b[188:162];
27'b000000000000000000010000000:
_461_ = b[215:189];
27'b000000000000000000100000000:
_461_ = b[242:216];
27'b000000000000000001000000000:
_461_ = b[269:243];
27'b000000000000000010000000000:
_461_ = b[296:270];
27'b000000000000000100000000000:
_461_ = b[323:297];
27'b000000000000001000000000000:
_461_ = b[350:324];
27'b000000000000010000000000000:
_461_ = b[377:351];
27'b000000000000100000000000000:
_461_ = b[404:378];
27'b000000000001000000000000000:
_461_ = b[431:405];
27'b000000000010000000000000000:
_461_ = b[458:432];
27'b000000000100000000000000000:
_461_ = b[485:459];
27'b000000001000000000000000000:
_461_ = b[512:486];
27'b000000010000000000000000000:
_461_ = b[539:513];
27'b000000100000000000000000000:
_461_ = b[566:540];
27'b000001000000000000000000000:
_461_ = b[593:567];
27'b000010000000000000000000000:
_461_ = b[620:594];
27'b000100000000000000000000000:
_461_ = b[647:621];
27'b001000000000000000000000000:
_461_ = b[674:648];
27'b010000000000000000000000000:
_461_ = b[701:675];
27'b100000000000000000000000000:
_461_ = b[728:702];
27'b000000000000000000000000000:
_461_ = a;
default:
_461_ = 27'bx;
endcase
endfunction
assign ap_NS_fsm = _461_(27'hxxxxxxx, { 25'h0000000, _046_, 702'h00000020000008000002000000800000200000080000020000008000002000000800000200000080000020000008000002000000800000200000080000020000008000002000000800000200000080000020000000000001 }, { _160_, _186_, _185_, _184_, _183_, _182_, _181_, _180_, _179_, _178_, _177_, _176_, _175_, _174_, _173_, _172_, _171_, _170_, _169_, _168_, _167_, _166_, _165_, _164_, _163_, _162_, _161_ });
assign _161_ = ap_CS_fsm == 27'h4000000;
assign _162_ = ap_CS_fsm == 26'h2000000;
assign _163_ = ap_CS_fsm == 25'h1000000;
assign _164_ = ap_CS_fsm == 24'h800000;
assign _165_ = ap_CS_fsm == 23'h400000;
assign _166_ = ap_CS_fsm == 22'h200000;
assign _167_ = ap_CS_fsm == 21'h100000;
assign _168_ = ap_CS_fsm == 20'h80000;
assign _169_ = ap_CS_fsm == 19'h40000;
assign _170_ = ap_CS_fsm == 18'h20000;
assign _171_ = ap_CS_fsm == 17'h10000;
assign _172_ = ap_CS_fsm == 16'h8000;
assign _173_ = ap_CS_fsm == 15'h4000;
assign _174_ = ap_CS_fsm == 14'h2000;
assign _175_ = ap_CS_fsm == 13'h1000;
assign _176_ = ap_CS_fsm == 12'h800;
assign _177_ = ap_CS_fsm == 11'h400;
assign _178_ = ap_CS_fsm == 10'h200;
assign _179_ = ap_CS_fsm == 9'h100;
assign _180_ = ap_CS_fsm == 8'h80;
assign _181_ = ap_CS_fsm == 7'h40;
assign _182_ = ap_CS_fsm == 6'h20;
assign _183_ = ap_CS_fsm == 5'h10;
assign _184_ = ap_CS_fsm == 4'h8;
assign _185_ = ap_CS_fsm == 3'h4;
assign _186_ = ap_CS_fsm == 2'h2;
assign op_29_ap_vld = ap_CS_fsm[26] ? 1'h1 : 1'h0;
assign ap_idle = _049_ ? 1'h1 : 1'h0;
assign _042_ = ap_CS_fsm[21] ? grp_fu_735_p2[34:3] : tmp_5_reg_1128;
assign _038_ = ap_CS_fsm[11] ? { op_3[3], op_3 } : sext_ln703_reg_983;
assign _036_ = ap_CS_fsm[15] ? select_ln353_fu_581_p3 : select_ln353_reg_1045;
assign _035_ = ap_CS_fsm[2] ? select_ln340_fu_307_p3 : select_ln340_reg_864;
assign _033_ = ap_CS_fsm[3] ? ret_V_9_fu_328_p3 : ret_V_9_reg_869;
assign _028_ = ap_CS_fsm[23] ? grp_fu_766_p2[33:2] : ret_V_36_cast_reg_1153;
assign _026_ = ap_CS_fsm[23] ? grp_fu_766_p2 : ret_V_32_reg_1148;
assign _027_ = ap_CS_fsm[14] ? grp_fu_549_p2[32:1] : ret_V_33_cast_reg_1038;
assign _024_ = ap_CS_fsm[14] ? grp_fu_549_p2 : ret_V_30_reg_1033;
assign _032_ = ap_CS_fsm[14] ? grp_fu_529_p2 : ret_V_8_reg_1028;
assign _043_ = ap_CS_fsm[7] ? grp_fu_404_p2[16:5] : tmp_8_reg_936;
assign _022_ = ap_CS_fsm[7] ? grp_fu_404_p2 : ret_V_28_reg_931;
assign _030_ = ap_CS_fsm[7] ? grp_fu_384_p2 : ret_V_5_reg_926;
assign _039_ = ap_CS_fsm[8] ? { tmp_8_reg_936[11], tmp_8_reg_936[11], tmp_8_reg_936[11], tmp_8_reg_936[11], tmp_8_reg_936[11], tmp_8_reg_936[11], tmp_8_reg_936[11], tmp_8_reg_936[11], tmp_8_reg_936[11], tmp_8_reg_936[11], tmp_8_reg_936[11], tmp_8_reg_936[11], tmp_8_reg_936[11], tmp_8_reg_936[11], tmp_8_reg_936[11], tmp_8_reg_936[11], tmp_8_reg_936[11], tmp_8_reg_936[11], tmp_8_reg_936[11], tmp_8_reg_936[11], tmp_8_reg_936 } : sext_ln831_reg_946;
assign _019_ = ap_CS_fsm[8] ? ret_V_24_fu_442_p3 : ret_V_24_reg_941;
assign _021_ = ap_CS_fsm[5] ? grp_fu_341_p2 : ret_V_27_reg_901;
assign _029_ = ap_CS_fsm[5] ? ret_V_23_fu_359_p2[7:2] : ret_V_3_reg_889;
assign _018_ = ap_CS_fsm[5] ? ret_V_23_fu_359_p2[7:2] : ret_V_23_reg_884[7:2];
assign _015_ = ap_CS_fsm[0] ? r_fu_219_p2[3:2] : p_Result_s_16_reg_840;
assign _041_ = ap_CS_fsm[0] ? r_fu_219_p2[1] : tmp_3_reg_834;
assign _045_ = ap_CS_fsm[0] ? r_fu_219_p2[1:0] : trunc_ln731_reg_828;
assign _040_ = ap_CS_fsm[0] ? op_4[3] : tmp_2_reg_822;
assign _014_ = ap_CS_fsm[19] ? grp_fu_713_p2 : op_27_V_reg_1113;
assign _016_ = ap_CS_fsm[19] ? grp_fu_708_p2 : ret_V_13_reg_1108;
assign _013_ = ap_CS_fsm[12] ? grp_fu_514_p2 : op_24_V_reg_1008;
assign _031_ = ap_CS_fsm[12] ? grp_fu_506_p2[4:1] : ret_V_8_cast_reg_1001;
assign _020_ = ap_CS_fsm[12] ? grp_fu_506_p2 : ret_V_25_reg_995;
assign _010_ = ap_CS_fsm[22] ? icmp_ln851_2_fu_776_p2 : icmp_ln851_2_reg_1143;
assign _009_ = ap_CS_fsm[6] ? icmp_ln851_1_fu_414_p2 : icmp_ln851_1_reg_921;
assign _011_ = ap_CS_fsm[6] ? icmp_ln851_fu_379_p2 : icmp_ln851_reg_906;
assign _007_ = ap_CS_fsm[1] ? icmp_ln786_1_fu_282_p2 : icmp_ln786_1_reg_858;
assign _008_ = ap_CS_fsm[1] ? icmp_ln786_fu_276_p2 : icmp_ln786_reg_852;
assign _006_ = ap_CS_fsm[1] ? icmp_ln785_fu_270_p2 : icmp_ln785_reg_846;
assign _004_ = ap_CS_fsm[10] ? grp_fu_469_p2 : add_ln69_reg_978;
assign _023_ = ap_CS_fsm[10] ? ret_V_29_fu_495_p3 : ret_V_29_reg_973;
assign _034_ = ap_CS_fsm[10] ? select_ln1192_fu_475_p3[4:1] : select_ln1192_reg_968[4:1];
assign _003_ = ap_CS_fsm[17] ? grp_fu_629_p2 : add_ln69_2_reg_1098;
assign _025_ = ap_CS_fsm[17] ? ret_V_31_fu_698_p3 : ret_V_31_reg_1093;
assign _037_ = ap_CS_fsm[17] ? select_ln703_fu_674_p3 : select_ln703_reg_1088;
assign _012_ = ap_CS_fsm[17] ? grp_fu_620_p2[4:1] : op_14_V_reg_1083;
assign _002_ = _048_ ? grp_fu_452_p2 : add_ln691_reg_953;
assign _001_ = _047_ ? grp_fu_792_p2 : add_ln691_2_reg_1160;
assign _000_ = ap_CS_fsm[16] ? grp_fu_588_p2 : add_ln691_1_reg_1073;
assign _044_ = ap_CS_fsm[16] ? ret_V_21_fu_600_p2[1] : tmp_reg_1061;
assign _017_ = ap_CS_fsm[16] ? ret_V_21_fu_600_p2 : ret_V_21_reg_1055;
assign _005_ = ap_rst ? 27'h0000001 : ap_NS_fsm;
assign icmp_ln785_fu_270_p2 = _156_ ? 1'h1 : 1'h0;
assign icmp_ln786_1_fu_282_p2 = _157_ ? 1'h1 : 1'h0;
assign icmp_ln786_fu_276_p2 = _052_ ? 1'h1 : 1'h0;
assign icmp_ln851_1_fu_414_p2 = _158_ ? 1'h1 : 1'h0;
assign icmp_ln851_2_fu_776_p2 = _159_ ? 1'h1 : 1'h0;
assign icmp_ln851_fu_379_p2 = _053_ ? 1'h1 : 1'h0;
assign op_29 = ret_V_32_reg_1148[34] ? select_ln850_6_fu_804_p3 : ret_V_36_cast_reg_1153;
assign ret_V_22_fu_657_p3 = ret_V_21_reg_1055[4] ? select_ln850_fu_650_p3 : tmp_reg_1061;
assign ret_V_24_fu_442_p3 = ret_V_23_reg_884[7] ? select_ln850_1_fu_437_p3 : ret_V_3_reg_889;
assign ret_V_29_fu_495_p3 = ret_V_28_reg_931[16] ? select_ln850_4_fu_490_p3 : sext_ln831_reg_946;
assign ret_V_31_fu_698_p3 = ret_V_30_reg_1033[33] ? select_ln850_5_fu_692_p3 : ret_V_33_cast_reg_1038;
assign ret_V_9_fu_328_p3 = or_ln785_fu_322_p2 ? select_ln340_reg_864 : trunc_ln731_reg_828;
assign select_ln1192_fu_475_p3 = op_0 ? 5'h00 : 5'h1e;
assign select_ln340_fu_307_p3 = and_ln340_fu_301_p2 ? trunc_ln731_reg_828 : 2'h0;
assign select_ln353_fu_581_p3 = ret_V_25_reg_995[4] ? select_ln850_3_fu_575_p3 : ret_V_8_cast_reg_1001;
assign select_ln703_fu_674_p3 = ret_V_22_fu_657_p3 ? 5'h1f : 5'h00;
assign select_ln850_1_fu_437_p3 = icmp_ln851_reg_906 ? ret_V_3_reg_889 : ret_V_5_reg_926;
assign select_ln850_3_fu_575_p3 = ret_V_25_reg_995[0] ? ret_V_8_reg_1028 : ret_V_8_cast_reg_1001;
assign select_ln850_4_fu_490_p3 = icmp_ln851_1_reg_921 ? add_ln691_reg_953 : sext_ln831_reg_946;
assign select_ln850_5_fu_692_p3 = op_15[0] ? add_ln691_1_reg_1073 : ret_V_33_cast_reg_1038;
assign select_ln850_6_fu_804_p3 = icmp_ln851_2_reg_1143 ? add_ln691_2_reg_1160 : ret_V_36_cast_reg_1153;
assign select_ln850_fu_650_p3 = ret_V_21_reg_1055[0] ? ret_V_fu_645_p2 : tmp_reg_1061;
assign ret_V_21_fu_600_p2 = sext_ln703_reg_983 ^ { op_4, 1'h0 };
assign and_ln_fu_255_p3 = { tmp_3_reg_834, 3'h0 };
assign ap_CS_fsm_state1 = ap_CS_fsm[0];
assign ap_CS_fsm_state10 = ap_CS_fsm[9];
assign ap_CS_fsm_state11 = ap_CS_fsm[10];
assign ap_CS_fsm_state12 = ap_CS_fsm[11];
assign ap_CS_fsm_state13 = ap_CS_fsm[12];
assign ap_CS_fsm_state14 = ap_CS_fsm[13];
assign ap_CS_fsm_state15 = ap_CS_fsm[14];
assign ap_CS_fsm_state16 = ap_CS_fsm[15];
assign ap_CS_fsm_state17 = ap_CS_fsm[16];
assign ap_CS_fsm_state18 = ap_CS_fsm[17];
assign ap_CS_fsm_state19 = ap_CS_fsm[18];
assign ap_CS_fsm_state2 = ap_CS_fsm[1];
assign ap_CS_fsm_state20 = ap_CS_fsm[19];
assign ap_CS_fsm_state21 = ap_CS_fsm[20];
assign ap_CS_fsm_state22 = ap_CS_fsm[21];
assign ap_CS_fsm_state23 = ap_CS_fsm[22];
assign ap_CS_fsm_state24 = ap_CS_fsm[23];
assign ap_CS_fsm_state25 = ap_CS_fsm[24];
assign ap_CS_fsm_state26 = ap_CS_fsm[25];
assign ap_CS_fsm_state27 = ap_CS_fsm[26];
assign ap_CS_fsm_state3 = ap_CS_fsm[2];
assign ap_CS_fsm_state4 = ap_CS_fsm[3];
assign ap_CS_fsm_state5 = ap_CS_fsm[4];
assign ap_CS_fsm_state6 = ap_CS_fsm[5];
assign ap_CS_fsm_state7 = ap_CS_fsm[6];
assign ap_CS_fsm_state8 = ap_CS_fsm[7];
assign ap_CS_fsm_state9 = ap_CS_fsm[8];
assign ap_done = op_29_ap_vld;
assign ap_ready = op_29_ap_vld;
assign grp_fu_341_p0 = { ret_V_9_reg_869[1], ret_V_9_reg_869 };
assign grp_fu_341_p1 = { op_10[1], op_10 };
assign grp_fu_404_p0 = { ret_V_27_reg_901[2], ret_V_27_reg_901[2], ret_V_27_reg_901[2], ret_V_27_reg_901[2], ret_V_27_reg_901[2], ret_V_27_reg_901[2], ret_V_27_reg_901[2], ret_V_27_reg_901[2], ret_V_27_reg_901[2], ret_V_27_reg_901, 5'h00 };
assign grp_fu_404_p1 = { op_11[15], op_11 };
assign grp_fu_452_p0 = { tmp_8_reg_936[11], tmp_8_reg_936[11], tmp_8_reg_936[11], tmp_8_reg_936[11], tmp_8_reg_936[11], tmp_8_reg_936[11], tmp_8_reg_936[11], tmp_8_reg_936[11], tmp_8_reg_936[11], tmp_8_reg_936[11], tmp_8_reg_936[11], tmp_8_reg_936[11], tmp_8_reg_936[11], tmp_8_reg_936[11], tmp_8_reg_936[11], tmp_8_reg_936[11], tmp_8_reg_936[11], tmp_8_reg_936[11], tmp_8_reg_936[11], tmp_8_reg_936[11], tmp_8_reg_936 };
assign grp_fu_469_p0 = { 1'h0, ret_V_24_reg_941[5], ret_V_24_reg_941[5], ret_V_24_reg_941 };
assign grp_fu_469_p1 = { 7'h00, op_13 };
assign grp_fu_506_p1 = { op_3[3], op_3 };
assign grp_fu_514_p0 = { 23'h000000, add_ln69_reg_978 };
assign grp_fu_549_p0 = { op_24_V_reg_1008[31], op_24_V_reg_1008, 1'h0 };
assign grp_fu_549_p1 = { op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15 };
assign grp_fu_620_p0 = { select_ln353_reg_1045, 1'h0 };
assign grp_fu_629_p0 = { op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17 };
assign grp_fu_708_p0 = { op_14_V_reg_1083[3], op_14_V_reg_1083 };
assign grp_fu_735_p0 = { op_27_V_reg_1113, 3'h0 };
assign grp_fu_735_p1 = { ret_V_13_reg_1108[4], ret_V_13_reg_1108[4], ret_V_13_reg_1108[4], ret_V_13_reg_1108[4], ret_V_13_reg_1108[4], ret_V_13_reg_1108[4], ret_V_13_reg_1108[4], ret_V_13_reg_1108[4], ret_V_13_reg_1108[4], ret_V_13_reg_1108[4], ret_V_13_reg_1108[4], ret_V_13_reg_1108[4], ret_V_13_reg_1108[4], ret_V_13_reg_1108[4], ret_V_13_reg_1108[4], ret_V_13_reg_1108[4], ret_V_13_reg_1108[4], ret_V_13_reg_1108[4], ret_V_13_reg_1108[4], ret_V_13_reg_1108[4], ret_V_13_reg_1108[4], ret_V_13_reg_1108[4], ret_V_13_reg_1108[4], ret_V_13_reg_1108[4], ret_V_13_reg_1108[4], ret_V_13_reg_1108[4], ret_V_13_reg_1108[4], ret_V_13_reg_1108, 3'h0 };
assign grp_fu_766_p0 = { tmp_5_reg_1128[31], tmp_5_reg_1128, 2'h0 };
assign grp_fu_766_p1 = { op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19 };
assign lhs_fu_347_p3 = { op_5, 2'h0 };
assign op_18_V_fu_717_p3 = { ret_V_13_reg_1108, 3'h0 };
assign or_ln786_fu_287_p2 = or_ln786_1_fu_314_p2;
assign or_ln_fu_262_p4 = { tmp_3_reg_834, 1'h0, p_Result_s_16_reg_840 };
assign p_Result_1_fu_430_p3 = ret_V_23_reg_884[7];
assign p_Result_2_fu_565_p3 = ret_V_25_reg_995[4];
assign p_Result_3_fu_483_p3 = ret_V_28_reg_931[16];
assign p_Result_4_fu_682_p3 = ret_V_30_reg_1033[33];
assign p_Result_5_fu_797_p3 = ret_V_32_reg_1148[34];
assign p_Result_s_fu_635_p3 = ret_V_21_reg_1055[4];
assign rhs_5_fu_538_p3 = { op_24_V_reg_1008, 1'h0 };
assign rhs_8_fu_755_p3 = { tmp_5_reg_1128, 2'h0 };
assign rhs_fu_593_p3 = { op_4, 1'h0 };
assign sext_ln1192_1_fu_389_p0 = op_11;
assign sext_ln1194_fu_355_p1 = { op_5[3], op_5[3], op_5, 2'h0 };
assign sext_ln69_1_fu_458_p1 = { ret_V_24_reg_941[5], ret_V_24_reg_941[5], ret_V_24_reg_941 };
assign sext_ln703_2_fu_534_p0 = op_15;
assign sext_ln703_3_fu_751_p0 = op_19;
assign sext_ln703_fu_502_p1 = { op_3[3], op_3 };
assign sext_ln831_fu_449_p1 = { tmp_8_reg_936[11], tmp_8_reg_936[11], tmp_8_reg_936[11], tmp_8_reg_936[11], tmp_8_reg_936[11], tmp_8_reg_936[11], tmp_8_reg_936[11], tmp_8_reg_936[11], tmp_8_reg_936[11], tmp_8_reg_936[11], tmp_8_reg_936[11], tmp_8_reg_936[11], tmp_8_reg_936[11], tmp_8_reg_936[11], tmp_8_reg_936[11], tmp_8_reg_936[11], tmp_8_reg_936[11], tmp_8_reg_936[11], tmp_8_reg_936[11], tmp_8_reg_936[11], tmp_8_reg_936 };
assign tmp_4_fu_393_p3 = { ret_V_27_reg_901, 5'h00 };
assign trunc_ln731_fu_233_p1 = r_fu_219_p2[1:0];
assign trunc_ln851_1_fu_375_p1 = ret_V_23_fu_359_p2[1:0];
assign trunc_ln851_2_fu_572_p1 = ret_V_25_reg_995[0];
assign trunc_ln851_3_fu_410_p0 = op_11;
assign trunc_ln851_3_fu_410_p1 = op_11[4:0];
assign trunc_ln851_4_fu_689_p0 = op_15;
assign trunc_ln851_4_fu_689_p1 = op_15[0];
assign trunc_ln851_5_fu_772_p0 = op_19;
assign trunc_ln851_5_fu_772_p1 = op_19[1:0];
assign trunc_ln851_fu_642_p1 = ret_V_21_reg_1055[0];
assign \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.ain_s0  = \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.a ;
assign \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.bin_s0  = \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.b ;
assign \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.s  = { \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.fas_s2 , \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.sum_s1  };
assign \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.u2.a  = \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.ain_s1 ;
assign \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.u2.b  = \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.bin_s1 ;
assign \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.u2.cin  = \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.carry_s1 ;
assign \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.facout_s2  = \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.u2.cout ;
assign \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.fas_s2  = \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.u2.s ;
assign \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.u1.a  = \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.a [3:0];
assign \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.u1.b  = \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.b [3:0];
assign \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.u1.cin  = 1'h0;
assign \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.facout_s1  = \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.u1.cout ;
assign \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.fas_s1  = \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.u1.s ;
assign \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.a  = \add_9ns_9ns_9_2_1_U5.din0 ;
assign \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.b  = \add_9ns_9ns_9_2_1_U5.din1 ;
assign \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.ce  = \add_9ns_9ns_9_2_1_U5.ce ;
assign \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.clk  = \add_9ns_9ns_9_2_1_U5.clk ;
assign \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.reset  = \add_9ns_9ns_9_2_1_U5.reset ;
assign \add_9ns_9ns_9_2_1_U5.dout  = \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.s ;
assign \add_9ns_9ns_9_2_1_U5.ce  = 1'h1;
assign \add_9ns_9ns_9_2_1_U5.clk  = ap_clk;
assign \add_9ns_9ns_9_2_1_U5.din0  = { 1'h0, ret_V_24_reg_941[5], ret_V_24_reg_941[5], ret_V_24_reg_941 };
assign \add_9ns_9ns_9_2_1_U5.din1  = { 7'h00, op_13 };
assign grp_fu_469_p2 = \add_9ns_9ns_9_2_1_U5.dout ;
assign \add_9ns_9ns_9_2_1_U5.reset  = ap_rst;
assign \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.ain_s0  = \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.a ;
assign \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.bin_s0  = \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.b ;
assign \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.s  = { \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.fas_s2 , \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.sum_s1  };
assign \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.u2.a  = \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.ain_s1 ;
assign \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.u2.b  = \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.bin_s1 ;
assign \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.u2.cin  = \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.carry_s1 ;
assign \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.facout_s2  = \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.u2.cout ;
assign \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.fas_s2  = \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.u2.s ;
assign \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.u1.a  = \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.a [2:0];
assign \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.u1.b  = \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.b [2:0];
assign \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.u1.cin  = 1'h0;
assign \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.facout_s1  = \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.u1.cout ;
assign \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.fas_s1  = \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.u1.s ;
assign \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.a  = \add_6ns_6ns_6_2_1_U2.din0 ;
assign \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.b  = \add_6ns_6ns_6_2_1_U2.din1 ;
assign \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.ce  = \add_6ns_6ns_6_2_1_U2.ce ;
assign \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.clk  = \add_6ns_6ns_6_2_1_U2.clk ;
assign \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.reset  = \add_6ns_6ns_6_2_1_U2.reset ;
assign \add_6ns_6ns_6_2_1_U2.dout  = \add_6ns_6ns_6_2_1_U2.top_add_6ns_6ns_6_2_1_Adder_1_U.s ;
assign \add_6ns_6ns_6_2_1_U2.ce  = 1'h1;
assign \add_6ns_6ns_6_2_1_U2.clk  = ap_clk;
assign \add_6ns_6ns_6_2_1_U2.din0  = ret_V_3_reg_889;
assign \add_6ns_6ns_6_2_1_U2.din1  = 6'h01;
assign grp_fu_384_p2 = \add_6ns_6ns_6_2_1_U2.dout ;
assign \add_6ns_6ns_6_2_1_U2.reset  = ap_rst;
assign \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.ain_s0  = \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.a ;
assign \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.bin_s0  = \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.b ;
assign \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.s  = { \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.fas_s2 , \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.sum_s1  };
assign \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.u2.a  = \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.ain_s1 ;
assign \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.u2.b  = \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.bin_s1 ;
assign \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.u2.cin  = \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.carry_s1 ;
assign \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.facout_s2  = \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.u2.cout ;
assign \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.fas_s2  = \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.u2.s ;
assign \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.u1.a  = \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.a [1:0];
assign \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.u1.b  = \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.b [1:0];
assign \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.u1.cin  = 1'h0;
assign \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.facout_s1  = \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.u1.cout ;
assign \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.fas_s1  = \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.u1.s ;
assign \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.a  = \add_5s_5ns_5_2_1_U13.din0 ;
assign \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.b  = \add_5s_5ns_5_2_1_U13.din1 ;
assign \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.ce  = \add_5s_5ns_5_2_1_U13.ce ;
assign \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.clk  = \add_5s_5ns_5_2_1_U13.clk ;
assign \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.reset  = \add_5s_5ns_5_2_1_U13.reset ;
assign \add_5s_5ns_5_2_1_U13.dout  = \add_5s_5ns_5_2_1_U13.top_add_5s_5ns_5_2_1_Adder_9_U.s ;
assign \add_5s_5ns_5_2_1_U13.ce  = 1'h1;
assign \add_5s_5ns_5_2_1_U13.clk  = ap_clk;
assign \add_5s_5ns_5_2_1_U13.din0  = { op_14_V_reg_1083[3], op_14_V_reg_1083 };
assign \add_5s_5ns_5_2_1_U13.din1  = select_ln703_reg_1088;
assign grp_fu_708_p2 = \add_5s_5ns_5_2_1_U13.dout ;
assign \add_5s_5ns_5_2_1_U13.reset  = ap_rst;
assign \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.ain_s0  = \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.a ;
assign \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.bin_s0  = \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.b ;
assign \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.s  = { \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.fas_s2 , \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.sum_s1  };
assign \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.u2.a  = \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.ain_s1 ;
assign \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.u2.b  = \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.bin_s1 ;
assign \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.u2.cin  = \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.carry_s1 ;
assign \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.facout_s2  = \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.u2.cout ;
assign \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.fas_s2  = \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.u2.s ;
assign \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.u1.a  = \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.a [1:0];
assign \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.u1.b  = \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.b [1:0];
assign \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.u1.cin  = 1'h0;
assign \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.facout_s1  = \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.u1.cout ;
assign \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.fas_s1  = \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.u1.s ;
assign \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.a  = \add_5ns_5s_5_2_1_U6.din0 ;
assign \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.b  = \add_5ns_5s_5_2_1_U6.din1 ;
assign \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.ce  = \add_5ns_5s_5_2_1_U6.ce ;
assign \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.clk  = \add_5ns_5s_5_2_1_U6.clk ;
assign \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.reset  = \add_5ns_5s_5_2_1_U6.reset ;
assign \add_5ns_5s_5_2_1_U6.dout  = \add_5ns_5s_5_2_1_U6.top_add_5ns_5s_5_2_1_Adder_5_U.s ;
assign \add_5ns_5s_5_2_1_U6.ce  = 1'h1;
assign \add_5ns_5s_5_2_1_U6.clk  = ap_clk;
assign \add_5ns_5s_5_2_1_U6.din0  = select_ln1192_reg_968;
assign \add_5ns_5s_5_2_1_U6.din1  = { op_3[3], op_3 };
assign grp_fu_506_p2 = \add_5ns_5s_5_2_1_U6.dout ;
assign \add_5ns_5s_5_2_1_U6.reset  = ap_rst;
assign \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.ain_s0  = \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.a ;
assign \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.bin_s0  = \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.b ;
assign \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.s  = { \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.fas_s2 , \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.sum_s1  };
assign \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.u2.a  = \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.ain_s1 ;
assign \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.u2.b  = \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.bin_s1 ;
assign \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.u2.cin  = \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.carry_s1 ;
assign \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.facout_s2  = \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.u2.cout ;
assign \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.fas_s2  = \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.u2.s ;
assign \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.u1.a  = \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.a [1:0];
assign \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.u1.b  = \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.b [1:0];
assign \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.u1.cin  = 1'h0;
assign \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.facout_s1  = \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.u1.cout ;
assign \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.fas_s1  = \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.u1.s ;
assign \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.a  = \add_5ns_5s_5_2_1_U11.din0 ;
assign \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.b  = \add_5ns_5s_5_2_1_U11.din1 ;
assign \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.ce  = \add_5ns_5s_5_2_1_U11.ce ;
assign \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.clk  = \add_5ns_5s_5_2_1_U11.clk ;
assign \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.reset  = \add_5ns_5s_5_2_1_U11.reset ;
assign \add_5ns_5s_5_2_1_U11.dout  = \add_5ns_5s_5_2_1_U11.top_add_5ns_5s_5_2_1_Adder_5_U.s ;
assign \add_5ns_5s_5_2_1_U11.ce  = 1'h1;
assign \add_5ns_5s_5_2_1_U11.clk  = ap_clk;
assign \add_5ns_5s_5_2_1_U11.din0  = { select_ln353_reg_1045, 1'h0 };
assign \add_5ns_5s_5_2_1_U11.din1  = sext_ln703_reg_983;
assign grp_fu_620_p2 = \add_5ns_5s_5_2_1_U11.dout ;
assign \add_5ns_5s_5_2_1_U11.reset  = ap_rst;
assign \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.ain_s0  = \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.a ;
assign \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.bin_s0  = \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.b ;
assign \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.s  = { \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.fas_s2 , \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.sum_s1  };
assign \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.u2.a  = \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.ain_s1 ;
assign \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.u2.b  = \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.bin_s1 ;
assign \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.u2.cin  = \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.carry_s1 ;
assign \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.facout_s2  = \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.u2.cout ;
assign \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.fas_s2  = \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.u2.s ;
assign \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.u1.a  = \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.a [1:0];
assign \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.u1.b  = \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.b [1:0];
assign \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.u1.cin  = 1'h0;
assign \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.facout_s1  = \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.u1.cout ;
assign \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.fas_s1  = \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.u1.s ;
assign \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.a  = \add_4ns_4ns_4_2_1_U8.din0 ;
assign \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.b  = \add_4ns_4ns_4_2_1_U8.din1 ;
assign \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.ce  = \add_4ns_4ns_4_2_1_U8.ce ;
assign \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.clk  = \add_4ns_4ns_4_2_1_U8.clk ;
assign \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.reset  = \add_4ns_4ns_4_2_1_U8.reset ;
assign \add_4ns_4ns_4_2_1_U8.dout  = \add_4ns_4ns_4_2_1_U8.top_add_4ns_4ns_4_2_1_Adder_7_U.s ;
assign \add_4ns_4ns_4_2_1_U8.ce  = 1'h1;
assign \add_4ns_4ns_4_2_1_U8.clk  = ap_clk;
assign \add_4ns_4ns_4_2_1_U8.din0  = ret_V_8_cast_reg_1001;
assign \add_4ns_4ns_4_2_1_U8.din1  = 4'h1;
assign grp_fu_529_p2 = \add_4ns_4ns_4_2_1_U8.dout ;
assign \add_4ns_4ns_4_2_1_U8.reset  = ap_rst;
assign \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.ain_s0  = \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.a ;
assign \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.bin_s0  = \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.b ;
assign \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.s  = { \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.fas_s2 , \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.sum_s1  };
assign \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.u2.a  = \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.ain_s1 ;
assign \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.u2.b  = \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.bin_s1 ;
assign \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.u2.cin  = \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.carry_s1 ;
assign \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.facout_s2  = \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.u2.cout ;
assign \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.fas_s2  = \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.u2.s ;
assign \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.u1.a  = \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.a [0];
assign \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.u1.b  = \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.b [0];
assign \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.u1.cin  = 1'h0;
assign \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.facout_s1  = \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.u1.cout ;
assign \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.fas_s1  = \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.u1.s ;
assign \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.a  = \add_3s_3s_3_2_1_U1.din0 ;
assign \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.b  = \add_3s_3s_3_2_1_U1.din1 ;
assign \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.ce  = \add_3s_3s_3_2_1_U1.ce ;
assign \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.clk  = \add_3s_3s_3_2_1_U1.clk ;
assign \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.reset  = \add_3s_3s_3_2_1_U1.reset ;
assign \add_3s_3s_3_2_1_U1.dout  = \add_3s_3s_3_2_1_U1.top_add_3s_3s_3_2_1_Adder_0_U.s ;
assign \add_3s_3s_3_2_1_U1.ce  = 1'h1;
assign \add_3s_3s_3_2_1_U1.clk  = ap_clk;
assign \add_3s_3s_3_2_1_U1.din0  = { ret_V_9_reg_869[1], ret_V_9_reg_869 };
assign \add_3s_3s_3_2_1_U1.din1  = { op_10[1], op_10 };
assign grp_fu_341_p2 = \add_3s_3s_3_2_1_U1.dout ;
assign \add_3s_3s_3_2_1_U1.reset  = ap_rst;
assign \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.ain_s0  = \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.a ;
assign \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.bin_s0  = \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.b ;
assign \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.s  = { \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.fas_s2 , \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.sum_s1  };
assign \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.u2.a  = \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.ain_s1 ;
assign \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.u2.b  = \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.bin_s1 ;
assign \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.u2.cin  = \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.carry_s1 ;
assign \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.facout_s2  = \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.u2.cout ;
assign \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.fas_s2  = \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.u2.s ;
assign \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.u1.a  = \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.a [16:0];
assign \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.u1.b  = \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.b [16:0];
assign \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.u1.cin  = 1'h0;
assign \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.facout_s1  = \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.u1.cout ;
assign \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.fas_s1  = \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.u1.s ;
assign \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.a  = \add_35s_35s_35_2_1_U16.din0 ;
assign \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.b  = \add_35s_35s_35_2_1_U16.din1 ;
assign \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.ce  = \add_35s_35s_35_2_1_U16.ce ;
assign \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.clk  = \add_35s_35s_35_2_1_U16.clk ;
assign \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.reset  = \add_35s_35s_35_2_1_U16.reset ;
assign \add_35s_35s_35_2_1_U16.dout  = \add_35s_35s_35_2_1_U16.top_add_35s_35s_35_2_1_Adder_11_U.s ;
assign \add_35s_35s_35_2_1_U16.ce  = 1'h1;
assign \add_35s_35s_35_2_1_U16.clk  = ap_clk;
assign \add_35s_35s_35_2_1_U16.din0  = { tmp_5_reg_1128[31], tmp_5_reg_1128, 2'h0 };
assign \add_35s_35s_35_2_1_U16.din1  = { op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19[3], op_19 };
assign grp_fu_766_p2 = \add_35s_35s_35_2_1_U16.dout ;
assign \add_35s_35s_35_2_1_U16.reset  = ap_rst;
assign \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.ain_s0  = \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.a ;
assign \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.bin_s0  = \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.b ;
assign \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.s  = { \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.fas_s2 , \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.sum_s1  };
assign \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.u2.a  = \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.ain_s1 ;
assign \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.u2.b  = \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.bin_s1 ;
assign \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.u2.cin  = \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.carry_s1 ;
assign \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.facout_s2  = \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.u2.cout ;
assign \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.fas_s2  = \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.u2.s ;
assign \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.u1.a  = \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.a [16:0];
assign \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.u1.b  = \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.b [16:0];
assign \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.u1.cin  = 1'h0;
assign \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.facout_s1  = \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.u1.cout ;
assign \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.fas_s1  = \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.u1.s ;
assign \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.a  = \add_35ns_35s_35_2_1_U15.din0 ;
assign \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.b  = \add_35ns_35s_35_2_1_U15.din1 ;
assign \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.ce  = \add_35ns_35s_35_2_1_U15.ce ;
assign \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.clk  = \add_35ns_35s_35_2_1_U15.clk ;
assign \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.reset  = \add_35ns_35s_35_2_1_U15.reset ;
assign \add_35ns_35s_35_2_1_U15.dout  = \add_35ns_35s_35_2_1_U15.top_add_35ns_35s_35_2_1_Adder_10_U.s ;
assign \add_35ns_35s_35_2_1_U15.ce  = 1'h1;
assign \add_35ns_35s_35_2_1_U15.clk  = ap_clk;
assign \add_35ns_35s_35_2_1_U15.din0  = { op_27_V_reg_1113, 3'h0 };
assign \add_35ns_35s_35_2_1_U15.din1  = { ret_V_13_reg_1108[4], ret_V_13_reg_1108[4], ret_V_13_reg_1108[4], ret_V_13_reg_1108[4], ret_V_13_reg_1108[4], ret_V_13_reg_1108[4], ret_V_13_reg_1108[4], ret_V_13_reg_1108[4], ret_V_13_reg_1108[4], ret_V_13_reg_1108[4], ret_V_13_reg_1108[4], ret_V_13_reg_1108[4], ret_V_13_reg_1108[4], ret_V_13_reg_1108[4], ret_V_13_reg_1108[4], ret_V_13_reg_1108[4], ret_V_13_reg_1108[4], ret_V_13_reg_1108[4], ret_V_13_reg_1108[4], ret_V_13_reg_1108[4], ret_V_13_reg_1108[4], ret_V_13_reg_1108[4], ret_V_13_reg_1108[4], ret_V_13_reg_1108[4], ret_V_13_reg_1108[4], ret_V_13_reg_1108[4], ret_V_13_reg_1108[4], ret_V_13_reg_1108, 3'h0 };
assign grp_fu_735_p2 = \add_35ns_35s_35_2_1_U15.dout ;
assign \add_35ns_35s_35_2_1_U15.reset  = ap_rst;
assign \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.ain_s0  = \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.a ;
assign \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.bin_s0  = \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.b ;
assign \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.s  = { \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.fas_s2 , \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.sum_s1  };
assign \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.u2.a  = \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.ain_s1 ;
assign \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.u2.b  = \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.bin_s1 ;
assign \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.u2.cin  = \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.carry_s1 ;
assign \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.facout_s2  = \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.u2.cout ;
assign \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.fas_s2  = \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.u2.s ;
assign \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.u1.a  = \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.a [16:0];
assign \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.u1.b  = \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.b [16:0];
assign \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.u1.cin  = 1'h0;
assign \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.facout_s1  = \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.u1.cout ;
assign \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.fas_s1  = \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.u1.s ;
assign \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.a  = \add_34s_34s_34_2_1_U9.din0 ;
assign \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.b  = \add_34s_34s_34_2_1_U9.din1 ;
assign \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.ce  = \add_34s_34s_34_2_1_U9.ce ;
assign \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.clk  = \add_34s_34s_34_2_1_U9.clk ;
assign \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.reset  = \add_34s_34s_34_2_1_U9.reset ;
assign \add_34s_34s_34_2_1_U9.dout  = \add_34s_34s_34_2_1_U9.top_add_34s_34s_34_2_1_Adder_8_U.s ;
assign \add_34s_34s_34_2_1_U9.ce  = 1'h1;
assign \add_34s_34s_34_2_1_U9.clk  = ap_clk;
assign \add_34s_34s_34_2_1_U9.din0  = { op_24_V_reg_1008[31], op_24_V_reg_1008, 1'h0 };
assign \add_34s_34s_34_2_1_U9.din1  = { op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15 };
assign grp_fu_549_p2 = \add_34s_34s_34_2_1_U9.dout ;
assign \add_34s_34s_34_2_1_U9.reset  = ap_rst;
assign \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.ain_s0  = \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.a ;
assign \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.bin_s0  = \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.b ;
assign \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.s  = { \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.fas_s2 , \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.sum_s1  };
assign \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.u2.a  = \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.ain_s1 ;
assign \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.u2.b  = \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.bin_s1 ;
assign \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.u2.cin  = \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.carry_s1 ;
assign \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.facout_s2  = \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.u2.cout ;
assign \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.fas_s2  = \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.u2.s ;
assign \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.u1.a  = \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.a [15:0];
assign \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.u1.b  = \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.b [15:0];
assign \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.u1.cin  = 1'h0;
assign \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.facout_s1  = \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.u1.cout ;
assign \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.fas_s1  = \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.u1.s ;
assign \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.a  = \add_32s_32ns_32_2_1_U4.din0 ;
assign \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.b  = \add_32s_32ns_32_2_1_U4.din1 ;
assign \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.ce  = \add_32s_32ns_32_2_1_U4.ce ;
assign \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.clk  = \add_32s_32ns_32_2_1_U4.clk ;
assign \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.reset  = \add_32s_32ns_32_2_1_U4.reset ;
assign \add_32s_32ns_32_2_1_U4.dout  = \add_32s_32ns_32_2_1_U4.top_add_32s_32ns_32_2_1_Adder_3_U.s ;
assign \add_32s_32ns_32_2_1_U4.ce  = 1'h1;
assign \add_32s_32ns_32_2_1_U4.clk  = ap_clk;
assign \add_32s_32ns_32_2_1_U4.din0  = { tmp_8_reg_936[11], tmp_8_reg_936[11], tmp_8_reg_936[11], tmp_8_reg_936[11], tmp_8_reg_936[11], tmp_8_reg_936[11], tmp_8_reg_936[11], tmp_8_reg_936[11], tmp_8_reg_936[11], tmp_8_reg_936[11], tmp_8_reg_936[11], tmp_8_reg_936[11], tmp_8_reg_936[11], tmp_8_reg_936[11], tmp_8_reg_936[11], tmp_8_reg_936[11], tmp_8_reg_936[11], tmp_8_reg_936[11], tmp_8_reg_936[11], tmp_8_reg_936[11], tmp_8_reg_936 };
assign \add_32s_32ns_32_2_1_U4.din1  = 32'd1;
assign grp_fu_452_p2 = \add_32s_32ns_32_2_1_U4.dout ;
assign \add_32s_32ns_32_2_1_U4.reset  = ap_rst;
assign \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.ain_s0  = \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.a ;
assign \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.bin_s0  = \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.b ;
assign \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.s  = { \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.fas_s2 , \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.sum_s1  };
assign \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.u2.a  = \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.ain_s1 ;
assign \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.u2.b  = \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.bin_s1 ;
assign \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.u2.cin  = \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.carry_s1 ;
assign \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.facout_s2  = \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.u2.cout ;
assign \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.fas_s2  = \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.u2.s ;
assign \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.u1.a  = \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.a [15:0];
assign \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.u1.b  = \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.b [15:0];
assign \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.u1.cin  = 1'h0;
assign \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.facout_s1  = \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.u1.cout ;
assign \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.fas_s1  = \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.u1.s ;
assign \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.a  = \add_32s_32ns_32_2_1_U12.din0 ;
assign \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.b  = \add_32s_32ns_32_2_1_U12.din1 ;
assign \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.ce  = \add_32s_32ns_32_2_1_U12.ce ;
assign \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.clk  = \add_32s_32ns_32_2_1_U12.clk ;
assign \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.reset  = \add_32s_32ns_32_2_1_U12.reset ;
assign \add_32s_32ns_32_2_1_U12.dout  = \add_32s_32ns_32_2_1_U12.top_add_32s_32ns_32_2_1_Adder_3_U.s ;
assign \add_32s_32ns_32_2_1_U12.ce  = 1'h1;
assign \add_32s_32ns_32_2_1_U12.clk  = ap_clk;
assign \add_32s_32ns_32_2_1_U12.din0  = { op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17[3], op_17 };
assign \add_32s_32ns_32_2_1_U12.din1  = op_16;
assign grp_fu_629_p2 = \add_32s_32ns_32_2_1_U12.dout ;
assign \add_32s_32ns_32_2_1_U12.reset  = ap_rst;
assign \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s0  = \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.a ;
assign \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s0  = \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.b ;
assign \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.s  = { \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s2 , \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.sum_s1  };
assign \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.a  = \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s1 ;
assign \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.b  = \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s1 ;
assign \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cin  = \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.carry_s1 ;
assign \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s2  = \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cout ;
assign \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s2  = \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.s ;
assign \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.a  = \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.a [15:0];
assign \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.b  = \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.b [15:0];
assign \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cin  = 1'h0;
assign \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s1  = \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cout ;
assign \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s1  = \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.s ;
assign \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.a  = \add_32ns_32ns_32_2_1_U7.din0 ;
assign \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.b  = \add_32ns_32ns_32_2_1_U7.din1 ;
assign \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  = \add_32ns_32ns_32_2_1_U7.ce ;
assign \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.clk  = \add_32ns_32ns_32_2_1_U7.clk ;
assign \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.reset  = \add_32ns_32ns_32_2_1_U7.reset ;
assign \add_32ns_32ns_32_2_1_U7.dout  = \add_32ns_32ns_32_2_1_U7.top_add_32ns_32ns_32_2_1_Adder_6_U.s ;
assign \add_32ns_32ns_32_2_1_U7.ce  = 1'h1;
assign \add_32ns_32ns_32_2_1_U7.clk  = ap_clk;
assign \add_32ns_32ns_32_2_1_U7.din0  = { 23'h000000, add_ln69_reg_978 };
assign \add_32ns_32ns_32_2_1_U7.din1  = ret_V_29_reg_973;
assign grp_fu_514_p2 = \add_32ns_32ns_32_2_1_U7.dout ;
assign \add_32ns_32ns_32_2_1_U7.reset  = ap_rst;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s0  = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.a ;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s0  = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.b ;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.s  = { \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s2 , \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.sum_s1  };
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.a  = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s1 ;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.b  = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s1 ;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cin  = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.carry_s1 ;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s2  = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cout ;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s2  = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.s ;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.a  = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.a [15:0];
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.b  = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.b [15:0];
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cin  = 1'h0;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s1  = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cout ;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s1  = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.s ;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.a  = \add_32ns_32ns_32_2_1_U17.din0 ;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.b  = \add_32ns_32ns_32_2_1_U17.din1 ;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  = \add_32ns_32ns_32_2_1_U17.ce ;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.clk  = \add_32ns_32ns_32_2_1_U17.clk ;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.reset  = \add_32ns_32ns_32_2_1_U17.reset ;
assign \add_32ns_32ns_32_2_1_U17.dout  = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_6_U.s ;
assign \add_32ns_32ns_32_2_1_U17.ce  = 1'h1;
assign \add_32ns_32ns_32_2_1_U17.clk  = ap_clk;
assign \add_32ns_32ns_32_2_1_U17.din0  = ret_V_36_cast_reg_1153;
assign \add_32ns_32ns_32_2_1_U17.din1  = 32'd1;
assign grp_fu_792_p2 = \add_32ns_32ns_32_2_1_U17.dout ;
assign \add_32ns_32ns_32_2_1_U17.reset  = ap_rst;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s0  = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.a ;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s0  = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.b ;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.s  = { \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s2 , \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.sum_s1  };
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.a  = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s1 ;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.b  = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s1 ;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cin  = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.carry_s1 ;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s2  = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cout ;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s2  = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.s ;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.a  = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.a [15:0];
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.b  = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.b [15:0];
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cin  = 1'h0;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s1  = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cout ;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s1  = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.s ;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.a  = \add_32ns_32ns_32_2_1_U14.din0 ;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.b  = \add_32ns_32ns_32_2_1_U14.din1 ;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  = \add_32ns_32ns_32_2_1_U14.ce ;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.clk  = \add_32ns_32ns_32_2_1_U14.clk ;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.reset  = \add_32ns_32ns_32_2_1_U14.reset ;
assign \add_32ns_32ns_32_2_1_U14.dout  = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_6_U.s ;
assign \add_32ns_32ns_32_2_1_U14.ce  = 1'h1;
assign \add_32ns_32ns_32_2_1_U14.clk  = ap_clk;
assign \add_32ns_32ns_32_2_1_U14.din0  = add_ln69_2_reg_1098;
assign \add_32ns_32ns_32_2_1_U14.din1  = ret_V_31_reg_1093;
assign grp_fu_713_p2 = \add_32ns_32ns_32_2_1_U14.dout ;
assign \add_32ns_32ns_32_2_1_U14.reset  = ap_rst;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s0  = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.a ;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s0  = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.b ;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.s  = { \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s2 , \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.sum_s1  };
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.a  = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.ain_s1 ;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.b  = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.bin_s1 ;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cin  = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.carry_s1 ;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s2  = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.cout ;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s2  = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.u2.s ;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.a  = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.a [15:0];
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.b  = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.b [15:0];
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cin  = 1'h0;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.facout_s1  = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.cout ;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.fas_s1  = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.u1.s ;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.a  = \add_32ns_32ns_32_2_1_U10.din0 ;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.b  = \add_32ns_32ns_32_2_1_U10.din1 ;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.ce  = \add_32ns_32ns_32_2_1_U10.ce ;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.clk  = \add_32ns_32ns_32_2_1_U10.clk ;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.reset  = \add_32ns_32ns_32_2_1_U10.reset ;
assign \add_32ns_32ns_32_2_1_U10.dout  = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_6_U.s ;
assign \add_32ns_32ns_32_2_1_U10.ce  = 1'h1;
assign \add_32ns_32ns_32_2_1_U10.clk  = ap_clk;
assign \add_32ns_32ns_32_2_1_U10.din0  = ret_V_33_cast_reg_1038;
assign \add_32ns_32ns_32_2_1_U10.din1  = 32'd1;
assign grp_fu_588_p2 = \add_32ns_32ns_32_2_1_U10.dout ;
assign \add_32ns_32ns_32_2_1_U10.reset  = ap_rst;
assign \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.ain_s0  = \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.a ;
assign \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.bin_s0  = \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.b ;
assign \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.s  = { \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.fas_s2 , \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.sum_s1  };
assign \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.u2.a  = \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.ain_s1 ;
assign \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.u2.b  = \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.bin_s1 ;
assign \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.u2.cin  = \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.carry_s1 ;
assign \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.facout_s2  = \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.u2.cout ;
assign \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.fas_s2  = \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.u2.s ;
assign \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.u1.a  = \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.a [7:0];
assign \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.u1.b  = \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.b [7:0];
assign \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.u1.cin  = 1'h0;
assign \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.facout_s1  = \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.u1.cout ;
assign \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.fas_s1  = \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.u1.s ;
assign \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.a  = \add_17s_17s_17_2_1_U3.din0 ;
assign \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.b  = \add_17s_17s_17_2_1_U3.din1 ;
assign \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.ce  = \add_17s_17s_17_2_1_U3.ce ;
assign \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.clk  = \add_17s_17s_17_2_1_U3.clk ;
assign \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.reset  = \add_17s_17s_17_2_1_U3.reset ;
assign \add_17s_17s_17_2_1_U3.dout  = \add_17s_17s_17_2_1_U3.top_add_17s_17s_17_2_1_Adder_2_U.s ;
assign \add_17s_17s_17_2_1_U3.ce  = 1'h1;
assign \add_17s_17s_17_2_1_U3.clk  = ap_clk;
assign \add_17s_17s_17_2_1_U3.din0  = { ret_V_27_reg_901[2], ret_V_27_reg_901[2], ret_V_27_reg_901[2], ret_V_27_reg_901[2], ret_V_27_reg_901[2], ret_V_27_reg_901[2], ret_V_27_reg_901[2], ret_V_27_reg_901[2], ret_V_27_reg_901[2], ret_V_27_reg_901, 5'h00 };
assign \add_17s_17s_17_2_1_U3.din1  = { op_11[15], op_11 };
assign grp_fu_404_p2 = \add_17s_17s_17_2_1_U3.dout ;
assign \add_17s_17s_17_2_1_U3.reset  = ap_rst;
endmodule


// Product machine:
module top_A_times_top_B (ap_start, op_0, op_10, op_11, op_13, op_15, op_16, op_17, op_19, op_3, op_4, op_5, op_9, ap_clk, unsafe_signal);
input ap_start;
input op_0;
input [1:0] op_10;
input [15:0] op_11;
input [1:0] op_13;
input [3:0] op_15;
input [31:0] op_16;
input [3:0] op_17;
input [3:0] op_19;
input [3:0] op_3;
input [3:0] op_4;
input [3:0] op_5;
input [7:0] op_9;
input ap_clk;
output unsafe_signal;
reg _setup;
initial _setup = 1'b0;
always @ (posedge ap_clk) _setup <= 1'b1;
reg ap_start_internal;
always @ (posedge ap_clk) if (!_setup) ap_start_internal <= ap_start;
reg op_0_internal;
always @ (posedge ap_clk) if (!_setup) op_0_internal <= op_0;
reg [1:0] op_10_internal;
always @ (posedge ap_clk) if (!_setup) op_10_internal <= op_10;
reg [15:0] op_11_internal;
always @ (posedge ap_clk) if (!_setup) op_11_internal <= op_11;
reg [1:0] op_13_internal;
always @ (posedge ap_clk) if (!_setup) op_13_internal <= op_13;
reg [3:0] op_15_internal;
always @ (posedge ap_clk) if (!_setup) op_15_internal <= op_15;
reg [31:0] op_16_internal;
always @ (posedge ap_clk) if (!_setup) op_16_internal <= op_16;
reg [3:0] op_17_internal;
always @ (posedge ap_clk) if (!_setup) op_17_internal <= op_17;
reg [3:0] op_19_internal;
always @ (posedge ap_clk) if (!_setup) op_19_internal <= op_19;
reg [3:0] op_3_internal;
always @ (posedge ap_clk) if (!_setup) op_3_internal <= op_3;
reg [3:0] op_4_internal;
always @ (posedge ap_clk) if (!_setup) op_4_internal <= op_4;
reg [3:0] op_5_internal;
always @ (posedge ap_clk) if (!_setup) op_5_internal <= op_5;
reg [7:0] op_9_internal;
always @ (posedge ap_clk) if (!_setup) op_9_internal <= op_9;
wire ap_done_A;
wire ap_done_B;
wire ap_done_eq;
assign ap_done_eq = ap_done_A == ap_done_B;
wire ap_idle_A;
wire ap_idle_B;
wire ap_idle_eq;
assign ap_idle_eq = ap_idle_A == ap_idle_B;
wire ap_ready_A;
wire ap_ready_B;
wire ap_ready_eq;
assign ap_ready_eq = ap_ready_A == ap_ready_B;
wire [31:0] op_29_A;
wire [31:0] op_29_B;
wire op_29_eq;
assign op_29_eq = op_29_A == op_29_B;
wire op_29_ap_vld_A;
wire op_29_ap_vld_B;
wire clk_enable_A;
wire clk_enable_B;
assign clk_enable_A = _setup & (~op_29_ap_vld_A | op_29_ap_vld_B);
assign clk_enable_B = _setup;
wire divergent;
assign divergent = ~(ap_done_eq & ap_idle_eq & ap_ready_eq & op_29_eq);
assign unsafe_signal = op_29_ap_vld_A & op_29_ap_vld_B & divergent;
top_A instance_A (
    .ap_clk(ap_clk),
    .clk_enable(clk_enable_A),
    .ap_start(ap_start_internal),
    .op_0(op_0_internal),
    .op_10(op_10_internal),
    .op_11(op_11_internal),
    .op_13(op_13_internal),
    .op_15(op_15_internal),
    .op_16(op_16_internal),
    .op_17(op_17_internal),
    .op_19(op_19_internal),
    .op_3(op_3_internal),
    .op_4(op_4_internal),
    .op_5(op_5_internal),
    .op_9(op_9_internal),
    .ap_done(ap_done_A),
    .ap_idle(ap_idle_A),
    .ap_ready(ap_ready_A),
    .op_29(op_29_A),
    .op_29_ap_vld(op_29_ap_vld_A)
);
top_B instance_B (
    .ap_clk(ap_clk),
    .clk_enable(clk_enable_B),
    .ap_start(ap_start_internal),
    .op_0(op_0_internal),
    .op_10(op_10_internal),
    .op_11(op_11_internal),
    .op_13(op_13_internal),
    .op_15(op_15_internal),
    .op_16(op_16_internal),
    .op_17(op_17_internal),
    .op_19(op_19_internal),
    .op_3(op_3_internal),
    .op_4(op_4_internal),
    .op_5(op_5_internal),
    .op_9(op_9_internal),
    .ap_done(ap_done_B),
    .ap_idle(ap_idle_B),
    .ap_ready(ap_ready_B),
    .op_29(op_29_B),
    .op_29_ap_vld(op_29_ap_vld_B)
);
endmodule
