// Processed by function `construct_kairos` in `verilog_tricks.py`.
// Machine A:
// Processed by function `add_clk_enable_signal` in `verilog_tricks.py`.
// Processed by function `remove_reset_signal` in `verilog_tricks.py`.
module top_A (
  ap_clk,
  ap_start,
  ap_done,
  ap_idle,
  ap_ready,
  op_0,
  op_2,
  op_3,
  op_5,
  op_6,
  op_7,
  op_12,
  op_15,
  op_16,
  op_18,
  op_19,
  op_30,
  op_30_ap_vld,
clk_enable
);
input clk_enable;


input ap_clk;
wire ap_rst;
assign ap_rst = op_30_ap_vld;
input ap_start;
input op_0;
input op_12;
input [3:0] op_15;
input [15:0] op_16;
input [3:0] op_18;
input [3:0] op_19;
input op_2;
input [3:0] op_3;
input [1:0] op_5;
input [7:0] op_6;
input [3:0] op_7;
output ap_done;
output ap_idle;
output ap_ready;
output [31:0] op_30;
output op_30_ap_vld;


reg Range1_all_ones_reg_1583;
reg Range1_all_zeros_reg_1590;
reg Range2_all_ones_reg_1578;
reg \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.ain_s1 ;
reg \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.bin_s1 ;
reg \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.carry_s1 ;
reg \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.sum_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.ain_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.bin_s1 ;
reg \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.carry_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.sum_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.ain_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.bin_s1 ;
reg \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.carry_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.sum_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.ain_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.bin_s1 ;
reg \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.carry_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.sum_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.ain_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.bin_s1 ;
reg \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.carry_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.sum_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.ain_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.bin_s1 ;
reg \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.carry_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.sum_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.ain_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.bin_s1 ;
reg \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.carry_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.sum_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_11_U.ain_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_11_U.bin_s1 ;
reg \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_11_U.carry_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_11_U.sum_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_11_U.ain_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_11_U.bin_s1 ;
reg \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_11_U.carry_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_11_U.sum_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_11_U.ain_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_11_U.bin_s1 ;
reg \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_11_U.carry_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_11_U.sum_s1 ;
reg [16:0] \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_10_U.ain_s1 ;
reg [16:0] \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_10_U.bin_s1 ;
reg \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_10_U.carry_s1 ;
reg [16:0] \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_10_U.sum_s1 ;
reg [16:0] \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_10_U.ain_s1 ;
reg [16:0] \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_10_U.bin_s1 ;
reg \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_10_U.carry_s1 ;
reg [16:0] \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_10_U.sum_s1 ;
reg [16:0] \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_10_U.ain_s1 ;
reg [16:0] \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_10_U.bin_s1 ;
reg \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_10_U.carry_s1 ;
reg [16:0] \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_10_U.sum_s1 ;
reg [17:0] \add_35s_35s_35_2_1_U23.top_add_35s_35s_35_2_1_Adder_12_U.ain_s1 ;
reg [17:0] \add_35s_35s_35_2_1_U23.top_add_35s_35s_35_2_1_Adder_12_U.bin_s1 ;
reg \add_35s_35s_35_2_1_U23.top_add_35s_35s_35_2_1_Adder_12_U.carry_s1 ;
reg [16:0] \add_35s_35s_35_2_1_U23.top_add_35s_35s_35_2_1_Adder_12_U.sum_s1 ;
reg [1:0] \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.ain_s1 ;
reg [1:0] \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.bin_s1 ;
reg \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.carry_s1 ;
reg [1:0] \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.sum_s1 ;
reg [1:0] \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.ain_s1 ;
reg [1:0] \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.bin_s1 ;
reg \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.carry_s1 ;
reg [1:0] \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.sum_s1 ;
reg [2:0] \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.ain_s1 ;
reg [2:0] \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.bin_s1 ;
reg \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.carry_s1 ;
reg [1:0] \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.sum_s1 ;
reg [2:0] \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_5_U.ain_s1 ;
reg [2:0] \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_5_U.bin_s1 ;
reg \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_5_U.carry_s1 ;
reg [2:0] \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_5_U.sum_s1 ;
reg [2:0] \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.ain_s1 ;
reg [2:0] \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.bin_s1 ;
reg \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.carry_s1 ;
reg [2:0] \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.sum_s1 ;
reg [3:0] \add_8s_8ns_8_2_1_U11.top_add_8s_8ns_8_2_1_Adder_8_U.ain_s1 ;
reg [3:0] \add_8s_8ns_8_2_1_U11.top_add_8s_8ns_8_2_1_Adder_8_U.bin_s1 ;
reg \add_8s_8ns_8_2_1_U11.top_add_8s_8ns_8_2_1_Adder_8_U.carry_s1 ;
reg [3:0] \add_8s_8ns_8_2_1_U11.top_add_8s_8ns_8_2_1_Adder_8_U.sum_s1 ;
reg [3:0] \add_8s_8s_8_2_1_U10.top_add_8s_8s_8_2_1_Adder_7_U.ain_s1 ;
reg [3:0] \add_8s_8s_8_2_1_U10.top_add_8s_8s_8_2_1_Adder_7_U.bin_s1 ;
reg \add_8s_8s_8_2_1_U10.top_add_8s_8s_8_2_1_Adder_7_U.carry_s1 ;
reg [3:0] \add_8s_8s_8_2_1_U10.top_add_8s_8s_8_2_1_Adder_7_U.sum_s1 ;
reg [4:0] \add_9s_9ns_9_2_1_U5.top_add_9s_9ns_9_2_1_Adder_3_U.ain_s1 ;
reg [4:0] \add_9s_9ns_9_2_1_U5.top_add_9s_9ns_9_2_1_Adder_3_U.bin_s1 ;
reg \add_9s_9ns_9_2_1_U5.top_add_9s_9ns_9_2_1_Adder_3_U.carry_s1 ;
reg [3:0] \add_9s_9ns_9_2_1_U5.top_add_9s_9ns_9_2_1_Adder_3_U.sum_s1 ;
reg [4:0] \add_9s_9s_9_2_1_U8.top_add_9s_9s_9_2_1_Adder_6_U.ain_s1 ;
reg [4:0] \add_9s_9s_9_2_1_U8.top_add_9s_9s_9_2_1_Adder_6_U.bin_s1 ;
reg \add_9s_9s_9_2_1_U8.top_add_9s_9s_9_2_1_Adder_6_U.carry_s1 ;
reg [3:0] \add_9s_9s_9_2_1_U8.top_add_9s_9s_9_2_1_Adder_6_U.sum_s1 ;
reg [31:0] add_ln691_1_reg_1828;
reg [31:0] add_ln691_2_reg_1938;
reg [31:0] add_ln691_3_reg_1975;
reg [31:0] add_ln691_4_reg_2027;
reg [7:0] add_ln691_reg_1790;
reg and_ln406_reg_1573;
reg and_ln408_reg_1768;
reg and_ln785_1_reg_1687;
reg and_ln786_reg_1673;
reg [56:0] ap_CS_fsm = 57'h000000000000001;
reg carry_2_reg_1654;
reg carry_reg_1859;
reg deleted_zeros_reg_1661;
reg icmp_ln1497_reg_1886;
reg icmp_ln768_reg_1495;
reg icmp_ln786_reg_1500;
reg icmp_ln790_reg_1505;
reg icmp_ln851_1_reg_1617;
reg icmp_ln851_2_reg_2010;
reg icmp_ln851_reg_1419;
reg lhs_V_2_reg_1864;
reg [15:0] \mul_16ns_4s_20_7_1_U4.top_mul_16ns_4s_20_7_1_Mul_DSP_0_U.a_reg0 ;
reg [3:0] \mul_16ns_4s_20_7_1_U4.top_mul_16ns_4s_20_7_1_Mul_DSP_0_U.b_reg0 ;
reg [19:0] \mul_16ns_4s_20_7_1_U4.top_mul_16ns_4s_20_7_1_Mul_DSP_0_U.buff0 ;
reg [19:0] \mul_16ns_4s_20_7_1_U4.top_mul_16ns_4s_20_7_1_Mul_DSP_0_U.buff1 ;
reg [19:0] \mul_16ns_4s_20_7_1_U4.top_mul_16ns_4s_20_7_1_Mul_DSP_0_U.buff2 ;
reg [19:0] \mul_16ns_4s_20_7_1_U4.top_mul_16ns_4s_20_7_1_Mul_DSP_0_U.buff3 ;
reg [19:0] \mul_16ns_4s_20_7_1_U4.top_mul_16ns_4s_20_7_1_Mul_DSP_0_U.buff4 ;
reg newsignbit_reg_1879;
reg [5:0] op_10_V_reg_1795;
reg [31:0] op_23_V_reg_1874;
reg [31:0] op_28_V_reg_1995;
reg [7:0] op_8_V_reg_1521;
reg [3:0] op_9_V_reg_1722;
reg or_ln340_reg_1681;
reg or_ln384_reg_1516;
reg overflow_reg_1510;
reg p_Result_21_reg_1853;
reg p_Result_22_reg_1733;
reg p_Result_23_reg_1472;
reg p_Result_24_reg_1478;
reg p_Result_25_reg_1533;
reg p_Result_27_reg_1546;
reg p_Result_28_reg_1631;
reg p_Result_29_reg_1551;
reg [12:0] p_Result_6_reg_1557;
reg [13:0] p_Result_7_reg_1562;
reg [3:0] p_Val2_6_reg_1541;
reg [3:0] p_Val2_7_reg_1622;
reg [19:0] r_V_1_reg_1526;
reg r_reg_1753;
reg [4:0] ret_V_20_reg_1424;
reg [1:0] ret_V_21_reg_1441;
reg [31:0] ret_V_24_cast_reg_1821;
reg [8:0] ret_V_24_reg_1595;
reg [7:0] ret_V_25_reg_1758;
reg [33:0] ret_V_26_reg_1816;
reg [31:0] ret_V_27_reg_1833;
reg [31:0] ret_V_28_reg_1896;
reg [31:0] ret_V_29_reg_1906;
reg [1:0] ret_V_2_reg_1436;
reg [31:0] ret_V_30_cast_reg_1931;
reg [33:0] ret_V_30_reg_1926;
reg [33:0] ret_V_31_reg_1963;
reg [31:0] ret_V_32_cast_reg_1968;
reg [31:0] ret_V_32_reg_1985;
reg [34:0] ret_V_33_reg_2015;
reg [31:0] ret_V_34_cast_reg_2020;
reg [31:0] ret_V_34_reg_2032;
reg [5:0] ret_V_7_reg_1600;
reg [5:0] ret_V_9_reg_1638;
reg [1:0] ret_V_reg_1429;
reg [16:0] ret_reg_1467;
reg sel_tmp11_reg_1697;
reg [31:0] select_ln1192_reg_1901;
reg [16:0] select_ln1347_reg_1447;
reg [3:0] select_ln340_1_reg_1692;
reg [31:0] select_ln353_2_reg_1943;
reg [7:0] select_ln353_reg_1801;
reg [31:0] select_ln69_reg_1838;
reg [4:0] select_ln703_reg_1402;
reg [5:0] select_ln850_4_reg_1649;
reg [7:0] sext_ln850_reg_1773;
reg signbit_3_reg_1869;
reg [8:0] \sub_17ns_17ns_17_2_1_U3.top_sub_17ns_17ns_17_2_1_Adder_2_U.ain_s1 ;
reg [8:0] \sub_17ns_17ns_17_2_1_U3.top_sub_17ns_17ns_17_2_1_Adder_2_U.bin_s1 ;
reg \sub_17ns_17ns_17_2_1_U3.top_sub_17ns_17ns_17_2_1_Adder_2_U.carry_s1 ;
reg [7:0] \sub_17ns_17ns_17_2_1_U3.top_sub_17ns_17ns_17_2_1_Adder_2_U.sum_s1 ;
reg [11:0] tmp_2_reg_1484;
reg [6:0] tmp_3_reg_1763;
reg [4:0] trunc_ln2_reg_1728;
reg trunc_ln415_reg_1848;
reg [2:0] trunc_ln718_reg_1738;
reg [3:0] trunc_ln790_reg_1490;
reg [2:0] trunc_ln851_1_reg_1607;
reg xor_ln1497_reg_1980;
reg xor_ln416_reg_1643;
reg xor_ln785_3_reg_1667;
wire _000_;
wire _001_;
wire _002_;
wire [31:0] _003_;
wire [31:0] _004_;
wire [31:0] _005_;
wire [31:0] _006_;
wire [7:0] _007_;
wire _008_;
wire _009_;
wire _010_;
wire _011_;
wire [56:0] _012_;
wire _013_;
wire _014_;
wire _015_;
wire _016_;
wire _017_;
wire _018_;
wire _019_;
wire _020_;
wire _021_;
wire _022_;
wire _023_;
wire _024_;
wire [5:0] _025_;
wire [31:0] _026_;
wire [31:0] _027_;
wire [7:0] _028_;
wire [3:0] _029_;
wire _030_;
wire _031_;
wire _032_;
wire _033_;
wire _034_;
wire _035_;
wire _036_;
wire _037_;
wire _038_;
wire _039_;
wire _040_;
wire [12:0] _041_;
wire [13:0] _042_;
wire [3:0] _043_;
wire [3:0] _044_;
wire [19:0] _045_;
wire _046_;
wire [4:0] _047_;
wire [1:0] _048_;
wire [31:0] _049_;
wire [8:0] _050_;
wire [7:0] _051_;
wire [33:0] _052_;
wire [31:0] _053_;
wire [31:0] _054_;
wire [31:0] _055_;
wire [1:0] _056_;
wire [31:0] _057_;
wire [33:0] _058_;
wire [33:0] _059_;
wire [31:0] _060_;
wire [31:0] _061_;
wire [34:0] _062_;
wire [31:0] _063_;
wire [31:0] _064_;
wire [5:0] _065_;
wire [5:0] _066_;
wire [1:0] _067_;
wire [16:0] _068_;
wire _069_;
wire [31:0] _070_;
wire [16:0] _071_;
wire [3:0] _072_;
wire [31:0] _073_;
wire [7:0] _074_;
wire [31:0] _075_;
wire [1:0] _076_;
wire [5:0] _077_;
wire [7:0] _078_;
wire _079_;
wire [11:0] _080_;
wire [6:0] _081_;
wire [4:0] _082_;
wire _083_;
wire [2:0] _084_;
wire [3:0] _085_;
wire [2:0] _086_;
wire _087_;
wire _088_;
wire _089_;
wire [1:0] _090_;
wire _091_;
wire _092_;
wire _093_;
wire _094_;
wire _095_;
wire _096_;
wire _097_;
wire _098_;
wire _099_;
wire _100_;
wire _101_;
wire _102_;
wire _103_;
wire _104_;
wire _105_;
wire _106_;
wire _107_;
wire _108_;
wire [1:0] _109_;
wire [1:0] _110_;
wire [15:0] _111_;
wire [15:0] _112_;
wire _113_;
wire [15:0] _114_;
wire [16:0] _115_;
wire [16:0] _116_;
wire [15:0] _117_;
wire [15:0] _118_;
wire _119_;
wire [15:0] _120_;
wire [16:0] _121_;
wire [16:0] _122_;
wire [15:0] _123_;
wire [15:0] _124_;
wire _125_;
wire [15:0] _126_;
wire [16:0] _127_;
wire [16:0] _128_;
wire [15:0] _129_;
wire [15:0] _130_;
wire _131_;
wire [15:0] _132_;
wire [16:0] _133_;
wire [16:0] _134_;
wire [15:0] _135_;
wire [15:0] _136_;
wire _137_;
wire [15:0] _138_;
wire [16:0] _139_;
wire [16:0] _140_;
wire [15:0] _141_;
wire [15:0] _142_;
wire _143_;
wire [15:0] _144_;
wire [16:0] _145_;
wire [16:0] _146_;
wire [15:0] _147_;
wire [15:0] _148_;
wire _149_;
wire [15:0] _150_;
wire [16:0] _151_;
wire [16:0] _152_;
wire [15:0] _153_;
wire [15:0] _154_;
wire _155_;
wire [15:0] _156_;
wire [16:0] _157_;
wire [16:0] _158_;
wire [15:0] _159_;
wire [15:0] _160_;
wire _161_;
wire [15:0] _162_;
wire [16:0] _163_;
wire [16:0] _164_;
wire [16:0] _165_;
wire [16:0] _166_;
wire _167_;
wire [16:0] _168_;
wire [17:0] _169_;
wire [17:0] _170_;
wire [16:0] _171_;
wire [16:0] _172_;
wire _173_;
wire [16:0] _174_;
wire [17:0] _175_;
wire [17:0] _176_;
wire [16:0] _177_;
wire [16:0] _178_;
wire _179_;
wire [16:0] _180_;
wire [17:0] _181_;
wire [17:0] _182_;
wire [17:0] _183_;
wire [17:0] _184_;
wire _185_;
wire [16:0] _186_;
wire [17:0] _187_;
wire [18:0] _188_;
wire [1:0] _189_;
wire [1:0] _190_;
wire _191_;
wire [1:0] _192_;
wire [2:0] _193_;
wire [2:0] _194_;
wire [1:0] _195_;
wire [1:0] _196_;
wire _197_;
wire [1:0] _198_;
wire [2:0] _199_;
wire [2:0] _200_;
wire [2:0] _201_;
wire [2:0] _202_;
wire _203_;
wire [1:0] _204_;
wire [2:0] _205_;
wire [3:0] _206_;
wire [2:0] _207_;
wire [2:0] _208_;
wire _209_;
wire [2:0] _210_;
wire [3:0] _211_;
wire [3:0] _212_;
wire [2:0] _213_;
wire [2:0] _214_;
wire _215_;
wire [2:0] _216_;
wire [3:0] _217_;
wire [3:0] _218_;
wire [3:0] _219_;
wire [3:0] _220_;
wire _221_;
wire [3:0] _222_;
wire [4:0] _223_;
wire [4:0] _224_;
wire [3:0] _225_;
wire [3:0] _226_;
wire _227_;
wire [3:0] _228_;
wire [4:0] _229_;
wire [4:0] _230_;
wire [4:0] _231_;
wire [4:0] _232_;
wire _233_;
wire [3:0] _234_;
wire [4:0] _235_;
wire [5:0] _236_;
wire [4:0] _237_;
wire [4:0] _238_;
wire _239_;
wire [3:0] _240_;
wire [4:0] _241_;
wire [5:0] _242_;
wire [15:0] _243_;
wire [3:0] _244_;
wire [19:0] _245_;
wire [19:0] _246_;
wire [19:0] _247_;
wire [19:0] _248_;
wire [19:0] _249_;
wire [8:0] _250_;
wire [8:0] _251_;
wire _252_;
wire [7:0] _253_;
wire [8:0] _254_;
wire [9:0] _255_;
wire _256_;
wire _257_;
wire _258_;
wire _259_;
wire _260_;
wire _261_;
wire _262_;
wire _263_;
wire _264_;
wire _265_;
wire _266_;
wire _267_;
wire _268_;
wire _269_;
wire _270_;
wire _271_;
wire _272_;
wire _273_;
wire _274_;
wire _275_;
wire _276_;
wire _277_;
wire _278_;
wire _279_;
wire _280_;
wire _281_;
wire _282_;
wire _283_;
wire _284_;
wire _285_;
wire _286_;
wire _287_;
wire _288_;
wire _289_;
wire _290_;
wire _291_;
wire _292_;
wire _293_;
wire _294_;
wire _295_;
wire _296_;
wire _297_;
wire _298_;
wire _299_;
wire _300_;
wire _301_;
wire _302_;
wire _303_;
wire _304_;
wire _305_;
wire _306_;
wire _307_;
wire _308_;
wire _309_;
wire _310_;
wire _311_;
wire _312_;
wire _313_;
wire _314_;
wire _315_;
wire _316_;
wire _317_;
wire _318_;
wire _319_;
wire Range1_all_ones_fu_549_p2;
wire Range1_all_zeros_fu_554_p2;
wire Range2_all_ones_fu_544_p2;
wire \add_2ns_2ns_2_2_1_U2.ce ;
wire \add_2ns_2ns_2_2_1_U2.clk ;
wire [1:0] \add_2ns_2ns_2_2_1_U2.din0 ;
wire [1:0] \add_2ns_2ns_2_2_1_U2.din1 ;
wire [1:0] \add_2ns_2ns_2_2_1_U2.dout ;
wire \add_2ns_2ns_2_2_1_U2.reset ;
wire [1:0] \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.a ;
wire [1:0] \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.ain_s0 ;
wire [1:0] \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.b ;
wire [1:0] \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.bin_s0 ;
wire \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.ce ;
wire \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.clk ;
wire \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.facout_s1 ;
wire \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.facout_s2 ;
wire \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.fas_s1 ;
wire \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.fas_s2 ;
wire \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.reset ;
wire [1:0] \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.s ;
wire \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.a ;
wire \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.b ;
wire \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.cin ;
wire \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.cout ;
wire \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.s ;
wire \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.a ;
wire \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.b ;
wire \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.cin ;
wire \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.cout ;
wire \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.s ;
wire \add_32ns_32ns_32_2_1_U14.ce ;
wire \add_32ns_32ns_32_2_1_U14.clk ;
wire [31:0] \add_32ns_32ns_32_2_1_U14.din0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U14.din1 ;
wire [31:0] \add_32ns_32ns_32_2_1_U14.dout ;
wire \add_32ns_32ns_32_2_1_U14.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.a ;
wire [31:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.ain_s0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.b ;
wire [31:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.bin_s0 ;
wire \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.ce ;
wire \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.clk ;
wire \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.facout_s1 ;
wire \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.facout_s2 ;
wire [15:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.fas_s1 ;
wire [15:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.fas_s2 ;
wire \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.b ;
wire \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.cin ;
wire \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.b ;
wire \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.cin ;
wire \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.s ;
wire \add_32ns_32ns_32_2_1_U15.ce ;
wire \add_32ns_32ns_32_2_1_U15.clk ;
wire [31:0] \add_32ns_32ns_32_2_1_U15.din0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U15.din1 ;
wire [31:0] \add_32ns_32ns_32_2_1_U15.dout ;
wire \add_32ns_32ns_32_2_1_U15.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.a ;
wire [31:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.ain_s0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.b ;
wire [31:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.bin_s0 ;
wire \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.ce ;
wire \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.clk ;
wire \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.facout_s1 ;
wire \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.facout_s2 ;
wire [15:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.fas_s1 ;
wire [15:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.fas_s2 ;
wire \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.b ;
wire \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.cin ;
wire \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.b ;
wire \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.cin ;
wire \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.s ;
wire \add_32ns_32ns_32_2_1_U16.ce ;
wire \add_32ns_32ns_32_2_1_U16.clk ;
wire [31:0] \add_32ns_32ns_32_2_1_U16.din0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U16.din1 ;
wire [31:0] \add_32ns_32ns_32_2_1_U16.dout ;
wire \add_32ns_32ns_32_2_1_U16.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.a ;
wire [31:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.ain_s0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.b ;
wire [31:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.bin_s0 ;
wire \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.ce ;
wire \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.clk ;
wire \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.facout_s1 ;
wire \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.facout_s2 ;
wire [15:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.fas_s1 ;
wire [15:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.fas_s2 ;
wire \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.b ;
wire \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.cin ;
wire \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.b ;
wire \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.cin ;
wire \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.s ;
wire \add_32ns_32ns_32_2_1_U17.ce ;
wire \add_32ns_32ns_32_2_1_U17.clk ;
wire [31:0] \add_32ns_32ns_32_2_1_U17.din0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U17.din1 ;
wire [31:0] \add_32ns_32ns_32_2_1_U17.dout ;
wire \add_32ns_32ns_32_2_1_U17.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.a ;
wire [31:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.ain_s0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.b ;
wire [31:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.bin_s0 ;
wire \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.ce ;
wire \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.clk ;
wire \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.facout_s1 ;
wire \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.facout_s2 ;
wire [15:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.fas_s1 ;
wire [15:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.fas_s2 ;
wire \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.b ;
wire \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.cin ;
wire \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.b ;
wire \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.cin ;
wire \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.s ;
wire \add_32ns_32ns_32_2_1_U19.ce ;
wire \add_32ns_32ns_32_2_1_U19.clk ;
wire [31:0] \add_32ns_32ns_32_2_1_U19.din0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U19.din1 ;
wire [31:0] \add_32ns_32ns_32_2_1_U19.dout ;
wire \add_32ns_32ns_32_2_1_U19.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.a ;
wire [31:0] \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.ain_s0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.b ;
wire [31:0] \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.bin_s0 ;
wire \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.ce ;
wire \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.clk ;
wire \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.facout_s1 ;
wire \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.facout_s2 ;
wire [15:0] \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.fas_s1 ;
wire [15:0] \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.fas_s2 ;
wire \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.b ;
wire \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.cin ;
wire \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.b ;
wire \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.cin ;
wire \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.s ;
wire \add_32ns_32ns_32_2_1_U21.ce ;
wire \add_32ns_32ns_32_2_1_U21.clk ;
wire [31:0] \add_32ns_32ns_32_2_1_U21.din0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U21.din1 ;
wire [31:0] \add_32ns_32ns_32_2_1_U21.dout ;
wire \add_32ns_32ns_32_2_1_U21.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.a ;
wire [31:0] \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.ain_s0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.b ;
wire [31:0] \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.bin_s0 ;
wire \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.ce ;
wire \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.clk ;
wire \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.facout_s1 ;
wire \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.facout_s2 ;
wire [15:0] \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.fas_s1 ;
wire [15:0] \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.fas_s2 ;
wire \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.b ;
wire \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.cin ;
wire \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.b ;
wire \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.cin ;
wire \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.s ;
wire \add_32ns_32ns_32_2_1_U22.ce ;
wire \add_32ns_32ns_32_2_1_U22.clk ;
wire [31:0] \add_32ns_32ns_32_2_1_U22.din0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U22.din1 ;
wire [31:0] \add_32ns_32ns_32_2_1_U22.dout ;
wire \add_32ns_32ns_32_2_1_U22.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_11_U.a ;
wire [31:0] \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_11_U.ain_s0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_11_U.b ;
wire [31:0] \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_11_U.bin_s0 ;
wire \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_11_U.ce ;
wire \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_11_U.clk ;
wire \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_11_U.facout_s1 ;
wire \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_11_U.facout_s2 ;
wire [15:0] \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_11_U.fas_s1 ;
wire [15:0] \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_11_U.fas_s2 ;
wire \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_11_U.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_11_U.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.b ;
wire \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.cin ;
wire \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.b ;
wire \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.cin ;
wire \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.s ;
wire \add_32ns_32ns_32_2_1_U24.ce ;
wire \add_32ns_32ns_32_2_1_U24.clk ;
wire [31:0] \add_32ns_32ns_32_2_1_U24.din0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U24.din1 ;
wire [31:0] \add_32ns_32ns_32_2_1_U24.dout ;
wire \add_32ns_32ns_32_2_1_U24.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_11_U.a ;
wire [31:0] \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_11_U.ain_s0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_11_U.b ;
wire [31:0] \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_11_U.bin_s0 ;
wire \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_11_U.ce ;
wire \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_11_U.clk ;
wire \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_11_U.facout_s1 ;
wire \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_11_U.facout_s2 ;
wire [15:0] \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_11_U.fas_s1 ;
wire [15:0] \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_11_U.fas_s2 ;
wire \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_11_U.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_11_U.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.b ;
wire \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.cin ;
wire \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.b ;
wire \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.cin ;
wire \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.s ;
wire \add_32ns_32ns_32_2_1_U25.ce ;
wire \add_32ns_32ns_32_2_1_U25.clk ;
wire [31:0] \add_32ns_32ns_32_2_1_U25.din0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U25.din1 ;
wire [31:0] \add_32ns_32ns_32_2_1_U25.dout ;
wire \add_32ns_32ns_32_2_1_U25.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_11_U.a ;
wire [31:0] \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_11_U.ain_s0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_11_U.b ;
wire [31:0] \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_11_U.bin_s0 ;
wire \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_11_U.ce ;
wire \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_11_U.clk ;
wire \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_11_U.facout_s1 ;
wire \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_11_U.facout_s2 ;
wire [15:0] \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_11_U.fas_s1 ;
wire [15:0] \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_11_U.fas_s2 ;
wire \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_11_U.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_11_U.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.b ;
wire \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.cin ;
wire \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.b ;
wire \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.cin ;
wire \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.s ;
wire \add_34s_34s_34_2_1_U13.ce ;
wire \add_34s_34s_34_2_1_U13.clk ;
wire [33:0] \add_34s_34s_34_2_1_U13.din0 ;
wire [33:0] \add_34s_34s_34_2_1_U13.din1 ;
wire [33:0] \add_34s_34s_34_2_1_U13.dout ;
wire \add_34s_34s_34_2_1_U13.reset ;
wire [33:0] \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_10_U.a ;
wire [33:0] \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_10_U.ain_s0 ;
wire [33:0] \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_10_U.b ;
wire [33:0] \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_10_U.bin_s0 ;
wire \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_10_U.ce ;
wire \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_10_U.clk ;
wire \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_10_U.facout_s1 ;
wire \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_10_U.facout_s2 ;
wire [16:0] \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_10_U.fas_s1 ;
wire [16:0] \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_10_U.fas_s2 ;
wire \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_10_U.reset ;
wire [33:0] \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_10_U.s ;
wire [16:0] \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_10_U.u1.a ;
wire [16:0] \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_10_U.u1.b ;
wire \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_10_U.u1.cin ;
wire \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_10_U.u1.cout ;
wire [16:0] \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_10_U.u1.s ;
wire [16:0] \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_10_U.u2.a ;
wire [16:0] \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_10_U.u2.b ;
wire \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_10_U.u2.cin ;
wire \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_10_U.u2.cout ;
wire [16:0] \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_10_U.u2.s ;
wire \add_34s_34s_34_2_1_U18.ce ;
wire \add_34s_34s_34_2_1_U18.clk ;
wire [33:0] \add_34s_34s_34_2_1_U18.din0 ;
wire [33:0] \add_34s_34s_34_2_1_U18.din1 ;
wire [33:0] \add_34s_34s_34_2_1_U18.dout ;
wire \add_34s_34s_34_2_1_U18.reset ;
wire [33:0] \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_10_U.a ;
wire [33:0] \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_10_U.ain_s0 ;
wire [33:0] \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_10_U.b ;
wire [33:0] \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_10_U.bin_s0 ;
wire \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_10_U.ce ;
wire \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_10_U.clk ;
wire \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_10_U.facout_s1 ;
wire \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_10_U.facout_s2 ;
wire [16:0] \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_10_U.fas_s1 ;
wire [16:0] \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_10_U.fas_s2 ;
wire \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_10_U.reset ;
wire [33:0] \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_10_U.s ;
wire [16:0] \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_10_U.u1.a ;
wire [16:0] \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_10_U.u1.b ;
wire \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_10_U.u1.cin ;
wire \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_10_U.u1.cout ;
wire [16:0] \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_10_U.u1.s ;
wire [16:0] \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_10_U.u2.a ;
wire [16:0] \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_10_U.u2.b ;
wire \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_10_U.u2.cin ;
wire \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_10_U.u2.cout ;
wire [16:0] \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_10_U.u2.s ;
wire \add_34s_34s_34_2_1_U20.ce ;
wire \add_34s_34s_34_2_1_U20.clk ;
wire [33:0] \add_34s_34s_34_2_1_U20.din0 ;
wire [33:0] \add_34s_34s_34_2_1_U20.din1 ;
wire [33:0] \add_34s_34s_34_2_1_U20.dout ;
wire \add_34s_34s_34_2_1_U20.reset ;
wire [33:0] \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_10_U.a ;
wire [33:0] \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_10_U.ain_s0 ;
wire [33:0] \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_10_U.b ;
wire [33:0] \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_10_U.bin_s0 ;
wire \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_10_U.ce ;
wire \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_10_U.clk ;
wire \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_10_U.facout_s1 ;
wire \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_10_U.facout_s2 ;
wire [16:0] \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_10_U.fas_s1 ;
wire [16:0] \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_10_U.fas_s2 ;
wire \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_10_U.reset ;
wire [33:0] \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_10_U.s ;
wire [16:0] \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_10_U.u1.a ;
wire [16:0] \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_10_U.u1.b ;
wire \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_10_U.u1.cin ;
wire \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_10_U.u1.cout ;
wire [16:0] \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_10_U.u1.s ;
wire [16:0] \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_10_U.u2.a ;
wire [16:0] \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_10_U.u2.b ;
wire \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_10_U.u2.cin ;
wire \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_10_U.u2.cout ;
wire [16:0] \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_10_U.u2.s ;
wire \add_35s_35s_35_2_1_U23.ce ;
wire \add_35s_35s_35_2_1_U23.clk ;
wire [34:0] \add_35s_35s_35_2_1_U23.din0 ;
wire [34:0] \add_35s_35s_35_2_1_U23.din1 ;
wire [34:0] \add_35s_35s_35_2_1_U23.dout ;
wire \add_35s_35s_35_2_1_U23.reset ;
wire [34:0] \add_35s_35s_35_2_1_U23.top_add_35s_35s_35_2_1_Adder_12_U.a ;
wire [34:0] \add_35s_35s_35_2_1_U23.top_add_35s_35s_35_2_1_Adder_12_U.ain_s0 ;
wire [34:0] \add_35s_35s_35_2_1_U23.top_add_35s_35s_35_2_1_Adder_12_U.b ;
wire [34:0] \add_35s_35s_35_2_1_U23.top_add_35s_35s_35_2_1_Adder_12_U.bin_s0 ;
wire \add_35s_35s_35_2_1_U23.top_add_35s_35s_35_2_1_Adder_12_U.ce ;
wire \add_35s_35s_35_2_1_U23.top_add_35s_35s_35_2_1_Adder_12_U.clk ;
wire \add_35s_35s_35_2_1_U23.top_add_35s_35s_35_2_1_Adder_12_U.facout_s1 ;
wire \add_35s_35s_35_2_1_U23.top_add_35s_35s_35_2_1_Adder_12_U.facout_s2 ;
wire [16:0] \add_35s_35s_35_2_1_U23.top_add_35s_35s_35_2_1_Adder_12_U.fas_s1 ;
wire [17:0] \add_35s_35s_35_2_1_U23.top_add_35s_35s_35_2_1_Adder_12_U.fas_s2 ;
wire \add_35s_35s_35_2_1_U23.top_add_35s_35s_35_2_1_Adder_12_U.reset ;
wire [34:0] \add_35s_35s_35_2_1_U23.top_add_35s_35s_35_2_1_Adder_12_U.s ;
wire [16:0] \add_35s_35s_35_2_1_U23.top_add_35s_35s_35_2_1_Adder_12_U.u1.a ;
wire [16:0] \add_35s_35s_35_2_1_U23.top_add_35s_35s_35_2_1_Adder_12_U.u1.b ;
wire \add_35s_35s_35_2_1_U23.top_add_35s_35s_35_2_1_Adder_12_U.u1.cin ;
wire \add_35s_35s_35_2_1_U23.top_add_35s_35s_35_2_1_Adder_12_U.u1.cout ;
wire [16:0] \add_35s_35s_35_2_1_U23.top_add_35s_35s_35_2_1_Adder_12_U.u1.s ;
wire [17:0] \add_35s_35s_35_2_1_U23.top_add_35s_35s_35_2_1_Adder_12_U.u2.a ;
wire [17:0] \add_35s_35s_35_2_1_U23.top_add_35s_35s_35_2_1_Adder_12_U.u2.b ;
wire \add_35s_35s_35_2_1_U23.top_add_35s_35s_35_2_1_Adder_12_U.u2.cin ;
wire \add_35s_35s_35_2_1_U23.top_add_35s_35s_35_2_1_Adder_12_U.u2.cout ;
wire [17:0] \add_35s_35s_35_2_1_U23.top_add_35s_35s_35_2_1_Adder_12_U.u2.s ;
wire \add_4ns_4ns_4_2_1_U6.ce ;
wire \add_4ns_4ns_4_2_1_U6.clk ;
wire [3:0] \add_4ns_4ns_4_2_1_U6.din0 ;
wire [3:0] \add_4ns_4ns_4_2_1_U6.din1 ;
wire [3:0] \add_4ns_4ns_4_2_1_U6.dout ;
wire \add_4ns_4ns_4_2_1_U6.reset ;
wire [3:0] \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.a ;
wire [3:0] \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.ain_s0 ;
wire [3:0] \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.b ;
wire [3:0] \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.bin_s0 ;
wire \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.ce ;
wire \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.clk ;
wire \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.facout_s1 ;
wire \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.facout_s2 ;
wire [1:0] \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.fas_s1 ;
wire [1:0] \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.fas_s2 ;
wire \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.reset ;
wire [3:0] \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.s ;
wire [1:0] \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.u1.a ;
wire [1:0] \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.u1.b ;
wire \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.u1.cin ;
wire \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.u1.cout ;
wire [1:0] \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.u1.s ;
wire [1:0] \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.u2.a ;
wire [1:0] \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.u2.b ;
wire \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.u2.cin ;
wire \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.u2.cout ;
wire [1:0] \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.u2.s ;
wire \add_4ns_4ns_4_2_1_U9.ce ;
wire \add_4ns_4ns_4_2_1_U9.clk ;
wire [3:0] \add_4ns_4ns_4_2_1_U9.din0 ;
wire [3:0] \add_4ns_4ns_4_2_1_U9.din1 ;
wire [3:0] \add_4ns_4ns_4_2_1_U9.dout ;
wire \add_4ns_4ns_4_2_1_U9.reset ;
wire [3:0] \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.a ;
wire [3:0] \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.ain_s0 ;
wire [3:0] \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.b ;
wire [3:0] \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.bin_s0 ;
wire \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.ce ;
wire \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.clk ;
wire \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.facout_s1 ;
wire \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.facout_s2 ;
wire [1:0] \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.fas_s1 ;
wire [1:0] \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.fas_s2 ;
wire \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.reset ;
wire [3:0] \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.s ;
wire [1:0] \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.u1.a ;
wire [1:0] \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.u1.b ;
wire \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.u1.cin ;
wire \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.u1.cout ;
wire [1:0] \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.u1.s ;
wire [1:0] \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.u2.a ;
wire [1:0] \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.u2.b ;
wire \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.u2.cin ;
wire \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.u2.cout ;
wire [1:0] \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.u2.s ;
wire \add_5ns_5s_5_2_1_U1.ce ;
wire \add_5ns_5s_5_2_1_U1.clk ;
wire [4:0] \add_5ns_5s_5_2_1_U1.din0 ;
wire [4:0] \add_5ns_5s_5_2_1_U1.din1 ;
wire [4:0] \add_5ns_5s_5_2_1_U1.dout ;
wire \add_5ns_5s_5_2_1_U1.reset ;
wire [4:0] \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.a ;
wire [4:0] \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.ain_s0 ;
wire [4:0] \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.b ;
wire [4:0] \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.bin_s0 ;
wire \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.ce ;
wire \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.clk ;
wire \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.facout_s1 ;
wire \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.facout_s2 ;
wire [1:0] \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.fas_s1 ;
wire [2:0] \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.fas_s2 ;
wire \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.reset ;
wire [4:0] \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.s ;
wire [1:0] \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.u1.a ;
wire [1:0] \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.u1.b ;
wire \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.u1.cin ;
wire \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.u1.cout ;
wire [1:0] \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.u1.s ;
wire [2:0] \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.u2.a ;
wire [2:0] \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.u2.b ;
wire \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.u2.cin ;
wire \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.u2.cout ;
wire [2:0] \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.u2.s ;
wire \add_6ns_6ns_6_2_1_U7.ce ;
wire \add_6ns_6ns_6_2_1_U7.clk ;
wire [5:0] \add_6ns_6ns_6_2_1_U7.din0 ;
wire [5:0] \add_6ns_6ns_6_2_1_U7.din1 ;
wire [5:0] \add_6ns_6ns_6_2_1_U7.dout ;
wire \add_6ns_6ns_6_2_1_U7.reset ;
wire [5:0] \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_5_U.a ;
wire [5:0] \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_5_U.ain_s0 ;
wire [5:0] \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_5_U.b ;
wire [5:0] \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_5_U.bin_s0 ;
wire \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_5_U.ce ;
wire \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_5_U.clk ;
wire \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_5_U.facout_s1 ;
wire \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_5_U.facout_s2 ;
wire [2:0] \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_5_U.fas_s1 ;
wire [2:0] \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_5_U.fas_s2 ;
wire \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_5_U.reset ;
wire [5:0] \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_5_U.s ;
wire [2:0] \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_5_U.u1.a ;
wire [2:0] \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_5_U.u1.b ;
wire \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_5_U.u1.cin ;
wire \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_5_U.u1.cout ;
wire [2:0] \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_5_U.u1.s ;
wire [2:0] \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_5_U.u2.a ;
wire [2:0] \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_5_U.u2.b ;
wire \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_5_U.u2.cin ;
wire \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_5_U.u2.cout ;
wire [2:0] \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_5_U.u2.s ;
wire \add_6s_6ns_6_2_1_U12.ce ;
wire \add_6s_6ns_6_2_1_U12.clk ;
wire [5:0] \add_6s_6ns_6_2_1_U12.din0 ;
wire [5:0] \add_6s_6ns_6_2_1_U12.din1 ;
wire [5:0] \add_6s_6ns_6_2_1_U12.dout ;
wire \add_6s_6ns_6_2_1_U12.reset ;
wire [5:0] \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.a ;
wire [5:0] \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.ain_s0 ;
wire [5:0] \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.b ;
wire [5:0] \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.bin_s0 ;
wire \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.ce ;
wire \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.clk ;
wire \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.facout_s1 ;
wire \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.facout_s2 ;
wire [2:0] \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.fas_s1 ;
wire [2:0] \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.fas_s2 ;
wire \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.reset ;
wire [5:0] \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.s ;
wire [2:0] \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.u1.a ;
wire [2:0] \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.u1.b ;
wire \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.u1.cin ;
wire \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.u1.cout ;
wire [2:0] \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.u1.s ;
wire [2:0] \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.u2.a ;
wire [2:0] \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.u2.b ;
wire \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.u2.cin ;
wire \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.u2.cout ;
wire [2:0] \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.u2.s ;
wire \add_8s_8ns_8_2_1_U11.ce ;
wire \add_8s_8ns_8_2_1_U11.clk ;
wire [7:0] \add_8s_8ns_8_2_1_U11.din0 ;
wire [7:0] \add_8s_8ns_8_2_1_U11.din1 ;
wire [7:0] \add_8s_8ns_8_2_1_U11.dout ;
wire \add_8s_8ns_8_2_1_U11.reset ;
wire [7:0] \add_8s_8ns_8_2_1_U11.top_add_8s_8ns_8_2_1_Adder_8_U.a ;
wire [7:0] \add_8s_8ns_8_2_1_U11.top_add_8s_8ns_8_2_1_Adder_8_U.ain_s0 ;
wire [7:0] \add_8s_8ns_8_2_1_U11.top_add_8s_8ns_8_2_1_Adder_8_U.b ;
wire [7:0] \add_8s_8ns_8_2_1_U11.top_add_8s_8ns_8_2_1_Adder_8_U.bin_s0 ;
wire \add_8s_8ns_8_2_1_U11.top_add_8s_8ns_8_2_1_Adder_8_U.ce ;
wire \add_8s_8ns_8_2_1_U11.top_add_8s_8ns_8_2_1_Adder_8_U.clk ;
wire \add_8s_8ns_8_2_1_U11.top_add_8s_8ns_8_2_1_Adder_8_U.facout_s1 ;
wire \add_8s_8ns_8_2_1_U11.top_add_8s_8ns_8_2_1_Adder_8_U.facout_s2 ;
wire [3:0] \add_8s_8ns_8_2_1_U11.top_add_8s_8ns_8_2_1_Adder_8_U.fas_s1 ;
wire [3:0] \add_8s_8ns_8_2_1_U11.top_add_8s_8ns_8_2_1_Adder_8_U.fas_s2 ;
wire \add_8s_8ns_8_2_1_U11.top_add_8s_8ns_8_2_1_Adder_8_U.reset ;
wire [7:0] \add_8s_8ns_8_2_1_U11.top_add_8s_8ns_8_2_1_Adder_8_U.s ;
wire [3:0] \add_8s_8ns_8_2_1_U11.top_add_8s_8ns_8_2_1_Adder_8_U.u1.a ;
wire [3:0] \add_8s_8ns_8_2_1_U11.top_add_8s_8ns_8_2_1_Adder_8_U.u1.b ;
wire \add_8s_8ns_8_2_1_U11.top_add_8s_8ns_8_2_1_Adder_8_U.u1.cin ;
wire \add_8s_8ns_8_2_1_U11.top_add_8s_8ns_8_2_1_Adder_8_U.u1.cout ;
wire [3:0] \add_8s_8ns_8_2_1_U11.top_add_8s_8ns_8_2_1_Adder_8_U.u1.s ;
wire [3:0] \add_8s_8ns_8_2_1_U11.top_add_8s_8ns_8_2_1_Adder_8_U.u2.a ;
wire [3:0] \add_8s_8ns_8_2_1_U11.top_add_8s_8ns_8_2_1_Adder_8_U.u2.b ;
wire \add_8s_8ns_8_2_1_U11.top_add_8s_8ns_8_2_1_Adder_8_U.u2.cin ;
wire \add_8s_8ns_8_2_1_U11.top_add_8s_8ns_8_2_1_Adder_8_U.u2.cout ;
wire [3:0] \add_8s_8ns_8_2_1_U11.top_add_8s_8ns_8_2_1_Adder_8_U.u2.s ;
wire \add_8s_8s_8_2_1_U10.ce ;
wire \add_8s_8s_8_2_1_U10.clk ;
wire [7:0] \add_8s_8s_8_2_1_U10.din0 ;
wire [7:0] \add_8s_8s_8_2_1_U10.din1 ;
wire [7:0] \add_8s_8s_8_2_1_U10.dout ;
wire \add_8s_8s_8_2_1_U10.reset ;
wire [7:0] \add_8s_8s_8_2_1_U10.top_add_8s_8s_8_2_1_Adder_7_U.a ;
wire [7:0] \add_8s_8s_8_2_1_U10.top_add_8s_8s_8_2_1_Adder_7_U.ain_s0 ;
wire [7:0] \add_8s_8s_8_2_1_U10.top_add_8s_8s_8_2_1_Adder_7_U.b ;
wire [7:0] \add_8s_8s_8_2_1_U10.top_add_8s_8s_8_2_1_Adder_7_U.bin_s0 ;
wire \add_8s_8s_8_2_1_U10.top_add_8s_8s_8_2_1_Adder_7_U.ce ;
wire \add_8s_8s_8_2_1_U10.top_add_8s_8s_8_2_1_Adder_7_U.clk ;
wire \add_8s_8s_8_2_1_U10.top_add_8s_8s_8_2_1_Adder_7_U.facout_s1 ;
wire \add_8s_8s_8_2_1_U10.top_add_8s_8s_8_2_1_Adder_7_U.facout_s2 ;
wire [3:0] \add_8s_8s_8_2_1_U10.top_add_8s_8s_8_2_1_Adder_7_U.fas_s1 ;
wire [3:0] \add_8s_8s_8_2_1_U10.top_add_8s_8s_8_2_1_Adder_7_U.fas_s2 ;
wire \add_8s_8s_8_2_1_U10.top_add_8s_8s_8_2_1_Adder_7_U.reset ;
wire [7:0] \add_8s_8s_8_2_1_U10.top_add_8s_8s_8_2_1_Adder_7_U.s ;
wire [3:0] \add_8s_8s_8_2_1_U10.top_add_8s_8s_8_2_1_Adder_7_U.u1.a ;
wire [3:0] \add_8s_8s_8_2_1_U10.top_add_8s_8s_8_2_1_Adder_7_U.u1.b ;
wire \add_8s_8s_8_2_1_U10.top_add_8s_8s_8_2_1_Adder_7_U.u1.cin ;
wire \add_8s_8s_8_2_1_U10.top_add_8s_8s_8_2_1_Adder_7_U.u1.cout ;
wire [3:0] \add_8s_8s_8_2_1_U10.top_add_8s_8s_8_2_1_Adder_7_U.u1.s ;
wire [3:0] \add_8s_8s_8_2_1_U10.top_add_8s_8s_8_2_1_Adder_7_U.u2.a ;
wire [3:0] \add_8s_8s_8_2_1_U10.top_add_8s_8s_8_2_1_Adder_7_U.u2.b ;
wire \add_8s_8s_8_2_1_U10.top_add_8s_8s_8_2_1_Adder_7_U.u2.cin ;
wire \add_8s_8s_8_2_1_U10.top_add_8s_8s_8_2_1_Adder_7_U.u2.cout ;
wire [3:0] \add_8s_8s_8_2_1_U10.top_add_8s_8s_8_2_1_Adder_7_U.u2.s ;
wire \add_9s_9ns_9_2_1_U5.ce ;
wire \add_9s_9ns_9_2_1_U5.clk ;
wire [8:0] \add_9s_9ns_9_2_1_U5.din0 ;
wire [8:0] \add_9s_9ns_9_2_1_U5.din1 ;
wire [8:0] \add_9s_9ns_9_2_1_U5.dout ;
wire \add_9s_9ns_9_2_1_U5.reset ;
wire [8:0] \add_9s_9ns_9_2_1_U5.top_add_9s_9ns_9_2_1_Adder_3_U.a ;
wire [8:0] \add_9s_9ns_9_2_1_U5.top_add_9s_9ns_9_2_1_Adder_3_U.ain_s0 ;
wire [8:0] \add_9s_9ns_9_2_1_U5.top_add_9s_9ns_9_2_1_Adder_3_U.b ;
wire [8:0] \add_9s_9ns_9_2_1_U5.top_add_9s_9ns_9_2_1_Adder_3_U.bin_s0 ;
wire \add_9s_9ns_9_2_1_U5.top_add_9s_9ns_9_2_1_Adder_3_U.ce ;
wire \add_9s_9ns_9_2_1_U5.top_add_9s_9ns_9_2_1_Adder_3_U.clk ;
wire \add_9s_9ns_9_2_1_U5.top_add_9s_9ns_9_2_1_Adder_3_U.facout_s1 ;
wire \add_9s_9ns_9_2_1_U5.top_add_9s_9ns_9_2_1_Adder_3_U.facout_s2 ;
wire [3:0] \add_9s_9ns_9_2_1_U5.top_add_9s_9ns_9_2_1_Adder_3_U.fas_s1 ;
wire [4:0] \add_9s_9ns_9_2_1_U5.top_add_9s_9ns_9_2_1_Adder_3_U.fas_s2 ;
wire \add_9s_9ns_9_2_1_U5.top_add_9s_9ns_9_2_1_Adder_3_U.reset ;
wire [8:0] \add_9s_9ns_9_2_1_U5.top_add_9s_9ns_9_2_1_Adder_3_U.s ;
wire [3:0] \add_9s_9ns_9_2_1_U5.top_add_9s_9ns_9_2_1_Adder_3_U.u1.a ;
wire [3:0] \add_9s_9ns_9_2_1_U5.top_add_9s_9ns_9_2_1_Adder_3_U.u1.b ;
wire \add_9s_9ns_9_2_1_U5.top_add_9s_9ns_9_2_1_Adder_3_U.u1.cin ;
wire \add_9s_9ns_9_2_1_U5.top_add_9s_9ns_9_2_1_Adder_3_U.u1.cout ;
wire [3:0] \add_9s_9ns_9_2_1_U5.top_add_9s_9ns_9_2_1_Adder_3_U.u1.s ;
wire [4:0] \add_9s_9ns_9_2_1_U5.top_add_9s_9ns_9_2_1_Adder_3_U.u2.a ;
wire [4:0] \add_9s_9ns_9_2_1_U5.top_add_9s_9ns_9_2_1_Adder_3_U.u2.b ;
wire \add_9s_9ns_9_2_1_U5.top_add_9s_9ns_9_2_1_Adder_3_U.u2.cin ;
wire \add_9s_9ns_9_2_1_U5.top_add_9s_9ns_9_2_1_Adder_3_U.u2.cout ;
wire [4:0] \add_9s_9ns_9_2_1_U5.top_add_9s_9ns_9_2_1_Adder_3_U.u2.s ;
wire \add_9s_9s_9_2_1_U8.ce ;
wire \add_9s_9s_9_2_1_U8.clk ;
wire [8:0] \add_9s_9s_9_2_1_U8.din0 ;
wire [8:0] \add_9s_9s_9_2_1_U8.din1 ;
wire [8:0] \add_9s_9s_9_2_1_U8.dout ;
wire \add_9s_9s_9_2_1_U8.reset ;
wire [8:0] \add_9s_9s_9_2_1_U8.top_add_9s_9s_9_2_1_Adder_6_U.a ;
wire [8:0] \add_9s_9s_9_2_1_U8.top_add_9s_9s_9_2_1_Adder_6_U.ain_s0 ;
wire [8:0] \add_9s_9s_9_2_1_U8.top_add_9s_9s_9_2_1_Adder_6_U.b ;
wire [8:0] \add_9s_9s_9_2_1_U8.top_add_9s_9s_9_2_1_Adder_6_U.bin_s0 ;
wire \add_9s_9s_9_2_1_U8.top_add_9s_9s_9_2_1_Adder_6_U.ce ;
wire \add_9s_9s_9_2_1_U8.top_add_9s_9s_9_2_1_Adder_6_U.clk ;
wire \add_9s_9s_9_2_1_U8.top_add_9s_9s_9_2_1_Adder_6_U.facout_s1 ;
wire \add_9s_9s_9_2_1_U8.top_add_9s_9s_9_2_1_Adder_6_U.facout_s2 ;
wire [3:0] \add_9s_9s_9_2_1_U8.top_add_9s_9s_9_2_1_Adder_6_U.fas_s1 ;
wire [4:0] \add_9s_9s_9_2_1_U8.top_add_9s_9s_9_2_1_Adder_6_U.fas_s2 ;
wire \add_9s_9s_9_2_1_U8.top_add_9s_9s_9_2_1_Adder_6_U.reset ;
wire [8:0] \add_9s_9s_9_2_1_U8.top_add_9s_9s_9_2_1_Adder_6_U.s ;
wire [3:0] \add_9s_9s_9_2_1_U8.top_add_9s_9s_9_2_1_Adder_6_U.u1.a ;
wire [3:0] \add_9s_9s_9_2_1_U8.top_add_9s_9s_9_2_1_Adder_6_U.u1.b ;
wire \add_9s_9s_9_2_1_U8.top_add_9s_9s_9_2_1_Adder_6_U.u1.cin ;
wire \add_9s_9s_9_2_1_U8.top_add_9s_9s_9_2_1_Adder_6_U.u1.cout ;
wire [3:0] \add_9s_9s_9_2_1_U8.top_add_9s_9s_9_2_1_Adder_6_U.u1.s ;
wire [4:0] \add_9s_9s_9_2_1_U8.top_add_9s_9s_9_2_1_Adder_6_U.u2.a ;
wire [4:0] \add_9s_9s_9_2_1_U8.top_add_9s_9s_9_2_1_Adder_6_U.u2.b ;
wire \add_9s_9s_9_2_1_U8.top_add_9s_9s_9_2_1_Adder_6_U.u2.cin ;
wire \add_9s_9s_9_2_1_U8.top_add_9s_9s_9_2_1_Adder_6_U.u2.cout ;
wire [4:0] \add_9s_9s_9_2_1_U8.top_add_9s_9s_9_2_1_Adder_6_U.u2.s ;
wire and_ln340_fu_768_p2;
wire and_ln406_fu_538_p2;
wire and_ln408_fu_889_p2;
wire and_ln780_fu_637_p2;
wire and_ln781_fu_658_p2;
wire and_ln785_1_fu_703_p2;
wire and_ln785_2_fu_759_p2;
wire and_ln785_fu_694_p2;
wire and_ln786_fu_653_p2;
wire and_ln850_fu_1027_p2;
wire ap_CS_fsm_state1;
wire ap_CS_fsm_state10;
wire ap_CS_fsm_state11;
wire ap_CS_fsm_state12;
wire ap_CS_fsm_state13;
wire ap_CS_fsm_state14;
wire ap_CS_fsm_state15;
wire ap_CS_fsm_state16;
wire ap_CS_fsm_state17;
wire ap_CS_fsm_state18;
wire ap_CS_fsm_state19;
wire ap_CS_fsm_state2;
wire ap_CS_fsm_state20;
wire ap_CS_fsm_state21;
wire ap_CS_fsm_state22;
wire ap_CS_fsm_state23;
wire ap_CS_fsm_state24;
wire ap_CS_fsm_state25;
wire ap_CS_fsm_state26;
wire ap_CS_fsm_state27;
wire ap_CS_fsm_state28;
wire ap_CS_fsm_state29;
wire ap_CS_fsm_state3;
wire ap_CS_fsm_state30;
wire ap_CS_fsm_state31;
wire ap_CS_fsm_state32;
wire ap_CS_fsm_state33;
wire ap_CS_fsm_state34;
wire ap_CS_fsm_state35;
wire ap_CS_fsm_state36;
wire ap_CS_fsm_state37;
wire ap_CS_fsm_state38;
wire ap_CS_fsm_state39;
wire ap_CS_fsm_state4;
wire ap_CS_fsm_state40;
wire ap_CS_fsm_state41;
wire ap_CS_fsm_state42;
wire ap_CS_fsm_state43;
wire ap_CS_fsm_state44;
wire ap_CS_fsm_state45;
wire ap_CS_fsm_state46;
wire ap_CS_fsm_state47;
wire ap_CS_fsm_state48;
wire ap_CS_fsm_state49;
wire ap_CS_fsm_state5;
wire ap_CS_fsm_state50;
wire ap_CS_fsm_state51;
wire ap_CS_fsm_state52;
wire ap_CS_fsm_state53;
wire ap_CS_fsm_state54;
wire ap_CS_fsm_state55;
wire ap_CS_fsm_state56;
wire ap_CS_fsm_state57;
wire ap_CS_fsm_state6;
wire ap_CS_fsm_state7;
wire ap_CS_fsm_state8;
wire ap_CS_fsm_state9;
wire [56:0] ap_NS_fsm;
wire ap_clk;
wire ap_done;
wire ap_idle;
wire ap_ready;
wire ap_rst;
wire ap_start;
wire carry_2_fu_623_p2;
wire deleted_ones_fu_642_p3;
wire deleted_zeros_fu_627_p3;
wire [31:0] grp_fu_1003_p2;
wire [31:0] grp_fu_1147_p1;
wire [31:0] grp_fu_1147_p2;
wire [31:0] grp_fu_1187_p2;
wire [33:0] grp_fu_1206_p0;
wire [33:0] grp_fu_1206_p1;
wire [33:0] grp_fu_1206_p2;
wire [31:0] grp_fu_1222_p2;
wire [33:0] grp_fu_1265_p0;
wire [33:0] grp_fu_1265_p1;
wire [33:0] grp_fu_1265_p2;
wire [31:0] grp_fu_1281_p2;
wire [31:0] grp_fu_1317_p1;
wire [31:0] grp_fu_1317_p2;
wire [34:0] grp_fu_1337_p0;
wire [34:0] grp_fu_1337_p1;
wire [34:0] grp_fu_1337_p2;
wire [31:0] grp_fu_1363_p2;
wire [31:0] grp_fu_1391_p1;
wire [31:0] grp_fu_1391_p2;
wire [4:0] grp_fu_265_p1;
wire [4:0] grp_fu_265_p2;
wire [1:0] grp_fu_286_p2;
wire [16:0] grp_fu_324_p1;
wire [16:0] grp_fu_324_p2;
wire [15:0] grp_fu_336_p0;
wire [19:0] grp_fu_336_p00;
wire [19:0] grp_fu_336_p2;
wire [8:0] grp_fu_517_p0;
wire [8:0] grp_fu_517_p2;
wire [3:0] grp_fu_576_p1;
wire [3:0] grp_fu_576_p2;
wire [5:0] grp_fu_586_p2;
wire [8:0] grp_fu_809_p0;
wire [8:0] grp_fu_809_p1;
wire [8:0] grp_fu_809_p2;
wire [3:0] grp_fu_815_p0;
wire [3:0] grp_fu_815_p1;
wire [3:0] grp_fu_815_p2;
wire [7:0] grp_fu_868_p0;
wire [7:0] grp_fu_868_p1;
wire [7:0] grp_fu_868_p2;
wire [7:0] grp_fu_896_p0;
wire [7:0] grp_fu_896_p2;
wire [5:0] grp_fu_908_p0;
wire [5:0] grp_fu_908_p1;
wire [5:0] grp_fu_908_p2;
wire [33:0] grp_fu_951_p0;
wire [33:0] grp_fu_951_p1;
wire [33:0] grp_fu_951_p2;
wire [31:0] grp_fu_967_p2;
wire icmp_ln1497_fu_1138_p2;
wire icmp_ln768_fu_372_p2;
wire icmp_ln786_fu_377_p2;
wire icmp_ln790_fu_389_p2;
wire icmp_ln851_1_fu_581_p2;
wire icmp_ln851_2_fu_1347_p2;
wire icmp_ln851_fu_270_p2;
wire lhs_V_2_fu_1093_p2;
wire [3:0] lhs_fu_785_p1;
wire [5:0] lhs_fu_785_p3;
wire \mul_16ns_4s_20_7_1_U4.ce ;
wire \mul_16ns_4s_20_7_1_U4.clk ;
wire [15:0] \mul_16ns_4s_20_7_1_U4.din0 ;
wire [3:0] \mul_16ns_4s_20_7_1_U4.din1 ;
wire [19:0] \mul_16ns_4s_20_7_1_U4.dout ;
wire \mul_16ns_4s_20_7_1_U4.reset ;
wire [15:0] \mul_16ns_4s_20_7_1_U4.top_mul_16ns_4s_20_7_1_Mul_DSP_0_U.a ;
wire [3:0] \mul_16ns_4s_20_7_1_U4.top_mul_16ns_4s_20_7_1_Mul_DSP_0_U.b ;
wire \mul_16ns_4s_20_7_1_U4.top_mul_16ns_4s_20_7_1_Mul_DSP_0_U.ce ;
wire \mul_16ns_4s_20_7_1_U4.top_mul_16ns_4s_20_7_1_Mul_DSP_0_U.clk ;
wire [19:0] \mul_16ns_4s_20_7_1_U4.top_mul_16ns_4s_20_7_1_Mul_DSP_0_U.p ;
wire [19:0] \mul_16ns_4s_20_7_1_U4.top_mul_16ns_4s_20_7_1_Mul_DSP_0_U.tmp_product ;
wire neg_src_2_fu_1152_p2;
wire neg_src_fu_668_p2;
wire newsignbit_fu_1123_p2;
wire op_0;
wire [1:0] op_11_V_fu_1127_p3;
wire op_12;
wire op_14_V_fu_1174_p2;
wire [3:0] op_15;
wire [15:0] op_16;
wire [3:0] op_18;
wire [3:0] op_19;
wire op_2;
wire [3:0] op_3;
wire [31:0] op_30;
wire op_30_ap_vld;
wire [1:0] op_5;
wire [7:0] op_6;
wire [3:0] op_7;
wire [7:0] op_8_V_fu_453_p3;
wire [3:0] op_9_V_fu_826_p3;
wire or_ln340_1_fu_748_p2;
wire or_ln340_2_fu_773_p2;
wire or_ln340_fu_688_p2;
wire or_ln384_fu_430_p2;
wire or_ln406_fu_533_p2;
wire or_ln785_1_fu_678_p2;
wire or_ln785_2_fu_698_p2;
wire or_ln785_fu_395_p2;
wire or_ln788_1_fu_420_p2;
wire or_ln788_fu_415_p2;
wire overflow_1_fu_683_p2;
wire overflow_fu_404_p2;
wire [3:0] p_Result_14_fu_739_p4;
wire p_Result_15_fu_604_p3;
wire p_Result_16_fu_914_p3;
wire p_Result_17_fu_972_p3;
wire p_Result_18_fu_1227_p3;
wire p_Result_19_fu_1291_p3;
wire [1:0] p_Result_1_fu_1015_p1;
wire p_Result_1_fu_1015_p3;
wire p_Result_20_fu_1368_p3;
wire p_Result_26_fu_523_p3;
wire [6:0] p_Result_3_fu_382_p3;
wire p_Result_s_fu_291_p3;
wire [7:0] p_Val2_4_fu_438_p3;
wire [2:0] p_Val2_8_fu_734_p2;
wire r_1_fu_530_p1;
wire [1:0] r_V_fu_1053_p2;
wire [1:0] r_V_fu_1053_p3;
wire r_fu_874_p2;
wire [1:0] ret_V_21_fu_303_p3;
wire ret_V_22_fu_1033_p2;
wire [31:0] ret_V_27_fu_988_p3;
wire [31:0] ret_V_32_fu_1307_p3;
wire [31:0] ret_V_34_fu_1380_p3;
wire [1:0] ret_V_4_fu_1007_p1;
wire ret_V_4_fu_1007_p3;
wire [6:0] rhs_2_fu_857_p3;
wire [32:0] rhs_6_fu_1195_p3;
wire [32:0] rhs_7_fu_1254_p3;
wire [33:0] rhs_9_fu_1326_p3;
wire sel_tmp11_fu_779_p2;
wire [31:0] select_ln1192_fu_1179_p3;
wire [16:0] select_ln1347_fu_310_p3;
wire [3:0] select_ln340_1_fu_752_p3;
wire select_ln340_fu_1161_p3;
wire [31:0] select_ln353_2_fu_1243_p3;
wire [7:0] select_ln353_fu_930_p3;
wire [7:0] select_ln384_fu_446_p3;
wire [31:0] select_ln69_fu_995_p3;
wire [4:0] select_ln703_fu_249_p3;
wire [3:0] select_ln785_fu_821_p3;
wire [5:0] select_ln850_2_fu_611_p3;
wire [31:0] select_ln850_3_fu_982_p3;
wire [5:0] select_ln850_4_fu_616_p3;
wire [31:0] select_ln850_5_fu_1301_p3;
wire [31:0] select_ln850_6_fu_1375_p3;
wire [7:0] select_ln850_7_fu_924_p3;
wire [31:0] select_ln850_8_fu_1237_p3;
wire [1:0] select_ln850_fu_298_p3;
wire [1:0] sext_ln1299_1_fu_1039_p0;
wire [17:0] sext_ln1299_1_fu_1039_p1;
wire [1:0] sext_ln1299_2_fu_1043_p0;
wire [5:0] sext_ln1299_2_fu_1043_p1;
wire [1:0] sext_ln1299_fu_1120_p0;
wire [2:0] sext_ln1299_fu_1120_p1;
wire [15:0] sext_ln1347_fu_317_p1;
wire [16:0] sext_ln1499_fu_1106_p1;
wire [7:0] sext_ln703_1_fu_796_p0;
wire [3:0] sext_ln703_4_fu_1191_p0;
wire [15:0] sext_ln703_5_fu_1250_p0;
wire [3:0] sext_ln703_6_fu_1322_p0;
wire [3:0] sext_ln703_fu_257_p0;
wire [7:0] sext_ln850_fu_893_p1;
wire [3:0] shl_ln1192_fu_804_p0;
wire [1:0] shl_ln1299_fu_1047_p0;
wire [1:0] shl_ln1299_fu_1047_p2;
wire [4:0] shl_ln1_fu_1081_p3;
wire signbit_3_fu_1114_p2;
wire \sub_17ns_17ns_17_2_1_U3.ce ;
wire \sub_17ns_17ns_17_2_1_U3.clk ;
wire [16:0] \sub_17ns_17ns_17_2_1_U3.din0 ;
wire [16:0] \sub_17ns_17ns_17_2_1_U3.din1 ;
wire [16:0] \sub_17ns_17ns_17_2_1_U3.dout ;
wire \sub_17ns_17ns_17_2_1_U3.reset ;
wire [16:0] \sub_17ns_17ns_17_2_1_U3.top_sub_17ns_17ns_17_2_1_Adder_2_U.a ;
wire [16:0] \sub_17ns_17ns_17_2_1_U3.top_sub_17ns_17ns_17_2_1_Adder_2_U.ain_s0 ;
wire [16:0] \sub_17ns_17ns_17_2_1_U3.top_sub_17ns_17ns_17_2_1_Adder_2_U.b ;
wire [16:0] \sub_17ns_17ns_17_2_1_U3.top_sub_17ns_17ns_17_2_1_Adder_2_U.bin_s0 ;
wire \sub_17ns_17ns_17_2_1_U3.top_sub_17ns_17ns_17_2_1_Adder_2_U.ce ;
wire \sub_17ns_17ns_17_2_1_U3.top_sub_17ns_17ns_17_2_1_Adder_2_U.clk ;
wire \sub_17ns_17ns_17_2_1_U3.top_sub_17ns_17ns_17_2_1_Adder_2_U.facout_s1 ;
wire \sub_17ns_17ns_17_2_1_U3.top_sub_17ns_17ns_17_2_1_Adder_2_U.facout_s2 ;
wire [7:0] \sub_17ns_17ns_17_2_1_U3.top_sub_17ns_17ns_17_2_1_Adder_2_U.fas_s1 ;
wire [8:0] \sub_17ns_17ns_17_2_1_U3.top_sub_17ns_17ns_17_2_1_Adder_2_U.fas_s2 ;
wire \sub_17ns_17ns_17_2_1_U3.top_sub_17ns_17ns_17_2_1_Adder_2_U.reset ;
wire [16:0] \sub_17ns_17ns_17_2_1_U3.top_sub_17ns_17ns_17_2_1_Adder_2_U.s ;
wire [7:0] \sub_17ns_17ns_17_2_1_U3.top_sub_17ns_17ns_17_2_1_Adder_2_U.u1.a ;
wire [7:0] \sub_17ns_17ns_17_2_1_U3.top_sub_17ns_17ns_17_2_1_Adder_2_U.u1.b ;
wire \sub_17ns_17ns_17_2_1_U3.top_sub_17ns_17ns_17_2_1_Adder_2_U.u1.cin ;
wire \sub_17ns_17ns_17_2_1_U3.top_sub_17ns_17ns_17_2_1_Adder_2_U.u1.cout ;
wire [7:0] \sub_17ns_17ns_17_2_1_U3.top_sub_17ns_17ns_17_2_1_Adder_2_U.u1.s ;
wire [8:0] \sub_17ns_17ns_17_2_1_U3.top_sub_17ns_17ns_17_2_1_Adder_2_U.u2.a ;
wire [8:0] \sub_17ns_17ns_17_2_1_U3.top_sub_17ns_17ns_17_2_1_Adder_2_U.u2.b ;
wire \sub_17ns_17ns_17_2_1_U3.top_sub_17ns_17ns_17_2_1_Adder_2_U.u2.cin ;
wire \sub_17ns_17ns_17_2_1_U3.top_sub_17ns_17ns_17_2_1_Adder_2_U.u2.cout ;
wire [8:0] \sub_17ns_17ns_17_2_1_U3.top_sub_17ns_17ns_17_2_1_Adder_2_U.u2.s ;
wire tmp_1_fu_715_p3;
wire [2:0] tmp_7_fu_1099_p3;
wire [8:0] tmp_8_fu_940_p3;
wire tmp_fu_708_p3;
wire [7:0] trunc_ln1192_1_fu_800_p0;
wire [3:0] trunc_ln1192_fu_261_p0;
wire [2:0] trunc_ln1192_fu_261_p1;
wire trunc_ln415_fu_1061_p1;
wire [2:0] trunc_ln718_fu_850_p1;
wire [4:0] trunc_ln731_fu_435_p1;
wire [3:0] trunc_ln790_fu_368_p1;
wire [2:0] trunc_ln851_1_fu_569_p1;
wire trunc_ln851_2_fu_921_p1;
wire trunc_ln851_3_fu_979_p1;
wire [3:0] trunc_ln851_4_fu_1234_p0;
wire trunc_ln851_4_fu_1234_p1;
wire [15:0] trunc_ln851_5_fu_1298_p0;
wire trunc_ln851_5_fu_1298_p1;
wire [3:0] trunc_ln851_6_fu_1343_p0;
wire [1:0] trunc_ln851_6_fu_1343_p1;
wire [1:0] trunc_ln851_fu_1023_p0;
wire trunc_ln851_fu_1023_p1;
wire underflow_fu_425_p2;
wire xor_ln1497_fu_1286_p2;
wire xor_ln340_fu_1168_p2;
wire xor_ln365_1_fu_728_p2;
wire xor_ln365_fu_722_p2;
wire xor_ln416_fu_599_p2;
wire xor_ln780_fu_632_p2;
wire xor_ln781_fu_662_p2;
wire xor_ln785_1_fu_399_p2;
wire xor_ln785_2_fu_673_p2;
wire xor_ln785_3_fu_648_p2;
wire xor_ln785_fu_1156_p2;
wire xor_ln786_1_fu_763_p2;
wire xor_ln786_fu_410_p2;
wire [2:0] zext_ln1497_fu_1134_p1;
wire [17:0] zext_ln1499_1_fu_1110_p1;
wire [5:0] zext_ln1499_fu_1089_p1;


assign _091_ = icmp_ln851_2_reg_2010 & ap_CS_fsm[53];
assign _092_ = ap_CS_fsm[4] & _096_;
assign _093_ = ap_CS_fsm[20] & _097_;
assign _094_ = _098_ & ap_CS_fsm[0];
assign _095_ = ap_start & ap_CS_fsm[0];
assign and_ln340_fu_768_p2 = xor_ln786_1_fu_763_p2 & or_ln340_reg_1681;
assign and_ln406_fu_538_p2 = r_V_1_reg_1526[1] & or_ln406_fu_533_p2;
assign and_ln408_fu_889_p2 = r_reg_1753 & p_Result_22_reg_1733;
assign and_ln780_fu_637_p2 = xor_ln780_fu_632_p2 & Range2_all_ones_reg_1578;
assign and_ln781_fu_658_p2 = carry_2_reg_1654 & Range1_all_ones_reg_1583;
assign and_ln785_1_fu_703_p2 = or_ln785_2_fu_698_p2 & and_ln786_reg_1673;
assign and_ln785_2_fu_759_p2 = xor_ln785_3_reg_1667 & and_ln786_reg_1673;
assign and_ln785_fu_694_p2 = xor_ln416_reg_1643 & deleted_zeros_reg_1661;
assign and_ln786_fu_653_p2 = p_Result_28_reg_1631 & deleted_ones_fu_642_p3;
assign and_ln850_fu_1027_p2 = op_5[0] & op_5[1];
assign carry_2_fu_623_p2 = xor_ln416_reg_1643 & p_Result_27_reg_1546;
assign neg_src_2_fu_1152_p2 = p_Result_21_reg_1853 & newsignbit_reg_1879;
assign neg_src_fu_668_p2 = xor_ln781_fu_662_p2 & p_Result_25_reg_1533;
assign op_14_V_fu_1174_p2 = xor_ln340_fu_1168_p2 & newsignbit_reg_1879;
assign overflow_1_fu_683_p2 = xor_ln785_3_reg_1667 & or_ln785_1_fu_678_p2;
assign overflow_fu_404_p2 = xor_ln785_1_fu_399_p2 & or_ln785_fu_395_p2;
assign sel_tmp11_fu_779_p2 = xor_ln365_1_fu_728_p2 & or_ln340_2_fu_773_p2;
assign underflow_fu_425_p2 = p_Result_23_reg_1472 & or_ln788_1_fu_420_p2;
assign xor_ln786_1_fu_763_p2 = ~ and_ln786_reg_1673;
assign xor_ln780_fu_632_p2 = ~ p_Result_29_reg_1551;
assign xor_ln781_fu_662_p2 = ~ and_ln781_fu_658_p2;
assign xor_ln785_fu_1156_p2 = ~ p_Result_21_reg_1853;
assign xor_ln340_fu_1168_p2 = ~ select_ln340_fu_1161_p3;
assign xor_ln785_2_fu_673_p2 = ~ deleted_zeros_reg_1661;
assign xor_ln786_fu_410_p2 = ~ p_Result_24_reg_1478;
assign xor_ln785_1_fu_399_p2 = ~ p_Result_23_reg_1472;
assign xor_ln365_1_fu_728_p2 = ~ xor_ln365_fu_722_p2;
assign xor_ln1497_fu_1286_p2 = ~ icmp_ln1497_reg_1886;
assign xor_ln416_fu_599_p2 = ~ p_Result_28_reg_1631;
assign xor_ln785_3_fu_648_p2 = ~ p_Result_25_reg_1533;
assign p_Val2_8_fu_734_p2 = ~ p_Val2_7_reg_1622[2:0];
assign _096_ = ~ icmp_ln851_reg_1419;
assign _097_ = ~ and_ln785_1_reg_1687;
assign _098_ = ~ ap_start;
assign _099_ = p_Result_7_reg_1562 == 14'h3fff;
assign _100_ = ! p_Result_7_reg_1562;
assign _101_ = p_Result_6_reg_1557 == 13'h1fff;
assign _102_ = ! { trunc_ln790_reg_1490, 3'h0 };
assign _103_ = ! trunc_ln851_1_reg_1607;
assign _104_ = ! op_3[2:0];
always @(posedge \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.clk )
\add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.bin_s1  <= _106_;
always @(posedge \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.clk )
\add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.ain_s1  <= _105_;
always @(posedge \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.clk )
\add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.sum_s1  <= _108_;
always @(posedge \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.clk )
\add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.carry_s1  <= _107_;
assign _106_ = \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.ce  ? \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.b [1] : \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.bin_s1 ;
assign _105_ = \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.ce  ? \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.a [1] : \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.ain_s1 ;
assign _107_ = \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.ce  ? \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.facout_s1  : \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.carry_s1 ;
assign _108_ = \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.ce  ? \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.fas_s1  : \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.sum_s1 ;
assign _109_ = \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.a  + \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.b ;
assign { \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.cout , \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.s  } = _109_ + \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.cin ;
assign _110_ = \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.a  + \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.b ;
assign { \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.cout , \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.s  } = _110_ + \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.cin ;
always @(posedge \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.clk )
\add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.bin_s1  <= _112_;
always @(posedge \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.clk )
\add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.ain_s1  <= _111_;
always @(posedge \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.clk )
\add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.sum_s1  <= _114_;
always @(posedge \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.clk )
\add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.carry_s1  <= _113_;
assign _112_ = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.ce  ? \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.b [31:16] : \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.bin_s1 ;
assign _111_ = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.ce  ? \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.a [31:16] : \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.ain_s1 ;
assign _113_ = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.ce  ? \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.facout_s1  : \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.carry_s1 ;
assign _114_ = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.ce  ? \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.fas_s1  : \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.sum_s1 ;
assign _115_ = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.a  + \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.b ;
assign { \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.cout , \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.s  } = _115_ + \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.cin ;
assign _116_ = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.a  + \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.b ;
assign { \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.cout , \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.s  } = _116_ + \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.cin ;
always @(posedge \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.clk )
\add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.bin_s1  <= _118_;
always @(posedge \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.clk )
\add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.ain_s1  <= _117_;
always @(posedge \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.clk )
\add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.sum_s1  <= _120_;
always @(posedge \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.clk )
\add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.carry_s1  <= _119_;
assign _118_ = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.ce  ? \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.b [31:16] : \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.bin_s1 ;
assign _117_ = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.ce  ? \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.a [31:16] : \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.ain_s1 ;
assign _119_ = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.ce  ? \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.facout_s1  : \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.carry_s1 ;
assign _120_ = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.ce  ? \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.fas_s1  : \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.sum_s1 ;
assign _121_ = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.a  + \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.b ;
assign { \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.cout , \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.s  } = _121_ + \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.cin ;
assign _122_ = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.a  + \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.b ;
assign { \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.cout , \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.s  } = _122_ + \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.cin ;
always @(posedge \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.clk )
\add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.bin_s1  <= _124_;
always @(posedge \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.clk )
\add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.ain_s1  <= _123_;
always @(posedge \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.clk )
\add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.sum_s1  <= _126_;
always @(posedge \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.clk )
\add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.carry_s1  <= _125_;
assign _124_ = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.ce  ? \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.b [31:16] : \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.bin_s1 ;
assign _123_ = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.ce  ? \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.a [31:16] : \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.ain_s1 ;
assign _125_ = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.ce  ? \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.facout_s1  : \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.carry_s1 ;
assign _126_ = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.ce  ? \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.fas_s1  : \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.sum_s1 ;
assign _127_ = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.a  + \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.b ;
assign { \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.cout , \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.s  } = _127_ + \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.cin ;
assign _128_ = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.a  + \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.b ;
assign { \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.cout , \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.s  } = _128_ + \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.cin ;
always @(posedge \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.clk )
\add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.bin_s1  <= _130_;
always @(posedge \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.clk )
\add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.ain_s1  <= _129_;
always @(posedge \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.clk )
\add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.sum_s1  <= _132_;
always @(posedge \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.clk )
\add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.carry_s1  <= _131_;
assign _130_ = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.ce  ? \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.b [31:16] : \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.bin_s1 ;
assign _129_ = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.ce  ? \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.a [31:16] : \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.ain_s1 ;
assign _131_ = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.ce  ? \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.facout_s1  : \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.carry_s1 ;
assign _132_ = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.ce  ? \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.fas_s1  : \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.sum_s1 ;
assign _133_ = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.a  + \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.b ;
assign { \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.cout , \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.s  } = _133_ + \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.cin ;
assign _134_ = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.a  + \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.b ;
assign { \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.cout , \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.s  } = _134_ + \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.cin ;
always @(posedge \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.clk )
\add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.bin_s1  <= _136_;
always @(posedge \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.clk )
\add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.ain_s1  <= _135_;
always @(posedge \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.clk )
\add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.sum_s1  <= _138_;
always @(posedge \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.clk )
\add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.carry_s1  <= _137_;
assign _136_ = \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.ce  ? \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.b [31:16] : \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.bin_s1 ;
assign _135_ = \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.ce  ? \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.a [31:16] : \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.ain_s1 ;
assign _137_ = \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.ce  ? \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.facout_s1  : \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.carry_s1 ;
assign _138_ = \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.ce  ? \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.fas_s1  : \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.sum_s1 ;
assign _139_ = \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.a  + \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.b ;
assign { \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.cout , \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.s  } = _139_ + \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.cin ;
assign _140_ = \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.a  + \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.b ;
assign { \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.cout , \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.s  } = _140_ + \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.cin ;
always @(posedge \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.clk )
\add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.bin_s1  <= _142_;
always @(posedge \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.clk )
\add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.ain_s1  <= _141_;
always @(posedge \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.clk )
\add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.sum_s1  <= _144_;
always @(posedge \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.clk )
\add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.carry_s1  <= _143_;
assign _142_ = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.ce  ? \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.b [31:16] : \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.bin_s1 ;
assign _141_ = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.ce  ? \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.a [31:16] : \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.ain_s1 ;
assign _143_ = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.ce  ? \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.facout_s1  : \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.carry_s1 ;
assign _144_ = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.ce  ? \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.fas_s1  : \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.sum_s1 ;
assign _145_ = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.a  + \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.b ;
assign { \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.cout , \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.s  } = _145_ + \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.cin ;
assign _146_ = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.a  + \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.b ;
assign { \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.cout , \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.s  } = _146_ + \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.cin ;
always @(posedge \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_11_U.clk )
\add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_11_U.bin_s1  <= _148_;
always @(posedge \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_11_U.clk )
\add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_11_U.ain_s1  <= _147_;
always @(posedge \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_11_U.clk )
\add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_11_U.sum_s1  <= _150_;
always @(posedge \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_11_U.clk )
\add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_11_U.carry_s1  <= _149_;
assign _148_ = \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_11_U.ce  ? \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_11_U.b [31:16] : \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_11_U.bin_s1 ;
assign _147_ = \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_11_U.ce  ? \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_11_U.a [31:16] : \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_11_U.ain_s1 ;
assign _149_ = \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_11_U.ce  ? \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_11_U.facout_s1  : \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_11_U.carry_s1 ;
assign _150_ = \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_11_U.ce  ? \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_11_U.fas_s1  : \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_11_U.sum_s1 ;
assign _151_ = \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.a  + \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.b ;
assign { \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.cout , \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.s  } = _151_ + \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.cin ;
assign _152_ = \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.a  + \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.b ;
assign { \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.cout , \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.s  } = _152_ + \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.cin ;
always @(posedge \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_11_U.clk )
\add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_11_U.bin_s1  <= _154_;
always @(posedge \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_11_U.clk )
\add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_11_U.ain_s1  <= _153_;
always @(posedge \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_11_U.clk )
\add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_11_U.sum_s1  <= _156_;
always @(posedge \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_11_U.clk )
\add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_11_U.carry_s1  <= _155_;
assign _154_ = \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_11_U.ce  ? \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_11_U.b [31:16] : \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_11_U.bin_s1 ;
assign _153_ = \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_11_U.ce  ? \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_11_U.a [31:16] : \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_11_U.ain_s1 ;
assign _155_ = \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_11_U.ce  ? \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_11_U.facout_s1  : \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_11_U.carry_s1 ;
assign _156_ = \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_11_U.ce  ? \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_11_U.fas_s1  : \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_11_U.sum_s1 ;
assign _157_ = \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.a  + \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.b ;
assign { \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.cout , \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.s  } = _157_ + \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.cin ;
assign _158_ = \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.a  + \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.b ;
assign { \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.cout , \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.s  } = _158_ + \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.cin ;
always @(posedge \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_11_U.clk )
\add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_11_U.bin_s1  <= _160_;
always @(posedge \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_11_U.clk )
\add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_11_U.ain_s1  <= _159_;
always @(posedge \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_11_U.clk )
\add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_11_U.sum_s1  <= _162_;
always @(posedge \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_11_U.clk )
\add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_11_U.carry_s1  <= _161_;
assign _160_ = \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_11_U.ce  ? \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_11_U.b [31:16] : \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_11_U.bin_s1 ;
assign _159_ = \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_11_U.ce  ? \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_11_U.a [31:16] : \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_11_U.ain_s1 ;
assign _161_ = \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_11_U.ce  ? \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_11_U.facout_s1  : \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_11_U.carry_s1 ;
assign _162_ = \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_11_U.ce  ? \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_11_U.fas_s1  : \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_11_U.sum_s1 ;
assign _163_ = \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.a  + \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.b ;
assign { \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.cout , \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.s  } = _163_ + \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.cin ;
assign _164_ = \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.a  + \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.b ;
assign { \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.cout , \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.s  } = _164_ + \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.cin ;
always @(posedge \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_10_U.clk )
\add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_10_U.bin_s1  <= _166_;
always @(posedge \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_10_U.clk )
\add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_10_U.ain_s1  <= _165_;
always @(posedge \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_10_U.clk )
\add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_10_U.sum_s1  <= _168_;
always @(posedge \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_10_U.clk )
\add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_10_U.carry_s1  <= _167_;
assign _166_ = \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_10_U.ce  ? \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_10_U.b [33:17] : \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_10_U.bin_s1 ;
assign _165_ = \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_10_U.ce  ? \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_10_U.a [33:17] : \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_10_U.ain_s1 ;
assign _167_ = \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_10_U.ce  ? \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_10_U.facout_s1  : \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_10_U.carry_s1 ;
assign _168_ = \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_10_U.ce  ? \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_10_U.fas_s1  : \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_10_U.sum_s1 ;
assign _169_ = \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_10_U.u1.a  + \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_10_U.u1.b ;
assign { \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_10_U.u1.cout , \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_10_U.u1.s  } = _169_ + \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_10_U.u1.cin ;
assign _170_ = \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_10_U.u2.a  + \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_10_U.u2.b ;
assign { \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_10_U.u2.cout , \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_10_U.u2.s  } = _170_ + \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_10_U.u2.cin ;
always @(posedge \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_10_U.clk )
\add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_10_U.bin_s1  <= _172_;
always @(posedge \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_10_U.clk )
\add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_10_U.ain_s1  <= _171_;
always @(posedge \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_10_U.clk )
\add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_10_U.sum_s1  <= _174_;
always @(posedge \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_10_U.clk )
\add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_10_U.carry_s1  <= _173_;
assign _172_ = \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_10_U.ce  ? \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_10_U.b [33:17] : \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_10_U.bin_s1 ;
assign _171_ = \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_10_U.ce  ? \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_10_U.a [33:17] : \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_10_U.ain_s1 ;
assign _173_ = \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_10_U.ce  ? \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_10_U.facout_s1  : \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_10_U.carry_s1 ;
assign _174_ = \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_10_U.ce  ? \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_10_U.fas_s1  : \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_10_U.sum_s1 ;
assign _175_ = \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_10_U.u1.a  + \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_10_U.u1.b ;
assign { \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_10_U.u1.cout , \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_10_U.u1.s  } = _175_ + \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_10_U.u1.cin ;
assign _176_ = \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_10_U.u2.a  + \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_10_U.u2.b ;
assign { \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_10_U.u2.cout , \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_10_U.u2.s  } = _176_ + \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_10_U.u2.cin ;
always @(posedge \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_10_U.clk )
\add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_10_U.bin_s1  <= _178_;
always @(posedge \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_10_U.clk )
\add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_10_U.ain_s1  <= _177_;
always @(posedge \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_10_U.clk )
\add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_10_U.sum_s1  <= _180_;
always @(posedge \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_10_U.clk )
\add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_10_U.carry_s1  <= _179_;
assign _178_ = \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_10_U.ce  ? \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_10_U.b [33:17] : \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_10_U.bin_s1 ;
assign _177_ = \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_10_U.ce  ? \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_10_U.a [33:17] : \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_10_U.ain_s1 ;
assign _179_ = \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_10_U.ce  ? \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_10_U.facout_s1  : \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_10_U.carry_s1 ;
assign _180_ = \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_10_U.ce  ? \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_10_U.fas_s1  : \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_10_U.sum_s1 ;
assign _181_ = \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_10_U.u1.a  + \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_10_U.u1.b ;
assign { \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_10_U.u1.cout , \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_10_U.u1.s  } = _181_ + \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_10_U.u1.cin ;
assign _182_ = \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_10_U.u2.a  + \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_10_U.u2.b ;
assign { \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_10_U.u2.cout , \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_10_U.u2.s  } = _182_ + \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_10_U.u2.cin ;
always @(posedge \add_35s_35s_35_2_1_U23.top_add_35s_35s_35_2_1_Adder_12_U.clk )
\add_35s_35s_35_2_1_U23.top_add_35s_35s_35_2_1_Adder_12_U.bin_s1  <= _184_;
always @(posedge \add_35s_35s_35_2_1_U23.top_add_35s_35s_35_2_1_Adder_12_U.clk )
\add_35s_35s_35_2_1_U23.top_add_35s_35s_35_2_1_Adder_12_U.ain_s1  <= _183_;
always @(posedge \add_35s_35s_35_2_1_U23.top_add_35s_35s_35_2_1_Adder_12_U.clk )
\add_35s_35s_35_2_1_U23.top_add_35s_35s_35_2_1_Adder_12_U.sum_s1  <= _186_;
always @(posedge \add_35s_35s_35_2_1_U23.top_add_35s_35s_35_2_1_Adder_12_U.clk )
\add_35s_35s_35_2_1_U23.top_add_35s_35s_35_2_1_Adder_12_U.carry_s1  <= _185_;
assign _184_ = \add_35s_35s_35_2_1_U23.top_add_35s_35s_35_2_1_Adder_12_U.ce  ? \add_35s_35s_35_2_1_U23.top_add_35s_35s_35_2_1_Adder_12_U.b [34:17] : \add_35s_35s_35_2_1_U23.top_add_35s_35s_35_2_1_Adder_12_U.bin_s1 ;
assign _183_ = \add_35s_35s_35_2_1_U23.top_add_35s_35s_35_2_1_Adder_12_U.ce  ? \add_35s_35s_35_2_1_U23.top_add_35s_35s_35_2_1_Adder_12_U.a [34:17] : \add_35s_35s_35_2_1_U23.top_add_35s_35s_35_2_1_Adder_12_U.ain_s1 ;
assign _185_ = \add_35s_35s_35_2_1_U23.top_add_35s_35s_35_2_1_Adder_12_U.ce  ? \add_35s_35s_35_2_1_U23.top_add_35s_35s_35_2_1_Adder_12_U.facout_s1  : \add_35s_35s_35_2_1_U23.top_add_35s_35s_35_2_1_Adder_12_U.carry_s1 ;
assign _186_ = \add_35s_35s_35_2_1_U23.top_add_35s_35s_35_2_1_Adder_12_U.ce  ? \add_35s_35s_35_2_1_U23.top_add_35s_35s_35_2_1_Adder_12_U.fas_s1  : \add_35s_35s_35_2_1_U23.top_add_35s_35s_35_2_1_Adder_12_U.sum_s1 ;
assign _187_ = \add_35s_35s_35_2_1_U23.top_add_35s_35s_35_2_1_Adder_12_U.u1.a  + \add_35s_35s_35_2_1_U23.top_add_35s_35s_35_2_1_Adder_12_U.u1.b ;
assign { \add_35s_35s_35_2_1_U23.top_add_35s_35s_35_2_1_Adder_12_U.u1.cout , \add_35s_35s_35_2_1_U23.top_add_35s_35s_35_2_1_Adder_12_U.u1.s  } = _187_ + \add_35s_35s_35_2_1_U23.top_add_35s_35s_35_2_1_Adder_12_U.u1.cin ;
assign _188_ = \add_35s_35s_35_2_1_U23.top_add_35s_35s_35_2_1_Adder_12_U.u2.a  + \add_35s_35s_35_2_1_U23.top_add_35s_35s_35_2_1_Adder_12_U.u2.b ;
assign { \add_35s_35s_35_2_1_U23.top_add_35s_35s_35_2_1_Adder_12_U.u2.cout , \add_35s_35s_35_2_1_U23.top_add_35s_35s_35_2_1_Adder_12_U.u2.s  } = _188_ + \add_35s_35s_35_2_1_U23.top_add_35s_35s_35_2_1_Adder_12_U.u2.cin ;
always @(posedge \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.clk )
\add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.bin_s1  <= _190_;
always @(posedge \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.clk )
\add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.ain_s1  <= _189_;
always @(posedge \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.clk )
\add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.sum_s1  <= _192_;
always @(posedge \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.clk )
\add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.carry_s1  <= _191_;
assign _190_ = \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.ce  ? \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.b [3:2] : \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.bin_s1 ;
assign _189_ = \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.ce  ? \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.a [3:2] : \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.ain_s1 ;
assign _191_ = \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.ce  ? \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.facout_s1  : \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.carry_s1 ;
assign _192_ = \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.ce  ? \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.fas_s1  : \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.sum_s1 ;
assign _193_ = \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.u1.a  + \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.u1.b ;
assign { \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.u1.cout , \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.u1.s  } = _193_ + \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.u1.cin ;
assign _194_ = \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.u2.a  + \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.u2.b ;
assign { \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.u2.cout , \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.u2.s  } = _194_ + \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.u2.cin ;
always @(posedge \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.clk )
\add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.bin_s1  <= _196_;
always @(posedge \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.clk )
\add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.ain_s1  <= _195_;
always @(posedge \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.clk )
\add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.sum_s1  <= _198_;
always @(posedge \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.clk )
\add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.carry_s1  <= _197_;
assign _196_ = \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.ce  ? \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.b [3:2] : \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.bin_s1 ;
assign _195_ = \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.ce  ? \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.a [3:2] : \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.ain_s1 ;
assign _197_ = \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.ce  ? \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.facout_s1  : \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.carry_s1 ;
assign _198_ = \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.ce  ? \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.fas_s1  : \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.sum_s1 ;
assign _199_ = \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.u1.a  + \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.u1.b ;
assign { \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.u1.cout , \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.u1.s  } = _199_ + \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.u1.cin ;
assign _200_ = \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.u2.a  + \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.u2.b ;
assign { \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.u2.cout , \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.u2.s  } = _200_ + \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.u2.cin ;
always @(posedge \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.clk )
\add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.bin_s1  <= _202_;
always @(posedge \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.clk )
\add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.ain_s1  <= _201_;
always @(posedge \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.clk )
\add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.sum_s1  <= _204_;
always @(posedge \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.clk )
\add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.carry_s1  <= _203_;
assign _202_ = \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.ce  ? \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.b [4:2] : \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.bin_s1 ;
assign _201_ = \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.ce  ? \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.a [4:2] : \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.ain_s1 ;
assign _203_ = \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.ce  ? \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.facout_s1  : \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.carry_s1 ;
assign _204_ = \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.ce  ? \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.fas_s1  : \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.sum_s1 ;
assign _205_ = \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.u1.a  + \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.u1.b ;
assign { \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.u1.cout , \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.u1.s  } = _205_ + \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.u1.cin ;
assign _206_ = \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.u2.a  + \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.u2.b ;
assign { \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.u2.cout , \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.u2.s  } = _206_ + \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.u2.cin ;
always @(posedge \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_5_U.clk )
\add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_5_U.bin_s1  <= _208_;
always @(posedge \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_5_U.clk )
\add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_5_U.ain_s1  <= _207_;
always @(posedge \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_5_U.clk )
\add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_5_U.sum_s1  <= _210_;
always @(posedge \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_5_U.clk )
\add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_5_U.carry_s1  <= _209_;
assign _208_ = \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_5_U.ce  ? \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_5_U.b [5:3] : \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_5_U.bin_s1 ;
assign _207_ = \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_5_U.ce  ? \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_5_U.a [5:3] : \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_5_U.ain_s1 ;
assign _209_ = \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_5_U.ce  ? \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_5_U.facout_s1  : \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_5_U.carry_s1 ;
assign _210_ = \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_5_U.ce  ? \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_5_U.fas_s1  : \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_5_U.sum_s1 ;
assign _211_ = \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_5_U.u1.a  + \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_5_U.u1.b ;
assign { \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_5_U.u1.cout , \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_5_U.u1.s  } = _211_ + \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_5_U.u1.cin ;
assign _212_ = \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_5_U.u2.a  + \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_5_U.u2.b ;
assign { \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_5_U.u2.cout , \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_5_U.u2.s  } = _212_ + \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_5_U.u2.cin ;
always @(posedge \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.clk )
\add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.bin_s1  <= _214_;
always @(posedge \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.clk )
\add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.ain_s1  <= _213_;
always @(posedge \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.clk )
\add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.sum_s1  <= _216_;
always @(posedge \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.clk )
\add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.carry_s1  <= _215_;
assign _214_ = \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.ce  ? \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.b [5:3] : \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.bin_s1 ;
assign _213_ = \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.ce  ? \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.a [5:3] : \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.ain_s1 ;
assign _215_ = \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.ce  ? \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.facout_s1  : \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.carry_s1 ;
assign _216_ = \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.ce  ? \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.fas_s1  : \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.sum_s1 ;
assign _217_ = \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.u1.a  + \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.u1.b ;
assign { \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.u1.cout , \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.u1.s  } = _217_ + \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.u1.cin ;
assign _218_ = \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.u2.a  + \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.u2.b ;
assign { \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.u2.cout , \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.u2.s  } = _218_ + \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.u2.cin ;
always @(posedge \add_8s_8ns_8_2_1_U11.top_add_8s_8ns_8_2_1_Adder_8_U.clk )
\add_8s_8ns_8_2_1_U11.top_add_8s_8ns_8_2_1_Adder_8_U.bin_s1  <= _220_;
always @(posedge \add_8s_8ns_8_2_1_U11.top_add_8s_8ns_8_2_1_Adder_8_U.clk )
\add_8s_8ns_8_2_1_U11.top_add_8s_8ns_8_2_1_Adder_8_U.ain_s1  <= _219_;
always @(posedge \add_8s_8ns_8_2_1_U11.top_add_8s_8ns_8_2_1_Adder_8_U.clk )
\add_8s_8ns_8_2_1_U11.top_add_8s_8ns_8_2_1_Adder_8_U.sum_s1  <= _222_;
always @(posedge \add_8s_8ns_8_2_1_U11.top_add_8s_8ns_8_2_1_Adder_8_U.clk )
\add_8s_8ns_8_2_1_U11.top_add_8s_8ns_8_2_1_Adder_8_U.carry_s1  <= _221_;
assign _220_ = \add_8s_8ns_8_2_1_U11.top_add_8s_8ns_8_2_1_Adder_8_U.ce  ? \add_8s_8ns_8_2_1_U11.top_add_8s_8ns_8_2_1_Adder_8_U.b [7:4] : \add_8s_8ns_8_2_1_U11.top_add_8s_8ns_8_2_1_Adder_8_U.bin_s1 ;
assign _219_ = \add_8s_8ns_8_2_1_U11.top_add_8s_8ns_8_2_1_Adder_8_U.ce  ? \add_8s_8ns_8_2_1_U11.top_add_8s_8ns_8_2_1_Adder_8_U.a [7:4] : \add_8s_8ns_8_2_1_U11.top_add_8s_8ns_8_2_1_Adder_8_U.ain_s1 ;
assign _221_ = \add_8s_8ns_8_2_1_U11.top_add_8s_8ns_8_2_1_Adder_8_U.ce  ? \add_8s_8ns_8_2_1_U11.top_add_8s_8ns_8_2_1_Adder_8_U.facout_s1  : \add_8s_8ns_8_2_1_U11.top_add_8s_8ns_8_2_1_Adder_8_U.carry_s1 ;
assign _222_ = \add_8s_8ns_8_2_1_U11.top_add_8s_8ns_8_2_1_Adder_8_U.ce  ? \add_8s_8ns_8_2_1_U11.top_add_8s_8ns_8_2_1_Adder_8_U.fas_s1  : \add_8s_8ns_8_2_1_U11.top_add_8s_8ns_8_2_1_Adder_8_U.sum_s1 ;
assign _223_ = \add_8s_8ns_8_2_1_U11.top_add_8s_8ns_8_2_1_Adder_8_U.u1.a  + \add_8s_8ns_8_2_1_U11.top_add_8s_8ns_8_2_1_Adder_8_U.u1.b ;
assign { \add_8s_8ns_8_2_1_U11.top_add_8s_8ns_8_2_1_Adder_8_U.u1.cout , \add_8s_8ns_8_2_1_U11.top_add_8s_8ns_8_2_1_Adder_8_U.u1.s  } = _223_ + \add_8s_8ns_8_2_1_U11.top_add_8s_8ns_8_2_1_Adder_8_U.u1.cin ;
assign _224_ = \add_8s_8ns_8_2_1_U11.top_add_8s_8ns_8_2_1_Adder_8_U.u2.a  + \add_8s_8ns_8_2_1_U11.top_add_8s_8ns_8_2_1_Adder_8_U.u2.b ;
assign { \add_8s_8ns_8_2_1_U11.top_add_8s_8ns_8_2_1_Adder_8_U.u2.cout , \add_8s_8ns_8_2_1_U11.top_add_8s_8ns_8_2_1_Adder_8_U.u2.s  } = _224_ + \add_8s_8ns_8_2_1_U11.top_add_8s_8ns_8_2_1_Adder_8_U.u2.cin ;
always @(posedge \add_8s_8s_8_2_1_U10.top_add_8s_8s_8_2_1_Adder_7_U.clk )
\add_8s_8s_8_2_1_U10.top_add_8s_8s_8_2_1_Adder_7_U.bin_s1  <= _226_;
always @(posedge \add_8s_8s_8_2_1_U10.top_add_8s_8s_8_2_1_Adder_7_U.clk )
\add_8s_8s_8_2_1_U10.top_add_8s_8s_8_2_1_Adder_7_U.ain_s1  <= _225_;
always @(posedge \add_8s_8s_8_2_1_U10.top_add_8s_8s_8_2_1_Adder_7_U.clk )
\add_8s_8s_8_2_1_U10.top_add_8s_8s_8_2_1_Adder_7_U.sum_s1  <= _228_;
always @(posedge \add_8s_8s_8_2_1_U10.top_add_8s_8s_8_2_1_Adder_7_U.clk )
\add_8s_8s_8_2_1_U10.top_add_8s_8s_8_2_1_Adder_7_U.carry_s1  <= _227_;
assign _226_ = \add_8s_8s_8_2_1_U10.top_add_8s_8s_8_2_1_Adder_7_U.ce  ? \add_8s_8s_8_2_1_U10.top_add_8s_8s_8_2_1_Adder_7_U.b [7:4] : \add_8s_8s_8_2_1_U10.top_add_8s_8s_8_2_1_Adder_7_U.bin_s1 ;
assign _225_ = \add_8s_8s_8_2_1_U10.top_add_8s_8s_8_2_1_Adder_7_U.ce  ? \add_8s_8s_8_2_1_U10.top_add_8s_8s_8_2_1_Adder_7_U.a [7:4] : \add_8s_8s_8_2_1_U10.top_add_8s_8s_8_2_1_Adder_7_U.ain_s1 ;
assign _227_ = \add_8s_8s_8_2_1_U10.top_add_8s_8s_8_2_1_Adder_7_U.ce  ? \add_8s_8s_8_2_1_U10.top_add_8s_8s_8_2_1_Adder_7_U.facout_s1  : \add_8s_8s_8_2_1_U10.top_add_8s_8s_8_2_1_Adder_7_U.carry_s1 ;
assign _228_ = \add_8s_8s_8_2_1_U10.top_add_8s_8s_8_2_1_Adder_7_U.ce  ? \add_8s_8s_8_2_1_U10.top_add_8s_8s_8_2_1_Adder_7_U.fas_s1  : \add_8s_8s_8_2_1_U10.top_add_8s_8s_8_2_1_Adder_7_U.sum_s1 ;
assign _229_ = \add_8s_8s_8_2_1_U10.top_add_8s_8s_8_2_1_Adder_7_U.u1.a  + \add_8s_8s_8_2_1_U10.top_add_8s_8s_8_2_1_Adder_7_U.u1.b ;
assign { \add_8s_8s_8_2_1_U10.top_add_8s_8s_8_2_1_Adder_7_U.u1.cout , \add_8s_8s_8_2_1_U10.top_add_8s_8s_8_2_1_Adder_7_U.u1.s  } = _229_ + \add_8s_8s_8_2_1_U10.top_add_8s_8s_8_2_1_Adder_7_U.u1.cin ;
assign _230_ = \add_8s_8s_8_2_1_U10.top_add_8s_8s_8_2_1_Adder_7_U.u2.a  + \add_8s_8s_8_2_1_U10.top_add_8s_8s_8_2_1_Adder_7_U.u2.b ;
assign { \add_8s_8s_8_2_1_U10.top_add_8s_8s_8_2_1_Adder_7_U.u2.cout , \add_8s_8s_8_2_1_U10.top_add_8s_8s_8_2_1_Adder_7_U.u2.s  } = _230_ + \add_8s_8s_8_2_1_U10.top_add_8s_8s_8_2_1_Adder_7_U.u2.cin ;
always @(posedge \add_9s_9ns_9_2_1_U5.top_add_9s_9ns_9_2_1_Adder_3_U.clk )
\add_9s_9ns_9_2_1_U5.top_add_9s_9ns_9_2_1_Adder_3_U.bin_s1  <= _232_;
always @(posedge \add_9s_9ns_9_2_1_U5.top_add_9s_9ns_9_2_1_Adder_3_U.clk )
\add_9s_9ns_9_2_1_U5.top_add_9s_9ns_9_2_1_Adder_3_U.ain_s1  <= _231_;
always @(posedge \add_9s_9ns_9_2_1_U5.top_add_9s_9ns_9_2_1_Adder_3_U.clk )
\add_9s_9ns_9_2_1_U5.top_add_9s_9ns_9_2_1_Adder_3_U.sum_s1  <= _234_;
always @(posedge \add_9s_9ns_9_2_1_U5.top_add_9s_9ns_9_2_1_Adder_3_U.clk )
\add_9s_9ns_9_2_1_U5.top_add_9s_9ns_9_2_1_Adder_3_U.carry_s1  <= _233_;
assign _232_ = \add_9s_9ns_9_2_1_U5.top_add_9s_9ns_9_2_1_Adder_3_U.ce  ? \add_9s_9ns_9_2_1_U5.top_add_9s_9ns_9_2_1_Adder_3_U.b [8:4] : \add_9s_9ns_9_2_1_U5.top_add_9s_9ns_9_2_1_Adder_3_U.bin_s1 ;
assign _231_ = \add_9s_9ns_9_2_1_U5.top_add_9s_9ns_9_2_1_Adder_3_U.ce  ? \add_9s_9ns_9_2_1_U5.top_add_9s_9ns_9_2_1_Adder_3_U.a [8:4] : \add_9s_9ns_9_2_1_U5.top_add_9s_9ns_9_2_1_Adder_3_U.ain_s1 ;
assign _233_ = \add_9s_9ns_9_2_1_U5.top_add_9s_9ns_9_2_1_Adder_3_U.ce  ? \add_9s_9ns_9_2_1_U5.top_add_9s_9ns_9_2_1_Adder_3_U.facout_s1  : \add_9s_9ns_9_2_1_U5.top_add_9s_9ns_9_2_1_Adder_3_U.carry_s1 ;
assign _234_ = \add_9s_9ns_9_2_1_U5.top_add_9s_9ns_9_2_1_Adder_3_U.ce  ? \add_9s_9ns_9_2_1_U5.top_add_9s_9ns_9_2_1_Adder_3_U.fas_s1  : \add_9s_9ns_9_2_1_U5.top_add_9s_9ns_9_2_1_Adder_3_U.sum_s1 ;
assign _235_ = \add_9s_9ns_9_2_1_U5.top_add_9s_9ns_9_2_1_Adder_3_U.u1.a  + \add_9s_9ns_9_2_1_U5.top_add_9s_9ns_9_2_1_Adder_3_U.u1.b ;
assign { \add_9s_9ns_9_2_1_U5.top_add_9s_9ns_9_2_1_Adder_3_U.u1.cout , \add_9s_9ns_9_2_1_U5.top_add_9s_9ns_9_2_1_Adder_3_U.u1.s  } = _235_ + \add_9s_9ns_9_2_1_U5.top_add_9s_9ns_9_2_1_Adder_3_U.u1.cin ;
assign _236_ = \add_9s_9ns_9_2_1_U5.top_add_9s_9ns_9_2_1_Adder_3_U.u2.a  + \add_9s_9ns_9_2_1_U5.top_add_9s_9ns_9_2_1_Adder_3_U.u2.b ;
assign { \add_9s_9ns_9_2_1_U5.top_add_9s_9ns_9_2_1_Adder_3_U.u2.cout , \add_9s_9ns_9_2_1_U5.top_add_9s_9ns_9_2_1_Adder_3_U.u2.s  } = _236_ + \add_9s_9ns_9_2_1_U5.top_add_9s_9ns_9_2_1_Adder_3_U.u2.cin ;
always @(posedge \add_9s_9s_9_2_1_U8.top_add_9s_9s_9_2_1_Adder_6_U.clk )
\add_9s_9s_9_2_1_U8.top_add_9s_9s_9_2_1_Adder_6_U.bin_s1  <= _238_;
always @(posedge \add_9s_9s_9_2_1_U8.top_add_9s_9s_9_2_1_Adder_6_U.clk )
\add_9s_9s_9_2_1_U8.top_add_9s_9s_9_2_1_Adder_6_U.ain_s1  <= _237_;
always @(posedge \add_9s_9s_9_2_1_U8.top_add_9s_9s_9_2_1_Adder_6_U.clk )
\add_9s_9s_9_2_1_U8.top_add_9s_9s_9_2_1_Adder_6_U.sum_s1  <= _240_;
always @(posedge \add_9s_9s_9_2_1_U8.top_add_9s_9s_9_2_1_Adder_6_U.clk )
\add_9s_9s_9_2_1_U8.top_add_9s_9s_9_2_1_Adder_6_U.carry_s1  <= _239_;
assign _238_ = \add_9s_9s_9_2_1_U8.top_add_9s_9s_9_2_1_Adder_6_U.ce  ? \add_9s_9s_9_2_1_U8.top_add_9s_9s_9_2_1_Adder_6_U.b [8:4] : \add_9s_9s_9_2_1_U8.top_add_9s_9s_9_2_1_Adder_6_U.bin_s1 ;
assign _237_ = \add_9s_9s_9_2_1_U8.top_add_9s_9s_9_2_1_Adder_6_U.ce  ? \add_9s_9s_9_2_1_U8.top_add_9s_9s_9_2_1_Adder_6_U.a [8:4] : \add_9s_9s_9_2_1_U8.top_add_9s_9s_9_2_1_Adder_6_U.ain_s1 ;
assign _239_ = \add_9s_9s_9_2_1_U8.top_add_9s_9s_9_2_1_Adder_6_U.ce  ? \add_9s_9s_9_2_1_U8.top_add_9s_9s_9_2_1_Adder_6_U.facout_s1  : \add_9s_9s_9_2_1_U8.top_add_9s_9s_9_2_1_Adder_6_U.carry_s1 ;
assign _240_ = \add_9s_9s_9_2_1_U8.top_add_9s_9s_9_2_1_Adder_6_U.ce  ? \add_9s_9s_9_2_1_U8.top_add_9s_9s_9_2_1_Adder_6_U.fas_s1  : \add_9s_9s_9_2_1_U8.top_add_9s_9s_9_2_1_Adder_6_U.sum_s1 ;
assign _241_ = \add_9s_9s_9_2_1_U8.top_add_9s_9s_9_2_1_Adder_6_U.u1.a  + \add_9s_9s_9_2_1_U8.top_add_9s_9s_9_2_1_Adder_6_U.u1.b ;
assign { \add_9s_9s_9_2_1_U8.top_add_9s_9s_9_2_1_Adder_6_U.u1.cout , \add_9s_9s_9_2_1_U8.top_add_9s_9s_9_2_1_Adder_6_U.u1.s  } = _241_ + \add_9s_9s_9_2_1_U8.top_add_9s_9s_9_2_1_Adder_6_U.u1.cin ;
assign _242_ = \add_9s_9s_9_2_1_U8.top_add_9s_9s_9_2_1_Adder_6_U.u2.a  + \add_9s_9s_9_2_1_U8.top_add_9s_9s_9_2_1_Adder_6_U.u2.b ;
assign { \add_9s_9s_9_2_1_U8.top_add_9s_9s_9_2_1_Adder_6_U.u2.cout , \add_9s_9s_9_2_1_U8.top_add_9s_9s_9_2_1_Adder_6_U.u2.s  } = _242_ + \add_9s_9s_9_2_1_U8.top_add_9s_9s_9_2_1_Adder_6_U.u2.cin ;
assign \mul_16ns_4s_20_7_1_U4.top_mul_16ns_4s_20_7_1_Mul_DSP_0_U.tmp_product  = $signed({ 1'h0, \mul_16ns_4s_20_7_1_U4.top_mul_16ns_4s_20_7_1_Mul_DSP_0_U.a_reg0  }) * $signed(\mul_16ns_4s_20_7_1_U4.top_mul_16ns_4s_20_7_1_Mul_DSP_0_U.b_reg0 );
always @(posedge \mul_16ns_4s_20_7_1_U4.top_mul_16ns_4s_20_7_1_Mul_DSP_0_U.clk )
\mul_16ns_4s_20_7_1_U4.top_mul_16ns_4s_20_7_1_Mul_DSP_0_U.a_reg0  <= _243_;
always @(posedge \mul_16ns_4s_20_7_1_U4.top_mul_16ns_4s_20_7_1_Mul_DSP_0_U.clk )
\mul_16ns_4s_20_7_1_U4.top_mul_16ns_4s_20_7_1_Mul_DSP_0_U.b_reg0  <= _244_;
always @(posedge \mul_16ns_4s_20_7_1_U4.top_mul_16ns_4s_20_7_1_Mul_DSP_0_U.clk )
\mul_16ns_4s_20_7_1_U4.top_mul_16ns_4s_20_7_1_Mul_DSP_0_U.buff0  <= _245_;
always @(posedge \mul_16ns_4s_20_7_1_U4.top_mul_16ns_4s_20_7_1_Mul_DSP_0_U.clk )
\mul_16ns_4s_20_7_1_U4.top_mul_16ns_4s_20_7_1_Mul_DSP_0_U.buff1  <= _246_;
always @(posedge \mul_16ns_4s_20_7_1_U4.top_mul_16ns_4s_20_7_1_Mul_DSP_0_U.clk )
\mul_16ns_4s_20_7_1_U4.top_mul_16ns_4s_20_7_1_Mul_DSP_0_U.buff2  <= _247_;
always @(posedge \mul_16ns_4s_20_7_1_U4.top_mul_16ns_4s_20_7_1_Mul_DSP_0_U.clk )
\mul_16ns_4s_20_7_1_U4.top_mul_16ns_4s_20_7_1_Mul_DSP_0_U.buff3  <= _248_;
always @(posedge \mul_16ns_4s_20_7_1_U4.top_mul_16ns_4s_20_7_1_Mul_DSP_0_U.clk )
\mul_16ns_4s_20_7_1_U4.top_mul_16ns_4s_20_7_1_Mul_DSP_0_U.buff4  <= _249_;
assign _249_ = \mul_16ns_4s_20_7_1_U4.top_mul_16ns_4s_20_7_1_Mul_DSP_0_U.ce  ? \mul_16ns_4s_20_7_1_U4.top_mul_16ns_4s_20_7_1_Mul_DSP_0_U.buff3  : \mul_16ns_4s_20_7_1_U4.top_mul_16ns_4s_20_7_1_Mul_DSP_0_U.buff4 ;
assign _248_ = \mul_16ns_4s_20_7_1_U4.top_mul_16ns_4s_20_7_1_Mul_DSP_0_U.ce  ? \mul_16ns_4s_20_7_1_U4.top_mul_16ns_4s_20_7_1_Mul_DSP_0_U.buff2  : \mul_16ns_4s_20_7_1_U4.top_mul_16ns_4s_20_7_1_Mul_DSP_0_U.buff3 ;
assign _247_ = \mul_16ns_4s_20_7_1_U4.top_mul_16ns_4s_20_7_1_Mul_DSP_0_U.ce  ? \mul_16ns_4s_20_7_1_U4.top_mul_16ns_4s_20_7_1_Mul_DSP_0_U.buff1  : \mul_16ns_4s_20_7_1_U4.top_mul_16ns_4s_20_7_1_Mul_DSP_0_U.buff2 ;
assign _246_ = \mul_16ns_4s_20_7_1_U4.top_mul_16ns_4s_20_7_1_Mul_DSP_0_U.ce  ? \mul_16ns_4s_20_7_1_U4.top_mul_16ns_4s_20_7_1_Mul_DSP_0_U.buff0  : \mul_16ns_4s_20_7_1_U4.top_mul_16ns_4s_20_7_1_Mul_DSP_0_U.buff1 ;
assign _245_ = \mul_16ns_4s_20_7_1_U4.top_mul_16ns_4s_20_7_1_Mul_DSP_0_U.ce  ? \mul_16ns_4s_20_7_1_U4.top_mul_16ns_4s_20_7_1_Mul_DSP_0_U.tmp_product  : \mul_16ns_4s_20_7_1_U4.top_mul_16ns_4s_20_7_1_Mul_DSP_0_U.buff0 ;
assign _244_ = \mul_16ns_4s_20_7_1_U4.top_mul_16ns_4s_20_7_1_Mul_DSP_0_U.ce  ? \mul_16ns_4s_20_7_1_U4.top_mul_16ns_4s_20_7_1_Mul_DSP_0_U.b  : \mul_16ns_4s_20_7_1_U4.top_mul_16ns_4s_20_7_1_Mul_DSP_0_U.b_reg0 ;
assign _243_ = \mul_16ns_4s_20_7_1_U4.top_mul_16ns_4s_20_7_1_Mul_DSP_0_U.ce  ? \mul_16ns_4s_20_7_1_U4.top_mul_16ns_4s_20_7_1_Mul_DSP_0_U.a  : \mul_16ns_4s_20_7_1_U4.top_mul_16ns_4s_20_7_1_Mul_DSP_0_U.a_reg0 ;
assign \sub_17ns_17ns_17_2_1_U3.top_sub_17ns_17ns_17_2_1_Adder_2_U.bin_s0  = ~ \sub_17ns_17ns_17_2_1_U3.top_sub_17ns_17ns_17_2_1_Adder_2_U.b ;
always @(posedge \sub_17ns_17ns_17_2_1_U3.top_sub_17ns_17ns_17_2_1_Adder_2_U.clk )
\sub_17ns_17ns_17_2_1_U3.top_sub_17ns_17ns_17_2_1_Adder_2_U.bin_s1  <= _251_;
always @(posedge \sub_17ns_17ns_17_2_1_U3.top_sub_17ns_17ns_17_2_1_Adder_2_U.clk )
\sub_17ns_17ns_17_2_1_U3.top_sub_17ns_17ns_17_2_1_Adder_2_U.ain_s1  <= _250_;
always @(posedge \sub_17ns_17ns_17_2_1_U3.top_sub_17ns_17ns_17_2_1_Adder_2_U.clk )
\sub_17ns_17ns_17_2_1_U3.top_sub_17ns_17ns_17_2_1_Adder_2_U.sum_s1  <= _253_;
always @(posedge \sub_17ns_17ns_17_2_1_U3.top_sub_17ns_17ns_17_2_1_Adder_2_U.clk )
\sub_17ns_17ns_17_2_1_U3.top_sub_17ns_17ns_17_2_1_Adder_2_U.carry_s1  <= _252_;
assign _251_ = \sub_17ns_17ns_17_2_1_U3.top_sub_17ns_17ns_17_2_1_Adder_2_U.ce  ? \sub_17ns_17ns_17_2_1_U3.top_sub_17ns_17ns_17_2_1_Adder_2_U.bin_s0 [16:8] : \sub_17ns_17ns_17_2_1_U3.top_sub_17ns_17ns_17_2_1_Adder_2_U.bin_s1 ;
assign _250_ = \sub_17ns_17ns_17_2_1_U3.top_sub_17ns_17ns_17_2_1_Adder_2_U.ce  ? \sub_17ns_17ns_17_2_1_U3.top_sub_17ns_17ns_17_2_1_Adder_2_U.a [16:8] : \sub_17ns_17ns_17_2_1_U3.top_sub_17ns_17ns_17_2_1_Adder_2_U.ain_s1 ;
assign _252_ = \sub_17ns_17ns_17_2_1_U3.top_sub_17ns_17ns_17_2_1_Adder_2_U.ce  ? \sub_17ns_17ns_17_2_1_U3.top_sub_17ns_17ns_17_2_1_Adder_2_U.facout_s1  : \sub_17ns_17ns_17_2_1_U3.top_sub_17ns_17ns_17_2_1_Adder_2_U.carry_s1 ;
assign _253_ = \sub_17ns_17ns_17_2_1_U3.top_sub_17ns_17ns_17_2_1_Adder_2_U.ce  ? \sub_17ns_17ns_17_2_1_U3.top_sub_17ns_17ns_17_2_1_Adder_2_U.fas_s1  : \sub_17ns_17ns_17_2_1_U3.top_sub_17ns_17ns_17_2_1_Adder_2_U.sum_s1 ;
assign _254_ = \sub_17ns_17ns_17_2_1_U3.top_sub_17ns_17ns_17_2_1_Adder_2_U.u1.a  + \sub_17ns_17ns_17_2_1_U3.top_sub_17ns_17ns_17_2_1_Adder_2_U.u1.b ;
assign { \sub_17ns_17ns_17_2_1_U3.top_sub_17ns_17ns_17_2_1_Adder_2_U.u1.cout , \sub_17ns_17ns_17_2_1_U3.top_sub_17ns_17ns_17_2_1_Adder_2_U.u1.s  } = _254_ + \sub_17ns_17ns_17_2_1_U3.top_sub_17ns_17ns_17_2_1_Adder_2_U.u1.cin ;
assign _255_ = \sub_17ns_17ns_17_2_1_U3.top_sub_17ns_17ns_17_2_1_Adder_2_U.u2.a  + \sub_17ns_17ns_17_2_1_U3.top_sub_17ns_17ns_17_2_1_Adder_2_U.u2.b ;
assign { \sub_17ns_17ns_17_2_1_U3.top_sub_17ns_17ns_17_2_1_Adder_2_U.u2.cout , \sub_17ns_17ns_17_2_1_U3.top_sub_17ns_17ns_17_2_1_Adder_2_U.u2.s  } = _255_ + \sub_17ns_17ns_17_2_1_U3.top_sub_17ns_17ns_17_2_1_Adder_2_U.u2.cin ;
assign _256_ = $signed({ 1'h0, signbit_3_reg_1869, 1'h0 }) < $signed(op_5);
assign _257_ = | tmp_2_reg_1484;
assign _258_ = tmp_2_reg_1484 != 12'hfff;
assign _259_ = | op_18[1:0];
assign _260_ = { op_5[1], op_5[1], op_5[1], op_5[1], op_5 } != { op_7, 1'h0 };
assign _261_ = | trunc_ln718_reg_1738;
assign _262_ = { ret_V_21_reg_1441[1], ret_V_21_reg_1441[1], ret_V_21_reg_1441[1], ret_V_21_reg_1441[1], ret_V_21_reg_1441[1], ret_V_21_reg_1441[1], ret_V_21_reg_1441[1], ret_V_21_reg_1441[1], ret_V_21_reg_1441[1], ret_V_21_reg_1441[1], ret_V_21_reg_1441[1], ret_V_21_reg_1441[1], ret_V_21_reg_1441[1], ret_V_21_reg_1441[1], ret_V_21_reg_1441, 1'h0 } != { op_5[1], op_5[1], op_5[1], op_5[1], op_5[1], op_5[1], op_5[1], op_5[1], op_5[1], op_5[1], op_5[1], op_5[1], op_5[1], op_5[1], op_5[1], op_5[1], op_5 };
assign or_ln340_1_fu_748_p2 = or_ln340_reg_1681 | and_ln786_reg_1673;
assign or_ln340_2_fu_773_p2 = and_ln785_2_fu_759_p2 | and_ln340_fu_768_p2;
assign or_ln340_fu_688_p2 = overflow_1_fu_683_p2 | neg_src_fu_668_p2;
assign or_ln384_fu_430_p2 = underflow_fu_425_p2 | overflow_reg_1510;
assign or_ln406_fu_533_p2 = r_V_1_reg_1526[0] | p_Result_25_reg_1533;
assign or_ln785_1_fu_678_p2 = xor_ln785_2_fu_673_p2 | p_Result_28_reg_1631;
assign or_ln785_2_fu_698_p2 = p_Result_25_reg_1533 | and_ln785_fu_694_p2;
assign or_ln785_fu_395_p2 = p_Result_24_reg_1478 | icmp_ln768_reg_1495;
assign or_ln788_1_fu_420_p2 = or_ln788_fu_415_p2 | icmp_ln786_reg_1500;
assign or_ln788_fu_415_p2 = xor_ln786_fu_410_p2 | icmp_ln790_reg_1505;
always @(posedge ap_clk)
select_ln703_reg_1402[2:0] <= 3'h0;
always @(posedge ap_clk)
xor_ln416_reg_1643 <= _088_;
always @(posedge ap_clk)
select_ln850_4_reg_1649 <= _077_;
always @(posedge ap_clk)
select_ln703_reg_1402[4:3] <= _076_;
always @(posedge ap_clk)
select_ln353_2_reg_1943 <= _073_;
always @(posedge ap_clk)
select_ln340_1_reg_1692 <= _072_;
always @(posedge ap_clk)
sel_tmp11_reg_1697 <= _069_;
always @(posedge ap_clk)
ret_V_34_reg_2032 <= _064_;
always @(posedge ap_clk)
ret_V_33_reg_2015 <= _062_;
always @(posedge ap_clk)
ret_V_34_cast_reg_2020 <= _063_;
always @(posedge ap_clk)
xor_ln1497_reg_1980 <= _087_;
always @(posedge ap_clk)
ret_V_32_reg_1985 <= _061_;
always @(posedge ap_clk)
ret_V_31_reg_1963 <= _059_;
always @(posedge ap_clk)
ret_V_32_cast_reg_1968 <= _060_;
always @(posedge ap_clk)
ret_V_30_reg_1926 <= _058_;
always @(posedge ap_clk)
ret_V_30_cast_reg_1931 <= _057_;
always @(posedge ap_clk)
ret_V_2_reg_1436 <= _056_;
always @(posedge ap_clk)
ret_V_29_reg_1906 <= _055_;
always @(posedge ap_clk)
ret_V_28_reg_1896 <= _054_;
always @(posedge ap_clk)
select_ln1192_reg_1901 <= _070_;
always @(posedge ap_clk)
ret_V_27_reg_1833 <= _053_;
always @(posedge ap_clk)
select_ln69_reg_1838 <= _075_;
always @(posedge ap_clk)
ret_V_26_reg_1816 <= _052_;
always @(posedge ap_clk)
ret_V_24_cast_reg_1821 <= _049_;
always @(posedge ap_clk)
ret_V_21_reg_1441 <= _048_;
always @(posedge ap_clk)
select_ln1347_reg_1447 <= _071_;
always @(posedge ap_clk)
ret_V_20_reg_1424 <= _047_;
always @(posedge ap_clk)
ret_V_reg_1429 <= _067_;
always @(posedge ap_clk)
r_reg_1753 <= _046_;
always @(posedge ap_clk)
ret_V_25_reg_1758 <= _051_;
always @(posedge ap_clk)
tmp_3_reg_1763 <= _081_;
always @(posedge ap_clk)
p_Val2_7_reg_1622 <= _044_;
always @(posedge ap_clk)
p_Result_28_reg_1631 <= _039_;
always @(posedge ap_clk)
ret_V_9_reg_1638 <= _066_;
always @(posedge ap_clk)
r_V_1_reg_1526 <= _045_;
always @(posedge ap_clk)
p_Result_25_reg_1533 <= _037_;
always @(posedge ap_clk)
p_Val2_6_reg_1541 <= _043_;
always @(posedge ap_clk)
p_Result_27_reg_1546 <= _038_;
always @(posedge ap_clk)
p_Result_29_reg_1551 <= _040_;
always @(posedge ap_clk)
p_Result_6_reg_1557 <= _041_;
always @(posedge ap_clk)
p_Result_7_reg_1562 <= _042_;
always @(posedge ap_clk)
ret_reg_1467 <= _068_;
always @(posedge ap_clk)
p_Result_23_reg_1472 <= _035_;
always @(posedge ap_clk)
p_Result_24_reg_1478 <= _036_;
always @(posedge ap_clk)
tmp_2_reg_1484 <= _080_;
always @(posedge ap_clk)
trunc_ln790_reg_1490 <= _085_;
always @(posedge ap_clk)
trunc_ln2_reg_1728 <= _082_;
always @(posedge ap_clk)
p_Result_22_reg_1733 <= _034_;
always @(posedge ap_clk)
trunc_ln718_reg_1738 <= _084_;
always @(posedge ap_clk)
overflow_reg_1510 <= _032_;
always @(posedge ap_clk)
or_ln384_reg_1516 <= _031_;
always @(posedge ap_clk)
op_9_V_reg_1722 <= _029_;
always @(posedge ap_clk)
op_8_V_reg_1521 <= _028_;
always @(posedge ap_clk)
op_28_V_reg_1995 <= _027_;
always @(posedge ap_clk)
op_10_V_reg_1795 <= _025_;
always @(posedge ap_clk)
select_ln353_reg_1801 <= _074_;
always @(posedge ap_clk)
icmp_ln851_reg_1419 <= _022_;
always @(posedge ap_clk)
icmp_ln851_2_reg_2010 <= _021_;
always @(posedge ap_clk)
icmp_ln851_1_reg_1617 <= _020_;
always @(posedge ap_clk)
icmp_ln768_reg_1495 <= _017_;
always @(posedge ap_clk)
icmp_ln786_reg_1500 <= _018_;
always @(posedge ap_clk)
icmp_ln790_reg_1505 <= _019_;
always @(posedge ap_clk)
newsignbit_reg_1879 <= _024_;
always @(posedge ap_clk)
icmp_ln1497_reg_1886 <= _016_;
always @(posedge ap_clk)
trunc_ln415_reg_1848 <= _083_;
always @(posedge ap_clk)
p_Result_21_reg_1853 <= _033_;
always @(posedge ap_clk)
carry_reg_1859 <= _014_;
always @(posedge ap_clk)
lhs_V_2_reg_1864 <= _023_;
always @(posedge ap_clk)
signbit_3_reg_1869 <= _079_;
always @(posedge ap_clk)
op_23_V_reg_1874 <= _026_;
always @(posedge ap_clk)
carry_2_reg_1654 <= _013_;
always @(posedge ap_clk)
deleted_zeros_reg_1661 <= _015_;
always @(posedge ap_clk)
xor_ln785_3_reg_1667 <= _089_;
always @(posedge ap_clk)
and_ln786_reg_1673 <= _011_;
always @(posedge ap_clk)
or_ln340_reg_1681 <= _030_;
always @(posedge ap_clk)
and_ln785_1_reg_1687 <= _010_;
always @(posedge ap_clk)
and_ln408_reg_1768 <= _009_;
always @(posedge ap_clk)
sext_ln850_reg_1773 <= _078_;
always @(posedge ap_clk)
add_ln691_reg_1790 <= _007_;
always @(posedge ap_clk)
add_ln691_4_reg_2027 <= _006_;
always @(posedge ap_clk)
add_ln691_3_reg_1975 <= _005_;
always @(posedge ap_clk)
add_ln691_2_reg_1938 <= _004_;
always @(posedge ap_clk)
add_ln691_1_reg_1828 <= _003_;
always @(posedge ap_clk)
and_ln406_reg_1573 <= _008_;
always @(posedge ap_clk)
Range2_all_ones_reg_1578 <= _002_;
always @(posedge ap_clk)
Range1_all_ones_reg_1583 <= _000_;
always @(posedge ap_clk)
Range1_all_zeros_reg_1590 <= _001_;
always @(posedge ap_clk)
ret_V_24_reg_1595 <= _050_;
always @(posedge ap_clk)
ret_V_7_reg_1600 <= _065_;
always @(posedge ap_clk)
trunc_ln851_1_reg_1607 <= _086_;
always @(posedge ap_clk)
ap_CS_fsm <= _012_;
assign _090_ = _095_ ? 2'h2 : 2'h1;
assign _263_ = ap_CS_fsm == 1'h1;
function [56:0] _779_;
input [56:0] a;
input [3248:0] b;
input [56:0] s;
case (s)
57'b000000000000000000000000000000000000000000000000000000001:
_779_ = b[56:0];
57'b000000000000000000000000000000000000000000000000000000010:
_779_ = b[113:57];
57'b000000000000000000000000000000000000000000000000000000100:
_779_ = b[170:114];
57'b000000000000000000000000000000000000000000000000000001000:
_779_ = b[227:171];
57'b000000000000000000000000000000000000000000000000000010000:
_779_ = b[284:228];
57'b000000000000000000000000000000000000000000000000000100000:
_779_ = b[341:285];
57'b000000000000000000000000000000000000000000000000001000000:
_779_ = b[398:342];
57'b000000000000000000000000000000000000000000000000010000000:
_779_ = b[455:399];
57'b000000000000000000000000000000000000000000000000100000000:
_779_ = b[512:456];
57'b000000000000000000000000000000000000000000000001000000000:
_779_ = b[569:513];
57'b000000000000000000000000000000000000000000000010000000000:
_779_ = b[626:570];
57'b000000000000000000000000000000000000000000000100000000000:
_779_ = b[683:627];
57'b000000000000000000000000000000000000000000001000000000000:
_779_ = b[740:684];
57'b000000000000000000000000000000000000000000010000000000000:
_779_ = b[797:741];
57'b000000000000000000000000000000000000000000100000000000000:
_779_ = b[854:798];
57'b000000000000000000000000000000000000000001000000000000000:
_779_ = b[911:855];
57'b000000000000000000000000000000000000000010000000000000000:
_779_ = b[968:912];
57'b000000000000000000000000000000000000000100000000000000000:
_779_ = b[1025:969];
57'b000000000000000000000000000000000000001000000000000000000:
_779_ = b[1082:1026];
57'b000000000000000000000000000000000000010000000000000000000:
_779_ = b[1139:1083];
57'b000000000000000000000000000000000000100000000000000000000:
_779_ = b[1196:1140];
57'b000000000000000000000000000000000001000000000000000000000:
_779_ = b[1253:1197];
57'b000000000000000000000000000000000010000000000000000000000:
_779_ = b[1310:1254];
57'b000000000000000000000000000000000100000000000000000000000:
_779_ = b[1367:1311];
57'b000000000000000000000000000000001000000000000000000000000:
_779_ = b[1424:1368];
57'b000000000000000000000000000000010000000000000000000000000:
_779_ = b[1481:1425];
57'b000000000000000000000000000000100000000000000000000000000:
_779_ = b[1538:1482];
57'b000000000000000000000000000001000000000000000000000000000:
_779_ = b[1595:1539];
57'b000000000000000000000000000010000000000000000000000000000:
_779_ = b[1652:1596];
57'b000000000000000000000000000100000000000000000000000000000:
_779_ = b[1709:1653];
57'b000000000000000000000000001000000000000000000000000000000:
_779_ = b[1766:1710];
57'b000000000000000000000000010000000000000000000000000000000:
_779_ = b[1823:1767];
57'b000000000000000000000000100000000000000000000000000000000:
_779_ = b[1880:1824];
57'b000000000000000000000001000000000000000000000000000000000:
_779_ = b[1937:1881];
57'b000000000000000000000010000000000000000000000000000000000:
_779_ = b[1994:1938];
57'b000000000000000000000100000000000000000000000000000000000:
_779_ = b[2051:1995];
57'b000000000000000000001000000000000000000000000000000000000:
_779_ = b[2108:2052];
57'b000000000000000000010000000000000000000000000000000000000:
_779_ = b[2165:2109];
57'b000000000000000000100000000000000000000000000000000000000:
_779_ = b[2222:2166];
57'b000000000000000001000000000000000000000000000000000000000:
_779_ = b[2279:2223];
57'b000000000000000010000000000000000000000000000000000000000:
_779_ = b[2336:2280];
57'b000000000000000100000000000000000000000000000000000000000:
_779_ = b[2393:2337];
57'b000000000000001000000000000000000000000000000000000000000:
_779_ = b[2450:2394];
57'b000000000000010000000000000000000000000000000000000000000:
_779_ = b[2507:2451];
57'b000000000000100000000000000000000000000000000000000000000:
_779_ = b[2564:2508];
57'b000000000001000000000000000000000000000000000000000000000:
_779_ = b[2621:2565];
57'b000000000010000000000000000000000000000000000000000000000:
_779_ = b[2678:2622];
57'b000000000100000000000000000000000000000000000000000000000:
_779_ = b[2735:2679];
57'b000000001000000000000000000000000000000000000000000000000:
_779_ = b[2792:2736];
57'b000000010000000000000000000000000000000000000000000000000:
_779_ = b[2849:2793];
57'b000000100000000000000000000000000000000000000000000000000:
_779_ = b[2906:2850];
57'b000001000000000000000000000000000000000000000000000000000:
_779_ = b[2963:2907];
57'b000010000000000000000000000000000000000000000000000000000:
_779_ = b[3020:2964];
57'b000100000000000000000000000000000000000000000000000000000:
_779_ = b[3077:3021];
57'b001000000000000000000000000000000000000000000000000000000:
_779_ = b[3134:3078];
57'b010000000000000000000000000000000000000000000000000000000:
_779_ = b[3191:3135];
57'b100000000000000000000000000000000000000000000000000000000:
_779_ = b[3248:3192];
57'b000000000000000000000000000000000000000000000000000000000:
_779_ = a;
default:
_779_ = 57'bx;
endcase
endfunction
assign ap_NS_fsm = _779_(57'hxxxxxxxxxxxxxxx, { 55'h00000000000000, _090_, 3192'h000000000000020000000000000200000000000002000000000000020000000000000200000000000002000000000000020000000000000200000000000002000000000000020000000000000200000000000002000000000000020000000000000200000000000002000000000000020000000000000200000000000002000000000000020000000000000200000000000002000000000000020000000000000200000000000002000000000000020000000000000200000000000002000000000000020000000000000200000000000002000000000000020000000000000200000000000002000000000000020000000000000200000000000002000000000000020000000000000200000000000002000000000000020000000000000200000000000002000000000000020000000000000200000000000002000000000000020000000000000200000000000002000000000000020000000000000200000000000002000000000000020000000000000200000000000002000000000000020000000000000000000000000001 }, { _263_, _319_, _318_, _317_, _316_, _315_, _314_, _313_, _312_, _311_, _310_, _309_, _308_, _307_, _306_, _305_, _304_, _303_, _302_, _301_, _300_, _299_, _298_, _297_, _296_, _295_, _294_, _293_, _292_, _291_, _290_, _289_, _288_, _287_, _286_, _285_, _284_, _283_, _282_, _281_, _280_, _279_, _278_, _277_, _276_, _275_, _274_, _273_, _272_, _271_, _270_, _269_, _268_, _267_, _266_, _265_, _264_ });
assign _264_ = ap_CS_fsm == 57'h100000000000000;
assign _265_ = ap_CS_fsm == 56'h80000000000000;
assign _266_ = ap_CS_fsm == 55'h40000000000000;
assign _267_ = ap_CS_fsm == 54'h20000000000000;
assign _268_ = ap_CS_fsm == 53'h10000000000000;
assign _269_ = ap_CS_fsm == 52'h8000000000000;
assign _270_ = ap_CS_fsm == 51'h4000000000000;
assign _271_ = ap_CS_fsm == 50'h2000000000000;
assign _272_ = ap_CS_fsm == 49'h1000000000000;
assign _273_ = ap_CS_fsm == 48'h800000000000;
assign _274_ = ap_CS_fsm == 47'h400000000000;
assign _275_ = ap_CS_fsm == 46'h200000000000;
assign _276_ = ap_CS_fsm == 45'h100000000000;
assign _277_ = ap_CS_fsm == 44'h80000000000;
assign _278_ = ap_CS_fsm == 43'h40000000000;
assign _279_ = ap_CS_fsm == 42'h20000000000;
assign _280_ = ap_CS_fsm == 41'h10000000000;
assign _281_ = ap_CS_fsm == 40'h8000000000;
assign _282_ = ap_CS_fsm == 39'h4000000000;
assign _283_ = ap_CS_fsm == 38'h2000000000;
assign _284_ = ap_CS_fsm == 37'h1000000000;
assign _285_ = ap_CS_fsm == 36'h800000000;
assign _286_ = ap_CS_fsm == 35'h400000000;
assign _287_ = ap_CS_fsm == 34'h200000000;
assign _288_ = ap_CS_fsm == 33'h100000000;
assign _289_ = ap_CS_fsm == 32'd2147483648;
assign _290_ = ap_CS_fsm == 31'h40000000;
assign _291_ = ap_CS_fsm == 30'h20000000;
assign _292_ = ap_CS_fsm == 29'h10000000;
assign _293_ = ap_CS_fsm == 28'h8000000;
assign _294_ = ap_CS_fsm == 27'h4000000;
assign _295_ = ap_CS_fsm == 26'h2000000;
assign _296_ = ap_CS_fsm == 25'h1000000;
assign _297_ = ap_CS_fsm == 24'h800000;
assign _298_ = ap_CS_fsm == 23'h400000;
assign _299_ = ap_CS_fsm == 22'h200000;
assign _300_ = ap_CS_fsm == 21'h100000;
assign _301_ = ap_CS_fsm == 20'h80000;
assign _302_ = ap_CS_fsm == 19'h40000;
assign _303_ = ap_CS_fsm == 18'h20000;
assign _304_ = ap_CS_fsm == 17'h10000;
assign _305_ = ap_CS_fsm == 16'h8000;
assign _306_ = ap_CS_fsm == 15'h4000;
assign _307_ = ap_CS_fsm == 14'h2000;
assign _308_ = ap_CS_fsm == 13'h1000;
assign _309_ = ap_CS_fsm == 12'h800;
assign _310_ = ap_CS_fsm == 11'h400;
assign _311_ = ap_CS_fsm == 10'h200;
assign _312_ = ap_CS_fsm == 9'h100;
assign _313_ = ap_CS_fsm == 8'h80;
assign _314_ = ap_CS_fsm == 7'h40;
assign _315_ = ap_CS_fsm == 6'h20;
assign _316_ = ap_CS_fsm == 5'h10;
assign _317_ = ap_CS_fsm == 4'h8;
assign _318_ = ap_CS_fsm == 3'h4;
assign _319_ = ap_CS_fsm == 2'h2;
assign op_30_ap_vld = ap_CS_fsm[56] ? 1'h1 : 1'h0;
assign ap_idle = _094_ ? 1'h1 : 1'h0;
assign _077_ = ap_CS_fsm[16] ? select_ln850_4_fu_616_p3 : select_ln850_4_reg_1649;
assign _088_ = ap_CS_fsm[16] ? xor_ln416_fu_599_p2 : xor_ln416_reg_1643;
assign _076_ = ap_CS_fsm[0] ? select_ln703_fu_249_p3[4:3] : select_ln703_reg_1402[4:3];
assign _073_ = ap_CS_fsm[42] ? select_ln353_2_fu_1243_p3 : select_ln353_2_reg_1943;
assign _072_ = _093_ ? select_ln340_1_fu_752_p3 : select_ln340_1_reg_1692;
assign _069_ = ap_CS_fsm[20] ? sel_tmp11_fu_779_p2 : sel_tmp11_reg_1697;
assign _064_ = ap_CS_fsm[54] ? ret_V_34_fu_1380_p3 : ret_V_34_reg_2032;
assign _063_ = ap_CS_fsm[51] ? grp_fu_1337_p2[33:2] : ret_V_34_cast_reg_2020;
assign _062_ = ap_CS_fsm[51] ? grp_fu_1337_p2 : ret_V_33_reg_2015;
assign _061_ = ap_CS_fsm[47] ? ret_V_32_fu_1307_p3 : ret_V_32_reg_1985;
assign _087_ = ap_CS_fsm[47] ? xor_ln1497_fu_1286_p2 : xor_ln1497_reg_1980;
assign _060_ = ap_CS_fsm[44] ? grp_fu_1265_p2[32:1] : ret_V_32_cast_reg_1968;
assign _059_ = ap_CS_fsm[44] ? grp_fu_1265_p2 : ret_V_31_reg_1963;
assign _057_ = ap_CS_fsm[39] ? grp_fu_1206_p2[32:1] : ret_V_30_cast_reg_1931;
assign _058_ = ap_CS_fsm[39] ? grp_fu_1206_p2 : ret_V_30_reg_1926;
assign _056_ = _092_ ? grp_fu_286_p2 : ret_V_2_reg_1436;
assign _055_ = ap_CS_fsm[37] ? grp_fu_1187_p2 : ret_V_29_reg_1906;
assign _070_ = ap_CS_fsm[35] ? select_ln1192_fu_1179_p3 : select_ln1192_reg_1901;
assign _054_ = ap_CS_fsm[35] ? grp_fu_1147_p2 : ret_V_28_reg_1896;
assign _075_ = ap_CS_fsm[31] ? select_ln69_fu_995_p3 : select_ln69_reg_1838;
assign _053_ = ap_CS_fsm[31] ? ret_V_27_fu_988_p3 : ret_V_27_reg_1833;
assign _049_ = ap_CS_fsm[28] ? grp_fu_951_p2[32:1] : ret_V_24_cast_reg_1821;
assign _052_ = ap_CS_fsm[28] ? grp_fu_951_p2 : ret_V_26_reg_1816;
assign _071_ = ap_CS_fsm[5] ? select_ln1347_fu_310_p3 : select_ln1347_reg_1447;
assign _048_ = ap_CS_fsm[5] ? ret_V_21_fu_303_p3 : ret_V_21_reg_1441;
assign _067_ = ap_CS_fsm[2] ? grp_fu_265_p2[4:3] : ret_V_reg_1429;
assign _047_ = ap_CS_fsm[2] ? grp_fu_265_p2 : ret_V_20_reg_1424;
assign _081_ = ap_CS_fsm[23] ? grp_fu_868_p2[7:1] : tmp_3_reg_1763;
assign _051_ = ap_CS_fsm[23] ? grp_fu_868_p2 : ret_V_25_reg_1758;
assign _046_ = ap_CS_fsm[23] ? r_fu_874_p2 : r_reg_1753;
assign _066_ = ap_CS_fsm[15] ? grp_fu_586_p2 : ret_V_9_reg_1638;
assign _039_ = ap_CS_fsm[15] ? grp_fu_576_p2[3] : p_Result_28_reg_1631;
assign _044_ = ap_CS_fsm[15] ? grp_fu_576_p2 : p_Val2_7_reg_1622;
assign _042_ = ap_CS_fsm[12] ? grp_fu_336_p2[19:6] : p_Result_7_reg_1562;
assign _041_ = ap_CS_fsm[12] ? grp_fu_336_p2[19:7] : p_Result_6_reg_1557;
assign _040_ = ap_CS_fsm[12] ? grp_fu_336_p2[6] : p_Result_29_reg_1551;
assign _038_ = ap_CS_fsm[12] ? grp_fu_336_p2[5] : p_Result_27_reg_1546;
assign _043_ = ap_CS_fsm[12] ? grp_fu_336_p2[5:2] : p_Val2_6_reg_1541;
assign _037_ = ap_CS_fsm[12] ? grp_fu_336_p2[19] : p_Result_25_reg_1533;
assign _045_ = ap_CS_fsm[12] ? grp_fu_336_p2 : r_V_1_reg_1526;
assign _085_ = ap_CS_fsm[7] ? grp_fu_324_p2[3:0] : trunc_ln790_reg_1490;
assign _080_ = ap_CS_fsm[7] ? grp_fu_324_p2[16:5] : tmp_2_reg_1484;
assign _036_ = ap_CS_fsm[7] ? grp_fu_324_p2[4] : p_Result_24_reg_1478;
assign _035_ = ap_CS_fsm[7] ? grp_fu_324_p2[16] : p_Result_23_reg_1472;
assign _068_ = ap_CS_fsm[7] ? grp_fu_324_p2 : ret_reg_1467;
assign _084_ = ap_CS_fsm[22] ? grp_fu_809_p2[2:0] : trunc_ln718_reg_1738;
assign _034_ = ap_CS_fsm[22] ? grp_fu_815_p2[3] : p_Result_22_reg_1733;
assign _082_ = ap_CS_fsm[22] ? grp_fu_809_p2[8:4] : trunc_ln2_reg_1728;
assign _032_ = ap_CS_fsm[9] ? overflow_fu_404_p2 : overflow_reg_1510;
assign _031_ = ap_CS_fsm[10] ? or_ln384_fu_430_p2 : or_ln384_reg_1516;
assign _029_ = ap_CS_fsm[21] ? op_9_V_fu_826_p3 : op_9_V_reg_1722;
assign _028_ = ap_CS_fsm[11] ? op_8_V_fu_453_p3 : op_8_V_reg_1521;
assign _027_ = ap_CS_fsm[49] ? grp_fu_1317_p2 : op_28_V_reg_1995;
assign _074_ = ap_CS_fsm[26] ? select_ln353_fu_930_p3 : select_ln353_reg_1801;
assign _025_ = ap_CS_fsm[26] ? grp_fu_908_p2 : op_10_V_reg_1795;
assign _022_ = ap_CS_fsm[1] ? icmp_ln851_fu_270_p2 : icmp_ln851_reg_1419;
assign _021_ = ap_CS_fsm[50] ? icmp_ln851_2_fu_1347_p2 : icmp_ln851_2_reg_2010;
assign _020_ = ap_CS_fsm[14] ? icmp_ln851_1_fu_581_p2 : icmp_ln851_1_reg_1617;
assign _019_ = ap_CS_fsm[8] ? icmp_ln790_fu_389_p2 : icmp_ln790_reg_1505;
assign _018_ = ap_CS_fsm[8] ? icmp_ln786_fu_377_p2 : icmp_ln786_reg_1500;
assign _017_ = ap_CS_fsm[8] ? icmp_ln768_fu_372_p2 : icmp_ln768_reg_1495;
assign _016_ = ap_CS_fsm[34] ? icmp_ln1497_fu_1138_p2 : icmp_ln1497_reg_1886;
assign _024_ = ap_CS_fsm[34] ? newsignbit_fu_1123_p2 : newsignbit_reg_1879;
assign _026_ = ap_CS_fsm[33] ? grp_fu_1003_p2 : op_23_V_reg_1874;
assign _079_ = ap_CS_fsm[33] ? signbit_3_fu_1114_p2 : signbit_3_reg_1869;
assign _023_ = ap_CS_fsm[33] ? lhs_V_2_fu_1093_p2 : lhs_V_2_reg_1864;
assign _014_ = ap_CS_fsm[33] ? r_V_fu_1053_p3[1] : carry_reg_1859;
assign _033_ = ap_CS_fsm[33] ? r_V_fu_1053_p3[1] : p_Result_21_reg_1853;
assign _083_ = ap_CS_fsm[33] ? r_V_fu_1053_p3[0] : trunc_ln415_reg_1848;
assign _013_ = ap_CS_fsm[17] ? carry_2_fu_623_p2 : carry_2_reg_1654;
assign _011_ = ap_CS_fsm[18] ? and_ln786_fu_653_p2 : and_ln786_reg_1673;
assign _089_ = ap_CS_fsm[18] ? xor_ln785_3_fu_648_p2 : xor_ln785_3_reg_1667;
assign _015_ = ap_CS_fsm[18] ? deleted_zeros_fu_627_p3 : deleted_zeros_reg_1661;
assign _010_ = ap_CS_fsm[19] ? and_ln785_1_fu_703_p2 : and_ln785_1_reg_1687;
assign _030_ = ap_CS_fsm[19] ? or_ln340_fu_688_p2 : or_ln340_reg_1681;
assign _078_ = ap_CS_fsm[24] ? { tmp_3_reg_1763[6], tmp_3_reg_1763 } : sext_ln850_reg_1773;
assign _009_ = ap_CS_fsm[24] ? and_ln408_fu_889_p2 : and_ln408_reg_1768;
assign _007_ = ap_CS_fsm[25] ? grp_fu_896_p2 : add_ln691_reg_1790;
assign _006_ = _091_ ? grp_fu_1363_p2 : add_ln691_4_reg_2027;
assign _005_ = ap_CS_fsm[46] ? grp_fu_1281_p2 : add_ln691_3_reg_1975;
assign _004_ = ap_CS_fsm[41] ? grp_fu_1222_p2 : add_ln691_2_reg_1938;
assign _003_ = ap_CS_fsm[30] ? grp_fu_967_p2 : add_ln691_1_reg_1828;
assign _086_ = ap_CS_fsm[13] ? grp_fu_517_p2[2:0] : trunc_ln851_1_reg_1607;
assign _065_ = ap_CS_fsm[13] ? grp_fu_517_p2[8:3] : ret_V_7_reg_1600;
assign _050_ = ap_CS_fsm[13] ? grp_fu_517_p2 : ret_V_24_reg_1595;
assign _001_ = ap_CS_fsm[13] ? Range1_all_zeros_fu_554_p2 : Range1_all_zeros_reg_1590;
assign _000_ = ap_CS_fsm[13] ? Range1_all_ones_fu_549_p2 : Range1_all_ones_reg_1583;
assign _002_ = ap_CS_fsm[13] ? Range2_all_ones_fu_544_p2 : Range2_all_ones_reg_1578;
assign _008_ = ap_CS_fsm[13] ? and_ln406_fu_538_p2 : and_ln406_reg_1573;
assign _012_ = ap_rst ? 57'h000000000000001 : ap_NS_fsm;
assign Range1_all_ones_fu_549_p2 = _099_ ? 1'h1 : 1'h0;
assign Range1_all_zeros_fu_554_p2 = _100_ ? 1'h1 : 1'h0;
assign Range2_all_ones_fu_544_p2 = _101_ ? 1'h1 : 1'h0;
assign deleted_ones_fu_642_p3 = carry_2_reg_1654 ? and_ln780_fu_637_p2 : Range1_all_ones_reg_1583;
assign deleted_zeros_fu_627_p3 = carry_2_reg_1654 ? Range1_all_ones_reg_1583 : Range1_all_zeros_reg_1590;
assign icmp_ln1497_fu_1138_p2 = _256_ ? 1'h1 : 1'h0;
assign icmp_ln768_fu_372_p2 = _257_ ? 1'h1 : 1'h0;
assign icmp_ln786_fu_377_p2 = _258_ ? 1'h1 : 1'h0;
assign icmp_ln790_fu_389_p2 = _102_ ? 1'h1 : 1'h0;
assign icmp_ln851_1_fu_581_p2 = _103_ ? 1'h1 : 1'h0;
assign icmp_ln851_2_fu_1347_p2 = _259_ ? 1'h1 : 1'h0;
assign icmp_ln851_fu_270_p2 = _104_ ? 1'h1 : 1'h0;
assign lhs_V_2_fu_1093_p2 = _260_ ? 1'h1 : 1'h0;
assign op_8_V_fu_453_p3 = or_ln384_reg_1516 ? select_ln384_fu_446_p3 : { ret_reg_1467[4:0], 3'h0 };
assign op_9_V_fu_826_p3 = sel_tmp11_reg_1697 ? p_Val2_7_reg_1622 : select_ln785_fu_821_p3;
assign r_V_fu_1053_p3 = ret_V_22_fu_1033_p2 ? { op_5[0], 1'h0 } : op_5;
assign r_fu_874_p2 = _261_ ? 1'h1 : 1'h0;
assign ret_V_21_fu_303_p3 = ret_V_20_reg_1424[4] ? select_ln850_fu_298_p3 : ret_V_reg_1429;
assign ret_V_27_fu_988_p3 = ret_V_26_reg_1816[33] ? select_ln850_3_fu_982_p3 : ret_V_24_cast_reg_1821;
assign ret_V_32_fu_1307_p3 = ret_V_31_reg_1963[33] ? select_ln850_5_fu_1301_p3 : ret_V_32_cast_reg_1968;
assign ret_V_34_fu_1380_p3 = ret_V_33_reg_2015[34] ? select_ln850_6_fu_1375_p3 : ret_V_34_cast_reg_2020;
assign select_ln1192_fu_1179_p3 = op_14_V_fu_1174_p2 ? 32'd4294967295 : 32'd0;
assign select_ln1347_fu_310_p3 = op_2 ? 17'h1ffff : 17'h00000;
assign select_ln340_1_fu_752_p3 = or_ln340_1_fu_748_p2 ? { p_Result_29_reg_1551, p_Val2_8_fu_734_p2 } : p_Val2_7_reg_1622;
assign select_ln340_fu_1161_p3 = newsignbit_reg_1879 ? xor_ln785_fu_1156_p2 : neg_src_2_fu_1152_p2;
assign select_ln353_2_fu_1243_p3 = ret_V_30_reg_1926[33] ? select_ln850_8_fu_1237_p3 : ret_V_30_cast_reg_1931;
assign select_ln353_fu_930_p3 = ret_V_25_reg_1758[7] ? select_ln850_7_fu_924_p3 : sext_ln850_reg_1773;
assign select_ln384_fu_446_p3 = overflow_reg_1510 ? 8'h7f : 8'h81;
assign select_ln69_fu_995_p3 = op_12 ? 32'd4294967295 : 32'd0;
assign select_ln703_fu_249_p3 = op_2 ? 5'h18 : 5'h00;
assign select_ln785_fu_821_p3 = and_ln785_1_reg_1687 ? p_Val2_7_reg_1622 : select_ln340_1_reg_1692;
assign select_ln850_2_fu_611_p3 = icmp_ln851_1_reg_1617 ? ret_V_7_reg_1600 : ret_V_9_reg_1638;
assign select_ln850_3_fu_982_p3 = op_10_V_reg_1795[0] ? add_ln691_1_reg_1828 : ret_V_24_cast_reg_1821;
assign select_ln850_4_fu_616_p3 = ret_V_24_reg_1595[8] ? select_ln850_2_fu_611_p3 : ret_V_7_reg_1600;
assign select_ln850_5_fu_1301_p3 = op_16[0] ? add_ln691_3_reg_1975 : ret_V_32_cast_reg_1968;
assign select_ln850_6_fu_1375_p3 = icmp_ln851_2_reg_2010 ? add_ln691_4_reg_2027 : ret_V_34_cast_reg_2020;
assign select_ln850_7_fu_924_p3 = op_9_V_reg_1722[0] ? add_ln691_reg_1790 : sext_ln850_reg_1773;
assign select_ln850_8_fu_1237_p3 = op_15[0] ? add_ln691_2_reg_1938 : ret_V_30_cast_reg_1931;
assign select_ln850_fu_298_p3 = icmp_ln851_reg_1419 ? ret_V_reg_1429 : ret_V_2_reg_1436;
assign signbit_3_fu_1114_p2 = _262_ ? 1'h1 : 1'h0;
assign newsignbit_fu_1123_p2 = trunc_ln415_reg_1848 ^ carry_reg_1859;
assign ret_V_22_fu_1033_p2 = op_5[1] ^ and_ln850_fu_1027_p2;
assign xor_ln365_fu_722_p2 = r_V_1_reg_1526[6] ^ p_Val2_7_reg_1622[3];
assign ap_CS_fsm_state1 = ap_CS_fsm[0];
assign ap_CS_fsm_state10 = ap_CS_fsm[9];
assign ap_CS_fsm_state11 = ap_CS_fsm[10];
assign ap_CS_fsm_state12 = ap_CS_fsm[11];
assign ap_CS_fsm_state13 = ap_CS_fsm[12];
assign ap_CS_fsm_state14 = ap_CS_fsm[13];
assign ap_CS_fsm_state15 = ap_CS_fsm[14];
assign ap_CS_fsm_state16 = ap_CS_fsm[15];
assign ap_CS_fsm_state17 = ap_CS_fsm[16];
assign ap_CS_fsm_state18 = ap_CS_fsm[17];
assign ap_CS_fsm_state19 = ap_CS_fsm[18];
assign ap_CS_fsm_state2 = ap_CS_fsm[1];
assign ap_CS_fsm_state20 = ap_CS_fsm[19];
assign ap_CS_fsm_state21 = ap_CS_fsm[20];
assign ap_CS_fsm_state22 = ap_CS_fsm[21];
assign ap_CS_fsm_state23 = ap_CS_fsm[22];
assign ap_CS_fsm_state24 = ap_CS_fsm[23];
assign ap_CS_fsm_state25 = ap_CS_fsm[24];
assign ap_CS_fsm_state26 = ap_CS_fsm[25];
assign ap_CS_fsm_state27 = ap_CS_fsm[26];
assign ap_CS_fsm_state28 = ap_CS_fsm[27];
assign ap_CS_fsm_state29 = ap_CS_fsm[28];
assign ap_CS_fsm_state3 = ap_CS_fsm[2];
assign ap_CS_fsm_state30 = ap_CS_fsm[29];
assign ap_CS_fsm_state31 = ap_CS_fsm[30];
assign ap_CS_fsm_state32 = ap_CS_fsm[31];
assign ap_CS_fsm_state33 = ap_CS_fsm[32];
assign ap_CS_fsm_state34 = ap_CS_fsm[33];
assign ap_CS_fsm_state35 = ap_CS_fsm[34];
assign ap_CS_fsm_state36 = ap_CS_fsm[35];
assign ap_CS_fsm_state37 = ap_CS_fsm[36];
assign ap_CS_fsm_state38 = ap_CS_fsm[37];
assign ap_CS_fsm_state39 = ap_CS_fsm[38];
assign ap_CS_fsm_state4 = ap_CS_fsm[3];
assign ap_CS_fsm_state40 = ap_CS_fsm[39];
assign ap_CS_fsm_state41 = ap_CS_fsm[40];
assign ap_CS_fsm_state42 = ap_CS_fsm[41];
assign ap_CS_fsm_state43 = ap_CS_fsm[42];
assign ap_CS_fsm_state44 = ap_CS_fsm[43];
assign ap_CS_fsm_state45 = ap_CS_fsm[44];
assign ap_CS_fsm_state46 = ap_CS_fsm[45];
assign ap_CS_fsm_state47 = ap_CS_fsm[46];
assign ap_CS_fsm_state48 = ap_CS_fsm[47];
assign ap_CS_fsm_state49 = ap_CS_fsm[48];
assign ap_CS_fsm_state5 = ap_CS_fsm[4];
assign ap_CS_fsm_state50 = ap_CS_fsm[49];
assign ap_CS_fsm_state51 = ap_CS_fsm[50];
assign ap_CS_fsm_state52 = ap_CS_fsm[51];
assign ap_CS_fsm_state53 = ap_CS_fsm[52];
assign ap_CS_fsm_state54 = ap_CS_fsm[53];
assign ap_CS_fsm_state55 = ap_CS_fsm[54];
assign ap_CS_fsm_state56 = ap_CS_fsm[55];
assign ap_CS_fsm_state57 = ap_CS_fsm[56];
assign ap_CS_fsm_state6 = ap_CS_fsm[5];
assign ap_CS_fsm_state7 = ap_CS_fsm[6];
assign ap_CS_fsm_state8 = ap_CS_fsm[7];
assign ap_CS_fsm_state9 = ap_CS_fsm[8];
assign ap_done = op_30_ap_vld;
assign ap_ready = op_30_ap_vld;
assign grp_fu_1147_p1 = { 31'h00000000, lhs_V_2_reg_1864 };
assign grp_fu_1206_p0 = { ret_V_29_reg_1906[31], ret_V_29_reg_1906, 1'h0 };
assign grp_fu_1206_p1 = { op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15 };
assign grp_fu_1265_p0 = { select_ln353_2_reg_1943[31], select_ln353_2_reg_1943, 1'h0 };
assign grp_fu_1265_p1 = { op_16[15], op_16[15], op_16[15], op_16[15], op_16[15], op_16[15], op_16[15], op_16[15], op_16[15], op_16[15], op_16[15], op_16[15], op_16[15], op_16[15], op_16[15], op_16[15], op_16[15], op_16[15], op_16 };
assign grp_fu_1317_p1 = { 31'h00000000, xor_ln1497_reg_1980 };
assign grp_fu_1337_p0 = { op_28_V_reg_1995[31], op_28_V_reg_1995, 2'h0 };
assign grp_fu_1337_p1 = { op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18 };
assign grp_fu_1391_p1 = { 28'h0000000, op_19 };
assign grp_fu_265_p1 = { op_3[3], op_3 };
assign grp_fu_324_p1 = { 1'h0, ret_V_21_reg_1441[1], ret_V_21_reg_1441[1], ret_V_21_reg_1441[1], ret_V_21_reg_1441[1], ret_V_21_reg_1441[1], ret_V_21_reg_1441[1], ret_V_21_reg_1441[1], ret_V_21_reg_1441[1], ret_V_21_reg_1441[1], ret_V_21_reg_1441[1], ret_V_21_reg_1441[1], ret_V_21_reg_1441[1], ret_V_21_reg_1441[1], ret_V_21_reg_1441[1], ret_V_21_reg_1441 };
assign grp_fu_336_p0 = { ret_V_21_reg_1441[1], ret_V_21_reg_1441[1], ret_V_21_reg_1441[1], ret_V_21_reg_1441[1], ret_V_21_reg_1441[1], ret_V_21_reg_1441[1], ret_V_21_reg_1441[1], ret_V_21_reg_1441[1], ret_V_21_reg_1441[1], ret_V_21_reg_1441[1], ret_V_21_reg_1441[1], ret_V_21_reg_1441[1], ret_V_21_reg_1441[1], ret_V_21_reg_1441[1], ret_V_21_reg_1441 };
assign grp_fu_336_p00 = { 4'h0, ret_V_21_reg_1441[1], ret_V_21_reg_1441[1], ret_V_21_reg_1441[1], ret_V_21_reg_1441[1], ret_V_21_reg_1441[1], ret_V_21_reg_1441[1], ret_V_21_reg_1441[1], ret_V_21_reg_1441[1], ret_V_21_reg_1441[1], ret_V_21_reg_1441[1], ret_V_21_reg_1441[1], ret_V_21_reg_1441[1], ret_V_21_reg_1441[1], ret_V_21_reg_1441[1], ret_V_21_reg_1441 };
assign grp_fu_517_p0 = { op_8_V_reg_1521[7], op_8_V_reg_1521 };
assign grp_fu_576_p1 = { 3'h0, and_ln406_reg_1573 };
assign grp_fu_809_p0 = { op_3[3], op_3[3], op_3[3], op_3, 2'h0 };
assign grp_fu_809_p1 = { op_6[7], op_6 };
assign grp_fu_815_p0 = { op_3[1:0], 2'h0 };
assign grp_fu_815_p1 = op_6[3:0];
assign grp_fu_868_p0 = { select_ln850_4_reg_1649[5], select_ln850_4_reg_1649, 1'h0 };
assign grp_fu_868_p1 = { op_9_V_reg_1722[3], op_9_V_reg_1722[3], op_9_V_reg_1722[3], op_9_V_reg_1722[3], op_9_V_reg_1722 };
assign grp_fu_896_p0 = { tmp_3_reg_1763[6], tmp_3_reg_1763 };
assign grp_fu_908_p0 = { trunc_ln2_reg_1728[4], trunc_ln2_reg_1728 };
assign grp_fu_908_p1 = { 5'h00, and_ln408_reg_1768 };
assign grp_fu_951_p0 = { select_ln353_reg_1801[7], select_ln353_reg_1801[7], select_ln353_reg_1801[7], select_ln353_reg_1801[7], select_ln353_reg_1801[7], select_ln353_reg_1801[7], select_ln353_reg_1801[7], select_ln353_reg_1801[7], select_ln353_reg_1801[7], select_ln353_reg_1801[7], select_ln353_reg_1801[7], select_ln353_reg_1801[7], select_ln353_reg_1801[7], select_ln353_reg_1801[7], select_ln353_reg_1801[7], select_ln353_reg_1801[7], select_ln353_reg_1801[7], select_ln353_reg_1801[7], select_ln353_reg_1801[7], select_ln353_reg_1801[7], select_ln353_reg_1801[7], select_ln353_reg_1801[7], select_ln353_reg_1801[7], select_ln353_reg_1801[7], select_ln353_reg_1801[7], select_ln353_reg_1801, 1'h0 };
assign grp_fu_951_p1 = { op_10_V_reg_1795[5], op_10_V_reg_1795[5], op_10_V_reg_1795[5], op_10_V_reg_1795[5], op_10_V_reg_1795[5], op_10_V_reg_1795[5], op_10_V_reg_1795[5], op_10_V_reg_1795[5], op_10_V_reg_1795[5], op_10_V_reg_1795[5], op_10_V_reg_1795[5], op_10_V_reg_1795[5], op_10_V_reg_1795[5], op_10_V_reg_1795[5], op_10_V_reg_1795[5], op_10_V_reg_1795[5], op_10_V_reg_1795[5], op_10_V_reg_1795[5], op_10_V_reg_1795[5], op_10_V_reg_1795[5], op_10_V_reg_1795[5], op_10_V_reg_1795[5], op_10_V_reg_1795[5], op_10_V_reg_1795[5], op_10_V_reg_1795[5], op_10_V_reg_1795[5], op_10_V_reg_1795[5], op_10_V_reg_1795[5], op_10_V_reg_1795 };
assign lhs_fu_785_p1 = op_3;
assign lhs_fu_785_p3 = { op_3, 2'h0 };
assign op_11_V_fu_1127_p3 = { signbit_3_reg_1869, 1'h0 };
assign op_30 = grp_fu_1391_p2;
assign p_Result_14_fu_739_p4 = { p_Result_29_reg_1551, p_Val2_8_fu_734_p2 };
assign p_Result_15_fu_604_p3 = ret_V_24_reg_1595[8];
assign p_Result_16_fu_914_p3 = ret_V_25_reg_1758[7];
assign p_Result_17_fu_972_p3 = ret_V_26_reg_1816[33];
assign p_Result_18_fu_1227_p3 = ret_V_30_reg_1926[33];
assign p_Result_19_fu_1291_p3 = ret_V_31_reg_1963[33];
assign p_Result_1_fu_1015_p1 = op_5;
assign p_Result_1_fu_1015_p3 = op_5[1];
assign p_Result_20_fu_1368_p3 = ret_V_33_reg_2015[34];
assign p_Result_26_fu_523_p3 = r_V_1_reg_1526[1];
assign p_Result_3_fu_382_p3 = { trunc_ln790_reg_1490, 3'h0 };
assign p_Result_s_fu_291_p3 = ret_V_20_reg_1424[4];
assign p_Val2_4_fu_438_p3 = { ret_reg_1467[4:0], 3'h0 };
assign r_1_fu_530_p1 = r_V_1_reg_1526[0];
assign r_V_fu_1053_p2 = op_5;
assign ret_V_4_fu_1007_p1 = op_5;
assign ret_V_4_fu_1007_p3 = op_5[1];
assign rhs_2_fu_857_p3 = { select_ln850_4_reg_1649, 1'h0 };
assign rhs_6_fu_1195_p3 = { ret_V_29_reg_1906, 1'h0 };
assign rhs_7_fu_1254_p3 = { select_ln353_2_reg_1943, 1'h0 };
assign rhs_9_fu_1326_p3 = { op_28_V_reg_1995, 2'h0 };
assign sext_ln1299_1_fu_1039_p0 = op_5;
assign sext_ln1299_1_fu_1039_p1 = { op_5[1], op_5[1], op_5[1], op_5[1], op_5[1], op_5[1], op_5[1], op_5[1], op_5[1], op_5[1], op_5[1], op_5[1], op_5[1], op_5[1], op_5[1], op_5[1], op_5 };
assign sext_ln1299_2_fu_1043_p0 = op_5;
assign sext_ln1299_2_fu_1043_p1 = { op_5[1], op_5[1], op_5[1], op_5[1], op_5 };
assign sext_ln1299_fu_1120_p0 = op_5;
assign sext_ln1299_fu_1120_p1 = { op_5[1], op_5 };
assign sext_ln1347_fu_317_p1 = { ret_V_21_reg_1441[1], ret_V_21_reg_1441[1], ret_V_21_reg_1441[1], ret_V_21_reg_1441[1], ret_V_21_reg_1441[1], ret_V_21_reg_1441[1], ret_V_21_reg_1441[1], ret_V_21_reg_1441[1], ret_V_21_reg_1441[1], ret_V_21_reg_1441[1], ret_V_21_reg_1441[1], ret_V_21_reg_1441[1], ret_V_21_reg_1441[1], ret_V_21_reg_1441[1], ret_V_21_reg_1441 };
assign sext_ln1499_fu_1106_p1 = { ret_V_21_reg_1441[1], ret_V_21_reg_1441[1], ret_V_21_reg_1441[1], ret_V_21_reg_1441[1], ret_V_21_reg_1441[1], ret_V_21_reg_1441[1], ret_V_21_reg_1441[1], ret_V_21_reg_1441[1], ret_V_21_reg_1441[1], ret_V_21_reg_1441[1], ret_V_21_reg_1441[1], ret_V_21_reg_1441[1], ret_V_21_reg_1441[1], ret_V_21_reg_1441[1], ret_V_21_reg_1441, 1'h0 };
assign sext_ln703_1_fu_796_p0 = op_6;
assign sext_ln703_4_fu_1191_p0 = op_15;
assign sext_ln703_5_fu_1250_p0 = op_16;
assign sext_ln703_6_fu_1322_p0 = op_18;
assign sext_ln703_fu_257_p0 = op_3;
assign sext_ln850_fu_893_p1 = { tmp_3_reg_1763[6], tmp_3_reg_1763 };
assign shl_ln1192_fu_804_p0 = op_3;
assign shl_ln1299_fu_1047_p0 = op_5;
assign shl_ln1299_fu_1047_p2 = { op_5[0], 1'h0 };
assign shl_ln1_fu_1081_p3 = { op_7, 1'h0 };
assign tmp_1_fu_715_p3 = p_Val2_7_reg_1622[3];
assign tmp_7_fu_1099_p3 = { ret_V_21_reg_1441, 1'h0 };
assign tmp_8_fu_940_p3 = { select_ln353_reg_1801, 1'h0 };
assign tmp_fu_708_p3 = r_V_1_reg_1526[6];
assign trunc_ln1192_1_fu_800_p0 = op_6;
assign trunc_ln1192_fu_261_p0 = op_3;
assign trunc_ln1192_fu_261_p1 = op_3[2:0];
assign trunc_ln415_fu_1061_p1 = r_V_fu_1053_p3[0];
assign trunc_ln718_fu_850_p1 = grp_fu_809_p2[2:0];
assign trunc_ln731_fu_435_p1 = ret_reg_1467[4:0];
assign trunc_ln790_fu_368_p1 = grp_fu_324_p2[3:0];
assign trunc_ln851_1_fu_569_p1 = grp_fu_517_p2[2:0];
assign trunc_ln851_2_fu_921_p1 = op_9_V_reg_1722[0];
assign trunc_ln851_3_fu_979_p1 = op_10_V_reg_1795[0];
assign trunc_ln851_4_fu_1234_p0 = op_15;
assign trunc_ln851_4_fu_1234_p1 = op_15[0];
assign trunc_ln851_5_fu_1298_p0 = op_16;
assign trunc_ln851_5_fu_1298_p1 = op_16[0];
assign trunc_ln851_6_fu_1343_p0 = op_18;
assign trunc_ln851_6_fu_1343_p1 = op_18[1:0];
assign trunc_ln851_fu_1023_p0 = op_5;
assign trunc_ln851_fu_1023_p1 = op_5[0];
assign zext_ln1497_fu_1134_p1 = { 1'h0, signbit_3_reg_1869, 1'h0 };
assign zext_ln1499_1_fu_1110_p1 = { 1'h0, ret_V_21_reg_1441[1], ret_V_21_reg_1441[1], ret_V_21_reg_1441[1], ret_V_21_reg_1441[1], ret_V_21_reg_1441[1], ret_V_21_reg_1441[1], ret_V_21_reg_1441[1], ret_V_21_reg_1441[1], ret_V_21_reg_1441[1], ret_V_21_reg_1441[1], ret_V_21_reg_1441[1], ret_V_21_reg_1441[1], ret_V_21_reg_1441[1], ret_V_21_reg_1441[1], ret_V_21_reg_1441, 1'h0 };
assign zext_ln1499_fu_1089_p1 = { 1'h0, op_7, 1'h0 };
assign \sub_17ns_17ns_17_2_1_U3.top_sub_17ns_17ns_17_2_1_Adder_2_U.ain_s0  = \sub_17ns_17ns_17_2_1_U3.top_sub_17ns_17ns_17_2_1_Adder_2_U.a ;
assign \sub_17ns_17ns_17_2_1_U3.top_sub_17ns_17ns_17_2_1_Adder_2_U.s  = { \sub_17ns_17ns_17_2_1_U3.top_sub_17ns_17ns_17_2_1_Adder_2_U.fas_s2 , \sub_17ns_17ns_17_2_1_U3.top_sub_17ns_17ns_17_2_1_Adder_2_U.sum_s1  };
assign \sub_17ns_17ns_17_2_1_U3.top_sub_17ns_17ns_17_2_1_Adder_2_U.u2.a  = \sub_17ns_17ns_17_2_1_U3.top_sub_17ns_17ns_17_2_1_Adder_2_U.ain_s1 ;
assign \sub_17ns_17ns_17_2_1_U3.top_sub_17ns_17ns_17_2_1_Adder_2_U.u2.b  = \sub_17ns_17ns_17_2_1_U3.top_sub_17ns_17ns_17_2_1_Adder_2_U.bin_s1 ;
assign \sub_17ns_17ns_17_2_1_U3.top_sub_17ns_17ns_17_2_1_Adder_2_U.u2.cin  = \sub_17ns_17ns_17_2_1_U3.top_sub_17ns_17ns_17_2_1_Adder_2_U.carry_s1 ;
assign \sub_17ns_17ns_17_2_1_U3.top_sub_17ns_17ns_17_2_1_Adder_2_U.facout_s2  = \sub_17ns_17ns_17_2_1_U3.top_sub_17ns_17ns_17_2_1_Adder_2_U.u2.cout ;
assign \sub_17ns_17ns_17_2_1_U3.top_sub_17ns_17ns_17_2_1_Adder_2_U.fas_s2  = \sub_17ns_17ns_17_2_1_U3.top_sub_17ns_17ns_17_2_1_Adder_2_U.u2.s ;
assign \sub_17ns_17ns_17_2_1_U3.top_sub_17ns_17ns_17_2_1_Adder_2_U.u1.a  = \sub_17ns_17ns_17_2_1_U3.top_sub_17ns_17ns_17_2_1_Adder_2_U.a [7:0];
assign \sub_17ns_17ns_17_2_1_U3.top_sub_17ns_17ns_17_2_1_Adder_2_U.u1.b  = \sub_17ns_17ns_17_2_1_U3.top_sub_17ns_17ns_17_2_1_Adder_2_U.bin_s0 [7:0];
assign \sub_17ns_17ns_17_2_1_U3.top_sub_17ns_17ns_17_2_1_Adder_2_U.u1.cin  = 1'h1;
assign \sub_17ns_17ns_17_2_1_U3.top_sub_17ns_17ns_17_2_1_Adder_2_U.facout_s1  = \sub_17ns_17ns_17_2_1_U3.top_sub_17ns_17ns_17_2_1_Adder_2_U.u1.cout ;
assign \sub_17ns_17ns_17_2_1_U3.top_sub_17ns_17ns_17_2_1_Adder_2_U.fas_s1  = \sub_17ns_17ns_17_2_1_U3.top_sub_17ns_17ns_17_2_1_Adder_2_U.u1.s ;
assign \sub_17ns_17ns_17_2_1_U3.top_sub_17ns_17ns_17_2_1_Adder_2_U.a  = \sub_17ns_17ns_17_2_1_U3.din0 ;
assign \sub_17ns_17ns_17_2_1_U3.top_sub_17ns_17ns_17_2_1_Adder_2_U.b  = \sub_17ns_17ns_17_2_1_U3.din1 ;
assign \sub_17ns_17ns_17_2_1_U3.top_sub_17ns_17ns_17_2_1_Adder_2_U.ce  = \sub_17ns_17ns_17_2_1_U3.ce ;
assign \sub_17ns_17ns_17_2_1_U3.top_sub_17ns_17ns_17_2_1_Adder_2_U.clk  = \sub_17ns_17ns_17_2_1_U3.clk ;
assign \sub_17ns_17ns_17_2_1_U3.top_sub_17ns_17ns_17_2_1_Adder_2_U.reset  = \sub_17ns_17ns_17_2_1_U3.reset ;
assign \sub_17ns_17ns_17_2_1_U3.dout  = \sub_17ns_17ns_17_2_1_U3.top_sub_17ns_17ns_17_2_1_Adder_2_U.s ;
assign \sub_17ns_17ns_17_2_1_U3.ce  = 1'h1;
assign \sub_17ns_17ns_17_2_1_U3.clk  = ap_clk;
assign \sub_17ns_17ns_17_2_1_U3.din0  = select_ln1347_reg_1447;
assign \sub_17ns_17ns_17_2_1_U3.din1  = { 1'h0, ret_V_21_reg_1441[1], ret_V_21_reg_1441[1], ret_V_21_reg_1441[1], ret_V_21_reg_1441[1], ret_V_21_reg_1441[1], ret_V_21_reg_1441[1], ret_V_21_reg_1441[1], ret_V_21_reg_1441[1], ret_V_21_reg_1441[1], ret_V_21_reg_1441[1], ret_V_21_reg_1441[1], ret_V_21_reg_1441[1], ret_V_21_reg_1441[1], ret_V_21_reg_1441[1], ret_V_21_reg_1441 };
assign grp_fu_324_p2 = \sub_17ns_17ns_17_2_1_U3.dout ;
assign \sub_17ns_17ns_17_2_1_U3.reset  = ap_rst;
assign \mul_16ns_4s_20_7_1_U4.top_mul_16ns_4s_20_7_1_Mul_DSP_0_U.p  = \mul_16ns_4s_20_7_1_U4.top_mul_16ns_4s_20_7_1_Mul_DSP_0_U.buff4 ;
assign \mul_16ns_4s_20_7_1_U4.top_mul_16ns_4s_20_7_1_Mul_DSP_0_U.a  = \mul_16ns_4s_20_7_1_U4.din0 ;
assign \mul_16ns_4s_20_7_1_U4.top_mul_16ns_4s_20_7_1_Mul_DSP_0_U.b  = \mul_16ns_4s_20_7_1_U4.din1 ;
assign \mul_16ns_4s_20_7_1_U4.top_mul_16ns_4s_20_7_1_Mul_DSP_0_U.ce  = \mul_16ns_4s_20_7_1_U4.ce ;
assign \mul_16ns_4s_20_7_1_U4.top_mul_16ns_4s_20_7_1_Mul_DSP_0_U.clk  = \mul_16ns_4s_20_7_1_U4.clk ;
assign \mul_16ns_4s_20_7_1_U4.dout  = \mul_16ns_4s_20_7_1_U4.top_mul_16ns_4s_20_7_1_Mul_DSP_0_U.p ;
assign \mul_16ns_4s_20_7_1_U4.ce  = 1'h1;
assign \mul_16ns_4s_20_7_1_U4.clk  = ap_clk;
assign \mul_16ns_4s_20_7_1_U4.din0  = { ret_V_21_reg_1441[1], ret_V_21_reg_1441[1], ret_V_21_reg_1441[1], ret_V_21_reg_1441[1], ret_V_21_reg_1441[1], ret_V_21_reg_1441[1], ret_V_21_reg_1441[1], ret_V_21_reg_1441[1], ret_V_21_reg_1441[1], ret_V_21_reg_1441[1], ret_V_21_reg_1441[1], ret_V_21_reg_1441[1], ret_V_21_reg_1441[1], ret_V_21_reg_1441[1], ret_V_21_reg_1441 };
assign \mul_16ns_4s_20_7_1_U4.din1  = op_3;
assign grp_fu_336_p2 = \mul_16ns_4s_20_7_1_U4.dout ;
assign \mul_16ns_4s_20_7_1_U4.reset  = ap_rst;
assign \add_9s_9s_9_2_1_U8.top_add_9s_9s_9_2_1_Adder_6_U.ain_s0  = \add_9s_9s_9_2_1_U8.top_add_9s_9s_9_2_1_Adder_6_U.a ;
assign \add_9s_9s_9_2_1_U8.top_add_9s_9s_9_2_1_Adder_6_U.bin_s0  = \add_9s_9s_9_2_1_U8.top_add_9s_9s_9_2_1_Adder_6_U.b ;
assign \add_9s_9s_9_2_1_U8.top_add_9s_9s_9_2_1_Adder_6_U.s  = { \add_9s_9s_9_2_1_U8.top_add_9s_9s_9_2_1_Adder_6_U.fas_s2 , \add_9s_9s_9_2_1_U8.top_add_9s_9s_9_2_1_Adder_6_U.sum_s1  };
assign \add_9s_9s_9_2_1_U8.top_add_9s_9s_9_2_1_Adder_6_U.u2.a  = \add_9s_9s_9_2_1_U8.top_add_9s_9s_9_2_1_Adder_6_U.ain_s1 ;
assign \add_9s_9s_9_2_1_U8.top_add_9s_9s_9_2_1_Adder_6_U.u2.b  = \add_9s_9s_9_2_1_U8.top_add_9s_9s_9_2_1_Adder_6_U.bin_s1 ;
assign \add_9s_9s_9_2_1_U8.top_add_9s_9s_9_2_1_Adder_6_U.u2.cin  = \add_9s_9s_9_2_1_U8.top_add_9s_9s_9_2_1_Adder_6_U.carry_s1 ;
assign \add_9s_9s_9_2_1_U8.top_add_9s_9s_9_2_1_Adder_6_U.facout_s2  = \add_9s_9s_9_2_1_U8.top_add_9s_9s_9_2_1_Adder_6_U.u2.cout ;
assign \add_9s_9s_9_2_1_U8.top_add_9s_9s_9_2_1_Adder_6_U.fas_s2  = \add_9s_9s_9_2_1_U8.top_add_9s_9s_9_2_1_Adder_6_U.u2.s ;
assign \add_9s_9s_9_2_1_U8.top_add_9s_9s_9_2_1_Adder_6_U.u1.a  = \add_9s_9s_9_2_1_U8.top_add_9s_9s_9_2_1_Adder_6_U.a [3:0];
assign \add_9s_9s_9_2_1_U8.top_add_9s_9s_9_2_1_Adder_6_U.u1.b  = \add_9s_9s_9_2_1_U8.top_add_9s_9s_9_2_1_Adder_6_U.b [3:0];
assign \add_9s_9s_9_2_1_U8.top_add_9s_9s_9_2_1_Adder_6_U.u1.cin  = 1'h0;
assign \add_9s_9s_9_2_1_U8.top_add_9s_9s_9_2_1_Adder_6_U.facout_s1  = \add_9s_9s_9_2_1_U8.top_add_9s_9s_9_2_1_Adder_6_U.u1.cout ;
assign \add_9s_9s_9_2_1_U8.top_add_9s_9s_9_2_1_Adder_6_U.fas_s1  = \add_9s_9s_9_2_1_U8.top_add_9s_9s_9_2_1_Adder_6_U.u1.s ;
assign \add_9s_9s_9_2_1_U8.top_add_9s_9s_9_2_1_Adder_6_U.a  = \add_9s_9s_9_2_1_U8.din0 ;
assign \add_9s_9s_9_2_1_U8.top_add_9s_9s_9_2_1_Adder_6_U.b  = \add_9s_9s_9_2_1_U8.din1 ;
assign \add_9s_9s_9_2_1_U8.top_add_9s_9s_9_2_1_Adder_6_U.ce  = \add_9s_9s_9_2_1_U8.ce ;
assign \add_9s_9s_9_2_1_U8.top_add_9s_9s_9_2_1_Adder_6_U.clk  = \add_9s_9s_9_2_1_U8.clk ;
assign \add_9s_9s_9_2_1_U8.top_add_9s_9s_9_2_1_Adder_6_U.reset  = \add_9s_9s_9_2_1_U8.reset ;
assign \add_9s_9s_9_2_1_U8.dout  = \add_9s_9s_9_2_1_U8.top_add_9s_9s_9_2_1_Adder_6_U.s ;
assign \add_9s_9s_9_2_1_U8.ce  = 1'h1;
assign \add_9s_9s_9_2_1_U8.clk  = ap_clk;
assign \add_9s_9s_9_2_1_U8.din0  = { op_3[3], op_3[3], op_3[3], op_3, 2'h0 };
assign \add_9s_9s_9_2_1_U8.din1  = { op_6[7], op_6 };
assign grp_fu_809_p2 = \add_9s_9s_9_2_1_U8.dout ;
assign \add_9s_9s_9_2_1_U8.reset  = ap_rst;
assign \add_9s_9ns_9_2_1_U5.top_add_9s_9ns_9_2_1_Adder_3_U.ain_s0  = \add_9s_9ns_9_2_1_U5.top_add_9s_9ns_9_2_1_Adder_3_U.a ;
assign \add_9s_9ns_9_2_1_U5.top_add_9s_9ns_9_2_1_Adder_3_U.bin_s0  = \add_9s_9ns_9_2_1_U5.top_add_9s_9ns_9_2_1_Adder_3_U.b ;
assign \add_9s_9ns_9_2_1_U5.top_add_9s_9ns_9_2_1_Adder_3_U.s  = { \add_9s_9ns_9_2_1_U5.top_add_9s_9ns_9_2_1_Adder_3_U.fas_s2 , \add_9s_9ns_9_2_1_U5.top_add_9s_9ns_9_2_1_Adder_3_U.sum_s1  };
assign \add_9s_9ns_9_2_1_U5.top_add_9s_9ns_9_2_1_Adder_3_U.u2.a  = \add_9s_9ns_9_2_1_U5.top_add_9s_9ns_9_2_1_Adder_3_U.ain_s1 ;
assign \add_9s_9ns_9_2_1_U5.top_add_9s_9ns_9_2_1_Adder_3_U.u2.b  = \add_9s_9ns_9_2_1_U5.top_add_9s_9ns_9_2_1_Adder_3_U.bin_s1 ;
assign \add_9s_9ns_9_2_1_U5.top_add_9s_9ns_9_2_1_Adder_3_U.u2.cin  = \add_9s_9ns_9_2_1_U5.top_add_9s_9ns_9_2_1_Adder_3_U.carry_s1 ;
assign \add_9s_9ns_9_2_1_U5.top_add_9s_9ns_9_2_1_Adder_3_U.facout_s2  = \add_9s_9ns_9_2_1_U5.top_add_9s_9ns_9_2_1_Adder_3_U.u2.cout ;
assign \add_9s_9ns_9_2_1_U5.top_add_9s_9ns_9_2_1_Adder_3_U.fas_s2  = \add_9s_9ns_9_2_1_U5.top_add_9s_9ns_9_2_1_Adder_3_U.u2.s ;
assign \add_9s_9ns_9_2_1_U5.top_add_9s_9ns_9_2_1_Adder_3_U.u1.a  = \add_9s_9ns_9_2_1_U5.top_add_9s_9ns_9_2_1_Adder_3_U.a [3:0];
assign \add_9s_9ns_9_2_1_U5.top_add_9s_9ns_9_2_1_Adder_3_U.u1.b  = \add_9s_9ns_9_2_1_U5.top_add_9s_9ns_9_2_1_Adder_3_U.b [3:0];
assign \add_9s_9ns_9_2_1_U5.top_add_9s_9ns_9_2_1_Adder_3_U.u1.cin  = 1'h0;
assign \add_9s_9ns_9_2_1_U5.top_add_9s_9ns_9_2_1_Adder_3_U.facout_s1  = \add_9s_9ns_9_2_1_U5.top_add_9s_9ns_9_2_1_Adder_3_U.u1.cout ;
assign \add_9s_9ns_9_2_1_U5.top_add_9s_9ns_9_2_1_Adder_3_U.fas_s1  = \add_9s_9ns_9_2_1_U5.top_add_9s_9ns_9_2_1_Adder_3_U.u1.s ;
assign \add_9s_9ns_9_2_1_U5.top_add_9s_9ns_9_2_1_Adder_3_U.a  = \add_9s_9ns_9_2_1_U5.din0 ;
assign \add_9s_9ns_9_2_1_U5.top_add_9s_9ns_9_2_1_Adder_3_U.b  = \add_9s_9ns_9_2_1_U5.din1 ;
assign \add_9s_9ns_9_2_1_U5.top_add_9s_9ns_9_2_1_Adder_3_U.ce  = \add_9s_9ns_9_2_1_U5.ce ;
assign \add_9s_9ns_9_2_1_U5.top_add_9s_9ns_9_2_1_Adder_3_U.clk  = \add_9s_9ns_9_2_1_U5.clk ;
assign \add_9s_9ns_9_2_1_U5.top_add_9s_9ns_9_2_1_Adder_3_U.reset  = \add_9s_9ns_9_2_1_U5.reset ;
assign \add_9s_9ns_9_2_1_U5.dout  = \add_9s_9ns_9_2_1_U5.top_add_9s_9ns_9_2_1_Adder_3_U.s ;
assign \add_9s_9ns_9_2_1_U5.ce  = 1'h1;
assign \add_9s_9ns_9_2_1_U5.clk  = ap_clk;
assign \add_9s_9ns_9_2_1_U5.din0  = { op_8_V_reg_1521[7], op_8_V_reg_1521 };
assign \add_9s_9ns_9_2_1_U5.din1  = 9'h008;
assign grp_fu_517_p2 = \add_9s_9ns_9_2_1_U5.dout ;
assign \add_9s_9ns_9_2_1_U5.reset  = ap_rst;
assign \add_8s_8s_8_2_1_U10.top_add_8s_8s_8_2_1_Adder_7_U.ain_s0  = \add_8s_8s_8_2_1_U10.top_add_8s_8s_8_2_1_Adder_7_U.a ;
assign \add_8s_8s_8_2_1_U10.top_add_8s_8s_8_2_1_Adder_7_U.bin_s0  = \add_8s_8s_8_2_1_U10.top_add_8s_8s_8_2_1_Adder_7_U.b ;
assign \add_8s_8s_8_2_1_U10.top_add_8s_8s_8_2_1_Adder_7_U.s  = { \add_8s_8s_8_2_1_U10.top_add_8s_8s_8_2_1_Adder_7_U.fas_s2 , \add_8s_8s_8_2_1_U10.top_add_8s_8s_8_2_1_Adder_7_U.sum_s1  };
assign \add_8s_8s_8_2_1_U10.top_add_8s_8s_8_2_1_Adder_7_U.u2.a  = \add_8s_8s_8_2_1_U10.top_add_8s_8s_8_2_1_Adder_7_U.ain_s1 ;
assign \add_8s_8s_8_2_1_U10.top_add_8s_8s_8_2_1_Adder_7_U.u2.b  = \add_8s_8s_8_2_1_U10.top_add_8s_8s_8_2_1_Adder_7_U.bin_s1 ;
assign \add_8s_8s_8_2_1_U10.top_add_8s_8s_8_2_1_Adder_7_U.u2.cin  = \add_8s_8s_8_2_1_U10.top_add_8s_8s_8_2_1_Adder_7_U.carry_s1 ;
assign \add_8s_8s_8_2_1_U10.top_add_8s_8s_8_2_1_Adder_7_U.facout_s2  = \add_8s_8s_8_2_1_U10.top_add_8s_8s_8_2_1_Adder_7_U.u2.cout ;
assign \add_8s_8s_8_2_1_U10.top_add_8s_8s_8_2_1_Adder_7_U.fas_s2  = \add_8s_8s_8_2_1_U10.top_add_8s_8s_8_2_1_Adder_7_U.u2.s ;
assign \add_8s_8s_8_2_1_U10.top_add_8s_8s_8_2_1_Adder_7_U.u1.a  = \add_8s_8s_8_2_1_U10.top_add_8s_8s_8_2_1_Adder_7_U.a [3:0];
assign \add_8s_8s_8_2_1_U10.top_add_8s_8s_8_2_1_Adder_7_U.u1.b  = \add_8s_8s_8_2_1_U10.top_add_8s_8s_8_2_1_Adder_7_U.b [3:0];
assign \add_8s_8s_8_2_1_U10.top_add_8s_8s_8_2_1_Adder_7_U.u1.cin  = 1'h0;
assign \add_8s_8s_8_2_1_U10.top_add_8s_8s_8_2_1_Adder_7_U.facout_s1  = \add_8s_8s_8_2_1_U10.top_add_8s_8s_8_2_1_Adder_7_U.u1.cout ;
assign \add_8s_8s_8_2_1_U10.top_add_8s_8s_8_2_1_Adder_7_U.fas_s1  = \add_8s_8s_8_2_1_U10.top_add_8s_8s_8_2_1_Adder_7_U.u1.s ;
assign \add_8s_8s_8_2_1_U10.top_add_8s_8s_8_2_1_Adder_7_U.a  = \add_8s_8s_8_2_1_U10.din0 ;
assign \add_8s_8s_8_2_1_U10.top_add_8s_8s_8_2_1_Adder_7_U.b  = \add_8s_8s_8_2_1_U10.din1 ;
assign \add_8s_8s_8_2_1_U10.top_add_8s_8s_8_2_1_Adder_7_U.ce  = \add_8s_8s_8_2_1_U10.ce ;
assign \add_8s_8s_8_2_1_U10.top_add_8s_8s_8_2_1_Adder_7_U.clk  = \add_8s_8s_8_2_1_U10.clk ;
assign \add_8s_8s_8_2_1_U10.top_add_8s_8s_8_2_1_Adder_7_U.reset  = \add_8s_8s_8_2_1_U10.reset ;
assign \add_8s_8s_8_2_1_U10.dout  = \add_8s_8s_8_2_1_U10.top_add_8s_8s_8_2_1_Adder_7_U.s ;
assign \add_8s_8s_8_2_1_U10.ce  = 1'h1;
assign \add_8s_8s_8_2_1_U10.clk  = ap_clk;
assign \add_8s_8s_8_2_1_U10.din0  = { select_ln850_4_reg_1649[5], select_ln850_4_reg_1649, 1'h0 };
assign \add_8s_8s_8_2_1_U10.din1  = { op_9_V_reg_1722[3], op_9_V_reg_1722[3], op_9_V_reg_1722[3], op_9_V_reg_1722[3], op_9_V_reg_1722 };
assign grp_fu_868_p2 = \add_8s_8s_8_2_1_U10.dout ;
assign \add_8s_8s_8_2_1_U10.reset  = ap_rst;
assign \add_8s_8ns_8_2_1_U11.top_add_8s_8ns_8_2_1_Adder_8_U.ain_s0  = \add_8s_8ns_8_2_1_U11.top_add_8s_8ns_8_2_1_Adder_8_U.a ;
assign \add_8s_8ns_8_2_1_U11.top_add_8s_8ns_8_2_1_Adder_8_U.bin_s0  = \add_8s_8ns_8_2_1_U11.top_add_8s_8ns_8_2_1_Adder_8_U.b ;
assign \add_8s_8ns_8_2_1_U11.top_add_8s_8ns_8_2_1_Adder_8_U.s  = { \add_8s_8ns_8_2_1_U11.top_add_8s_8ns_8_2_1_Adder_8_U.fas_s2 , \add_8s_8ns_8_2_1_U11.top_add_8s_8ns_8_2_1_Adder_8_U.sum_s1  };
assign \add_8s_8ns_8_2_1_U11.top_add_8s_8ns_8_2_1_Adder_8_U.u2.a  = \add_8s_8ns_8_2_1_U11.top_add_8s_8ns_8_2_1_Adder_8_U.ain_s1 ;
assign \add_8s_8ns_8_2_1_U11.top_add_8s_8ns_8_2_1_Adder_8_U.u2.b  = \add_8s_8ns_8_2_1_U11.top_add_8s_8ns_8_2_1_Adder_8_U.bin_s1 ;
assign \add_8s_8ns_8_2_1_U11.top_add_8s_8ns_8_2_1_Adder_8_U.u2.cin  = \add_8s_8ns_8_2_1_U11.top_add_8s_8ns_8_2_1_Adder_8_U.carry_s1 ;
assign \add_8s_8ns_8_2_1_U11.top_add_8s_8ns_8_2_1_Adder_8_U.facout_s2  = \add_8s_8ns_8_2_1_U11.top_add_8s_8ns_8_2_1_Adder_8_U.u2.cout ;
assign \add_8s_8ns_8_2_1_U11.top_add_8s_8ns_8_2_1_Adder_8_U.fas_s2  = \add_8s_8ns_8_2_1_U11.top_add_8s_8ns_8_2_1_Adder_8_U.u2.s ;
assign \add_8s_8ns_8_2_1_U11.top_add_8s_8ns_8_2_1_Adder_8_U.u1.a  = \add_8s_8ns_8_2_1_U11.top_add_8s_8ns_8_2_1_Adder_8_U.a [3:0];
assign \add_8s_8ns_8_2_1_U11.top_add_8s_8ns_8_2_1_Adder_8_U.u1.b  = \add_8s_8ns_8_2_1_U11.top_add_8s_8ns_8_2_1_Adder_8_U.b [3:0];
assign \add_8s_8ns_8_2_1_U11.top_add_8s_8ns_8_2_1_Adder_8_U.u1.cin  = 1'h0;
assign \add_8s_8ns_8_2_1_U11.top_add_8s_8ns_8_2_1_Adder_8_U.facout_s1  = \add_8s_8ns_8_2_1_U11.top_add_8s_8ns_8_2_1_Adder_8_U.u1.cout ;
assign \add_8s_8ns_8_2_1_U11.top_add_8s_8ns_8_2_1_Adder_8_U.fas_s1  = \add_8s_8ns_8_2_1_U11.top_add_8s_8ns_8_2_1_Adder_8_U.u1.s ;
assign \add_8s_8ns_8_2_1_U11.top_add_8s_8ns_8_2_1_Adder_8_U.a  = \add_8s_8ns_8_2_1_U11.din0 ;
assign \add_8s_8ns_8_2_1_U11.top_add_8s_8ns_8_2_1_Adder_8_U.b  = \add_8s_8ns_8_2_1_U11.din1 ;
assign \add_8s_8ns_8_2_1_U11.top_add_8s_8ns_8_2_1_Adder_8_U.ce  = \add_8s_8ns_8_2_1_U11.ce ;
assign \add_8s_8ns_8_2_1_U11.top_add_8s_8ns_8_2_1_Adder_8_U.clk  = \add_8s_8ns_8_2_1_U11.clk ;
assign \add_8s_8ns_8_2_1_U11.top_add_8s_8ns_8_2_1_Adder_8_U.reset  = \add_8s_8ns_8_2_1_U11.reset ;
assign \add_8s_8ns_8_2_1_U11.dout  = \add_8s_8ns_8_2_1_U11.top_add_8s_8ns_8_2_1_Adder_8_U.s ;
assign \add_8s_8ns_8_2_1_U11.ce  = 1'h1;
assign \add_8s_8ns_8_2_1_U11.clk  = ap_clk;
assign \add_8s_8ns_8_2_1_U11.din0  = { tmp_3_reg_1763[6], tmp_3_reg_1763 };
assign \add_8s_8ns_8_2_1_U11.din1  = 8'h01;
assign grp_fu_896_p2 = \add_8s_8ns_8_2_1_U11.dout ;
assign \add_8s_8ns_8_2_1_U11.reset  = ap_rst;
assign \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.ain_s0  = \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.a ;
assign \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.bin_s0  = \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.b ;
assign \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.s  = { \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.fas_s2 , \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.sum_s1  };
assign \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.u2.a  = \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.ain_s1 ;
assign \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.u2.b  = \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.bin_s1 ;
assign \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.u2.cin  = \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.carry_s1 ;
assign \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.facout_s2  = \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.u2.cout ;
assign \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.fas_s2  = \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.u2.s ;
assign \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.u1.a  = \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.a [2:0];
assign \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.u1.b  = \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.b [2:0];
assign \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.u1.cin  = 1'h0;
assign \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.facout_s1  = \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.u1.cout ;
assign \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.fas_s1  = \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.u1.s ;
assign \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.a  = \add_6s_6ns_6_2_1_U12.din0 ;
assign \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.b  = \add_6s_6ns_6_2_1_U12.din1 ;
assign \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.ce  = \add_6s_6ns_6_2_1_U12.ce ;
assign \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.clk  = \add_6s_6ns_6_2_1_U12.clk ;
assign \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.reset  = \add_6s_6ns_6_2_1_U12.reset ;
assign \add_6s_6ns_6_2_1_U12.dout  = \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.s ;
assign \add_6s_6ns_6_2_1_U12.ce  = 1'h1;
assign \add_6s_6ns_6_2_1_U12.clk  = ap_clk;
assign \add_6s_6ns_6_2_1_U12.din0  = { trunc_ln2_reg_1728[4], trunc_ln2_reg_1728 };
assign \add_6s_6ns_6_2_1_U12.din1  = { 5'h00, and_ln408_reg_1768 };
assign grp_fu_908_p2 = \add_6s_6ns_6_2_1_U12.dout ;
assign \add_6s_6ns_6_2_1_U12.reset  = ap_rst;
assign \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_5_U.ain_s0  = \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_5_U.a ;
assign \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_5_U.bin_s0  = \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_5_U.b ;
assign \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_5_U.s  = { \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_5_U.fas_s2 , \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_5_U.sum_s1  };
assign \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_5_U.u2.a  = \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_5_U.ain_s1 ;
assign \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_5_U.u2.b  = \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_5_U.bin_s1 ;
assign \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_5_U.u2.cin  = \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_5_U.carry_s1 ;
assign \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_5_U.facout_s2  = \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_5_U.u2.cout ;
assign \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_5_U.fas_s2  = \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_5_U.u2.s ;
assign \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_5_U.u1.a  = \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_5_U.a [2:0];
assign \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_5_U.u1.b  = \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_5_U.b [2:0];
assign \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_5_U.u1.cin  = 1'h0;
assign \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_5_U.facout_s1  = \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_5_U.u1.cout ;
assign \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_5_U.fas_s1  = \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_5_U.u1.s ;
assign \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_5_U.a  = \add_6ns_6ns_6_2_1_U7.din0 ;
assign \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_5_U.b  = \add_6ns_6ns_6_2_1_U7.din1 ;
assign \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_5_U.ce  = \add_6ns_6ns_6_2_1_U7.ce ;
assign \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_5_U.clk  = \add_6ns_6ns_6_2_1_U7.clk ;
assign \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_5_U.reset  = \add_6ns_6ns_6_2_1_U7.reset ;
assign \add_6ns_6ns_6_2_1_U7.dout  = \add_6ns_6ns_6_2_1_U7.top_add_6ns_6ns_6_2_1_Adder_5_U.s ;
assign \add_6ns_6ns_6_2_1_U7.ce  = 1'h1;
assign \add_6ns_6ns_6_2_1_U7.clk  = ap_clk;
assign \add_6ns_6ns_6_2_1_U7.din0  = ret_V_7_reg_1600;
assign \add_6ns_6ns_6_2_1_U7.din1  = 6'h01;
assign grp_fu_586_p2 = \add_6ns_6ns_6_2_1_U7.dout ;
assign \add_6ns_6ns_6_2_1_U7.reset  = ap_rst;
assign \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.ain_s0  = \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.a ;
assign \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.bin_s0  = \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.b ;
assign \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.s  = { \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.fas_s2 , \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.sum_s1  };
assign \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.u2.a  = \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.ain_s1 ;
assign \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.u2.b  = \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.bin_s1 ;
assign \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.u2.cin  = \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.carry_s1 ;
assign \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.facout_s2  = \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.u2.cout ;
assign \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.fas_s2  = \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.u2.s ;
assign \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.u1.a  = \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.a [1:0];
assign \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.u1.b  = \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.b [1:0];
assign \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.u1.cin  = 1'h0;
assign \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.facout_s1  = \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.u1.cout ;
assign \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.fas_s1  = \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.u1.s ;
assign \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.a  = \add_5ns_5s_5_2_1_U1.din0 ;
assign \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.b  = \add_5ns_5s_5_2_1_U1.din1 ;
assign \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.ce  = \add_5ns_5s_5_2_1_U1.ce ;
assign \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.clk  = \add_5ns_5s_5_2_1_U1.clk ;
assign \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.reset  = \add_5ns_5s_5_2_1_U1.reset ;
assign \add_5ns_5s_5_2_1_U1.dout  = \add_5ns_5s_5_2_1_U1.top_add_5ns_5s_5_2_1_Adder_0_U.s ;
assign \add_5ns_5s_5_2_1_U1.ce  = 1'h1;
assign \add_5ns_5s_5_2_1_U1.clk  = ap_clk;
assign \add_5ns_5s_5_2_1_U1.din0  = select_ln703_reg_1402;
assign \add_5ns_5s_5_2_1_U1.din1  = { op_3[3], op_3 };
assign grp_fu_265_p2 = \add_5ns_5s_5_2_1_U1.dout ;
assign \add_5ns_5s_5_2_1_U1.reset  = ap_rst;
assign \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.ain_s0  = \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.a ;
assign \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.bin_s0  = \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.b ;
assign \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.s  = { \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.fas_s2 , \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.sum_s1  };
assign \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.u2.a  = \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.ain_s1 ;
assign \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.u2.b  = \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.bin_s1 ;
assign \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.u2.cin  = \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.carry_s1 ;
assign \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.facout_s2  = \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.u2.cout ;
assign \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.fas_s2  = \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.u2.s ;
assign \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.u1.a  = \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.a [1:0];
assign \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.u1.b  = \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.b [1:0];
assign \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.u1.cin  = 1'h0;
assign \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.facout_s1  = \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.u1.cout ;
assign \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.fas_s1  = \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.u1.s ;
assign \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.a  = \add_4ns_4ns_4_2_1_U9.din0 ;
assign \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.b  = \add_4ns_4ns_4_2_1_U9.din1 ;
assign \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.ce  = \add_4ns_4ns_4_2_1_U9.ce ;
assign \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.clk  = \add_4ns_4ns_4_2_1_U9.clk ;
assign \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.reset  = \add_4ns_4ns_4_2_1_U9.reset ;
assign \add_4ns_4ns_4_2_1_U9.dout  = \add_4ns_4ns_4_2_1_U9.top_add_4ns_4ns_4_2_1_Adder_4_U.s ;
assign \add_4ns_4ns_4_2_1_U9.ce  = 1'h1;
assign \add_4ns_4ns_4_2_1_U9.clk  = ap_clk;
assign \add_4ns_4ns_4_2_1_U9.din0  = { op_3[1:0], 2'h0 };
assign \add_4ns_4ns_4_2_1_U9.din1  = op_6[3:0];
assign grp_fu_815_p2 = \add_4ns_4ns_4_2_1_U9.dout ;
assign \add_4ns_4ns_4_2_1_U9.reset  = ap_rst;
assign \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.ain_s0  = \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.a ;
assign \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.bin_s0  = \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.b ;
assign \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.s  = { \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.fas_s2 , \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.sum_s1  };
assign \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.u2.a  = \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.ain_s1 ;
assign \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.u2.b  = \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.bin_s1 ;
assign \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.u2.cin  = \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.carry_s1 ;
assign \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.facout_s2  = \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.u2.cout ;
assign \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.fas_s2  = \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.u2.s ;
assign \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.u1.a  = \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.a [1:0];
assign \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.u1.b  = \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.b [1:0];
assign \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.u1.cin  = 1'h0;
assign \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.facout_s1  = \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.u1.cout ;
assign \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.fas_s1  = \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.u1.s ;
assign \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.a  = \add_4ns_4ns_4_2_1_U6.din0 ;
assign \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.b  = \add_4ns_4ns_4_2_1_U6.din1 ;
assign \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.ce  = \add_4ns_4ns_4_2_1_U6.ce ;
assign \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.clk  = \add_4ns_4ns_4_2_1_U6.clk ;
assign \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.reset  = \add_4ns_4ns_4_2_1_U6.reset ;
assign \add_4ns_4ns_4_2_1_U6.dout  = \add_4ns_4ns_4_2_1_U6.top_add_4ns_4ns_4_2_1_Adder_4_U.s ;
assign \add_4ns_4ns_4_2_1_U6.ce  = 1'h1;
assign \add_4ns_4ns_4_2_1_U6.clk  = ap_clk;
assign \add_4ns_4ns_4_2_1_U6.din0  = p_Val2_6_reg_1541;
assign \add_4ns_4ns_4_2_1_U6.din1  = { 3'h0, and_ln406_reg_1573 };
assign grp_fu_576_p2 = \add_4ns_4ns_4_2_1_U6.dout ;
assign \add_4ns_4ns_4_2_1_U6.reset  = ap_rst;
assign \add_35s_35s_35_2_1_U23.top_add_35s_35s_35_2_1_Adder_12_U.ain_s0  = \add_35s_35s_35_2_1_U23.top_add_35s_35s_35_2_1_Adder_12_U.a ;
assign \add_35s_35s_35_2_1_U23.top_add_35s_35s_35_2_1_Adder_12_U.bin_s0  = \add_35s_35s_35_2_1_U23.top_add_35s_35s_35_2_1_Adder_12_U.b ;
assign \add_35s_35s_35_2_1_U23.top_add_35s_35s_35_2_1_Adder_12_U.s  = { \add_35s_35s_35_2_1_U23.top_add_35s_35s_35_2_1_Adder_12_U.fas_s2 , \add_35s_35s_35_2_1_U23.top_add_35s_35s_35_2_1_Adder_12_U.sum_s1  };
assign \add_35s_35s_35_2_1_U23.top_add_35s_35s_35_2_1_Adder_12_U.u2.a  = \add_35s_35s_35_2_1_U23.top_add_35s_35s_35_2_1_Adder_12_U.ain_s1 ;
assign \add_35s_35s_35_2_1_U23.top_add_35s_35s_35_2_1_Adder_12_U.u2.b  = \add_35s_35s_35_2_1_U23.top_add_35s_35s_35_2_1_Adder_12_U.bin_s1 ;
assign \add_35s_35s_35_2_1_U23.top_add_35s_35s_35_2_1_Adder_12_U.u2.cin  = \add_35s_35s_35_2_1_U23.top_add_35s_35s_35_2_1_Adder_12_U.carry_s1 ;
assign \add_35s_35s_35_2_1_U23.top_add_35s_35s_35_2_1_Adder_12_U.facout_s2  = \add_35s_35s_35_2_1_U23.top_add_35s_35s_35_2_1_Adder_12_U.u2.cout ;
assign \add_35s_35s_35_2_1_U23.top_add_35s_35s_35_2_1_Adder_12_U.fas_s2  = \add_35s_35s_35_2_1_U23.top_add_35s_35s_35_2_1_Adder_12_U.u2.s ;
assign \add_35s_35s_35_2_1_U23.top_add_35s_35s_35_2_1_Adder_12_U.u1.a  = \add_35s_35s_35_2_1_U23.top_add_35s_35s_35_2_1_Adder_12_U.a [16:0];
assign \add_35s_35s_35_2_1_U23.top_add_35s_35s_35_2_1_Adder_12_U.u1.b  = \add_35s_35s_35_2_1_U23.top_add_35s_35s_35_2_1_Adder_12_U.b [16:0];
assign \add_35s_35s_35_2_1_U23.top_add_35s_35s_35_2_1_Adder_12_U.u1.cin  = 1'h0;
assign \add_35s_35s_35_2_1_U23.top_add_35s_35s_35_2_1_Adder_12_U.facout_s1  = \add_35s_35s_35_2_1_U23.top_add_35s_35s_35_2_1_Adder_12_U.u1.cout ;
assign \add_35s_35s_35_2_1_U23.top_add_35s_35s_35_2_1_Adder_12_U.fas_s1  = \add_35s_35s_35_2_1_U23.top_add_35s_35s_35_2_1_Adder_12_U.u1.s ;
assign \add_35s_35s_35_2_1_U23.top_add_35s_35s_35_2_1_Adder_12_U.a  = \add_35s_35s_35_2_1_U23.din0 ;
assign \add_35s_35s_35_2_1_U23.top_add_35s_35s_35_2_1_Adder_12_U.b  = \add_35s_35s_35_2_1_U23.din1 ;
assign \add_35s_35s_35_2_1_U23.top_add_35s_35s_35_2_1_Adder_12_U.ce  = \add_35s_35s_35_2_1_U23.ce ;
assign \add_35s_35s_35_2_1_U23.top_add_35s_35s_35_2_1_Adder_12_U.clk  = \add_35s_35s_35_2_1_U23.clk ;
assign \add_35s_35s_35_2_1_U23.top_add_35s_35s_35_2_1_Adder_12_U.reset  = \add_35s_35s_35_2_1_U23.reset ;
assign \add_35s_35s_35_2_1_U23.dout  = \add_35s_35s_35_2_1_U23.top_add_35s_35s_35_2_1_Adder_12_U.s ;
assign \add_35s_35s_35_2_1_U23.ce  = 1'h1;
assign \add_35s_35s_35_2_1_U23.clk  = ap_clk;
assign \add_35s_35s_35_2_1_U23.din0  = { op_28_V_reg_1995[31], op_28_V_reg_1995, 2'h0 };
assign \add_35s_35s_35_2_1_U23.din1  = { op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18 };
assign grp_fu_1337_p2 = \add_35s_35s_35_2_1_U23.dout ;
assign \add_35s_35s_35_2_1_U23.reset  = ap_rst;
assign \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_10_U.ain_s0  = \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_10_U.a ;
assign \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_10_U.bin_s0  = \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_10_U.b ;
assign \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_10_U.s  = { \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_10_U.fas_s2 , \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_10_U.sum_s1  };
assign \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_10_U.u2.a  = \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_10_U.ain_s1 ;
assign \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_10_U.u2.b  = \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_10_U.bin_s1 ;
assign \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_10_U.u2.cin  = \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_10_U.carry_s1 ;
assign \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_10_U.facout_s2  = \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_10_U.u2.cout ;
assign \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_10_U.fas_s2  = \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_10_U.u2.s ;
assign \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_10_U.u1.a  = \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_10_U.a [16:0];
assign \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_10_U.u1.b  = \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_10_U.b [16:0];
assign \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_10_U.u1.cin  = 1'h0;
assign \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_10_U.facout_s1  = \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_10_U.u1.cout ;
assign \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_10_U.fas_s1  = \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_10_U.u1.s ;
assign \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_10_U.a  = \add_34s_34s_34_2_1_U20.din0 ;
assign \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_10_U.b  = \add_34s_34s_34_2_1_U20.din1 ;
assign \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_10_U.ce  = \add_34s_34s_34_2_1_U20.ce ;
assign \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_10_U.clk  = \add_34s_34s_34_2_1_U20.clk ;
assign \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_10_U.reset  = \add_34s_34s_34_2_1_U20.reset ;
assign \add_34s_34s_34_2_1_U20.dout  = \add_34s_34s_34_2_1_U20.top_add_34s_34s_34_2_1_Adder_10_U.s ;
assign \add_34s_34s_34_2_1_U20.ce  = 1'h1;
assign \add_34s_34s_34_2_1_U20.clk  = ap_clk;
assign \add_34s_34s_34_2_1_U20.din0  = { select_ln353_2_reg_1943[31], select_ln353_2_reg_1943, 1'h0 };
assign \add_34s_34s_34_2_1_U20.din1  = { op_16[15], op_16[15], op_16[15], op_16[15], op_16[15], op_16[15], op_16[15], op_16[15], op_16[15], op_16[15], op_16[15], op_16[15], op_16[15], op_16[15], op_16[15], op_16[15], op_16[15], op_16[15], op_16 };
assign grp_fu_1265_p2 = \add_34s_34s_34_2_1_U20.dout ;
assign \add_34s_34s_34_2_1_U20.reset  = ap_rst;
assign \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_10_U.ain_s0  = \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_10_U.a ;
assign \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_10_U.bin_s0  = \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_10_U.b ;
assign \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_10_U.s  = { \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_10_U.fas_s2 , \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_10_U.sum_s1  };
assign \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_10_U.u2.a  = \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_10_U.ain_s1 ;
assign \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_10_U.u2.b  = \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_10_U.bin_s1 ;
assign \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_10_U.u2.cin  = \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_10_U.carry_s1 ;
assign \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_10_U.facout_s2  = \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_10_U.u2.cout ;
assign \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_10_U.fas_s2  = \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_10_U.u2.s ;
assign \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_10_U.u1.a  = \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_10_U.a [16:0];
assign \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_10_U.u1.b  = \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_10_U.b [16:0];
assign \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_10_U.u1.cin  = 1'h0;
assign \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_10_U.facout_s1  = \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_10_U.u1.cout ;
assign \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_10_U.fas_s1  = \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_10_U.u1.s ;
assign \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_10_U.a  = \add_34s_34s_34_2_1_U18.din0 ;
assign \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_10_U.b  = \add_34s_34s_34_2_1_U18.din1 ;
assign \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_10_U.ce  = \add_34s_34s_34_2_1_U18.ce ;
assign \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_10_U.clk  = \add_34s_34s_34_2_1_U18.clk ;
assign \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_10_U.reset  = \add_34s_34s_34_2_1_U18.reset ;
assign \add_34s_34s_34_2_1_U18.dout  = \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_10_U.s ;
assign \add_34s_34s_34_2_1_U18.ce  = 1'h1;
assign \add_34s_34s_34_2_1_U18.clk  = ap_clk;
assign \add_34s_34s_34_2_1_U18.din0  = { ret_V_29_reg_1906[31], ret_V_29_reg_1906, 1'h0 };
assign \add_34s_34s_34_2_1_U18.din1  = { op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15 };
assign grp_fu_1206_p2 = \add_34s_34s_34_2_1_U18.dout ;
assign \add_34s_34s_34_2_1_U18.reset  = ap_rst;
assign \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_10_U.ain_s0  = \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_10_U.a ;
assign \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_10_U.bin_s0  = \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_10_U.b ;
assign \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_10_U.s  = { \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_10_U.fas_s2 , \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_10_U.sum_s1  };
assign \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_10_U.u2.a  = \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_10_U.ain_s1 ;
assign \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_10_U.u2.b  = \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_10_U.bin_s1 ;
assign \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_10_U.u2.cin  = \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_10_U.carry_s1 ;
assign \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_10_U.facout_s2  = \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_10_U.u2.cout ;
assign \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_10_U.fas_s2  = \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_10_U.u2.s ;
assign \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_10_U.u1.a  = \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_10_U.a [16:0];
assign \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_10_U.u1.b  = \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_10_U.b [16:0];
assign \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_10_U.u1.cin  = 1'h0;
assign \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_10_U.facout_s1  = \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_10_U.u1.cout ;
assign \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_10_U.fas_s1  = \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_10_U.u1.s ;
assign \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_10_U.a  = \add_34s_34s_34_2_1_U13.din0 ;
assign \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_10_U.b  = \add_34s_34s_34_2_1_U13.din1 ;
assign \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_10_U.ce  = \add_34s_34s_34_2_1_U13.ce ;
assign \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_10_U.clk  = \add_34s_34s_34_2_1_U13.clk ;
assign \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_10_U.reset  = \add_34s_34s_34_2_1_U13.reset ;
assign \add_34s_34s_34_2_1_U13.dout  = \add_34s_34s_34_2_1_U13.top_add_34s_34s_34_2_1_Adder_10_U.s ;
assign \add_34s_34s_34_2_1_U13.ce  = 1'h1;
assign \add_34s_34s_34_2_1_U13.clk  = ap_clk;
assign \add_34s_34s_34_2_1_U13.din0  = { select_ln353_reg_1801[7], select_ln353_reg_1801[7], select_ln353_reg_1801[7], select_ln353_reg_1801[7], select_ln353_reg_1801[7], select_ln353_reg_1801[7], select_ln353_reg_1801[7], select_ln353_reg_1801[7], select_ln353_reg_1801[7], select_ln353_reg_1801[7], select_ln353_reg_1801[7], select_ln353_reg_1801[7], select_ln353_reg_1801[7], select_ln353_reg_1801[7], select_ln353_reg_1801[7], select_ln353_reg_1801[7], select_ln353_reg_1801[7], select_ln353_reg_1801[7], select_ln353_reg_1801[7], select_ln353_reg_1801[7], select_ln353_reg_1801[7], select_ln353_reg_1801[7], select_ln353_reg_1801[7], select_ln353_reg_1801[7], select_ln353_reg_1801[7], select_ln353_reg_1801, 1'h0 };
assign \add_34s_34s_34_2_1_U13.din1  = { op_10_V_reg_1795[5], op_10_V_reg_1795[5], op_10_V_reg_1795[5], op_10_V_reg_1795[5], op_10_V_reg_1795[5], op_10_V_reg_1795[5], op_10_V_reg_1795[5], op_10_V_reg_1795[5], op_10_V_reg_1795[5], op_10_V_reg_1795[5], op_10_V_reg_1795[5], op_10_V_reg_1795[5], op_10_V_reg_1795[5], op_10_V_reg_1795[5], op_10_V_reg_1795[5], op_10_V_reg_1795[5], op_10_V_reg_1795[5], op_10_V_reg_1795[5], op_10_V_reg_1795[5], op_10_V_reg_1795[5], op_10_V_reg_1795[5], op_10_V_reg_1795[5], op_10_V_reg_1795[5], op_10_V_reg_1795[5], op_10_V_reg_1795[5], op_10_V_reg_1795[5], op_10_V_reg_1795[5], op_10_V_reg_1795[5], op_10_V_reg_1795 };
assign grp_fu_951_p2 = \add_34s_34s_34_2_1_U13.dout ;
assign \add_34s_34s_34_2_1_U13.reset  = ap_rst;
assign \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_11_U.ain_s0  = \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_11_U.a ;
assign \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_11_U.bin_s0  = \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_11_U.b ;
assign \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_11_U.s  = { \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_11_U.fas_s2 , \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_11_U.sum_s1  };
assign \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.a  = \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_11_U.ain_s1 ;
assign \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.b  = \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_11_U.bin_s1 ;
assign \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.cin  = \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_11_U.carry_s1 ;
assign \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_11_U.facout_s2  = \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.cout ;
assign \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_11_U.fas_s2  = \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.s ;
assign \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.a  = \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_11_U.a [15:0];
assign \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.b  = \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_11_U.b [15:0];
assign \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.cin  = 1'h0;
assign \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_11_U.facout_s1  = \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.cout ;
assign \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_11_U.fas_s1  = \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.s ;
assign \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_11_U.a  = \add_32ns_32ns_32_2_1_U25.din0 ;
assign \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_11_U.b  = \add_32ns_32ns_32_2_1_U25.din1 ;
assign \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_11_U.ce  = \add_32ns_32ns_32_2_1_U25.ce ;
assign \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_11_U.clk  = \add_32ns_32ns_32_2_1_U25.clk ;
assign \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_11_U.reset  = \add_32ns_32ns_32_2_1_U25.reset ;
assign \add_32ns_32ns_32_2_1_U25.dout  = \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_11_U.s ;
assign \add_32ns_32ns_32_2_1_U25.ce  = 1'h1;
assign \add_32ns_32ns_32_2_1_U25.clk  = ap_clk;
assign \add_32ns_32ns_32_2_1_U25.din0  = ret_V_34_reg_2032;
assign \add_32ns_32ns_32_2_1_U25.din1  = { 28'h0000000, op_19 };
assign grp_fu_1391_p2 = \add_32ns_32ns_32_2_1_U25.dout ;
assign \add_32ns_32ns_32_2_1_U25.reset  = ap_rst;
assign \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_11_U.ain_s0  = \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_11_U.a ;
assign \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_11_U.bin_s0  = \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_11_U.b ;
assign \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_11_U.s  = { \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_11_U.fas_s2 , \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_11_U.sum_s1  };
assign \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.a  = \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_11_U.ain_s1 ;
assign \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.b  = \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_11_U.bin_s1 ;
assign \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.cin  = \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_11_U.carry_s1 ;
assign \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_11_U.facout_s2  = \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.cout ;
assign \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_11_U.fas_s2  = \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.s ;
assign \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.a  = \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_11_U.a [15:0];
assign \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.b  = \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_11_U.b [15:0];
assign \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.cin  = 1'h0;
assign \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_11_U.facout_s1  = \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.cout ;
assign \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_11_U.fas_s1  = \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.s ;
assign \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_11_U.a  = \add_32ns_32ns_32_2_1_U24.din0 ;
assign \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_11_U.b  = \add_32ns_32ns_32_2_1_U24.din1 ;
assign \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_11_U.ce  = \add_32ns_32ns_32_2_1_U24.ce ;
assign \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_11_U.clk  = \add_32ns_32ns_32_2_1_U24.clk ;
assign \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_11_U.reset  = \add_32ns_32ns_32_2_1_U24.reset ;
assign \add_32ns_32ns_32_2_1_U24.dout  = \add_32ns_32ns_32_2_1_U24.top_add_32ns_32ns_32_2_1_Adder_11_U.s ;
assign \add_32ns_32ns_32_2_1_U24.ce  = 1'h1;
assign \add_32ns_32ns_32_2_1_U24.clk  = ap_clk;
assign \add_32ns_32ns_32_2_1_U24.din0  = ret_V_34_cast_reg_2020;
assign \add_32ns_32ns_32_2_1_U24.din1  = 32'd1;
assign grp_fu_1363_p2 = \add_32ns_32ns_32_2_1_U24.dout ;
assign \add_32ns_32ns_32_2_1_U24.reset  = ap_rst;
assign \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_11_U.ain_s0  = \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_11_U.a ;
assign \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_11_U.bin_s0  = \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_11_U.b ;
assign \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_11_U.s  = { \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_11_U.fas_s2 , \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_11_U.sum_s1  };
assign \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.a  = \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_11_U.ain_s1 ;
assign \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.b  = \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_11_U.bin_s1 ;
assign \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.cin  = \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_11_U.carry_s1 ;
assign \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_11_U.facout_s2  = \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.cout ;
assign \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_11_U.fas_s2  = \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.s ;
assign \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.a  = \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_11_U.a [15:0];
assign \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.b  = \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_11_U.b [15:0];
assign \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.cin  = 1'h0;
assign \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_11_U.facout_s1  = \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.cout ;
assign \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_11_U.fas_s1  = \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.s ;
assign \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_11_U.a  = \add_32ns_32ns_32_2_1_U22.din0 ;
assign \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_11_U.b  = \add_32ns_32ns_32_2_1_U22.din1 ;
assign \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_11_U.ce  = \add_32ns_32ns_32_2_1_U22.ce ;
assign \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_11_U.clk  = \add_32ns_32ns_32_2_1_U22.clk ;
assign \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_11_U.reset  = \add_32ns_32ns_32_2_1_U22.reset ;
assign \add_32ns_32ns_32_2_1_U22.dout  = \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_11_U.s ;
assign \add_32ns_32ns_32_2_1_U22.ce  = 1'h1;
assign \add_32ns_32ns_32_2_1_U22.clk  = ap_clk;
assign \add_32ns_32ns_32_2_1_U22.din0  = ret_V_32_reg_1985;
assign \add_32ns_32ns_32_2_1_U22.din1  = { 31'h00000000, xor_ln1497_reg_1980 };
assign grp_fu_1317_p2 = \add_32ns_32ns_32_2_1_U22.dout ;
assign \add_32ns_32ns_32_2_1_U22.reset  = ap_rst;
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.ain_s0  = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.a ;
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.bin_s0  = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.b ;
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.s  = { \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.fas_s2 , \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.sum_s1  };
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.a  = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.ain_s1 ;
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.b  = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.bin_s1 ;
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.cin  = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.carry_s1 ;
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.facout_s2  = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.cout ;
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.fas_s2  = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.s ;
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.a  = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.a [15:0];
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.b  = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.b [15:0];
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.cin  = 1'h0;
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.facout_s1  = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.cout ;
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.fas_s1  = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.s ;
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.a  = \add_32ns_32ns_32_2_1_U21.din0 ;
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.b  = \add_32ns_32ns_32_2_1_U21.din1 ;
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.ce  = \add_32ns_32ns_32_2_1_U21.ce ;
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.clk  = \add_32ns_32ns_32_2_1_U21.clk ;
assign \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.reset  = \add_32ns_32ns_32_2_1_U21.reset ;
assign \add_32ns_32ns_32_2_1_U21.dout  = \add_32ns_32ns_32_2_1_U21.top_add_32ns_32ns_32_2_1_Adder_11_U.s ;
assign \add_32ns_32ns_32_2_1_U21.ce  = 1'h1;
assign \add_32ns_32ns_32_2_1_U21.clk  = ap_clk;
assign \add_32ns_32ns_32_2_1_U21.din0  = ret_V_32_cast_reg_1968;
assign \add_32ns_32ns_32_2_1_U21.din1  = 32'd1;
assign grp_fu_1281_p2 = \add_32ns_32ns_32_2_1_U21.dout ;
assign \add_32ns_32ns_32_2_1_U21.reset  = ap_rst;
assign \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.ain_s0  = \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.a ;
assign \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.bin_s0  = \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.b ;
assign \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.s  = { \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.fas_s2 , \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.sum_s1  };
assign \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.a  = \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.ain_s1 ;
assign \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.b  = \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.bin_s1 ;
assign \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.cin  = \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.carry_s1 ;
assign \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.facout_s2  = \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.cout ;
assign \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.fas_s2  = \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.s ;
assign \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.a  = \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.a [15:0];
assign \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.b  = \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.b [15:0];
assign \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.cin  = 1'h0;
assign \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.facout_s1  = \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.cout ;
assign \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.fas_s1  = \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.s ;
assign \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.a  = \add_32ns_32ns_32_2_1_U19.din0 ;
assign \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.b  = \add_32ns_32ns_32_2_1_U19.din1 ;
assign \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.ce  = \add_32ns_32ns_32_2_1_U19.ce ;
assign \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.clk  = \add_32ns_32ns_32_2_1_U19.clk ;
assign \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.reset  = \add_32ns_32ns_32_2_1_U19.reset ;
assign \add_32ns_32ns_32_2_1_U19.dout  = \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.s ;
assign \add_32ns_32ns_32_2_1_U19.ce  = 1'h1;
assign \add_32ns_32ns_32_2_1_U19.clk  = ap_clk;
assign \add_32ns_32ns_32_2_1_U19.din0  = ret_V_30_cast_reg_1931;
assign \add_32ns_32ns_32_2_1_U19.din1  = 32'd1;
assign grp_fu_1222_p2 = \add_32ns_32ns_32_2_1_U19.dout ;
assign \add_32ns_32ns_32_2_1_U19.reset  = ap_rst;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.ain_s0  = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.a ;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.bin_s0  = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.b ;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.s  = { \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.fas_s2 , \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.sum_s1  };
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.a  = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.ain_s1 ;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.b  = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.bin_s1 ;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.cin  = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.carry_s1 ;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.facout_s2  = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.cout ;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.fas_s2  = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.s ;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.a  = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.a [15:0];
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.b  = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.b [15:0];
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.cin  = 1'h0;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.facout_s1  = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.cout ;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.fas_s1  = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.s ;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.a  = \add_32ns_32ns_32_2_1_U17.din0 ;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.b  = \add_32ns_32ns_32_2_1_U17.din1 ;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.ce  = \add_32ns_32ns_32_2_1_U17.ce ;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.clk  = \add_32ns_32ns_32_2_1_U17.clk ;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.reset  = \add_32ns_32ns_32_2_1_U17.reset ;
assign \add_32ns_32ns_32_2_1_U17.dout  = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.s ;
assign \add_32ns_32ns_32_2_1_U17.ce  = 1'h1;
assign \add_32ns_32ns_32_2_1_U17.clk  = ap_clk;
assign \add_32ns_32ns_32_2_1_U17.din0  = ret_V_28_reg_1896;
assign \add_32ns_32ns_32_2_1_U17.din1  = select_ln1192_reg_1901;
assign grp_fu_1187_p2 = \add_32ns_32ns_32_2_1_U17.dout ;
assign \add_32ns_32ns_32_2_1_U17.reset  = ap_rst;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.ain_s0  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.a ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.bin_s0  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.b ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.s  = { \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.fas_s2 , \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.sum_s1  };
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.a  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.ain_s1 ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.b  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.bin_s1 ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.cin  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.carry_s1 ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.facout_s2  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.cout ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.fas_s2  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.s ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.a  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.a [15:0];
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.b  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.b [15:0];
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.cin  = 1'h0;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.facout_s1  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.cout ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.fas_s1  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.s ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.a  = \add_32ns_32ns_32_2_1_U16.din0 ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.b  = \add_32ns_32ns_32_2_1_U16.din1 ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.ce  = \add_32ns_32ns_32_2_1_U16.ce ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.clk  = \add_32ns_32ns_32_2_1_U16.clk ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.reset  = \add_32ns_32ns_32_2_1_U16.reset ;
assign \add_32ns_32ns_32_2_1_U16.dout  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.s ;
assign \add_32ns_32ns_32_2_1_U16.ce  = 1'h1;
assign \add_32ns_32ns_32_2_1_U16.clk  = ap_clk;
assign \add_32ns_32ns_32_2_1_U16.din0  = op_23_V_reg_1874;
assign \add_32ns_32ns_32_2_1_U16.din1  = { 31'h00000000, lhs_V_2_reg_1864 };
assign grp_fu_1147_p2 = \add_32ns_32ns_32_2_1_U16.dout ;
assign \add_32ns_32ns_32_2_1_U16.reset  = ap_rst;
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.ain_s0  = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.a ;
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.bin_s0  = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.b ;
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.s  = { \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.fas_s2 , \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.sum_s1  };
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.a  = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.ain_s1 ;
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.b  = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.bin_s1 ;
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.cin  = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.carry_s1 ;
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.facout_s2  = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.cout ;
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.fas_s2  = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.s ;
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.a  = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.a [15:0];
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.b  = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.b [15:0];
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.cin  = 1'h0;
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.facout_s1  = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.cout ;
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.fas_s1  = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.s ;
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.a  = \add_32ns_32ns_32_2_1_U15.din0 ;
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.b  = \add_32ns_32ns_32_2_1_U15.din1 ;
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.ce  = \add_32ns_32ns_32_2_1_U15.ce ;
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.clk  = \add_32ns_32ns_32_2_1_U15.clk ;
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.reset  = \add_32ns_32ns_32_2_1_U15.reset ;
assign \add_32ns_32ns_32_2_1_U15.dout  = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.s ;
assign \add_32ns_32ns_32_2_1_U15.ce  = 1'h1;
assign \add_32ns_32ns_32_2_1_U15.clk  = ap_clk;
assign \add_32ns_32ns_32_2_1_U15.din0  = ret_V_27_reg_1833;
assign \add_32ns_32ns_32_2_1_U15.din1  = select_ln69_reg_1838;
assign grp_fu_1003_p2 = \add_32ns_32ns_32_2_1_U15.dout ;
assign \add_32ns_32ns_32_2_1_U15.reset  = ap_rst;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.ain_s0  = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.a ;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.bin_s0  = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.b ;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.s  = { \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.fas_s2 , \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.sum_s1  };
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.a  = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.ain_s1 ;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.b  = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.bin_s1 ;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.cin  = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.carry_s1 ;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.facout_s2  = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.cout ;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.fas_s2  = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.s ;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.a  = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.a [15:0];
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.b  = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.b [15:0];
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.cin  = 1'h0;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.facout_s1  = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.cout ;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.fas_s1  = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.s ;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.a  = \add_32ns_32ns_32_2_1_U14.din0 ;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.b  = \add_32ns_32ns_32_2_1_U14.din1 ;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.ce  = \add_32ns_32ns_32_2_1_U14.ce ;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.clk  = \add_32ns_32ns_32_2_1_U14.clk ;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.reset  = \add_32ns_32ns_32_2_1_U14.reset ;
assign \add_32ns_32ns_32_2_1_U14.dout  = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_11_U.s ;
assign \add_32ns_32ns_32_2_1_U14.ce  = 1'h1;
assign \add_32ns_32ns_32_2_1_U14.clk  = ap_clk;
assign \add_32ns_32ns_32_2_1_U14.din0  = ret_V_24_cast_reg_1821;
assign \add_32ns_32ns_32_2_1_U14.din1  = 32'd1;
assign grp_fu_967_p2 = \add_32ns_32ns_32_2_1_U14.dout ;
assign \add_32ns_32ns_32_2_1_U14.reset  = ap_rst;
assign \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.ain_s0  = \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.a ;
assign \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.bin_s0  = \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.b ;
assign \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.s  = { \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.fas_s2 , \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.sum_s1  };
assign \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.a  = \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.ain_s1 ;
assign \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.b  = \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.bin_s1 ;
assign \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.cin  = \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.carry_s1 ;
assign \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.facout_s2  = \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.cout ;
assign \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.fas_s2  = \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.s ;
assign \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.a  = \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.a [0];
assign \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.b  = \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.b [0];
assign \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.cin  = 1'h0;
assign \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.facout_s1  = \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.cout ;
assign \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.fas_s1  = \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.s ;
assign \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.a  = \add_2ns_2ns_2_2_1_U2.din0 ;
assign \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.b  = \add_2ns_2ns_2_2_1_U2.din1 ;
assign \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.ce  = \add_2ns_2ns_2_2_1_U2.ce ;
assign \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.clk  = \add_2ns_2ns_2_2_1_U2.clk ;
assign \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.reset  = \add_2ns_2ns_2_2_1_U2.reset ;
assign \add_2ns_2ns_2_2_1_U2.dout  = \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.s ;
assign \add_2ns_2ns_2_2_1_U2.ce  = 1'h1;
assign \add_2ns_2ns_2_2_1_U2.clk  = ap_clk;
assign \add_2ns_2ns_2_2_1_U2.din0  = ret_V_reg_1429;
assign \add_2ns_2ns_2_2_1_U2.din1  = 2'h1;
assign grp_fu_286_p2 = \add_2ns_2ns_2_2_1_U2.dout ;
assign \add_2ns_2ns_2_2_1_U2.reset  = ap_rst;
endmodule


// Machine B:
// Processed by function `add_clk_enable_signal` in `verilog_tricks.py`.
// Processed by function `remove_reset_signal` in `verilog_tricks.py`.
module top_B (
  ap_clk,
  ap_start,
  ap_done,
  ap_idle,
  ap_ready,
  op_0,
  op_2,
  op_3,
  op_5,
  op_6,
  op_7,
  op_12,
  op_15,
  op_16,
  op_18,
  op_19,
  op_30,
  op_30_ap_vld,
clk_enable
);
input clk_enable;


input ap_clk;
wire ap_rst;
assign ap_rst = op_30_ap_vld;
input ap_start;
input op_0;
input op_12;
input [3:0] op_15;
input [15:0] op_16;
input [3:0] op_18;
input [3:0] op_19;
input op_2;
input [3:0] op_3;
input [1:0] op_5;
input [7:0] op_6;
input [3:0] op_7;
output ap_done;
output ap_idle;
output ap_ready;
output [31:0] op_30;
output op_30_ap_vld;


reg [7:0] add_ln691_reg_1611;
reg and_ln785_1_reg_1574;
reg and_ln786_reg_1564;
reg [10:0] ap_CS_fsm = 11'h001;
reg icmp_ln1497_reg_1621;
reg icmp_ln851_2_reg_1687;
reg lhs_V_2_reg_1616;
reg [5:0] op_10_V_reg_1599;
reg [31:0] op_23_V_reg_1626;
reg [31:0] op_28_V_reg_1670;
reg [3:0] op_9_V_reg_1584;
reg or_ln340_reg_1569;
reg or_ln384_reg_1551;
reg overflow_reg_1546;
reg p_Result_25_reg_1511;
reg p_Result_27_reg_1519;
reg p_Result_29_reg_1524;
reg [12:0] p_Result_6_reg_1530;
reg [13:0] p_Result_7_reg_1535;
reg [3:0] p_Val2_7_reg_1556;
reg [19:0] r_V_1_reg_1503;
reg [1:0] ret_V_21_reg_1492;
reg [7:0] ret_V_25_reg_1589;
reg [31:0] ret_V_30_cast_reg_1646;
reg [33:0] ret_V_30_reg_1641;
reg [33:0] ret_V_31_reg_1658;
reg [31:0] ret_V_32_cast_reg_1663;
reg [34:0] ret_V_33_reg_1675;
reg [31:0] ret_V_34_cast_reg_1680;
reg [16:0] ret_reg_1541;
reg sel_tmp11_reg_1579;
reg [31:0] select_ln1192_reg_1631;
reg [15:0] sext_ln1347_reg_1498;
reg [7:0] sext_ln850_reg_1605;
reg [6:0] tmp_3_reg_1594;
wire [7:0] _000_;
wire _001_;
wire _002_;
wire [10:0] _003_;
wire _004_;
wire _005_;
wire _006_;
wire [5:0] _007_;
wire [31:0] _008_;
wire [31:0] _009_;
wire [3:0] _010_;
wire _011_;
wire _012_;
wire _013_;
wire _014_;
wire _015_;
wire _016_;
wire [12:0] _017_;
wire [13:0] _018_;
wire [3:0] _019_;
wire [19:0] _020_;
wire [1:0] _021_;
wire [7:0] _022_;
wire [31:0] _023_;
wire [33:0] _024_;
wire [33:0] _025_;
wire [31:0] _026_;
wire [34:0] _027_;
wire [31:0] _028_;
wire [16:0] _029_;
wire _030_;
wire [31:0] _031_;
wire [15:0] _032_;
wire [7:0] _033_;
wire [6:0] _034_;
wire [1:0] _035_;
wire _036_;
wire _037_;
wire _038_;
wire _039_;
wire _040_;
wire _041_;
wire _042_;
wire _043_;
wire _044_;
wire _045_;
wire _046_;
wire _047_;
wire _048_;
wire _049_;
wire _050_;
wire _051_;
wire _052_;
wire _053_;
wire _054_;
wire _055_;
wire _056_;
wire _057_;
wire _058_;
wire _059_;
wire _060_;
wire _061_;
wire _062_;
wire Range1_all_ones_fu_561_p2;
wire Range1_all_zeros_fu_566_p2;
wire Range2_all_ones_fu_556_p2;
wire [3:0] add_ln1192_1_fu_908_p2;
wire [31:0] add_ln691_1_fu_1209_p2;
wire [31:0] add_ln691_2_fu_1308_p2;
wire [31:0] add_ln691_3_fu_1374_p2;
wire [31:0] add_ln691_4_fu_1451_p2;
wire [7:0] add_ln691_fu_965_p2;
wire and_ln340_fu_706_p2;
wire and_ln406_fu_521_p2;
wire and_ln408_fu_946_p2;
wire and_ln780_fu_584_p2;
wire and_ln781_fu_598_p2;
wire and_ln785_1_fu_688_p2;
wire and_ln785_2_fu_694_p2;
wire and_ln785_fu_677_p2;
wire and_ln786_fu_638_p2;
wire and_ln850_fu_991_p2;
wire ap_CS_fsm_state1;
wire ap_CS_fsm_state10;
wire ap_CS_fsm_state11;
wire ap_CS_fsm_state2;
wire ap_CS_fsm_state3;
wire ap_CS_fsm_state4;
wire ap_CS_fsm_state5;
wire ap_CS_fsm_state6;
wire ap_CS_fsm_state7;
wire ap_CS_fsm_state8;
wire ap_CS_fsm_state9;
wire [10:0] ap_NS_fsm;
wire ap_clk;
wire ap_done;
wire ap_idle;
wire ap_ready;
wire ap_rst;
wire ap_start;
wire carry_2_fu_551_p2;
wire carry_fu_1041_p3;
wire deleted_ones_fu_590_p3;
wire deleted_zeros_fu_571_p3;
wire icmp_ln1497_fu_1138_p2;
wire icmp_ln768_fu_419_p2;
wire icmp_ln786_fu_449_p2;
wire icmp_ln790_fu_467_p2;
wire icmp_ln851_1_fu_818_p2;
wire icmp_ln851_2_fu_1438_p2;
wire icmp_ln851_fu_289_p2;
wire lhs_V_2_fu_1099_p2;
wire [3:0] lhs_fu_878_p1;
wire [5:0] lhs_fu_878_p3;
wire [15:0] \mul_16ns_4s_20_1_1_U1.din0 ;
wire [3:0] \mul_16ns_4s_20_1_1_U1.din1 ;
wire [19:0] \mul_16ns_4s_20_1_1_U1.dout ;
wire [15:0] \mul_16ns_4s_20_1_1_U1.top_mul_16ns_4s_20_1_1_Multiplier_0_U.a ;
wire [3:0] \mul_16ns_4s_20_1_1_U1.top_mul_16ns_4s_20_1_1_Multiplier_0_U.b ;
wire [19:0] \mul_16ns_4s_20_1_1_U1.top_mul_16ns_4s_20_1_1_Multiplier_0_U.p ;
wire neg_src_2_fu_1055_p2;
wire neg_src_fu_610_p2;
wire newsignbit_fu_1049_p2;
wire op_0;
wire [5:0] op_10_V_fu_956_p2;
wire [1:0] op_11_V_fu_1126_p3;
wire op_12;
wire op_14_V_fu_1081_p2;
wire [3:0] op_15;
wire [15:0] op_16;
wire [3:0] op_18;
wire [3:0] op_19;
wire op_2;
wire [31:0] op_23_V_fu_1239_p2;
wire [31:0] op_28_V_fu_1397_p2;
wire [3:0] op_3;
wire [31:0] op_30;
wire op_30_ap_vld;
wire [1:0] op_5;
wire [7:0] op_6;
wire [3:0] op_7;
wire [7:0] op_8_V_fu_742_p3;
wire [3:0] op_9_V_fu_780_p3;
wire or_ln340_1_fu_763_p2;
wire or_ln340_2_fu_712_p2;
wire or_ln340_fu_644_p2;
wire or_ln384_fu_491_p2;
wire or_ln406_fu_516_p2;
wire or_ln785_1_fu_621_p2;
wire or_ln785_2_fu_683_p2;
wire or_ln785_fu_425_p2;
wire or_ln788_1_fu_479_p2;
wire or_ln788_fu_473_p2;
wire overflow_1_fu_632_p2;
wire overflow_fu_437_p2;
wire [3:0] p_Result_14_fu_754_p4;
wire p_Result_15_fu_806_p3;
wire p_Result_16_fu_1144_p3;
wire p_Result_17_fu_1198_p3;
wire p_Result_18_fu_1298_p3;
wire p_Result_19_fu_1364_p3;
wire [1:0] p_Result_1_fu_979_p1;
wire p_Result_1_fu_979_p3;
wire p_Result_20_fu_1444_p3;
wire p_Result_21_fu_1033_p3;
wire p_Result_22_fu_928_p3;
wire p_Result_23_fu_393_p3;
wire p_Result_24_fu_401_p3;
wire p_Result_26_fu_506_p3;
wire p_Result_28_fu_537_p3;
wire [6:0] p_Result_3_fu_459_p3;
wire p_Result_s_fu_281_p3;
wire [7:0] p_Val2_4_fu_727_p3;
wire [3:0] p_Val2_6_fu_497_p4;
wire [3:0] p_Val2_7_fu_531_p2;
wire [2:0] p_Val2_8_fu_749_p2;
wire r_1_fu_513_p1;
wire [15:0] r_V_1_fu_327_p0;
wire [19:0] r_V_1_fu_327_p00;
wire [19:0] r_V_1_fu_327_p2;
wire [1:0] r_V_fu_1021_p2;
wire [1:0] r_V_fu_1021_p3;
wire r_fu_940_p2;
wire [4:0] ret_V_20_fu_265_p2;
wire [1:0] ret_V_21_fu_309_p3;
wire ret_V_22_fu_997_p2;
wire [8:0] ret_V_23_fu_902_p2;
wire [31:0] ret_V_24_cast_fu_1188_p4;
wire [8:0] ret_V_24_fu_790_p2;
wire [7:0] ret_V_25_fu_862_p2;
wire [33:0] ret_V_26_fu_1182_p2;
wire [31:0] ret_V_27_fu_1223_p3;
wire [31:0] ret_V_28_fu_1256_p2;
wire [31:0] ret_V_29_fu_1261_p2;
wire [1:0] ret_V_2_fu_295_p2;
wire [33:0] ret_V_30_fu_1282_p2;
wire [33:0] ret_V_31_fu_1343_p2;
wire [31:0] ret_V_32_fu_1386_p3;
wire [34:0] ret_V_33_fu_1418_p2;
wire [31:0] ret_V_34_fu_1462_p3;
wire [1:0] ret_V_4_fu_971_p1;
wire ret_V_4_fu_971_p3;
wire [5:0] ret_V_7_fu_796_p4;
wire [5:0] ret_V_9_fu_824_p2;
wire [1:0] ret_V_fu_271_p4;
wire [16:0] ret_fu_387_p2;
wire [6:0] rhs_2_fu_850_p3;
wire [32:0] rhs_6_fu_1270_p3;
wire [32:0] rhs_7_fu_1331_p3;
wire [33:0] rhs_9_fu_1407_p3;
wire sel_tmp11_fu_718_p2;
wire [31:0] select_ln1192_fu_1245_p3;
wire [16:0] select_ln1347_fu_377_p3;
wire [3:0] select_ln340_1_fu_767_p3;
wire select_ln340_fu_1067_p3;
wire [31:0] select_ln353_2_fu_1324_p3;
wire [7:0] select_ln353_fu_1163_p3;
wire [7:0] select_ln384_fu_735_p3;
wire [31:0] select_ln69_fu_1231_p3;
wire [4:0] select_ln703_fu_249_p3;
wire [3:0] select_ln785_fu_774_p3;
wire [5:0] select_ln850_2_fu_834_p3;
wire [31:0] select_ln850_3_fu_1215_p3;
wire [5:0] select_ln850_4_fu_842_p3;
wire [31:0] select_ln850_5_fu_1379_p3;
wire [31:0] select_ln850_6_fu_1456_p3;
wire [7:0] select_ln850_7_fu_1157_p3;
wire [31:0] select_ln850_8_fu_1317_p3;
wire [1:0] select_ln850_fu_301_p3;
wire [7:0] sext_ln1192_1_fu_830_p1;
wire [7:0] sext_ln1192_2_fu_858_p1;
wire [33:0] sext_ln1192_3_fu_1178_p1;
wire [33:0] sext_ln1192_4_fu_1278_p1;
wire [33:0] sext_ln1192_5_fu_1339_p1;
wire [34:0] sext_ln1192_6_fu_1414_p1;
wire [8:0] sext_ln1192_fu_885_p1;
wire [1:0] sext_ln1299_1_fu_1007_p0;
wire [17:0] sext_ln1299_1_fu_1007_p1;
wire [1:0] sext_ln1299_2_fu_1011_p0;
wire [5:0] sext_ln1299_2_fu_1011_p1;
wire [1:0] sext_ln1299_fu_1003_p0;
wire [2:0] sext_ln1299_fu_1003_p1;
wire [15:0] sext_ln1347_fu_317_p1;
wire [16:0] sext_ln1499_fu_1112_p1;
wire [7:0] sext_ln703_1_fu_889_p0;
wire [8:0] sext_ln703_1_fu_889_p1;
wire [8:0] sext_ln703_2_fu_786_p1;
wire [33:0] sext_ln703_3_fu_1154_p1;
wire [3:0] sext_ln703_4_fu_1266_p0;
wire [33:0] sext_ln703_4_fu_1266_p1;
wire [15:0] sext_ln703_5_fu_1313_p0;
wire [33:0] sext_ln703_5_fu_1313_p1;
wire [3:0] sext_ln703_6_fu_1403_p0;
wire [34:0] sext_ln703_6_fu_1403_p1;
wire [3:0] sext_ln703_fu_257_p0;
wire [4:0] sext_ln703_fu_257_p1;
wire [5:0] sext_ln713_fu_924_p1;
wire [7:0] sext_ln850_fu_962_p1;
wire [3:0] shl_ln1192_fu_897_p0;
wire [3:0] shl_ln1192_fu_897_p2;
wire [1:0] shl_ln1299_fu_1015_p0;
wire [1:0] shl_ln1299_fu_1015_p2;
wire [4:0] shl_ln1_fu_1087_p3;
wire signbit_3_fu_1120_p2;
wire tmp_1_fu_657_p3;
wire [11:0] tmp_2_fu_409_p4;
wire [2:0] tmp_7_fu_1105_p3;
wire [8:0] tmp_8_fu_1170_p3;
wire tmp_fu_650_p3;
wire [7:0] trunc_ln1192_1_fu_893_p0;
wire [3:0] trunc_ln1192_1_fu_893_p1;
wire [3:0] trunc_ln1192_fu_261_p0;
wire [2:0] trunc_ln1192_fu_261_p1;
wire [4:0] trunc_ln2_fu_914_p4;
wire trunc_ln415_fu_1029_p1;
wire [2:0] trunc_ln718_fu_936_p1;
wire [4:0] trunc_ln731_fu_724_p1;
wire [3:0] trunc_ln790_fu_455_p1;
wire [2:0] trunc_ln851_1_fu_814_p1;
wire trunc_ln851_2_fu_1151_p1;
wire trunc_ln851_3_fu_1206_p1;
wire [3:0] trunc_ln851_4_fu_1305_p0;
wire trunc_ln851_4_fu_1305_p1;
wire [15:0] trunc_ln851_5_fu_1371_p0;
wire trunc_ln851_5_fu_1371_p1;
wire [3:0] trunc_ln851_6_fu_1434_p0;
wire [1:0] trunc_ln851_6_fu_1434_p1;
wire [1:0] trunc_ln851_fu_987_p0;
wire trunc_ln851_fu_987_p1;
wire underflow_fu_485_p2;
wire xor_ln1497_fu_1359_p2;
wire xor_ln340_fu_1075_p2;
wire xor_ln365_1_fu_671_p2;
wire xor_ln365_fu_665_p2;
wire xor_ln416_fu_545_p2;
wire xor_ln780_fu_579_p2;
wire xor_ln781_fu_604_p2;
wire xor_ln785_1_fu_431_p2;
wire xor_ln785_2_fu_615_p2;
wire xor_ln785_3_fu_627_p2;
wire xor_ln785_fu_1061_p2;
wire xor_ln786_1_fu_700_p2;
wire xor_ln786_fu_443_p2;
wire [31:0] zext_ln1192_fu_1253_p1;
wire [16:0] zext_ln1347_fu_384_p1;
wire [2:0] zext_ln1497_fu_1134_p1;
wire [17:0] zext_ln1499_1_fu_1116_p1;
wire [5:0] zext_ln1499_fu_1095_p1;
wire [3:0] zext_ln415_1_fu_527_p1;
wire [5:0] zext_ln415_fu_952_p1;
wire [31:0] zext_ln69_1_fu_1469_p1;
wire [31:0] zext_ln69_fu_1393_p1;


assign add_ln1192_1_fu_908_p2 = { op_3[1:0], 2'h0 } + op_6[3:0];
assign add_ln691_1_fu_1209_p2 = { ret_V_26_fu_1182_p2[33], ret_V_26_fu_1182_p2[33], ret_V_26_fu_1182_p2[33], ret_V_26_fu_1182_p2[33], ret_V_26_fu_1182_p2[33], ret_V_26_fu_1182_p2[33], ret_V_26_fu_1182_p2[33], ret_V_26_fu_1182_p2[33], ret_V_26_fu_1182_p2[33], ret_V_26_fu_1182_p2[33], ret_V_26_fu_1182_p2[33], ret_V_26_fu_1182_p2[33], ret_V_26_fu_1182_p2[33], ret_V_26_fu_1182_p2[33], ret_V_26_fu_1182_p2[33], ret_V_26_fu_1182_p2[33], ret_V_26_fu_1182_p2[33], ret_V_26_fu_1182_p2[33], ret_V_26_fu_1182_p2[33], ret_V_26_fu_1182_p2[33], ret_V_26_fu_1182_p2[33], ret_V_26_fu_1182_p2[33], ret_V_26_fu_1182_p2[33], ret_V_26_fu_1182_p2[33], ret_V_26_fu_1182_p2[8:1] } + 1'h1;
assign add_ln691_2_fu_1308_p2 = ret_V_30_cast_reg_1646 + 1'h1;
assign add_ln691_3_fu_1374_p2 = ret_V_32_cast_reg_1663 + 1'h1;
assign add_ln691_4_fu_1451_p2 = ret_V_34_cast_reg_1680 + 1'h1;
assign add_ln691_fu_965_p2 = $signed(tmp_3_reg_1594) + $signed(2'h1);
assign op_10_V_fu_956_p2 = $signed(ret_V_23_fu_902_p2[8:4]) + $signed({ 1'h0, and_ln408_fu_946_p2 });
assign op_23_V_fu_1239_p2 = ret_V_27_fu_1223_p3 + select_ln69_fu_1231_p3;
assign op_28_V_fu_1397_p2 = ret_V_32_fu_1386_p3 + xor_ln1497_fu_1359_p2;
assign op_30 = ret_V_34_fu_1462_p3 + op_19;
assign p_Val2_7_fu_531_p2 = r_V_1_reg_1503[5:2] + and_ln406_fu_521_p2;
assign ret_V_20_fu_265_p2 = $signed(select_ln703_fu_249_p3) + $signed(op_3);
assign ret_V_23_fu_902_p2 = $signed({ op_3, 2'h0 }) + $signed(op_6);
assign ret_V_24_fu_790_p2 = $signed(op_8_V_fu_742_p3) + $signed(5'h08);
assign ret_V_25_fu_862_p2 = $signed({ select_ln850_4_fu_842_p3, 1'h0 }) + $signed(op_9_V_fu_780_p3);
assign { ret_V_26_fu_1182_p2[33], ret_V_26_fu_1182_p2[8:0] } = $signed({ select_ln353_fu_1163_p3, 1'h0 }) + $signed(op_10_V_reg_1599);
assign ret_V_28_fu_1256_p2 = op_23_V_reg_1626 + lhs_V_2_reg_1616;
assign ret_V_29_fu_1261_p2 = ret_V_28_fu_1256_p2 + select_ln1192_reg_1631;
assign ret_V_2_fu_295_p2 = ret_V_20_fu_265_p2[4:3] + 1'h1;
assign ret_V_30_fu_1282_p2 = $signed({ ret_V_29_fu_1261_p2, 1'h0 }) + $signed(op_15);
assign ret_V_31_fu_1343_p2 = $signed({ select_ln353_2_fu_1324_p3, 1'h0 }) + $signed(op_16);
assign ret_V_33_fu_1418_p2 = $signed({ op_28_V_reg_1670, 2'h0 }) + $signed(op_18);
assign ret_V_9_fu_824_p2 = ret_V_24_fu_790_p2[8:3] + 1'h1;
assign _036_ = ap_CS_fsm[0] & _038_;
assign _037_ = ap_CS_fsm[0] & ap_start;
assign and_ln340_fu_706_p2 = xor_ln786_1_fu_700_p2 & or_ln340_fu_644_p2;
assign and_ln406_fu_521_p2 = r_V_1_reg_1503[1] & or_ln406_fu_516_p2;
assign and_ln408_fu_946_p2 = r_fu_940_p2 & add_ln1192_1_fu_908_p2[3];
assign and_ln780_fu_584_p2 = xor_ln780_fu_579_p2 & Range2_all_ones_fu_556_p2;
assign and_ln781_fu_598_p2 = carry_2_fu_551_p2 & Range1_all_ones_fu_561_p2;
assign and_ln785_1_fu_688_p2 = or_ln785_2_fu_683_p2 & and_ln786_fu_638_p2;
assign and_ln785_2_fu_694_p2 = xor_ln785_3_fu_627_p2 & and_ln786_fu_638_p2;
assign and_ln785_fu_677_p2 = xor_ln416_fu_545_p2 & deleted_zeros_fu_571_p3;
assign and_ln786_fu_638_p2 = p_Val2_7_fu_531_p2[3] & deleted_ones_fu_590_p3;
assign and_ln850_fu_991_p2 = op_5[0] & op_5[1];
assign carry_2_fu_551_p2 = xor_ln416_fu_545_p2 & p_Result_27_reg_1519;
assign neg_src_2_fu_1055_p2 = r_V_fu_1021_p3[1] & newsignbit_fu_1049_p2;
assign neg_src_fu_610_p2 = xor_ln781_fu_604_p2 & p_Result_25_reg_1511;
assign op_14_V_fu_1081_p2 = xor_ln340_fu_1075_p2 & newsignbit_fu_1049_p2;
assign overflow_1_fu_632_p2 = xor_ln785_3_fu_627_p2 & or_ln785_1_fu_621_p2;
assign overflow_fu_437_p2 = xor_ln785_1_fu_431_p2 & or_ln785_fu_425_p2;
assign sel_tmp11_fu_718_p2 = xor_ln365_1_fu_671_p2 & or_ln340_2_fu_712_p2;
assign underflow_fu_485_p2 = ret_fu_387_p2[16] & or_ln788_1_fu_479_p2;
assign xor_ln416_fu_545_p2 = ~ p_Val2_7_fu_531_p2[3];
assign xor_ln781_fu_604_p2 = ~ and_ln781_fu_598_p2;
assign xor_ln785_2_fu_615_p2 = ~ deleted_zeros_fu_571_p3;
assign xor_ln785_3_fu_627_p2 = ~ p_Result_25_reg_1511;
assign xor_ln780_fu_579_p2 = ~ p_Result_29_reg_1524;
assign xor_ln786_1_fu_700_p2 = ~ and_ln786_fu_638_p2;
assign xor_ln785_fu_1061_p2 = ~ r_V_fu_1021_p3[1];
assign xor_ln340_fu_1075_p2 = ~ select_ln340_fu_1067_p3;
assign xor_ln1497_fu_1359_p2 = ~ icmp_ln1497_reg_1621;
assign xor_ln785_1_fu_431_p2 = ~ ret_fu_387_p2[16];
assign xor_ln786_fu_443_p2 = ~ ret_fu_387_p2[4];
assign xor_ln365_1_fu_671_p2 = ~ xor_ln365_fu_665_p2;
assign p_Val2_8_fu_749_p2 = ~ p_Val2_7_reg_1556[2:0];
assign _038_ = ~ ap_start;
assign _039_ = p_Result_7_reg_1535 == 14'h3fff;
assign _040_ = ! p_Result_7_reg_1535;
assign _041_ = p_Result_6_reg_1530 == 13'h1fff;
assign _042_ = ! { ret_fu_387_p2[3:0], 3'h0 };
assign _043_ = ! ret_V_24_fu_790_p2[2:0];
assign _044_ = ! op_3[2:0];
assign \mul_16ns_4s_20_1_1_U1.top_mul_16ns_4s_20_1_1_Multiplier_0_U.p  = $signed({ 1'h0, \mul_16ns_4s_20_1_1_U1.top_mul_16ns_4s_20_1_1_Multiplier_0_U.a  }) * $signed(\mul_16ns_4s_20_1_1_U1.top_mul_16ns_4s_20_1_1_Multiplier_0_U.b );
assign _045_ = $signed({ 1'h0, signbit_3_fu_1120_p2, 1'h0 }) < $signed(op_5);
assign _046_ = | ret_fu_387_p2[16:5];
assign _047_ = ret_fu_387_p2[16:5] != 12'hfff;
assign _048_ = | op_18[1:0];
assign _049_ = { op_5[1], op_5[1], op_5[1], op_5[1], op_5 } != { op_7, 1'h0 };
assign _050_ = | ret_V_23_fu_902_p2[2:0];
assign _051_ = { ret_V_21_reg_1492[1], ret_V_21_reg_1492[1], ret_V_21_reg_1492[1], ret_V_21_reg_1492[1], ret_V_21_reg_1492[1], ret_V_21_reg_1492[1], ret_V_21_reg_1492[1], ret_V_21_reg_1492[1], ret_V_21_reg_1492[1], ret_V_21_reg_1492[1], ret_V_21_reg_1492[1], ret_V_21_reg_1492[1], ret_V_21_reg_1492[1], ret_V_21_reg_1492[1], ret_V_21_reg_1492, 1'h0 } != { op_5[1], op_5[1], op_5[1], op_5[1], op_5[1], op_5[1], op_5[1], op_5[1], op_5[1], op_5[1], op_5[1], op_5[1], op_5[1], op_5[1], op_5[1], op_5[1], op_5 };
assign or_ln340_1_fu_763_p2 = or_ln340_reg_1569 | and_ln786_reg_1564;
assign or_ln340_2_fu_712_p2 = and_ln785_2_fu_694_p2 | and_ln340_fu_706_p2;
assign or_ln340_fu_644_p2 = overflow_1_fu_632_p2 | neg_src_fu_610_p2;
assign or_ln384_fu_491_p2 = underflow_fu_485_p2 | overflow_fu_437_p2;
assign or_ln406_fu_516_p2 = r_V_1_reg_1503[0] | p_Result_25_reg_1511;
assign or_ln785_1_fu_621_p2 = xor_ln785_2_fu_615_p2 | p_Val2_7_fu_531_p2[3];
assign or_ln785_2_fu_683_p2 = p_Result_25_reg_1511 | and_ln785_fu_677_p2;
assign or_ln785_fu_425_p2 = ret_fu_387_p2[4] | icmp_ln768_fu_419_p2;
assign or_ln788_1_fu_479_p2 = or_ln788_fu_473_p2 | icmp_ln786_fu_449_p2;
assign or_ln788_fu_473_p2 = xor_ln786_fu_443_p2 | icmp_ln790_fu_467_p2;
always @(posedge ap_clk)
ret_V_31_reg_1658 <= _025_;
always @(posedge ap_clk)
ret_V_32_cast_reg_1663 <= _026_;
always @(posedge ap_clk)
ret_V_30_reg_1641 <= _024_;
always @(posedge ap_clk)
ret_V_30_cast_reg_1646 <= _023_;
always @(posedge ap_clk)
ret_V_21_reg_1492 <= _021_;
always @(posedge ap_clk)
sext_ln1347_reg_1498 <= _032_;
always @(posedge ap_clk)
r_V_1_reg_1503 <= _020_;
always @(posedge ap_clk)
p_Result_25_reg_1511 <= _014_;
always @(posedge ap_clk)
p_Result_27_reg_1519 <= _015_;
always @(posedge ap_clk)
p_Result_29_reg_1524 <= _016_;
always @(posedge ap_clk)
p_Result_6_reg_1530 <= _017_;
always @(posedge ap_clk)
p_Result_7_reg_1535 <= _018_;
always @(posedge ap_clk)
op_9_V_reg_1584 <= _010_;
always @(posedge ap_clk)
ret_V_25_reg_1589 <= _022_;
always @(posedge ap_clk)
tmp_3_reg_1594 <= _034_;
always @(posedge ap_clk)
op_28_V_reg_1670 <= _009_;
always @(posedge ap_clk)
ret_V_33_reg_1675 <= _027_;
always @(posedge ap_clk)
ret_V_34_cast_reg_1680 <= _028_;
always @(posedge ap_clk)
icmp_ln851_2_reg_1687 <= _005_;
always @(posedge ap_clk)
lhs_V_2_reg_1616 <= _006_;
always @(posedge ap_clk)
icmp_ln1497_reg_1621 <= _004_;
always @(posedge ap_clk)
op_23_V_reg_1626 <= _008_;
always @(posedge ap_clk)
select_ln1192_reg_1631 <= _031_;
always @(posedge ap_clk)
ret_reg_1541 <= _029_;
always @(posedge ap_clk)
overflow_reg_1546 <= _013_;
always @(posedge ap_clk)
or_ln384_reg_1551 <= _012_;
always @(posedge ap_clk)
p_Val2_7_reg_1556 <= _019_;
always @(posedge ap_clk)
and_ln786_reg_1564 <= _002_;
always @(posedge ap_clk)
or_ln340_reg_1569 <= _011_;
always @(posedge ap_clk)
and_ln785_1_reg_1574 <= _001_;
always @(posedge ap_clk)
sel_tmp11_reg_1579 <= _030_;
always @(posedge ap_clk)
op_10_V_reg_1599 <= _007_;
always @(posedge ap_clk)
sext_ln850_reg_1605 <= _033_;
always @(posedge ap_clk)
add_ln691_reg_1611 <= _000_;
always @(posedge ap_clk)
ap_CS_fsm <= _003_;
assign _035_ = _037_ ? 2'h2 : 2'h1;
assign _052_ = ap_CS_fsm == 1'h1;
function [10:0] _181_;
input [10:0] a;
input [120:0] b;
input [10:0] s;
case (s)
11'b00000000001:
_181_ = b[10:0];
11'b00000000010:
_181_ = b[21:11];
11'b00000000100:
_181_ = b[32:22];
11'b00000001000:
_181_ = b[43:33];
11'b00000010000:
_181_ = b[54:44];
11'b00000100000:
_181_ = b[65:55];
11'b00001000000:
_181_ = b[76:66];
11'b00010000000:
_181_ = b[87:77];
11'b00100000000:
_181_ = b[98:88];
11'b01000000000:
_181_ = b[109:99];
11'b10000000000:
_181_ = b[120:110];
11'b00000000000:
_181_ = a;
default:
_181_ = 11'bx;
endcase
endfunction
assign ap_NS_fsm = _181_(11'hxxx, { 9'h000, _035_, 110'h0020080200802008020080200001 }, { _052_, _062_, _061_, _060_, _059_, _058_, _057_, _056_, _055_, _054_, _053_ });
assign _053_ = ap_CS_fsm == 11'h400;
assign _054_ = ap_CS_fsm == 10'h200;
assign _055_ = ap_CS_fsm == 9'h100;
assign _056_ = ap_CS_fsm == 8'h80;
assign _057_ = ap_CS_fsm == 7'h40;
assign _058_ = ap_CS_fsm == 6'h20;
assign _059_ = ap_CS_fsm == 5'h10;
assign _060_ = ap_CS_fsm == 4'h8;
assign _061_ = ap_CS_fsm == 3'h4;
assign _062_ = ap_CS_fsm == 2'h2;
assign op_30_ap_vld = ap_CS_fsm[10] ? 1'h1 : 1'h0;
assign ap_idle = _036_ ? 1'h1 : 1'h0;
assign _026_ = ap_CS_fsm[7] ? ret_V_31_fu_1343_p2[32:1] : ret_V_32_cast_reg_1663;
assign _025_ = ap_CS_fsm[7] ? ret_V_31_fu_1343_p2 : ret_V_31_reg_1658;
assign _023_ = ap_CS_fsm[6] ? ret_V_30_fu_1282_p2[32:1] : ret_V_30_cast_reg_1646;
assign _024_ = ap_CS_fsm[6] ? ret_V_30_fu_1282_p2 : ret_V_30_reg_1641;
assign _021_ = ap_CS_fsm[0] ? ret_V_21_fu_309_p3 : ret_V_21_reg_1492;
assign _018_ = ap_CS_fsm[1] ? r_V_1_fu_327_p2[19:6] : p_Result_7_reg_1535;
assign _017_ = ap_CS_fsm[1] ? r_V_1_fu_327_p2[19:7] : p_Result_6_reg_1530;
assign _016_ = ap_CS_fsm[1] ? r_V_1_fu_327_p2[6] : p_Result_29_reg_1524;
assign _015_ = ap_CS_fsm[1] ? r_V_1_fu_327_p2[5] : p_Result_27_reg_1519;
assign _014_ = ap_CS_fsm[1] ? r_V_1_fu_327_p2[19] : p_Result_25_reg_1511;
assign _020_ = ap_CS_fsm[1] ? r_V_1_fu_327_p2 : r_V_1_reg_1503;
assign _032_ = ap_CS_fsm[1] ? { ret_V_21_reg_1492[1], ret_V_21_reg_1492[1], ret_V_21_reg_1492[1], ret_V_21_reg_1492[1], ret_V_21_reg_1492[1], ret_V_21_reg_1492[1], ret_V_21_reg_1492[1], ret_V_21_reg_1492[1], ret_V_21_reg_1492[1], ret_V_21_reg_1492[1], ret_V_21_reg_1492[1], ret_V_21_reg_1492[1], ret_V_21_reg_1492[1], ret_V_21_reg_1492[1], ret_V_21_reg_1492 } : sext_ln1347_reg_1498;
assign _034_ = ap_CS_fsm[3] ? ret_V_25_fu_862_p2[7:1] : tmp_3_reg_1594;
assign _022_ = ap_CS_fsm[3] ? ret_V_25_fu_862_p2 : ret_V_25_reg_1589;
assign _010_ = ap_CS_fsm[3] ? op_9_V_fu_780_p3 : op_9_V_reg_1584;
assign _009_ = ap_CS_fsm[8] ? op_28_V_fu_1397_p2 : op_28_V_reg_1670;
assign _005_ = ap_CS_fsm[9] ? icmp_ln851_2_fu_1438_p2 : icmp_ln851_2_reg_1687;
assign _028_ = ap_CS_fsm[9] ? ret_V_33_fu_1418_p2[33:2] : ret_V_34_cast_reg_1680;
assign _027_ = ap_CS_fsm[9] ? ret_V_33_fu_1418_p2 : ret_V_33_reg_1675;
assign _031_ = ap_CS_fsm[5] ? select_ln1192_fu_1245_p3 : select_ln1192_reg_1631;
assign _008_ = ap_CS_fsm[5] ? op_23_V_fu_1239_p2 : op_23_V_reg_1626;
assign _004_ = ap_CS_fsm[5] ? icmp_ln1497_fu_1138_p2 : icmp_ln1497_reg_1621;
assign _006_ = ap_CS_fsm[5] ? lhs_V_2_fu_1099_p2 : lhs_V_2_reg_1616;
assign _030_ = ap_CS_fsm[2] ? sel_tmp11_fu_718_p2 : sel_tmp11_reg_1579;
assign _001_ = ap_CS_fsm[2] ? and_ln785_1_fu_688_p2 : and_ln785_1_reg_1574;
assign _011_ = ap_CS_fsm[2] ? or_ln340_fu_644_p2 : or_ln340_reg_1569;
assign _002_ = ap_CS_fsm[2] ? and_ln786_fu_638_p2 : and_ln786_reg_1564;
assign _019_ = ap_CS_fsm[2] ? p_Val2_7_fu_531_p2 : p_Val2_7_reg_1556;
assign _012_ = ap_CS_fsm[2] ? or_ln384_fu_491_p2 : or_ln384_reg_1551;
assign _013_ = ap_CS_fsm[2] ? overflow_fu_437_p2 : overflow_reg_1546;
assign _029_ = ap_CS_fsm[2] ? ret_fu_387_p2 : ret_reg_1541;
assign _000_ = ap_CS_fsm[4] ? add_ln691_fu_965_p2 : add_ln691_reg_1611;
assign _033_ = ap_CS_fsm[4] ? { tmp_3_reg_1594[6], tmp_3_reg_1594 } : sext_ln850_reg_1605;
assign _007_ = ap_CS_fsm[4] ? op_10_V_fu_956_p2 : op_10_V_reg_1599;
assign _003_ = ap_rst ? 11'h001 : ap_NS_fsm;
assign ret_fu_387_p2 = select_ln1347_fu_377_p3 - sext_ln1347_reg_1498;
assign Range1_all_ones_fu_561_p2 = _039_ ? 1'h1 : 1'h0;
assign Range1_all_zeros_fu_566_p2 = _040_ ? 1'h1 : 1'h0;
assign Range2_all_ones_fu_556_p2 = _041_ ? 1'h1 : 1'h0;
assign deleted_ones_fu_590_p3 = carry_2_fu_551_p2 ? and_ln780_fu_584_p2 : Range1_all_ones_fu_561_p2;
assign deleted_zeros_fu_571_p3 = carry_2_fu_551_p2 ? Range1_all_ones_fu_561_p2 : Range1_all_zeros_fu_566_p2;
assign icmp_ln1497_fu_1138_p2 = _045_ ? 1'h1 : 1'h0;
assign icmp_ln768_fu_419_p2 = _046_ ? 1'h1 : 1'h0;
assign icmp_ln786_fu_449_p2 = _047_ ? 1'h1 : 1'h0;
assign icmp_ln790_fu_467_p2 = _042_ ? 1'h1 : 1'h0;
assign icmp_ln851_1_fu_818_p2 = _043_ ? 1'h1 : 1'h0;
assign icmp_ln851_2_fu_1438_p2 = _048_ ? 1'h1 : 1'h0;
assign icmp_ln851_fu_289_p2 = _044_ ? 1'h1 : 1'h0;
assign lhs_V_2_fu_1099_p2 = _049_ ? 1'h1 : 1'h0;
assign op_8_V_fu_742_p3 = or_ln384_reg_1551 ? select_ln384_fu_735_p3 : { ret_reg_1541[4:0], 3'h0 };
assign op_9_V_fu_780_p3 = sel_tmp11_reg_1579 ? p_Val2_7_reg_1556 : select_ln785_fu_774_p3;
assign r_V_fu_1021_p3 = ret_V_22_fu_997_p2 ? { op_5[0], 1'h0 } : op_5;
assign r_fu_940_p2 = _050_ ? 1'h1 : 1'h0;
assign ret_V_21_fu_309_p3 = ret_V_20_fu_265_p2[4] ? select_ln850_fu_301_p3 : { 1'h0, ret_V_20_fu_265_p2[3] };
assign ret_V_27_fu_1223_p3 = ret_V_26_fu_1182_p2[33] ? select_ln850_3_fu_1215_p3 : { ret_V_26_fu_1182_p2[33], ret_V_26_fu_1182_p2[33], ret_V_26_fu_1182_p2[33], ret_V_26_fu_1182_p2[33], ret_V_26_fu_1182_p2[33], ret_V_26_fu_1182_p2[33], ret_V_26_fu_1182_p2[33], ret_V_26_fu_1182_p2[33], ret_V_26_fu_1182_p2[33], ret_V_26_fu_1182_p2[33], ret_V_26_fu_1182_p2[33], ret_V_26_fu_1182_p2[33], ret_V_26_fu_1182_p2[33], ret_V_26_fu_1182_p2[33], ret_V_26_fu_1182_p2[33], ret_V_26_fu_1182_p2[33], ret_V_26_fu_1182_p2[33], ret_V_26_fu_1182_p2[33], ret_V_26_fu_1182_p2[33], ret_V_26_fu_1182_p2[33], ret_V_26_fu_1182_p2[33], ret_V_26_fu_1182_p2[33], ret_V_26_fu_1182_p2[33], ret_V_26_fu_1182_p2[33], ret_V_26_fu_1182_p2[8:1] };
assign ret_V_32_fu_1386_p3 = ret_V_31_reg_1658[33] ? select_ln850_5_fu_1379_p3 : ret_V_32_cast_reg_1663;
assign ret_V_34_fu_1462_p3 = ret_V_33_reg_1675[34] ? select_ln850_6_fu_1456_p3 : ret_V_34_cast_reg_1680;
assign select_ln1192_fu_1245_p3 = op_14_V_fu_1081_p2 ? 32'd4294967295 : 32'd0;
assign select_ln1347_fu_377_p3 = op_2 ? 17'h1ffff : 17'h00000;
assign select_ln340_1_fu_767_p3 = or_ln340_1_fu_763_p2 ? { p_Result_29_reg_1524, p_Val2_8_fu_749_p2 } : p_Val2_7_reg_1556;
assign select_ln340_fu_1067_p3 = newsignbit_fu_1049_p2 ? xor_ln785_fu_1061_p2 : neg_src_2_fu_1055_p2;
assign select_ln353_2_fu_1324_p3 = ret_V_30_reg_1641[33] ? select_ln850_8_fu_1317_p3 : ret_V_30_cast_reg_1646;
assign select_ln353_fu_1163_p3 = ret_V_25_reg_1589[7] ? select_ln850_7_fu_1157_p3 : sext_ln850_reg_1605;
assign select_ln384_fu_735_p3 = overflow_reg_1546 ? 8'h7f : 8'h81;
assign select_ln69_fu_1231_p3 = op_12 ? 32'd4294967295 : 32'd0;
assign select_ln703_fu_249_p3 = op_2 ? 5'h18 : 5'h00;
assign select_ln785_fu_774_p3 = and_ln785_1_reg_1574 ? p_Val2_7_reg_1556 : select_ln340_1_fu_767_p3;
assign select_ln850_2_fu_834_p3 = icmp_ln851_1_fu_818_p2 ? { 1'h1, ret_V_24_fu_790_p2[7:3] } : ret_V_9_fu_824_p2;
assign select_ln850_3_fu_1215_p3 = op_10_V_reg_1599[0] ? add_ln691_1_fu_1209_p2 : { ret_V_26_fu_1182_p2[33], ret_V_26_fu_1182_p2[33], ret_V_26_fu_1182_p2[33], ret_V_26_fu_1182_p2[33], ret_V_26_fu_1182_p2[33], ret_V_26_fu_1182_p2[33], ret_V_26_fu_1182_p2[33], ret_V_26_fu_1182_p2[33], ret_V_26_fu_1182_p2[33], ret_V_26_fu_1182_p2[33], ret_V_26_fu_1182_p2[33], ret_V_26_fu_1182_p2[33], ret_V_26_fu_1182_p2[33], ret_V_26_fu_1182_p2[33], ret_V_26_fu_1182_p2[33], ret_V_26_fu_1182_p2[33], ret_V_26_fu_1182_p2[33], ret_V_26_fu_1182_p2[33], ret_V_26_fu_1182_p2[33], ret_V_26_fu_1182_p2[33], ret_V_26_fu_1182_p2[33], ret_V_26_fu_1182_p2[33], ret_V_26_fu_1182_p2[33], ret_V_26_fu_1182_p2[33], ret_V_26_fu_1182_p2[8:1] };
assign select_ln850_4_fu_842_p3 = ret_V_24_fu_790_p2[8] ? select_ln850_2_fu_834_p3 : { 1'h0, ret_V_24_fu_790_p2[7:3] };
assign select_ln850_5_fu_1379_p3 = op_16[0] ? add_ln691_3_fu_1374_p2 : ret_V_32_cast_reg_1663;
assign select_ln850_6_fu_1456_p3 = icmp_ln851_2_reg_1687 ? add_ln691_4_fu_1451_p2 : ret_V_34_cast_reg_1680;
assign select_ln850_7_fu_1157_p3 = op_9_V_reg_1584[0] ? add_ln691_reg_1611 : sext_ln850_reg_1605;
assign select_ln850_8_fu_1317_p3 = op_15[0] ? add_ln691_2_fu_1308_p2 : ret_V_30_cast_reg_1646;
assign select_ln850_fu_301_p3 = icmp_ln851_fu_289_p2 ? { 1'h1, ret_V_20_fu_265_p2[3] } : ret_V_2_fu_295_p2;
assign signbit_3_fu_1120_p2 = _051_ ? 1'h1 : 1'h0;
assign newsignbit_fu_1049_p2 = r_V_fu_1021_p3[0] ^ r_V_fu_1021_p3[1];
assign ret_V_22_fu_997_p2 = op_5[1] ^ and_ln850_fu_991_p2;
assign xor_ln365_fu_665_p2 = r_V_1_reg_1503[6] ^ p_Val2_7_fu_531_p2[3];
assign ap_CS_fsm_state1 = ap_CS_fsm[0];
assign ap_CS_fsm_state10 = ap_CS_fsm[9];
assign ap_CS_fsm_state11 = ap_CS_fsm[10];
assign ap_CS_fsm_state2 = ap_CS_fsm[1];
assign ap_CS_fsm_state3 = ap_CS_fsm[2];
assign ap_CS_fsm_state4 = ap_CS_fsm[3];
assign ap_CS_fsm_state5 = ap_CS_fsm[4];
assign ap_CS_fsm_state6 = ap_CS_fsm[5];
assign ap_CS_fsm_state7 = ap_CS_fsm[6];
assign ap_CS_fsm_state8 = ap_CS_fsm[7];
assign ap_CS_fsm_state9 = ap_CS_fsm[8];
assign ap_done = op_30_ap_vld;
assign ap_ready = op_30_ap_vld;
assign carry_fu_1041_p3 = r_V_fu_1021_p3[1];
assign lhs_fu_878_p1 = op_3;
assign lhs_fu_878_p3 = { op_3, 2'h0 };
assign op_11_V_fu_1126_p3 = { signbit_3_fu_1120_p2, 1'h0 };
assign p_Result_14_fu_754_p4 = { p_Result_29_reg_1524, p_Val2_8_fu_749_p2 };
assign p_Result_15_fu_806_p3 = ret_V_24_fu_790_p2[8];
assign p_Result_16_fu_1144_p3 = ret_V_25_reg_1589[7];
assign p_Result_17_fu_1198_p3 = ret_V_26_fu_1182_p2[33];
assign p_Result_18_fu_1298_p3 = ret_V_30_reg_1641[33];
assign p_Result_19_fu_1364_p3 = ret_V_31_reg_1658[33];
assign p_Result_1_fu_979_p1 = op_5;
assign p_Result_1_fu_979_p3 = op_5[1];
assign p_Result_20_fu_1444_p3 = ret_V_33_reg_1675[34];
assign p_Result_21_fu_1033_p3 = r_V_fu_1021_p3[1];
assign p_Result_22_fu_928_p3 = add_ln1192_1_fu_908_p2[3];
assign p_Result_23_fu_393_p3 = ret_fu_387_p2[16];
assign p_Result_24_fu_401_p3 = ret_fu_387_p2[4];
assign p_Result_26_fu_506_p3 = r_V_1_reg_1503[1];
assign p_Result_28_fu_537_p3 = p_Val2_7_fu_531_p2[3];
assign p_Result_3_fu_459_p3 = { ret_fu_387_p2[3:0], 3'h0 };
assign p_Result_s_fu_281_p3 = ret_V_20_fu_265_p2[4];
assign p_Val2_4_fu_727_p3 = { ret_reg_1541[4:0], 3'h0 };
assign p_Val2_6_fu_497_p4 = r_V_1_reg_1503[5:2];
assign r_1_fu_513_p1 = r_V_1_reg_1503[0];
assign r_V_1_fu_327_p0 = { ret_V_21_reg_1492[1], ret_V_21_reg_1492[1], ret_V_21_reg_1492[1], ret_V_21_reg_1492[1], ret_V_21_reg_1492[1], ret_V_21_reg_1492[1], ret_V_21_reg_1492[1], ret_V_21_reg_1492[1], ret_V_21_reg_1492[1], ret_V_21_reg_1492[1], ret_V_21_reg_1492[1], ret_V_21_reg_1492[1], ret_V_21_reg_1492[1], ret_V_21_reg_1492[1], ret_V_21_reg_1492 };
assign r_V_1_fu_327_p00 = { 4'h0, ret_V_21_reg_1492[1], ret_V_21_reg_1492[1], ret_V_21_reg_1492[1], ret_V_21_reg_1492[1], ret_V_21_reg_1492[1], ret_V_21_reg_1492[1], ret_V_21_reg_1492[1], ret_V_21_reg_1492[1], ret_V_21_reg_1492[1], ret_V_21_reg_1492[1], ret_V_21_reg_1492[1], ret_V_21_reg_1492[1], ret_V_21_reg_1492[1], ret_V_21_reg_1492[1], ret_V_21_reg_1492 };
assign r_V_fu_1021_p2 = op_5;
assign ret_V_24_cast_fu_1188_p4 = { ret_V_26_fu_1182_p2[33], ret_V_26_fu_1182_p2[33], ret_V_26_fu_1182_p2[33], ret_V_26_fu_1182_p2[33], ret_V_26_fu_1182_p2[33], ret_V_26_fu_1182_p2[33], ret_V_26_fu_1182_p2[33], ret_V_26_fu_1182_p2[33], ret_V_26_fu_1182_p2[33], ret_V_26_fu_1182_p2[33], ret_V_26_fu_1182_p2[33], ret_V_26_fu_1182_p2[33], ret_V_26_fu_1182_p2[33], ret_V_26_fu_1182_p2[33], ret_V_26_fu_1182_p2[33], ret_V_26_fu_1182_p2[33], ret_V_26_fu_1182_p2[33], ret_V_26_fu_1182_p2[33], ret_V_26_fu_1182_p2[33], ret_V_26_fu_1182_p2[33], ret_V_26_fu_1182_p2[33], ret_V_26_fu_1182_p2[33], ret_V_26_fu_1182_p2[33], ret_V_26_fu_1182_p2[33], ret_V_26_fu_1182_p2[8:1] };
assign ret_V_26_fu_1182_p2[32:9] = { ret_V_26_fu_1182_p2[33], ret_V_26_fu_1182_p2[33], ret_V_26_fu_1182_p2[33], ret_V_26_fu_1182_p2[33], ret_V_26_fu_1182_p2[33], ret_V_26_fu_1182_p2[33], ret_V_26_fu_1182_p2[33], ret_V_26_fu_1182_p2[33], ret_V_26_fu_1182_p2[33], ret_V_26_fu_1182_p2[33], ret_V_26_fu_1182_p2[33], ret_V_26_fu_1182_p2[33], ret_V_26_fu_1182_p2[33], ret_V_26_fu_1182_p2[33], ret_V_26_fu_1182_p2[33], ret_V_26_fu_1182_p2[33], ret_V_26_fu_1182_p2[33], ret_V_26_fu_1182_p2[33], ret_V_26_fu_1182_p2[33], ret_V_26_fu_1182_p2[33], ret_V_26_fu_1182_p2[33], ret_V_26_fu_1182_p2[33], ret_V_26_fu_1182_p2[33], ret_V_26_fu_1182_p2[33] };
assign ret_V_4_fu_971_p1 = op_5;
assign ret_V_4_fu_971_p3 = op_5[1];
assign ret_V_7_fu_796_p4 = ret_V_24_fu_790_p2[8:3];
assign ret_V_fu_271_p4 = ret_V_20_fu_265_p2[4:3];
assign rhs_2_fu_850_p3 = { select_ln850_4_fu_842_p3, 1'h0 };
assign rhs_6_fu_1270_p3 = { ret_V_29_fu_1261_p2, 1'h0 };
assign rhs_7_fu_1331_p3 = { select_ln353_2_fu_1324_p3, 1'h0 };
assign rhs_9_fu_1407_p3 = { op_28_V_reg_1670, 2'h0 };
assign sext_ln1192_1_fu_830_p1 = { op_9_V_fu_780_p3[3], op_9_V_fu_780_p3[3], op_9_V_fu_780_p3[3], op_9_V_fu_780_p3[3], op_9_V_fu_780_p3 };
assign sext_ln1192_2_fu_858_p1 = { select_ln850_4_fu_842_p3[5], select_ln850_4_fu_842_p3, 1'h0 };
assign sext_ln1192_3_fu_1178_p1 = { select_ln353_fu_1163_p3[7], select_ln353_fu_1163_p3[7], select_ln353_fu_1163_p3[7], select_ln353_fu_1163_p3[7], select_ln353_fu_1163_p3[7], select_ln353_fu_1163_p3[7], select_ln353_fu_1163_p3[7], select_ln353_fu_1163_p3[7], select_ln353_fu_1163_p3[7], select_ln353_fu_1163_p3[7], select_ln353_fu_1163_p3[7], select_ln353_fu_1163_p3[7], select_ln353_fu_1163_p3[7], select_ln353_fu_1163_p3[7], select_ln353_fu_1163_p3[7], select_ln353_fu_1163_p3[7], select_ln353_fu_1163_p3[7], select_ln353_fu_1163_p3[7], select_ln353_fu_1163_p3[7], select_ln353_fu_1163_p3[7], select_ln353_fu_1163_p3[7], select_ln353_fu_1163_p3[7], select_ln353_fu_1163_p3[7], select_ln353_fu_1163_p3[7], select_ln353_fu_1163_p3[7], select_ln353_fu_1163_p3, 1'h0 };
assign sext_ln1192_4_fu_1278_p1 = { ret_V_29_fu_1261_p2[31], ret_V_29_fu_1261_p2, 1'h0 };
assign sext_ln1192_5_fu_1339_p1 = { select_ln353_2_fu_1324_p3[31], select_ln353_2_fu_1324_p3, 1'h0 };
assign sext_ln1192_6_fu_1414_p1 = { op_28_V_reg_1670[31], op_28_V_reg_1670, 2'h0 };
assign sext_ln1192_fu_885_p1 = { op_3[3], op_3[3], op_3[3], op_3, 2'h0 };
assign sext_ln1299_1_fu_1007_p0 = op_5;
assign sext_ln1299_1_fu_1007_p1 = { op_5[1], op_5[1], op_5[1], op_5[1], op_5[1], op_5[1], op_5[1], op_5[1], op_5[1], op_5[1], op_5[1], op_5[1], op_5[1], op_5[1], op_5[1], op_5[1], op_5 };
assign sext_ln1299_2_fu_1011_p0 = op_5;
assign sext_ln1299_2_fu_1011_p1 = { op_5[1], op_5[1], op_5[1], op_5[1], op_5 };
assign sext_ln1299_fu_1003_p0 = op_5;
assign sext_ln1299_fu_1003_p1 = { op_5[1], op_5 };
assign sext_ln1347_fu_317_p1 = { ret_V_21_reg_1492[1], ret_V_21_reg_1492[1], ret_V_21_reg_1492[1], ret_V_21_reg_1492[1], ret_V_21_reg_1492[1], ret_V_21_reg_1492[1], ret_V_21_reg_1492[1], ret_V_21_reg_1492[1], ret_V_21_reg_1492[1], ret_V_21_reg_1492[1], ret_V_21_reg_1492[1], ret_V_21_reg_1492[1], ret_V_21_reg_1492[1], ret_V_21_reg_1492[1], ret_V_21_reg_1492 };
assign sext_ln1499_fu_1112_p1 = { ret_V_21_reg_1492[1], ret_V_21_reg_1492[1], ret_V_21_reg_1492[1], ret_V_21_reg_1492[1], ret_V_21_reg_1492[1], ret_V_21_reg_1492[1], ret_V_21_reg_1492[1], ret_V_21_reg_1492[1], ret_V_21_reg_1492[1], ret_V_21_reg_1492[1], ret_V_21_reg_1492[1], ret_V_21_reg_1492[1], ret_V_21_reg_1492[1], ret_V_21_reg_1492[1], ret_V_21_reg_1492, 1'h0 };
assign sext_ln703_1_fu_889_p0 = op_6;
assign sext_ln703_1_fu_889_p1 = { op_6[7], op_6 };
assign sext_ln703_2_fu_786_p1 = { op_8_V_fu_742_p3[7], op_8_V_fu_742_p3 };
assign sext_ln703_3_fu_1154_p1 = { op_10_V_reg_1599[5], op_10_V_reg_1599[5], op_10_V_reg_1599[5], op_10_V_reg_1599[5], op_10_V_reg_1599[5], op_10_V_reg_1599[5], op_10_V_reg_1599[5], op_10_V_reg_1599[5], op_10_V_reg_1599[5], op_10_V_reg_1599[5], op_10_V_reg_1599[5], op_10_V_reg_1599[5], op_10_V_reg_1599[5], op_10_V_reg_1599[5], op_10_V_reg_1599[5], op_10_V_reg_1599[5], op_10_V_reg_1599[5], op_10_V_reg_1599[5], op_10_V_reg_1599[5], op_10_V_reg_1599[5], op_10_V_reg_1599[5], op_10_V_reg_1599[5], op_10_V_reg_1599[5], op_10_V_reg_1599[5], op_10_V_reg_1599[5], op_10_V_reg_1599[5], op_10_V_reg_1599[5], op_10_V_reg_1599[5], op_10_V_reg_1599 };
assign sext_ln703_4_fu_1266_p0 = op_15;
assign sext_ln703_4_fu_1266_p1 = { op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15[3], op_15 };
assign sext_ln703_5_fu_1313_p0 = op_16;
assign sext_ln703_5_fu_1313_p1 = { op_16[15], op_16[15], op_16[15], op_16[15], op_16[15], op_16[15], op_16[15], op_16[15], op_16[15], op_16[15], op_16[15], op_16[15], op_16[15], op_16[15], op_16[15], op_16[15], op_16[15], op_16[15], op_16 };
assign sext_ln703_6_fu_1403_p0 = op_18;
assign sext_ln703_6_fu_1403_p1 = { op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18 };
assign sext_ln703_fu_257_p0 = op_3;
assign sext_ln703_fu_257_p1 = { op_3[3], op_3 };
assign sext_ln713_fu_924_p1 = { ret_V_23_fu_902_p2[8], ret_V_23_fu_902_p2[8:4] };
assign sext_ln850_fu_962_p1 = { tmp_3_reg_1594[6], tmp_3_reg_1594 };
assign shl_ln1192_fu_897_p0 = op_3;
assign shl_ln1192_fu_897_p2 = { op_3[1:0], 2'h0 };
assign shl_ln1299_fu_1015_p0 = op_5;
assign shl_ln1299_fu_1015_p2 = { op_5[0], 1'h0 };
assign shl_ln1_fu_1087_p3 = { op_7, 1'h0 };
assign tmp_1_fu_657_p3 = p_Val2_7_fu_531_p2[3];
assign tmp_2_fu_409_p4 = ret_fu_387_p2[16:5];
assign tmp_7_fu_1105_p3 = { ret_V_21_reg_1492, 1'h0 };
assign tmp_8_fu_1170_p3 = { select_ln353_fu_1163_p3, 1'h0 };
assign tmp_fu_650_p3 = r_V_1_reg_1503[6];
assign trunc_ln1192_1_fu_893_p0 = op_6;
assign trunc_ln1192_1_fu_893_p1 = op_6[3:0];
assign trunc_ln1192_fu_261_p0 = op_3;
assign trunc_ln1192_fu_261_p1 = op_3[2:0];
assign trunc_ln2_fu_914_p4 = ret_V_23_fu_902_p2[8:4];
assign trunc_ln415_fu_1029_p1 = r_V_fu_1021_p3[0];
assign trunc_ln718_fu_936_p1 = ret_V_23_fu_902_p2[2:0];
assign trunc_ln731_fu_724_p1 = ret_reg_1541[4:0];
assign trunc_ln790_fu_455_p1 = ret_fu_387_p2[3:0];
assign trunc_ln851_1_fu_814_p1 = ret_V_24_fu_790_p2[2:0];
assign trunc_ln851_2_fu_1151_p1 = op_9_V_reg_1584[0];
assign trunc_ln851_3_fu_1206_p1 = op_10_V_reg_1599[0];
assign trunc_ln851_4_fu_1305_p0 = op_15;
assign trunc_ln851_4_fu_1305_p1 = op_15[0];
assign trunc_ln851_5_fu_1371_p0 = op_16;
assign trunc_ln851_5_fu_1371_p1 = op_16[0];
assign trunc_ln851_6_fu_1434_p0 = op_18;
assign trunc_ln851_6_fu_1434_p1 = op_18[1:0];
assign trunc_ln851_fu_987_p0 = op_5;
assign trunc_ln851_fu_987_p1 = op_5[0];
assign zext_ln1192_fu_1253_p1 = { 31'h00000000, lhs_V_2_reg_1616 };
assign zext_ln1347_fu_384_p1 = { 1'h0, sext_ln1347_reg_1498 };
assign zext_ln1497_fu_1134_p1 = { 1'h0, signbit_3_fu_1120_p2, 1'h0 };
assign zext_ln1499_1_fu_1116_p1 = { 1'h0, ret_V_21_reg_1492[1], ret_V_21_reg_1492[1], ret_V_21_reg_1492[1], ret_V_21_reg_1492[1], ret_V_21_reg_1492[1], ret_V_21_reg_1492[1], ret_V_21_reg_1492[1], ret_V_21_reg_1492[1], ret_V_21_reg_1492[1], ret_V_21_reg_1492[1], ret_V_21_reg_1492[1], ret_V_21_reg_1492[1], ret_V_21_reg_1492[1], ret_V_21_reg_1492[1], ret_V_21_reg_1492, 1'h0 };
assign zext_ln1499_fu_1095_p1 = { 1'h0, op_7, 1'h0 };
assign zext_ln415_1_fu_527_p1 = { 3'h0, and_ln406_fu_521_p2 };
assign zext_ln415_fu_952_p1 = { 5'h00, and_ln408_fu_946_p2 };
assign zext_ln69_1_fu_1469_p1 = { 28'h0000000, op_19 };
assign zext_ln69_fu_1393_p1 = { 31'h00000000, xor_ln1497_fu_1359_p2 };
assign \mul_16ns_4s_20_1_1_U1.top_mul_16ns_4s_20_1_1_Multiplier_0_U.a  = \mul_16ns_4s_20_1_1_U1.din0 ;
assign \mul_16ns_4s_20_1_1_U1.top_mul_16ns_4s_20_1_1_Multiplier_0_U.b  = \mul_16ns_4s_20_1_1_U1.din1 ;
assign \mul_16ns_4s_20_1_1_U1.dout  = \mul_16ns_4s_20_1_1_U1.top_mul_16ns_4s_20_1_1_Multiplier_0_U.p ;
assign \mul_16ns_4s_20_1_1_U1.din0  = { ret_V_21_reg_1492[1], ret_V_21_reg_1492[1], ret_V_21_reg_1492[1], ret_V_21_reg_1492[1], ret_V_21_reg_1492[1], ret_V_21_reg_1492[1], ret_V_21_reg_1492[1], ret_V_21_reg_1492[1], ret_V_21_reg_1492[1], ret_V_21_reg_1492[1], ret_V_21_reg_1492[1], ret_V_21_reg_1492[1], ret_V_21_reg_1492[1], ret_V_21_reg_1492[1], ret_V_21_reg_1492 };
assign \mul_16ns_4s_20_1_1_U1.din1  = op_3;
assign r_V_1_fu_327_p2 = \mul_16ns_4s_20_1_1_U1.dout ;
endmodule


// Product machine:
module top_A_times_top_B (ap_start, op_0, op_12, op_15, op_16, op_18, op_19, op_2, op_3, op_5, op_6, op_7, ap_clk, unsafe_signal);
input ap_start;
input op_0;
input op_12;
input [3:0] op_15;
input [15:0] op_16;
input [3:0] op_18;
input [3:0] op_19;
input op_2;
input [3:0] op_3;
input [1:0] op_5;
input [7:0] op_6;
input [3:0] op_7;
input ap_clk;
output unsafe_signal;
reg _setup;
initial _setup = 1'b0;
always @ (posedge ap_clk) _setup <= 1'b1;
reg ap_start_internal;
always @ (posedge ap_clk) if (!_setup) ap_start_internal <= ap_start;
reg op_0_internal;
always @ (posedge ap_clk) if (!_setup) op_0_internal <= op_0;
reg op_12_internal;
always @ (posedge ap_clk) if (!_setup) op_12_internal <= op_12;
reg [3:0] op_15_internal;
always @ (posedge ap_clk) if (!_setup) op_15_internal <= op_15;
reg [15:0] op_16_internal;
always @ (posedge ap_clk) if (!_setup) op_16_internal <= op_16;
reg [3:0] op_18_internal;
always @ (posedge ap_clk) if (!_setup) op_18_internal <= op_18;
reg [3:0] op_19_internal;
always @ (posedge ap_clk) if (!_setup) op_19_internal <= op_19;
reg op_2_internal;
always @ (posedge ap_clk) if (!_setup) op_2_internal <= op_2;
reg [3:0] op_3_internal;
always @ (posedge ap_clk) if (!_setup) op_3_internal <= op_3;
reg [1:0] op_5_internal;
always @ (posedge ap_clk) if (!_setup) op_5_internal <= op_5;
reg [7:0] op_6_internal;
always @ (posedge ap_clk) if (!_setup) op_6_internal <= op_6;
reg [3:0] op_7_internal;
always @ (posedge ap_clk) if (!_setup) op_7_internal <= op_7;
wire ap_done_A;
wire ap_done_B;
wire ap_done_eq;
assign ap_done_eq = ap_done_A == ap_done_B;
wire ap_idle_A;
wire ap_idle_B;
wire ap_idle_eq;
assign ap_idle_eq = ap_idle_A == ap_idle_B;
wire ap_ready_A;
wire ap_ready_B;
wire ap_ready_eq;
assign ap_ready_eq = ap_ready_A == ap_ready_B;
wire [31:0] op_30_A;
wire [31:0] op_30_B;
wire op_30_eq;
assign op_30_eq = op_30_A == op_30_B;
wire op_30_ap_vld_A;
wire op_30_ap_vld_B;
wire clk_enable_A;
wire clk_enable_B;
assign clk_enable_A = _setup & (~op_30_ap_vld_A | op_30_ap_vld_B);
assign clk_enable_B = _setup;
wire divergent;
assign divergent = ~(ap_done_eq & ap_idle_eq & ap_ready_eq & op_30_eq);
assign unsafe_signal = op_30_ap_vld_A & op_30_ap_vld_B & divergent;
top_A instance_A (
    .ap_clk(ap_clk),
    .clk_enable(clk_enable_A),
    .ap_start(ap_start_internal),
    .op_0(op_0_internal),
    .op_12(op_12_internal),
    .op_15(op_15_internal),
    .op_16(op_16_internal),
    .op_18(op_18_internal),
    .op_19(op_19_internal),
    .op_2(op_2_internal),
    .op_3(op_3_internal),
    .op_5(op_5_internal),
    .op_6(op_6_internal),
    .op_7(op_7_internal),
    .ap_done(ap_done_A),
    .ap_idle(ap_idle_A),
    .ap_ready(ap_ready_A),
    .op_30(op_30_A),
    .op_30_ap_vld(op_30_ap_vld_A)
);
top_B instance_B (
    .ap_clk(ap_clk),
    .clk_enable(clk_enable_B),
    .ap_start(ap_start_internal),
    .op_0(op_0_internal),
    .op_12(op_12_internal),
    .op_15(op_15_internal),
    .op_16(op_16_internal),
    .op_18(op_18_internal),
    .op_19(op_19_internal),
    .op_2(op_2_internal),
    .op_3(op_3_internal),
    .op_5(op_5_internal),
    .op_6(op_6_internal),
    .op_7(op_7_internal),
    .ap_done(ap_done_B),
    .ap_idle(ap_idle_B),
    .ap_ready(ap_ready_B),
    .op_30(op_30_B),
    .op_30_ap_vld(op_30_ap_vld_B)
);
endmodule
