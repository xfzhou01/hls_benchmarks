// Processed by function `construct_kairos` in `verilog_tricks.py`.
// Machine A:
// Processed by function `add_clk_enable_signal` in `verilog_tricks.py`.
// Processed by function `remove_reset_signal` in `verilog_tricks.py`.
module top_A (
  ap_clk,
  ap_start,
  ap_done,
  ap_idle,
  ap_ready,
  op_0,
  op_1,
  op_4,
  op_5,
  op_6,
  op_11,
  op_18,
  op_27,
  op_27_ap_vld,
clk_enable
);
input clk_enable;


input ap_clk;
wire ap_rst;
assign ap_rst = op_27_ap_vld;
input ap_start;
input [7:0] op_0;
input [15:0] op_1;
input [1:0] op_11;
input [1:0] op_18;
input [7:0] op_4;
input [3:0] op_5;
input [1:0] op_6;
output ap_done;
output ap_idle;
output ap_ready;
output [31:0] op_27;
output op_27_ap_vld;


reg Range1_all_ones_reg_1903;
reg Range1_all_zeros_reg_1910;
reg Range2_all_ones_reg_1800;
reg [12:0] \add_26s_26ns_26_2_1_U9.top_add_26s_26ns_26_2_1_Adder_5_U.ain_s1 ;
reg [12:0] \add_26s_26ns_26_2_1_U9.top_add_26s_26ns_26_2_1_Adder_5_U.bin_s1 ;
reg \add_26s_26ns_26_2_1_U9.top_add_26s_26ns_26_2_1_Adder_5_U.carry_s1 ;
reg [12:0] \add_26s_26ns_26_2_1_U9.top_add_26s_26ns_26_2_1_Adder_5_U.sum_s1 ;
reg \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_4_U.ain_s1 ;
reg \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_4_U.bin_s1 ;
reg \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_4_U.carry_s1 ;
reg \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_4_U.sum_s1 ;
reg \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_4_U.ain_s1 ;
reg \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_4_U.bin_s1 ;
reg \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_4_U.carry_s1 ;
reg \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_4_U.sum_s1 ;
reg \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_4_U.ain_s1 ;
reg \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_4_U.bin_s1 ;
reg \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_4_U.carry_s1 ;
reg \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_4_U.sum_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s1 ;
reg \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.carry_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.sum_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s1 ;
reg \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_7_U.carry_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_7_U.sum_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s1 ;
reg \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_7_U.carry_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_7_U.sum_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s1 ;
reg \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_7_U.carry_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_7_U.sum_s1 ;
reg [15:0] \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.ain_s1 ;
reg [15:0] \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.bin_s1 ;
reg \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.carry_s1 ;
reg [15:0] \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.sum_s1 ;
reg [15:0] \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_9_U.ain_s1 ;
reg [15:0] \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_9_U.bin_s1 ;
reg \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_9_U.carry_s1 ;
reg [15:0] \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_9_U.sum_s1 ;
reg [16:0] \add_34s_34s_34_2_1_U12.top_add_34s_34s_34_2_1_Adder_6_U.ain_s1 ;
reg [16:0] \add_34s_34s_34_2_1_U12.top_add_34s_34s_34_2_1_Adder_6_U.bin_s1 ;
reg \add_34s_34s_34_2_1_U12.top_add_34s_34s_34_2_1_Adder_6_U.carry_s1 ;
reg [16:0] \add_34s_34s_34_2_1_U12.top_add_34s_34s_34_2_1_Adder_6_U.sum_s1 ;
reg [16:0] \add_34s_34s_34_2_1_U21.top_add_34s_34s_34_2_1_Adder_6_U.ain_s1 ;
reg [16:0] \add_34s_34s_34_2_1_U21.top_add_34s_34s_34_2_1_Adder_6_U.bin_s1 ;
reg \add_34s_34s_34_2_1_U21.top_add_34s_34s_34_2_1_Adder_6_U.carry_s1 ;
reg [16:0] \add_34s_34s_34_2_1_U21.top_add_34s_34s_34_2_1_Adder_6_U.sum_s1 ;
reg [16:0] \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_6_U.ain_s1 ;
reg [16:0] \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_6_U.bin_s1 ;
reg \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_6_U.carry_s1 ;
reg [16:0] \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_6_U.sum_s1 ;
reg [18:0] \add_37s_37s_37_2_1_U18.top_add_37s_37s_37_2_1_Adder_11_U.ain_s1 ;
reg [18:0] \add_37s_37s_37_2_1_U18.top_add_37s_37s_37_2_1_Adder_11_U.bin_s1 ;
reg \add_37s_37s_37_2_1_U18.top_add_37s_37s_37_2_1_Adder_11_U.carry_s1 ;
reg [17:0] \add_37s_37s_37_2_1_U18.top_add_37s_37s_37_2_1_Adder_11_U.sum_s1 ;
reg [1:0] \add_3s_3ns_3_2_1_U17.top_add_3s_3ns_3_2_1_Adder_10_U.ain_s1 ;
reg [1:0] \add_3s_3ns_3_2_1_U17.top_add_3s_3ns_3_2_1_Adder_10_U.bin_s1 ;
reg \add_3s_3ns_3_2_1_U17.top_add_3s_3ns_3_2_1_Adder_10_U.carry_s1 ;
reg \add_3s_3ns_3_2_1_U17.top_add_3s_3ns_3_2_1_Adder_10_U.sum_s1 ;
reg [1:0] \add_4ns_4ns_4_2_1_U3.top_add_4ns_4ns_4_2_1_Adder_2_U.ain_s1 ;
reg [1:0] \add_4ns_4ns_4_2_1_U3.top_add_4ns_4ns_4_2_1_Adder_2_U.bin_s1 ;
reg \add_4ns_4ns_4_2_1_U3.top_add_4ns_4ns_4_2_1_Adder_2_U.carry_s1 ;
reg [1:0] \add_4ns_4ns_4_2_1_U3.top_add_4ns_4ns_4_2_1_Adder_2_U.sum_s1 ;
reg [3:0] \add_7s_7ns_7_2_1_U10.top_add_7s_7ns_7_2_1_Adder_3_U.ain_s1 ;
reg [3:0] \add_7s_7ns_7_2_1_U10.top_add_7s_7ns_7_2_1_Adder_3_U.bin_s1 ;
reg \add_7s_7ns_7_2_1_U10.top_add_7s_7ns_7_2_1_Adder_3_U.carry_s1 ;
reg [2:0] \add_7s_7ns_7_2_1_U10.top_add_7s_7ns_7_2_1_Adder_3_U.sum_s1 ;
reg [3:0] \add_7s_7ns_7_2_1_U6.top_add_7s_7ns_7_2_1_Adder_3_U.ain_s1 ;
reg [3:0] \add_7s_7ns_7_2_1_U6.top_add_7s_7ns_7_2_1_Adder_3_U.bin_s1 ;
reg \add_7s_7ns_7_2_1_U6.top_add_7s_7ns_7_2_1_Adder_3_U.carry_s1 ;
reg [2:0] \add_7s_7ns_7_2_1_U6.top_add_7s_7ns_7_2_1_Adder_3_U.sum_s1 ;
reg [3:0] \add_8ns_8ns_8_2_1_U1.top_add_8ns_8ns_8_2_1_Adder_0_U.ain_s1 ;
reg [3:0] \add_8ns_8ns_8_2_1_U1.top_add_8ns_8ns_8_2_1_Adder_0_U.bin_s1 ;
reg \add_8ns_8ns_8_2_1_U1.top_add_8ns_8ns_8_2_1_Adder_0_U.carry_s1 ;
reg [3:0] \add_8ns_8ns_8_2_1_U1.top_add_8ns_8ns_8_2_1_Adder_0_U.sum_s1 ;
reg [31:0] add_ln691_1_reg_2018;
reg [31:0] add_ln691_2_reg_2199;
reg [31:0] add_ln691_3_reg_2237;
reg [31:0] add_ln691_4_reg_2279;
reg [6:0] add_ln691_reg_1948;
reg and_ln340_reg_2177;
reg and_ln410_reg_2138;
reg and_ln412_reg_1833;
reg and_ln414_1_reg_2087;
reg and_ln788_1_reg_1931;
reg [48:0] ap_CS_fsm = 49'h0000000000001;
reg [31:0] \ashr_32s_32s_32_7_1_U4.din1_cast_array[0] ;
reg [31:0] \ashr_32s_32s_32_7_1_U4.din1_cast_array[1] ;
reg [31:0] \ashr_32s_32s_32_7_1_U4.din1_cast_array[2] ;
reg [31:0] \ashr_32s_32s_32_7_1_U4.din1_cast_array[3] ;
reg [31:0] \ashr_32s_32s_32_7_1_U4.din1_cast_array[4] ;
reg [31:0] \ashr_32s_32s_32_7_1_U4.din1_cast_array[5] ;
reg [31:0] \ashr_32s_32s_32_7_1_U4.dout_array[0] ;
reg [31:0] \ashr_32s_32s_32_7_1_U4.dout_array[1] ;
reg [31:0] \ashr_32s_32s_32_7_1_U4.dout_array[2] ;
reg [31:0] \ashr_32s_32s_32_7_1_U4.dout_array[3] ;
reg [31:0] \ashr_32s_32s_32_7_1_U4.dout_array[4] ;
reg [31:0] \ashr_32s_32s_32_7_1_U4.dout_array[5] ;
reg [31:0] ashr_ln1497_reg_1667;
reg carry_1_reg_1896;
reg icmp_ln414_reg_2050;
reg icmp_ln785_reg_1705;
reg icmp_ln786_1_reg_1710;
reg icmp_ln786_reg_1726;
reg icmp_ln790_reg_1715;
reg icmp_ln851_1_reg_2008;
reg icmp_ln851_2_reg_1630;
reg icmp_ln851_3_reg_1848;
reg icmp_ln851_4_reg_2133;
reg icmp_ln851_reg_1575;
reg [3:0] \mul_4s_2s_6_7_1_U8.top_mul_4s_2s_6_7_1_Mul_DSP_0_U.a_reg0 ;
reg [1:0] \mul_4s_2s_6_7_1_U8.top_mul_4s_2s_6_7_1_Mul_DSP_0_U.b_reg0 ;
reg [5:0] \mul_4s_2s_6_7_1_U8.top_mul_4s_2s_6_7_1_Mul_DSP_0_U.buff0 ;
reg [5:0] \mul_4s_2s_6_7_1_U8.top_mul_4s_2s_6_7_1_Mul_DSP_0_U.buff1 ;
reg [5:0] \mul_4s_2s_6_7_1_U8.top_mul_4s_2s_6_7_1_Mul_DSP_0_U.buff2 ;
reg [5:0] \mul_4s_2s_6_7_1_U8.top_mul_4s_2s_6_7_1_Mul_DSP_0_U.buff3 ;
reg [5:0] \mul_4s_2s_6_7_1_U8.top_mul_4s_2s_6_7_1_Mul_DSP_0_U.buff4 ;
reg [3:0] op_12_V_reg_1789;
reg [1:0] op_14_V_reg_1953;
reg [1:0] op_17_V_reg_2204;
reg [3:0] op_19_V_reg_2193;
reg [31:0] op_23_V_reg_2097;
reg [31:0] op_26_V_reg_2252;
reg [7:0] op_2_V_reg_1741;
reg [3:0] or_ln1195_1_reg_1806;
reg [4:0] or_ln1195_reg_1794;
reg or_ln384_1_reg_1943;
reg or_ln384_reg_1731;
reg overflow_1_reg_1925;
reg overflow_reg_1720;
reg p_Result_23_reg_1682;
reg p_Result_24_reg_2076;
reg p_Result_26_reg_2187;
reg p_Result_27_reg_2034;
reg p_Result_28_reg_2149;
reg p_Result_29_reg_1812;
reg p_Result_32_reg_1879;
reg [4:0] p_Result_s_22_reg_1694;
reg [1:0] p_Val2_4_reg_2182;
reg [2:0] p_Val2_6_reg_2143;
reg [1:0] p_Val2_8_reg_1818;
reg [1:0] p_Val2_9_reg_1873;
reg [3:0] r_V_1_reg_2070;
reg [3:0] r_V_2_reg_2028;
reg [5:0] r_V_reg_1979;
reg [31:0] ret_V_19_cast_reg_2001;
reg [1:0] ret_V_19_reg_2023;
reg [7:0] ret_V_1_reg_1585;
reg [15:0] ret_V_20_reg_1608;
reg [3:0] ret_V_21_reg_1661;
reg [31:0] ret_V_22_cast_reg_2160;
reg [25:0] ret_V_22_reg_1915;
reg [33:0] ret_V_23_reg_1996;
reg [31:0] ret_V_24_reg_2045;
reg [31:0] ret_V_25_cast_reg_2230;
reg [36:0] ret_V_25_reg_2155;
reg [33:0] ret_V_26_reg_2225;
reg [31:0] ret_V_27_reg_2242;
reg [31:0] ret_V_28_cast_reg_2272;
reg [33:0] ret_V_28_reg_2267;
reg [7:0] ret_V_2_reg_1597;
reg [1:0] ret_V_3_cast_reg_1984;
reg [1:0] ret_V_3_reg_2013;
reg [6:0] ret_V_5_reg_1779;
reg [3:0] ret_V_7_reg_1640;
reg [3:0] ret_V_8_cast_reg_1613;
reg [6:0] ret_V_9_reg_2092;
reg [7:0] ret_V_reg_1568;
reg [1:0] ret_reg_1752;
reg rhs_1_reg_1590;
reg [31:0] select_ln1497_reg_1677;
reg [31:0] select_ln353_2_reg_2210;
reg [6:0] select_ln353_reg_1959;
reg [3:0] sext_ln745_reg_2172;
reg [6:0] sext_ln850_reg_1936;
reg [31:0] \shl_32s_32s_32_7_1_U5.din1_cast_array[0] ;
reg [31:0] \shl_32s_32s_32_7_1_U5.din1_cast_array[1] ;
reg [31:0] \shl_32s_32s_32_7_1_U5.din1_cast_array[2] ;
reg [31:0] \shl_32s_32s_32_7_1_U5.din1_cast_array[3] ;
reg [31:0] \shl_32s_32s_32_7_1_U5.din1_cast_array[4] ;
reg [31:0] \shl_32s_32s_32_7_1_U5.din1_cast_array[5] ;
reg [31:0] \shl_32s_32s_32_7_1_U5.dout_array[0] ;
reg [31:0] \shl_32s_32s_32_7_1_U5.dout_array[1] ;
reg [31:0] \shl_32s_32s_32_7_1_U5.dout_array[2] ;
reg [31:0] \shl_32s_32s_32_7_1_U5.dout_array[3] ;
reg [31:0] \shl_32s_32s_32_7_1_U5.dout_array[4] ;
reg [31:0] \shl_32s_32s_32_7_1_U5.dout_array[5] ;
reg \shl_4s_1ns_4_7_1_U11.din1_cast_array[0] ;
reg \shl_4s_1ns_4_7_1_U11.din1_cast_array[1] ;
reg \shl_4s_1ns_4_7_1_U11.din1_cast_array[2] ;
reg \shl_4s_1ns_4_7_1_U11.din1_cast_array[3] ;
reg \shl_4s_1ns_4_7_1_U11.din1_cast_array[4] ;
reg \shl_4s_1ns_4_7_1_U11.din1_cast_array[5] ;
reg [3:0] \shl_4s_1ns_4_7_1_U11.dout_array[0] ;
reg [3:0] \shl_4s_1ns_4_7_1_U11.dout_array[1] ;
reg [3:0] \shl_4s_1ns_4_7_1_U11.dout_array[2] ;
reg [3:0] \shl_4s_1ns_4_7_1_U11.dout_array[3] ;
reg [3:0] \shl_4s_1ns_4_7_1_U11.dout_array[4] ;
reg [3:0] \shl_4s_1ns_4_7_1_U11.dout_array[5] ;
reg [31:0] shl_ln1497_reg_1672;
reg signbit_reg_1784;
reg [3:0] \sub_7s_7ns_7_2_1_U15.top_sub_7s_7ns_7_2_1_Adder_8_U.ain_s1 ;
reg [3:0] \sub_7s_7ns_7_2_1_U15.top_sub_7s_7ns_7_2_1_Adder_8_U.bin_s1 ;
reg \sub_7s_7ns_7_2_1_U15.top_sub_7s_7ns_7_2_1_Adder_8_U.carry_s1 ;
reg [2:0] \sub_7s_7ns_7_2_1_U15.top_sub_7s_7ns_7_2_1_Adder_8_U.sum_s1 ;
reg [4:0] \sub_9ns_9s_9_2_1_U2.top_sub_9ns_9s_9_2_1_Adder_1_U.ain_s1 ;
reg [4:0] \sub_9ns_9s_9_2_1_U2.top_sub_9ns_9s_9_2_1_Adder_1_U.bin_s1 ;
reg \sub_9ns_9s_9_2_1_U2.top_sub_9ns_9s_9_2_1_Adder_1_U.carry_s1 ;
reg [3:0] \sub_9ns_9s_9_2_1_U2.top_sub_9ns_9s_9_2_1_Adder_1_U.sum_s1 ;
reg [8:0] sub_ln1497_reg_1635;
reg [4:0] tmp_1_reg_1858;
reg tmp_23_reg_1823;
reg tmp_4_reg_1688;
reg tmp_reg_1603;
reg [5:0] tmp_s_reg_1920;
reg trunc_ln1195_reg_1757;
reg [1:0] trunc_ln1_reg_2082;
reg [1:0] trunc_ln708_1_reg_2040;
reg [1:0] trunc_ln790_reg_1700;
reg [2:0] trunc_ln851_1_reg_1991;
reg [7:0] trunc_ln851_2_reg_1620;
reg [4:0] trunc_ln851_3_reg_1828;
reg [2:0] trunc_ln851_5_reg_2102;
reg [6:0] trunc_ln8_reg_1747;
reg ush_reg_1772;
reg xor_ln410_reg_2107;
wire _0000_;
wire _0001_;
wire _0002_;
wire [31:0] _0003_;
wire [31:0] _0004_;
wire [31:0] _0005_;
wire [31:0] _0006_;
wire [6:0] _0007_;
wire _0008_;
wire _0009_;
wire _0010_;
wire _0011_;
wire _0012_;
wire [48:0] _0013_;
wire [31:0] _0014_;
wire _0015_;
wire _0016_;
wire _0017_;
wire _0018_;
wire _0019_;
wire _0020_;
wire _0021_;
wire _0022_;
wire _0023_;
wire _0024_;
wire _0025_;
wire [3:0] _0026_;
wire [1:0] _0027_;
wire [1:0] _0028_;
wire [3:0] _0029_;
wire [31:0] _0030_;
wire [31:0] _0031_;
wire [7:0] _0032_;
wire [3:0] _0033_;
wire [4:0] _0034_;
wire _0035_;
wire _0036_;
wire _0037_;
wire _0038_;
wire _0039_;
wire _0040_;
wire _0041_;
wire _0042_;
wire _0043_;
wire _0044_;
wire _0045_;
wire [4:0] _0046_;
wire [1:0] _0047_;
wire [2:0] _0048_;
wire [1:0] _0049_;
wire [1:0] _0050_;
wire [3:0] _0051_;
wire [3:0] _0052_;
wire [5:0] _0053_;
wire [31:0] _0054_;
wire [1:0] _0055_;
wire [7:0] _0056_;
wire [15:0] _0057_;
wire [3:0] _0058_;
wire [31:0] _0059_;
wire [25:0] _0060_;
wire [33:0] _0061_;
wire [31:0] _0062_;
wire [31:0] _0063_;
wire [36:0] _0064_;
wire [33:0] _0065_;
wire [31:0] _0066_;
wire [31:0] _0067_;
wire [33:0] _0068_;
wire [7:0] _0069_;
wire [1:0] _0070_;
wire [1:0] _0071_;
wire [1:0] _0072_;
wire [3:0] _0073_;
wire [3:0] _0074_;
wire [6:0] _0075_;
wire [7:0] _0076_;
wire [1:0] _0077_;
wire _0078_;
wire [31:0] _0079_;
wire [31:0] _0080_;
wire [6:0] _0081_;
wire [3:0] _0082_;
wire [6:0] _0083_;
wire [31:0] _0084_;
wire _0085_;
wire [8:0] _0086_;
wire [4:0] _0087_;
wire _0088_;
wire _0089_;
wire _0090_;
wire [5:0] _0091_;
wire _0092_;
wire [1:0] _0093_;
wire [1:0] _0094_;
wire [1:0] _0095_;
wire [2:0] _0096_;
wire [7:0] _0097_;
wire [2:0] _0098_;
wire [6:0] _0099_;
wire _0100_;
wire _0101_;
wire [1:0] _0102_;
wire _0103_;
wire _0104_;
wire _0105_;
wire _0106_;
wire _0107_;
wire _0108_;
wire _0109_;
wire _0110_;
wire _0111_;
wire _0112_;
wire _0113_;
wire _0114_;
wire _0115_;
wire _0116_;
wire _0117_;
wire _0118_;
wire _0119_;
wire [12:0] _0120_;
wire [12:0] _0121_;
wire _0122_;
wire [12:0] _0123_;
wire [13:0] _0124_;
wire [13:0] _0125_;
wire _0126_;
wire _0127_;
wire _0128_;
wire _0129_;
wire [1:0] _0130_;
wire [1:0] _0131_;
wire _0132_;
wire _0133_;
wire _0134_;
wire _0135_;
wire [1:0] _0136_;
wire [1:0] _0137_;
wire _0138_;
wire _0139_;
wire _0140_;
wire _0141_;
wire [1:0] _0142_;
wire [1:0] _0143_;
wire [15:0] _0144_;
wire [15:0] _0145_;
wire _0146_;
wire [15:0] _0147_;
wire [16:0] _0148_;
wire [16:0] _0149_;
wire [15:0] _0150_;
wire [15:0] _0151_;
wire _0152_;
wire [15:0] _0153_;
wire [16:0] _0154_;
wire [16:0] _0155_;
wire [15:0] _0156_;
wire [15:0] _0157_;
wire _0158_;
wire [15:0] _0159_;
wire [16:0] _0160_;
wire [16:0] _0161_;
wire [15:0] _0162_;
wire [15:0] _0163_;
wire _0164_;
wire [15:0] _0165_;
wire [16:0] _0166_;
wire [16:0] _0167_;
wire [15:0] _0168_;
wire [15:0] _0169_;
wire _0170_;
wire [15:0] _0171_;
wire [16:0] _0172_;
wire [16:0] _0173_;
wire [15:0] _0174_;
wire [15:0] _0175_;
wire _0176_;
wire [15:0] _0177_;
wire [16:0] _0178_;
wire [16:0] _0179_;
wire [16:0] _0180_;
wire [16:0] _0181_;
wire _0182_;
wire [16:0] _0183_;
wire [17:0] _0184_;
wire [17:0] _0185_;
wire [16:0] _0186_;
wire [16:0] _0187_;
wire _0188_;
wire [16:0] _0189_;
wire [17:0] _0190_;
wire [17:0] _0191_;
wire [16:0] _0192_;
wire [16:0] _0193_;
wire _0194_;
wire [16:0] _0195_;
wire [17:0] _0196_;
wire [17:0] _0197_;
wire [18:0] _0198_;
wire [18:0] _0199_;
wire _0200_;
wire [17:0] _0201_;
wire [18:0] _0202_;
wire [19:0] _0203_;
wire [1:0] _0204_;
wire [1:0] _0205_;
wire _0206_;
wire _0207_;
wire [1:0] _0208_;
wire [2:0] _0209_;
wire [1:0] _0210_;
wire [1:0] _0211_;
wire _0212_;
wire [1:0] _0213_;
wire [2:0] _0214_;
wire [2:0] _0215_;
wire [3:0] _0216_;
wire [3:0] _0217_;
wire _0218_;
wire [2:0] _0219_;
wire [3:0] _0220_;
wire [4:0] _0221_;
wire [3:0] _0222_;
wire [3:0] _0223_;
wire _0224_;
wire [2:0] _0225_;
wire [3:0] _0226_;
wire [4:0] _0227_;
wire [3:0] _0228_;
wire [3:0] _0229_;
wire _0230_;
wire [3:0] _0231_;
wire [4:0] _0232_;
wire [4:0] _0233_;
wire [31:0] _0234_;
wire [31:0] _0235_;
wire [31:0] _0236_;
wire [31:0] _0237_;
wire [31:0] _0238_;
wire [31:0] _0239_;
wire [31:0] _0240_;
wire [31:0] _0241_;
wire [31:0] _0242_;
wire [31:0] _0243_;
wire [31:0] _0244_;
wire [31:0] _0245_;
wire [31:0] _0246_;
wire [31:0] _0247_;
wire [31:0] _0248_;
wire [31:0] _0249_;
wire [31:0] _0250_;
wire [31:0] _0251_;
wire [31:0] _0252_;
wire [31:0] _0253_;
wire [31:0] _0254_;
wire [31:0] _0255_;
wire [31:0] _0256_;
wire [31:0] _0257_;
wire [31:0] _0258_;
wire [31:0] _0259_;
wire [31:0] _0260_;
wire [31:0] _0261_;
wire [31:0] _0262_;
wire [31:0] _0263_;
wire [3:0] _0264_;
wire [1:0] _0265_;
wire [5:0] _0266_;
wire [5:0] _0267_;
wire [5:0] _0268_;
wire [5:0] _0269_;
wire [5:0] _0270_;
wire [31:0] _0271_;
wire [31:0] _0272_;
wire [31:0] _0273_;
wire [31:0] _0274_;
wire [31:0] _0275_;
wire [31:0] _0276_;
wire [31:0] _0277_;
wire [31:0] _0278_;
wire [31:0] _0279_;
wire [31:0] _0280_;
wire [31:0] _0281_;
wire [31:0] _0282_;
wire [31:0] _0283_;
wire [31:0] _0284_;
wire [31:0] _0285_;
wire [31:0] _0286_;
wire [31:0] _0287_;
wire [31:0] _0288_;
wire [31:0] _0289_;
wire [31:0] _0290_;
wire [31:0] _0291_;
wire [31:0] _0292_;
wire [31:0] _0293_;
wire [31:0] _0294_;
wire [31:0] _0295_;
wire [31:0] _0296_;
wire [31:0] _0297_;
wire [31:0] _0298_;
wire [31:0] _0299_;
wire [31:0] _0300_;
wire _0301_;
wire _0302_;
wire _0303_;
wire _0304_;
wire _0305_;
wire _0306_;
wire [3:0] _0307_;
wire [3:0] _0308_;
wire [3:0] _0309_;
wire [3:0] _0310_;
wire [3:0] _0311_;
wire [3:0] _0312_;
wire [3:0] _0313_;
wire _0314_;
wire [3:0] _0315_;
wire _0316_;
wire [3:0] _0317_;
wire _0318_;
wire [3:0] _0319_;
wire _0320_;
wire [3:0] _0321_;
wire _0322_;
wire [3:0] _0323_;
wire _0324_;
wire [3:0] _0325_;
wire [3:0] _0326_;
wire _0327_;
wire [2:0] _0328_;
wire [3:0] _0329_;
wire [4:0] _0330_;
wire [4:0] _0331_;
wire [4:0] _0332_;
wire _0333_;
wire [3:0] _0334_;
wire [4:0] _0335_;
wire [5:0] _0336_;
wire _0337_;
wire _0338_;
wire _0339_;
wire _0340_;
wire _0341_;
wire _0342_;
wire _0343_;
wire _0344_;
wire _0345_;
wire _0346_;
wire _0347_;
wire _0348_;
wire _0349_;
wire _0350_;
wire _0351_;
wire _0352_;
wire _0353_;
wire _0354_;
wire _0355_;
wire _0356_;
wire _0357_;
wire _0358_;
wire _0359_;
wire _0360_;
wire _0361_;
wire _0362_;
wire _0363_;
wire _0364_;
wire _0365_;
wire _0366_;
wire _0367_;
wire _0368_;
wire _0369_;
wire _0370_;
wire _0371_;
wire _0372_;
wire _0373_;
wire _0374_;
wire _0375_;
wire _0376_;
wire _0377_;
wire _0378_;
wire _0379_;
wire _0380_;
wire _0381_;
wire _0382_;
wire _0383_;
wire _0384_;
wire _0385_;
wire _0386_;
wire _0387_;
wire _0388_;
wire _0389_;
wire _0390_;
wire _0391_;
wire _0392_;
wire Range1_all_ones_fu_840_p2;
wire Range1_all_zeros_fu_846_p2;
wire [3:0] Range2_all_ones_fu_635_p1;
wire \add_26s_26ns_26_2_1_U9.ce ;
wire \add_26s_26ns_26_2_1_U9.clk ;
wire [25:0] \add_26s_26ns_26_2_1_U9.din0 ;
wire [25:0] \add_26s_26ns_26_2_1_U9.din1 ;
wire [25:0] \add_26s_26ns_26_2_1_U9.dout ;
wire \add_26s_26ns_26_2_1_U9.reset ;
wire [25:0] \add_26s_26ns_26_2_1_U9.top_add_26s_26ns_26_2_1_Adder_5_U.a ;
wire [25:0] \add_26s_26ns_26_2_1_U9.top_add_26s_26ns_26_2_1_Adder_5_U.ain_s0 ;
wire [25:0] \add_26s_26ns_26_2_1_U9.top_add_26s_26ns_26_2_1_Adder_5_U.b ;
wire [25:0] \add_26s_26ns_26_2_1_U9.top_add_26s_26ns_26_2_1_Adder_5_U.bin_s0 ;
wire \add_26s_26ns_26_2_1_U9.top_add_26s_26ns_26_2_1_Adder_5_U.ce ;
wire \add_26s_26ns_26_2_1_U9.top_add_26s_26ns_26_2_1_Adder_5_U.clk ;
wire \add_26s_26ns_26_2_1_U9.top_add_26s_26ns_26_2_1_Adder_5_U.facout_s1 ;
wire \add_26s_26ns_26_2_1_U9.top_add_26s_26ns_26_2_1_Adder_5_U.facout_s2 ;
wire [12:0] \add_26s_26ns_26_2_1_U9.top_add_26s_26ns_26_2_1_Adder_5_U.fas_s1 ;
wire [12:0] \add_26s_26ns_26_2_1_U9.top_add_26s_26ns_26_2_1_Adder_5_U.fas_s2 ;
wire \add_26s_26ns_26_2_1_U9.top_add_26s_26ns_26_2_1_Adder_5_U.reset ;
wire [25:0] \add_26s_26ns_26_2_1_U9.top_add_26s_26ns_26_2_1_Adder_5_U.s ;
wire [12:0] \add_26s_26ns_26_2_1_U9.top_add_26s_26ns_26_2_1_Adder_5_U.u1.a ;
wire [12:0] \add_26s_26ns_26_2_1_U9.top_add_26s_26ns_26_2_1_Adder_5_U.u1.b ;
wire \add_26s_26ns_26_2_1_U9.top_add_26s_26ns_26_2_1_Adder_5_U.u1.cin ;
wire \add_26s_26ns_26_2_1_U9.top_add_26s_26ns_26_2_1_Adder_5_U.u1.cout ;
wire [12:0] \add_26s_26ns_26_2_1_U9.top_add_26s_26ns_26_2_1_Adder_5_U.u1.s ;
wire [12:0] \add_26s_26ns_26_2_1_U9.top_add_26s_26ns_26_2_1_Adder_5_U.u2.a ;
wire [12:0] \add_26s_26ns_26_2_1_U9.top_add_26s_26ns_26_2_1_Adder_5_U.u2.b ;
wire \add_26s_26ns_26_2_1_U9.top_add_26s_26ns_26_2_1_Adder_5_U.u2.cin ;
wire \add_26s_26ns_26_2_1_U9.top_add_26s_26ns_26_2_1_Adder_5_U.u2.cout ;
wire [12:0] \add_26s_26ns_26_2_1_U9.top_add_26s_26ns_26_2_1_Adder_5_U.u2.s ;
wire \add_2ns_2ns_2_2_1_U13.ce ;
wire \add_2ns_2ns_2_2_1_U13.clk ;
wire [1:0] \add_2ns_2ns_2_2_1_U13.din0 ;
wire [1:0] \add_2ns_2ns_2_2_1_U13.din1 ;
wire [1:0] \add_2ns_2ns_2_2_1_U13.dout ;
wire \add_2ns_2ns_2_2_1_U13.reset ;
wire [1:0] \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_4_U.a ;
wire [1:0] \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_4_U.ain_s0 ;
wire [1:0] \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_4_U.b ;
wire [1:0] \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_4_U.bin_s0 ;
wire \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_4_U.ce ;
wire \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_4_U.clk ;
wire \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_4_U.facout_s1 ;
wire \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_4_U.facout_s2 ;
wire \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_4_U.fas_s1 ;
wire \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_4_U.fas_s2 ;
wire \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_4_U.reset ;
wire [1:0] \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_4_U.s ;
wire \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_4_U.u1.a ;
wire \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_4_U.u1.b ;
wire \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_4_U.u1.cin ;
wire \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_4_U.u1.cout ;
wire \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_4_U.u1.s ;
wire \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_4_U.u2.a ;
wire \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_4_U.u2.b ;
wire \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_4_U.u2.cin ;
wire \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_4_U.u2.cout ;
wire \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_4_U.u2.s ;
wire \add_2ns_2ns_2_2_1_U19.ce ;
wire \add_2ns_2ns_2_2_1_U19.clk ;
wire [1:0] \add_2ns_2ns_2_2_1_U19.din0 ;
wire [1:0] \add_2ns_2ns_2_2_1_U19.din1 ;
wire [1:0] \add_2ns_2ns_2_2_1_U19.dout ;
wire \add_2ns_2ns_2_2_1_U19.reset ;
wire [1:0] \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_4_U.a ;
wire [1:0] \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_4_U.ain_s0 ;
wire [1:0] \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_4_U.b ;
wire [1:0] \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_4_U.bin_s0 ;
wire \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_4_U.ce ;
wire \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_4_U.clk ;
wire \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_4_U.facout_s1 ;
wire \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_4_U.facout_s2 ;
wire \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_4_U.fas_s1 ;
wire \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_4_U.fas_s2 ;
wire \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_4_U.reset ;
wire [1:0] \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_4_U.s ;
wire \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_4_U.u1.a ;
wire \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_4_U.u1.b ;
wire \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_4_U.u1.cin ;
wire \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_4_U.u1.cout ;
wire \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_4_U.u1.s ;
wire \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_4_U.u2.a ;
wire \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_4_U.u2.b ;
wire \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_4_U.u2.cin ;
wire \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_4_U.u2.cout ;
wire \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_4_U.u2.s ;
wire \add_2ns_2ns_2_2_1_U7.ce ;
wire \add_2ns_2ns_2_2_1_U7.clk ;
wire [1:0] \add_2ns_2ns_2_2_1_U7.din0 ;
wire [1:0] \add_2ns_2ns_2_2_1_U7.din1 ;
wire [1:0] \add_2ns_2ns_2_2_1_U7.dout ;
wire \add_2ns_2ns_2_2_1_U7.reset ;
wire [1:0] \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_4_U.a ;
wire [1:0] \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_4_U.ain_s0 ;
wire [1:0] \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_4_U.b ;
wire [1:0] \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_4_U.bin_s0 ;
wire \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_4_U.ce ;
wire \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_4_U.clk ;
wire \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_4_U.facout_s1 ;
wire \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_4_U.facout_s2 ;
wire \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_4_U.fas_s1 ;
wire \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_4_U.fas_s2 ;
wire \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_4_U.reset ;
wire [1:0] \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_4_U.s ;
wire \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_4_U.u1.a ;
wire \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_4_U.u1.b ;
wire \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_4_U.u1.cin ;
wire \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_4_U.u1.cout ;
wire \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_4_U.u1.s ;
wire \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_4_U.u2.a ;
wire \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_4_U.u2.b ;
wire \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_4_U.u2.cin ;
wire \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_4_U.u2.cout ;
wire \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_4_U.u2.s ;
wire \add_32ns_32ns_32_2_1_U14.ce ;
wire \add_32ns_32ns_32_2_1_U14.clk ;
wire [31:0] \add_32ns_32ns_32_2_1_U14.din0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U14.din1 ;
wire [31:0] \add_32ns_32ns_32_2_1_U14.dout ;
wire \add_32ns_32ns_32_2_1_U14.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.a ;
wire [31:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.b ;
wire [31:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s0 ;
wire \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.ce ;
wire \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.clk ;
wire \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.facout_s1 ;
wire \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.facout_s2 ;
wire [15:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s1 ;
wire [15:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s2 ;
wire \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.b ;
wire \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cin ;
wire \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.b ;
wire \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cin ;
wire \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.s ;
wire \add_32ns_32ns_32_2_1_U20.ce ;
wire \add_32ns_32ns_32_2_1_U20.clk ;
wire [31:0] \add_32ns_32ns_32_2_1_U20.din0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U20.din1 ;
wire [31:0] \add_32ns_32ns_32_2_1_U20.dout ;
wire \add_32ns_32ns_32_2_1_U20.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_7_U.a ;
wire [31:0] \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_7_U.b ;
wire [31:0] \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s0 ;
wire \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_7_U.ce ;
wire \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_7_U.clk ;
wire \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_7_U.facout_s1 ;
wire \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_7_U.facout_s2 ;
wire [15:0] \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s1 ;
wire [15:0] \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s2 ;
wire \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_7_U.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_7_U.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.b ;
wire \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cin ;
wire \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.b ;
wire \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cin ;
wire \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.s ;
wire \add_32ns_32ns_32_2_1_U22.ce ;
wire \add_32ns_32ns_32_2_1_U22.clk ;
wire [31:0] \add_32ns_32ns_32_2_1_U22.din0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U22.din1 ;
wire [31:0] \add_32ns_32ns_32_2_1_U22.dout ;
wire \add_32ns_32ns_32_2_1_U22.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_7_U.a ;
wire [31:0] \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_7_U.b ;
wire [31:0] \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s0 ;
wire \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_7_U.ce ;
wire \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_7_U.clk ;
wire \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_7_U.facout_s1 ;
wire \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_7_U.facout_s2 ;
wire [15:0] \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s1 ;
wire [15:0] \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s2 ;
wire \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_7_U.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_7_U.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.b ;
wire \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cin ;
wire \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.b ;
wire \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cin ;
wire \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.s ;
wire \add_32ns_32ns_32_2_1_U25.ce ;
wire \add_32ns_32ns_32_2_1_U25.clk ;
wire [31:0] \add_32ns_32ns_32_2_1_U25.din0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U25.din1 ;
wire [31:0] \add_32ns_32ns_32_2_1_U25.dout ;
wire \add_32ns_32ns_32_2_1_U25.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_7_U.a ;
wire [31:0] \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_7_U.b ;
wire [31:0] \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s0 ;
wire \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_7_U.ce ;
wire \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_7_U.clk ;
wire \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_7_U.facout_s1 ;
wire \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_7_U.facout_s2 ;
wire [15:0] \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s1 ;
wire [15:0] \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s2 ;
wire \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_7_U.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_7_U.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.b ;
wire \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cin ;
wire \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.b ;
wire \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cin ;
wire \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.s ;
wire \add_32ns_32s_32_2_1_U16.ce ;
wire \add_32ns_32s_32_2_1_U16.clk ;
wire [31:0] \add_32ns_32s_32_2_1_U16.din0 ;
wire [31:0] \add_32ns_32s_32_2_1_U16.din1 ;
wire [31:0] \add_32ns_32s_32_2_1_U16.dout ;
wire \add_32ns_32s_32_2_1_U16.reset ;
wire [31:0] \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.a ;
wire [31:0] \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.ain_s0 ;
wire [31:0] \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.b ;
wire [31:0] \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.bin_s0 ;
wire \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.ce ;
wire \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.clk ;
wire \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.facout_s1 ;
wire \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.facout_s2 ;
wire [15:0] \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.fas_s1 ;
wire [15:0] \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.fas_s2 ;
wire \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.reset ;
wire [31:0] \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.s ;
wire [15:0] \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.u1.a ;
wire [15:0] \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.u1.b ;
wire \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.u1.cin ;
wire \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.u1.cout ;
wire [15:0] \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.u1.s ;
wire [15:0] \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.u2.a ;
wire [15:0] \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.u2.b ;
wire \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.u2.cin ;
wire \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.u2.cout ;
wire [15:0] \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.u2.s ;
wire \add_32ns_32s_32_2_1_U23.ce ;
wire \add_32ns_32s_32_2_1_U23.clk ;
wire [31:0] \add_32ns_32s_32_2_1_U23.din0 ;
wire [31:0] \add_32ns_32s_32_2_1_U23.din1 ;
wire [31:0] \add_32ns_32s_32_2_1_U23.dout ;
wire \add_32ns_32s_32_2_1_U23.reset ;
wire [31:0] \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_9_U.a ;
wire [31:0] \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_9_U.ain_s0 ;
wire [31:0] \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_9_U.b ;
wire [31:0] \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_9_U.bin_s0 ;
wire \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_9_U.ce ;
wire \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_9_U.clk ;
wire \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_9_U.facout_s1 ;
wire \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_9_U.facout_s2 ;
wire [15:0] \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_9_U.fas_s1 ;
wire [15:0] \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_9_U.fas_s2 ;
wire \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_9_U.reset ;
wire [31:0] \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_9_U.s ;
wire [15:0] \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_9_U.u1.a ;
wire [15:0] \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_9_U.u1.b ;
wire \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_9_U.u1.cin ;
wire \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_9_U.u1.cout ;
wire [15:0] \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_9_U.u1.s ;
wire [15:0] \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_9_U.u2.a ;
wire [15:0] \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_9_U.u2.b ;
wire \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_9_U.u2.cin ;
wire \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_9_U.u2.cout ;
wire [15:0] \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_9_U.u2.s ;
wire \add_34s_34s_34_2_1_U12.ce ;
wire \add_34s_34s_34_2_1_U12.clk ;
wire [33:0] \add_34s_34s_34_2_1_U12.din0 ;
wire [33:0] \add_34s_34s_34_2_1_U12.din1 ;
wire [33:0] \add_34s_34s_34_2_1_U12.dout ;
wire \add_34s_34s_34_2_1_U12.reset ;
wire [33:0] \add_34s_34s_34_2_1_U12.top_add_34s_34s_34_2_1_Adder_6_U.a ;
wire [33:0] \add_34s_34s_34_2_1_U12.top_add_34s_34s_34_2_1_Adder_6_U.ain_s0 ;
wire [33:0] \add_34s_34s_34_2_1_U12.top_add_34s_34s_34_2_1_Adder_6_U.b ;
wire [33:0] \add_34s_34s_34_2_1_U12.top_add_34s_34s_34_2_1_Adder_6_U.bin_s0 ;
wire \add_34s_34s_34_2_1_U12.top_add_34s_34s_34_2_1_Adder_6_U.ce ;
wire \add_34s_34s_34_2_1_U12.top_add_34s_34s_34_2_1_Adder_6_U.clk ;
wire \add_34s_34s_34_2_1_U12.top_add_34s_34s_34_2_1_Adder_6_U.facout_s1 ;
wire \add_34s_34s_34_2_1_U12.top_add_34s_34s_34_2_1_Adder_6_U.facout_s2 ;
wire [16:0] \add_34s_34s_34_2_1_U12.top_add_34s_34s_34_2_1_Adder_6_U.fas_s1 ;
wire [16:0] \add_34s_34s_34_2_1_U12.top_add_34s_34s_34_2_1_Adder_6_U.fas_s2 ;
wire \add_34s_34s_34_2_1_U12.top_add_34s_34s_34_2_1_Adder_6_U.reset ;
wire [33:0] \add_34s_34s_34_2_1_U12.top_add_34s_34s_34_2_1_Adder_6_U.s ;
wire [16:0] \add_34s_34s_34_2_1_U12.top_add_34s_34s_34_2_1_Adder_6_U.u1.a ;
wire [16:0] \add_34s_34s_34_2_1_U12.top_add_34s_34s_34_2_1_Adder_6_U.u1.b ;
wire \add_34s_34s_34_2_1_U12.top_add_34s_34s_34_2_1_Adder_6_U.u1.cin ;
wire \add_34s_34s_34_2_1_U12.top_add_34s_34s_34_2_1_Adder_6_U.u1.cout ;
wire [16:0] \add_34s_34s_34_2_1_U12.top_add_34s_34s_34_2_1_Adder_6_U.u1.s ;
wire [16:0] \add_34s_34s_34_2_1_U12.top_add_34s_34s_34_2_1_Adder_6_U.u2.a ;
wire [16:0] \add_34s_34s_34_2_1_U12.top_add_34s_34s_34_2_1_Adder_6_U.u2.b ;
wire \add_34s_34s_34_2_1_U12.top_add_34s_34s_34_2_1_Adder_6_U.u2.cin ;
wire \add_34s_34s_34_2_1_U12.top_add_34s_34s_34_2_1_Adder_6_U.u2.cout ;
wire [16:0] \add_34s_34s_34_2_1_U12.top_add_34s_34s_34_2_1_Adder_6_U.u2.s ;
wire \add_34s_34s_34_2_1_U21.ce ;
wire \add_34s_34s_34_2_1_U21.clk ;
wire [33:0] \add_34s_34s_34_2_1_U21.din0 ;
wire [33:0] \add_34s_34s_34_2_1_U21.din1 ;
wire [33:0] \add_34s_34s_34_2_1_U21.dout ;
wire \add_34s_34s_34_2_1_U21.reset ;
wire [33:0] \add_34s_34s_34_2_1_U21.top_add_34s_34s_34_2_1_Adder_6_U.a ;
wire [33:0] \add_34s_34s_34_2_1_U21.top_add_34s_34s_34_2_1_Adder_6_U.ain_s0 ;
wire [33:0] \add_34s_34s_34_2_1_U21.top_add_34s_34s_34_2_1_Adder_6_U.b ;
wire [33:0] \add_34s_34s_34_2_1_U21.top_add_34s_34s_34_2_1_Adder_6_U.bin_s0 ;
wire \add_34s_34s_34_2_1_U21.top_add_34s_34s_34_2_1_Adder_6_U.ce ;
wire \add_34s_34s_34_2_1_U21.top_add_34s_34s_34_2_1_Adder_6_U.clk ;
wire \add_34s_34s_34_2_1_U21.top_add_34s_34s_34_2_1_Adder_6_U.facout_s1 ;
wire \add_34s_34s_34_2_1_U21.top_add_34s_34s_34_2_1_Adder_6_U.facout_s2 ;
wire [16:0] \add_34s_34s_34_2_1_U21.top_add_34s_34s_34_2_1_Adder_6_U.fas_s1 ;
wire [16:0] \add_34s_34s_34_2_1_U21.top_add_34s_34s_34_2_1_Adder_6_U.fas_s2 ;
wire \add_34s_34s_34_2_1_U21.top_add_34s_34s_34_2_1_Adder_6_U.reset ;
wire [33:0] \add_34s_34s_34_2_1_U21.top_add_34s_34s_34_2_1_Adder_6_U.s ;
wire [16:0] \add_34s_34s_34_2_1_U21.top_add_34s_34s_34_2_1_Adder_6_U.u1.a ;
wire [16:0] \add_34s_34s_34_2_1_U21.top_add_34s_34s_34_2_1_Adder_6_U.u1.b ;
wire \add_34s_34s_34_2_1_U21.top_add_34s_34s_34_2_1_Adder_6_U.u1.cin ;
wire \add_34s_34s_34_2_1_U21.top_add_34s_34s_34_2_1_Adder_6_U.u1.cout ;
wire [16:0] \add_34s_34s_34_2_1_U21.top_add_34s_34s_34_2_1_Adder_6_U.u1.s ;
wire [16:0] \add_34s_34s_34_2_1_U21.top_add_34s_34s_34_2_1_Adder_6_U.u2.a ;
wire [16:0] \add_34s_34s_34_2_1_U21.top_add_34s_34s_34_2_1_Adder_6_U.u2.b ;
wire \add_34s_34s_34_2_1_U21.top_add_34s_34s_34_2_1_Adder_6_U.u2.cin ;
wire \add_34s_34s_34_2_1_U21.top_add_34s_34s_34_2_1_Adder_6_U.u2.cout ;
wire [16:0] \add_34s_34s_34_2_1_U21.top_add_34s_34s_34_2_1_Adder_6_U.u2.s ;
wire \add_34s_34s_34_2_1_U24.ce ;
wire \add_34s_34s_34_2_1_U24.clk ;
wire [33:0] \add_34s_34s_34_2_1_U24.din0 ;
wire [33:0] \add_34s_34s_34_2_1_U24.din1 ;
wire [33:0] \add_34s_34s_34_2_1_U24.dout ;
wire \add_34s_34s_34_2_1_U24.reset ;
wire [33:0] \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_6_U.a ;
wire [33:0] \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_6_U.ain_s0 ;
wire [33:0] \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_6_U.b ;
wire [33:0] \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_6_U.bin_s0 ;
wire \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_6_U.ce ;
wire \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_6_U.clk ;
wire \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_6_U.facout_s1 ;
wire \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_6_U.facout_s2 ;
wire [16:0] \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_6_U.fas_s1 ;
wire [16:0] \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_6_U.fas_s2 ;
wire \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_6_U.reset ;
wire [33:0] \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_6_U.s ;
wire [16:0] \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_6_U.u1.a ;
wire [16:0] \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_6_U.u1.b ;
wire \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_6_U.u1.cin ;
wire \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_6_U.u1.cout ;
wire [16:0] \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_6_U.u1.s ;
wire [16:0] \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_6_U.u2.a ;
wire [16:0] \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_6_U.u2.b ;
wire \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_6_U.u2.cin ;
wire \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_6_U.u2.cout ;
wire [16:0] \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_6_U.u2.s ;
wire \add_37s_37s_37_2_1_U18.ce ;
wire \add_37s_37s_37_2_1_U18.clk ;
wire [36:0] \add_37s_37s_37_2_1_U18.din0 ;
wire [36:0] \add_37s_37s_37_2_1_U18.din1 ;
wire [36:0] \add_37s_37s_37_2_1_U18.dout ;
wire \add_37s_37s_37_2_1_U18.reset ;
wire [36:0] \add_37s_37s_37_2_1_U18.top_add_37s_37s_37_2_1_Adder_11_U.a ;
wire [36:0] \add_37s_37s_37_2_1_U18.top_add_37s_37s_37_2_1_Adder_11_U.ain_s0 ;
wire [36:0] \add_37s_37s_37_2_1_U18.top_add_37s_37s_37_2_1_Adder_11_U.b ;
wire [36:0] \add_37s_37s_37_2_1_U18.top_add_37s_37s_37_2_1_Adder_11_U.bin_s0 ;
wire \add_37s_37s_37_2_1_U18.top_add_37s_37s_37_2_1_Adder_11_U.ce ;
wire \add_37s_37s_37_2_1_U18.top_add_37s_37s_37_2_1_Adder_11_U.clk ;
wire \add_37s_37s_37_2_1_U18.top_add_37s_37s_37_2_1_Adder_11_U.facout_s1 ;
wire \add_37s_37s_37_2_1_U18.top_add_37s_37s_37_2_1_Adder_11_U.facout_s2 ;
wire [17:0] \add_37s_37s_37_2_1_U18.top_add_37s_37s_37_2_1_Adder_11_U.fas_s1 ;
wire [18:0] \add_37s_37s_37_2_1_U18.top_add_37s_37s_37_2_1_Adder_11_U.fas_s2 ;
wire \add_37s_37s_37_2_1_U18.top_add_37s_37s_37_2_1_Adder_11_U.reset ;
wire [36:0] \add_37s_37s_37_2_1_U18.top_add_37s_37s_37_2_1_Adder_11_U.s ;
wire [17:0] \add_37s_37s_37_2_1_U18.top_add_37s_37s_37_2_1_Adder_11_U.u1.a ;
wire [17:0] \add_37s_37s_37_2_1_U18.top_add_37s_37s_37_2_1_Adder_11_U.u1.b ;
wire \add_37s_37s_37_2_1_U18.top_add_37s_37s_37_2_1_Adder_11_U.u1.cin ;
wire \add_37s_37s_37_2_1_U18.top_add_37s_37s_37_2_1_Adder_11_U.u1.cout ;
wire [17:0] \add_37s_37s_37_2_1_U18.top_add_37s_37s_37_2_1_Adder_11_U.u1.s ;
wire [18:0] \add_37s_37s_37_2_1_U18.top_add_37s_37s_37_2_1_Adder_11_U.u2.a ;
wire [18:0] \add_37s_37s_37_2_1_U18.top_add_37s_37s_37_2_1_Adder_11_U.u2.b ;
wire \add_37s_37s_37_2_1_U18.top_add_37s_37s_37_2_1_Adder_11_U.u2.cin ;
wire \add_37s_37s_37_2_1_U18.top_add_37s_37s_37_2_1_Adder_11_U.u2.cout ;
wire [18:0] \add_37s_37s_37_2_1_U18.top_add_37s_37s_37_2_1_Adder_11_U.u2.s ;
wire \add_3s_3ns_3_2_1_U17.ce ;
wire \add_3s_3ns_3_2_1_U17.clk ;
wire [2:0] \add_3s_3ns_3_2_1_U17.din0 ;
wire [2:0] \add_3s_3ns_3_2_1_U17.din1 ;
wire [2:0] \add_3s_3ns_3_2_1_U17.dout ;
wire \add_3s_3ns_3_2_1_U17.reset ;
wire [2:0] \add_3s_3ns_3_2_1_U17.top_add_3s_3ns_3_2_1_Adder_10_U.a ;
wire [2:0] \add_3s_3ns_3_2_1_U17.top_add_3s_3ns_3_2_1_Adder_10_U.ain_s0 ;
wire [2:0] \add_3s_3ns_3_2_1_U17.top_add_3s_3ns_3_2_1_Adder_10_U.b ;
wire [2:0] \add_3s_3ns_3_2_1_U17.top_add_3s_3ns_3_2_1_Adder_10_U.bin_s0 ;
wire \add_3s_3ns_3_2_1_U17.top_add_3s_3ns_3_2_1_Adder_10_U.ce ;
wire \add_3s_3ns_3_2_1_U17.top_add_3s_3ns_3_2_1_Adder_10_U.clk ;
wire \add_3s_3ns_3_2_1_U17.top_add_3s_3ns_3_2_1_Adder_10_U.facout_s1 ;
wire \add_3s_3ns_3_2_1_U17.top_add_3s_3ns_3_2_1_Adder_10_U.facout_s2 ;
wire \add_3s_3ns_3_2_1_U17.top_add_3s_3ns_3_2_1_Adder_10_U.fas_s1 ;
wire [1:0] \add_3s_3ns_3_2_1_U17.top_add_3s_3ns_3_2_1_Adder_10_U.fas_s2 ;
wire \add_3s_3ns_3_2_1_U17.top_add_3s_3ns_3_2_1_Adder_10_U.reset ;
wire [2:0] \add_3s_3ns_3_2_1_U17.top_add_3s_3ns_3_2_1_Adder_10_U.s ;
wire \add_3s_3ns_3_2_1_U17.top_add_3s_3ns_3_2_1_Adder_10_U.u1.a ;
wire \add_3s_3ns_3_2_1_U17.top_add_3s_3ns_3_2_1_Adder_10_U.u1.b ;
wire \add_3s_3ns_3_2_1_U17.top_add_3s_3ns_3_2_1_Adder_10_U.u1.cin ;
wire \add_3s_3ns_3_2_1_U17.top_add_3s_3ns_3_2_1_Adder_10_U.u1.cout ;
wire \add_3s_3ns_3_2_1_U17.top_add_3s_3ns_3_2_1_Adder_10_U.u1.s ;
wire [1:0] \add_3s_3ns_3_2_1_U17.top_add_3s_3ns_3_2_1_Adder_10_U.u2.a ;
wire [1:0] \add_3s_3ns_3_2_1_U17.top_add_3s_3ns_3_2_1_Adder_10_U.u2.b ;
wire \add_3s_3ns_3_2_1_U17.top_add_3s_3ns_3_2_1_Adder_10_U.u2.cin ;
wire \add_3s_3ns_3_2_1_U17.top_add_3s_3ns_3_2_1_Adder_10_U.u2.cout ;
wire [1:0] \add_3s_3ns_3_2_1_U17.top_add_3s_3ns_3_2_1_Adder_10_U.u2.s ;
wire \add_4ns_4ns_4_2_1_U3.ce ;
wire \add_4ns_4ns_4_2_1_U3.clk ;
wire [3:0] \add_4ns_4ns_4_2_1_U3.din0 ;
wire [3:0] \add_4ns_4ns_4_2_1_U3.din1 ;
wire [3:0] \add_4ns_4ns_4_2_1_U3.dout ;
wire \add_4ns_4ns_4_2_1_U3.reset ;
wire [3:0] \add_4ns_4ns_4_2_1_U3.top_add_4ns_4ns_4_2_1_Adder_2_U.a ;
wire [3:0] \add_4ns_4ns_4_2_1_U3.top_add_4ns_4ns_4_2_1_Adder_2_U.ain_s0 ;
wire [3:0] \add_4ns_4ns_4_2_1_U3.top_add_4ns_4ns_4_2_1_Adder_2_U.b ;
wire [3:0] \add_4ns_4ns_4_2_1_U3.top_add_4ns_4ns_4_2_1_Adder_2_U.bin_s0 ;
wire \add_4ns_4ns_4_2_1_U3.top_add_4ns_4ns_4_2_1_Adder_2_U.ce ;
wire \add_4ns_4ns_4_2_1_U3.top_add_4ns_4ns_4_2_1_Adder_2_U.clk ;
wire \add_4ns_4ns_4_2_1_U3.top_add_4ns_4ns_4_2_1_Adder_2_U.facout_s1 ;
wire \add_4ns_4ns_4_2_1_U3.top_add_4ns_4ns_4_2_1_Adder_2_U.facout_s2 ;
wire [1:0] \add_4ns_4ns_4_2_1_U3.top_add_4ns_4ns_4_2_1_Adder_2_U.fas_s1 ;
wire [1:0] \add_4ns_4ns_4_2_1_U3.top_add_4ns_4ns_4_2_1_Adder_2_U.fas_s2 ;
wire \add_4ns_4ns_4_2_1_U3.top_add_4ns_4ns_4_2_1_Adder_2_U.reset ;
wire [3:0] \add_4ns_4ns_4_2_1_U3.top_add_4ns_4ns_4_2_1_Adder_2_U.s ;
wire [1:0] \add_4ns_4ns_4_2_1_U3.top_add_4ns_4ns_4_2_1_Adder_2_U.u1.a ;
wire [1:0] \add_4ns_4ns_4_2_1_U3.top_add_4ns_4ns_4_2_1_Adder_2_U.u1.b ;
wire \add_4ns_4ns_4_2_1_U3.top_add_4ns_4ns_4_2_1_Adder_2_U.u1.cin ;
wire \add_4ns_4ns_4_2_1_U3.top_add_4ns_4ns_4_2_1_Adder_2_U.u1.cout ;
wire [1:0] \add_4ns_4ns_4_2_1_U3.top_add_4ns_4ns_4_2_1_Adder_2_U.u1.s ;
wire [1:0] \add_4ns_4ns_4_2_1_U3.top_add_4ns_4ns_4_2_1_Adder_2_U.u2.a ;
wire [1:0] \add_4ns_4ns_4_2_1_U3.top_add_4ns_4ns_4_2_1_Adder_2_U.u2.b ;
wire \add_4ns_4ns_4_2_1_U3.top_add_4ns_4ns_4_2_1_Adder_2_U.u2.cin ;
wire \add_4ns_4ns_4_2_1_U3.top_add_4ns_4ns_4_2_1_Adder_2_U.u2.cout ;
wire [1:0] \add_4ns_4ns_4_2_1_U3.top_add_4ns_4ns_4_2_1_Adder_2_U.u2.s ;
wire \add_7s_7ns_7_2_1_U10.ce ;
wire \add_7s_7ns_7_2_1_U10.clk ;
wire [6:0] \add_7s_7ns_7_2_1_U10.din0 ;
wire [6:0] \add_7s_7ns_7_2_1_U10.din1 ;
wire [6:0] \add_7s_7ns_7_2_1_U10.dout ;
wire \add_7s_7ns_7_2_1_U10.reset ;
wire [6:0] \add_7s_7ns_7_2_1_U10.top_add_7s_7ns_7_2_1_Adder_3_U.a ;
wire [6:0] \add_7s_7ns_7_2_1_U10.top_add_7s_7ns_7_2_1_Adder_3_U.ain_s0 ;
wire [6:0] \add_7s_7ns_7_2_1_U10.top_add_7s_7ns_7_2_1_Adder_3_U.b ;
wire [6:0] \add_7s_7ns_7_2_1_U10.top_add_7s_7ns_7_2_1_Adder_3_U.bin_s0 ;
wire \add_7s_7ns_7_2_1_U10.top_add_7s_7ns_7_2_1_Adder_3_U.ce ;
wire \add_7s_7ns_7_2_1_U10.top_add_7s_7ns_7_2_1_Adder_3_U.clk ;
wire \add_7s_7ns_7_2_1_U10.top_add_7s_7ns_7_2_1_Adder_3_U.facout_s1 ;
wire \add_7s_7ns_7_2_1_U10.top_add_7s_7ns_7_2_1_Adder_3_U.facout_s2 ;
wire [2:0] \add_7s_7ns_7_2_1_U10.top_add_7s_7ns_7_2_1_Adder_3_U.fas_s1 ;
wire [3:0] \add_7s_7ns_7_2_1_U10.top_add_7s_7ns_7_2_1_Adder_3_U.fas_s2 ;
wire \add_7s_7ns_7_2_1_U10.top_add_7s_7ns_7_2_1_Adder_3_U.reset ;
wire [6:0] \add_7s_7ns_7_2_1_U10.top_add_7s_7ns_7_2_1_Adder_3_U.s ;
wire [2:0] \add_7s_7ns_7_2_1_U10.top_add_7s_7ns_7_2_1_Adder_3_U.u1.a ;
wire [2:0] \add_7s_7ns_7_2_1_U10.top_add_7s_7ns_7_2_1_Adder_3_U.u1.b ;
wire \add_7s_7ns_7_2_1_U10.top_add_7s_7ns_7_2_1_Adder_3_U.u1.cin ;
wire \add_7s_7ns_7_2_1_U10.top_add_7s_7ns_7_2_1_Adder_3_U.u1.cout ;
wire [2:0] \add_7s_7ns_7_2_1_U10.top_add_7s_7ns_7_2_1_Adder_3_U.u1.s ;
wire [3:0] \add_7s_7ns_7_2_1_U10.top_add_7s_7ns_7_2_1_Adder_3_U.u2.a ;
wire [3:0] \add_7s_7ns_7_2_1_U10.top_add_7s_7ns_7_2_1_Adder_3_U.u2.b ;
wire \add_7s_7ns_7_2_1_U10.top_add_7s_7ns_7_2_1_Adder_3_U.u2.cin ;
wire \add_7s_7ns_7_2_1_U10.top_add_7s_7ns_7_2_1_Adder_3_U.u2.cout ;
wire [3:0] \add_7s_7ns_7_2_1_U10.top_add_7s_7ns_7_2_1_Adder_3_U.u2.s ;
wire \add_7s_7ns_7_2_1_U6.ce ;
wire \add_7s_7ns_7_2_1_U6.clk ;
wire [6:0] \add_7s_7ns_7_2_1_U6.din0 ;
wire [6:0] \add_7s_7ns_7_2_1_U6.din1 ;
wire [6:0] \add_7s_7ns_7_2_1_U6.dout ;
wire \add_7s_7ns_7_2_1_U6.reset ;
wire [6:0] \add_7s_7ns_7_2_1_U6.top_add_7s_7ns_7_2_1_Adder_3_U.a ;
wire [6:0] \add_7s_7ns_7_2_1_U6.top_add_7s_7ns_7_2_1_Adder_3_U.ain_s0 ;
wire [6:0] \add_7s_7ns_7_2_1_U6.top_add_7s_7ns_7_2_1_Adder_3_U.b ;
wire [6:0] \add_7s_7ns_7_2_1_U6.top_add_7s_7ns_7_2_1_Adder_3_U.bin_s0 ;
wire \add_7s_7ns_7_2_1_U6.top_add_7s_7ns_7_2_1_Adder_3_U.ce ;
wire \add_7s_7ns_7_2_1_U6.top_add_7s_7ns_7_2_1_Adder_3_U.clk ;
wire \add_7s_7ns_7_2_1_U6.top_add_7s_7ns_7_2_1_Adder_3_U.facout_s1 ;
wire \add_7s_7ns_7_2_1_U6.top_add_7s_7ns_7_2_1_Adder_3_U.facout_s2 ;
wire [2:0] \add_7s_7ns_7_2_1_U6.top_add_7s_7ns_7_2_1_Adder_3_U.fas_s1 ;
wire [3:0] \add_7s_7ns_7_2_1_U6.top_add_7s_7ns_7_2_1_Adder_3_U.fas_s2 ;
wire \add_7s_7ns_7_2_1_U6.top_add_7s_7ns_7_2_1_Adder_3_U.reset ;
wire [6:0] \add_7s_7ns_7_2_1_U6.top_add_7s_7ns_7_2_1_Adder_3_U.s ;
wire [2:0] \add_7s_7ns_7_2_1_U6.top_add_7s_7ns_7_2_1_Adder_3_U.u1.a ;
wire [2:0] \add_7s_7ns_7_2_1_U6.top_add_7s_7ns_7_2_1_Adder_3_U.u1.b ;
wire \add_7s_7ns_7_2_1_U6.top_add_7s_7ns_7_2_1_Adder_3_U.u1.cin ;
wire \add_7s_7ns_7_2_1_U6.top_add_7s_7ns_7_2_1_Adder_3_U.u1.cout ;
wire [2:0] \add_7s_7ns_7_2_1_U6.top_add_7s_7ns_7_2_1_Adder_3_U.u1.s ;
wire [3:0] \add_7s_7ns_7_2_1_U6.top_add_7s_7ns_7_2_1_Adder_3_U.u2.a ;
wire [3:0] \add_7s_7ns_7_2_1_U6.top_add_7s_7ns_7_2_1_Adder_3_U.u2.b ;
wire \add_7s_7ns_7_2_1_U6.top_add_7s_7ns_7_2_1_Adder_3_U.u2.cin ;
wire \add_7s_7ns_7_2_1_U6.top_add_7s_7ns_7_2_1_Adder_3_U.u2.cout ;
wire [3:0] \add_7s_7ns_7_2_1_U6.top_add_7s_7ns_7_2_1_Adder_3_U.u2.s ;
wire \add_8ns_8ns_8_2_1_U1.ce ;
wire \add_8ns_8ns_8_2_1_U1.clk ;
wire [7:0] \add_8ns_8ns_8_2_1_U1.din0 ;
wire [7:0] \add_8ns_8ns_8_2_1_U1.din1 ;
wire [7:0] \add_8ns_8ns_8_2_1_U1.dout ;
wire \add_8ns_8ns_8_2_1_U1.reset ;
wire [7:0] \add_8ns_8ns_8_2_1_U1.top_add_8ns_8ns_8_2_1_Adder_0_U.a ;
wire [7:0] \add_8ns_8ns_8_2_1_U1.top_add_8ns_8ns_8_2_1_Adder_0_U.ain_s0 ;
wire [7:0] \add_8ns_8ns_8_2_1_U1.top_add_8ns_8ns_8_2_1_Adder_0_U.b ;
wire [7:0] \add_8ns_8ns_8_2_1_U1.top_add_8ns_8ns_8_2_1_Adder_0_U.bin_s0 ;
wire \add_8ns_8ns_8_2_1_U1.top_add_8ns_8ns_8_2_1_Adder_0_U.ce ;
wire \add_8ns_8ns_8_2_1_U1.top_add_8ns_8ns_8_2_1_Adder_0_U.clk ;
wire \add_8ns_8ns_8_2_1_U1.top_add_8ns_8ns_8_2_1_Adder_0_U.facout_s1 ;
wire \add_8ns_8ns_8_2_1_U1.top_add_8ns_8ns_8_2_1_Adder_0_U.facout_s2 ;
wire [3:0] \add_8ns_8ns_8_2_1_U1.top_add_8ns_8ns_8_2_1_Adder_0_U.fas_s1 ;
wire [3:0] \add_8ns_8ns_8_2_1_U1.top_add_8ns_8ns_8_2_1_Adder_0_U.fas_s2 ;
wire \add_8ns_8ns_8_2_1_U1.top_add_8ns_8ns_8_2_1_Adder_0_U.reset ;
wire [7:0] \add_8ns_8ns_8_2_1_U1.top_add_8ns_8ns_8_2_1_Adder_0_U.s ;
wire [3:0] \add_8ns_8ns_8_2_1_U1.top_add_8ns_8ns_8_2_1_Adder_0_U.u1.a ;
wire [3:0] \add_8ns_8ns_8_2_1_U1.top_add_8ns_8ns_8_2_1_Adder_0_U.u1.b ;
wire \add_8ns_8ns_8_2_1_U1.top_add_8ns_8ns_8_2_1_Adder_0_U.u1.cin ;
wire \add_8ns_8ns_8_2_1_U1.top_add_8ns_8ns_8_2_1_Adder_0_U.u1.cout ;
wire [3:0] \add_8ns_8ns_8_2_1_U1.top_add_8ns_8ns_8_2_1_Adder_0_U.u1.s ;
wire [3:0] \add_8ns_8ns_8_2_1_U1.top_add_8ns_8ns_8_2_1_Adder_0_U.u2.a ;
wire [3:0] \add_8ns_8ns_8_2_1_U1.top_add_8ns_8ns_8_2_1_Adder_0_U.u2.b ;
wire \add_8ns_8ns_8_2_1_U1.top_add_8ns_8ns_8_2_1_Adder_0_U.u2.cin ;
wire \add_8ns_8ns_8_2_1_U1.top_add_8ns_8ns_8_2_1_Adder_0_U.u2.cout ;
wire [3:0] \add_8ns_8ns_8_2_1_U1.top_add_8ns_8ns_8_2_1_Adder_0_U.u2.s ;
wire and_ln340_fu_1356_p2;
wire and_ln410_fu_1296_p2;
wire and_ln412_fu_709_p2;
wire and_ln414_1_fu_1215_p2;
wire [1:0] and_ln414_fu_1145_p2;
wire and_ln780_fu_880_p2;
wire and_ln781_fu_936_p2;
wire [3:0] and_ln783_fu_1331_p2;
wire and_ln788_1_fu_922_p2;
wire and_ln788_fu_916_p2;
wire [7:0] and_ln_fu_469_p3;
wire ap_CS_fsm_state1;
wire ap_CS_fsm_state12;
wire ap_CS_fsm_state13;
wire ap_CS_fsm_state14;
wire ap_CS_fsm_state15;
wire ap_CS_fsm_state16;
wire ap_CS_fsm_state17;
wire ap_CS_fsm_state18;
wire ap_CS_fsm_state19;
wire ap_CS_fsm_state2;
wire ap_CS_fsm_state20;
wire ap_CS_fsm_state21;
wire ap_CS_fsm_state22;
wire ap_CS_fsm_state23;
wire ap_CS_fsm_state24;
wire ap_CS_fsm_state25;
wire ap_CS_fsm_state26;
wire ap_CS_fsm_state27;
wire ap_CS_fsm_state28;
wire ap_CS_fsm_state29;
wire ap_CS_fsm_state3;
wire ap_CS_fsm_state30;
wire ap_CS_fsm_state31;
wire ap_CS_fsm_state32;
wire ap_CS_fsm_state33;
wire ap_CS_fsm_state34;
wire ap_CS_fsm_state35;
wire ap_CS_fsm_state36;
wire ap_CS_fsm_state37;
wire ap_CS_fsm_state38;
wire ap_CS_fsm_state39;
wire ap_CS_fsm_state4;
wire ap_CS_fsm_state40;
wire ap_CS_fsm_state41;
wire ap_CS_fsm_state42;
wire ap_CS_fsm_state43;
wire ap_CS_fsm_state44;
wire ap_CS_fsm_state45;
wire ap_CS_fsm_state46;
wire ap_CS_fsm_state47;
wire ap_CS_fsm_state48;
wire ap_CS_fsm_state49;
wire ap_CS_fsm_state5;
wire ap_CS_fsm_state6;
wire [48:0] ap_NS_fsm;
wire ap_clk;
wire ap_done;
wire ap_idle;
wire ap_ready;
wire ap_rst;
wire ap_start;
wire \ashr_32s_32s_32_7_1_U4.ce ;
wire \ashr_32s_32s_32_7_1_U4.clk ;
wire [31:0] \ashr_32s_32s_32_7_1_U4.din0 ;
wire [31:0] \ashr_32s_32s_32_7_1_U4.din1 ;
wire [31:0] \ashr_32s_32s_32_7_1_U4.din1_cast ;
wire [31:0] \ashr_32s_32s_32_7_1_U4.din1_mask ;
wire [31:0] \ashr_32s_32s_32_7_1_U4.dout ;
wire \ashr_32s_32s_32_7_1_U4.reset ;
wire carry_1_fu_828_p2;
wire [7:0] conv_i847_fu_365_p0;
wire [31:0] conv_i847_fu_365_p1;
wire deleted_ones_fu_885_p3;
wire deleted_zeros_fu_862_p3;
wire [33:0] grp_fu_1015_p0;
wire [33:0] grp_fu_1015_p1;
wire [33:0] grp_fu_1015_p2;
wire [1:0] grp_fu_1050_p2;
wire [31:0] grp_fu_1055_p2;
wire [6:0] grp_fu_1183_p0;
wire [6:0] grp_fu_1183_p1;
wire [6:0] grp_fu_1183_p2;
wire [31:0] grp_fu_1192_p1;
wire [31:0] grp_fu_1192_p2;
wire [2:0] grp_fu_1234_p0;
wire [2:0] grp_fu_1234_p1;
wire [2:0] grp_fu_1234_p2;
wire [36:0] grp_fu_1262_p0;
wire [36:0] grp_fu_1262_p1;
wire [36:0] grp_fu_1262_p2;
wire [1:0] grp_fu_1323_p1;
wire [1:0] grp_fu_1323_p2;
wire [31:0] grp_fu_1361_p2;
wire [33:0] grp_fu_1449_p0;
wire [33:0] grp_fu_1449_p1;
wire [33:0] grp_fu_1449_p2;
wire [31:0] grp_fu_1465_p2;
wire [31:0] grp_fu_1497_p1;
wire [31:0] grp_fu_1497_p2;
wire [33:0] grp_fu_1516_p0;
wire [33:0] grp_fu_1516_p1;
wire [33:0] grp_fu_1516_p2;
wire [31:0] grp_fu_1532_p2;
wire [7:0] grp_fu_267_p0;
wire [7:0] grp_fu_267_p2;
wire [8:0] grp_fu_346_p1;
wire [8:0] grp_fu_346_p2;
wire [3:0] grp_fu_357_p2;
wire [31:0] grp_fu_368_p1;
wire [31:0] grp_fu_368_p2;
wire [31:0] grp_fu_377_p1;
wire [31:0] grp_fu_377_p2;
wire [6:0] grp_fu_730_p0;
wire [6:0] grp_fu_730_p1;
wire [6:0] grp_fu_730_p2;
wire [1:0] grp_fu_752_p1;
wire [1:0] grp_fu_752_p2;
wire [5:0] grp_fu_774_p2;
wire [25:0] grp_fu_810_p0;
wire [25:0] grp_fu_810_p1;
wire [25:0] grp_fu_810_p2;
wire [6:0] grp_fu_930_p0;
wire [6:0] grp_fu_930_p2;
wire [3:0] grp_fu_996_p1;
wire [3:0] grp_fu_996_p2;
wire icmp_ln414_fu_1167_p2;
wire icmp_ln785_fu_445_p2;
wire icmp_ln786_1_fu_451_p2;
wire icmp_ln786_fu_486_p2;
wire icmp_ln790_fu_463_p2;
wire icmp_ln851_1_fu_1045_p2;
wire icmp_ln851_2_fu_352_p2;
wire icmp_ln851_3_fu_743_p2;
wire icmp_ln851_4_fu_1275_p2;
wire icmp_ln851_fu_261_p2;
wire \mul_4s_2s_6_7_1_U8.ce ;
wire \mul_4s_2s_6_7_1_U8.clk ;
wire [3:0] \mul_4s_2s_6_7_1_U8.din0 ;
wire [1:0] \mul_4s_2s_6_7_1_U8.din1 ;
wire [5:0] \mul_4s_2s_6_7_1_U8.dout ;
wire \mul_4s_2s_6_7_1_U8.reset ;
wire [3:0] \mul_4s_2s_6_7_1_U8.top_mul_4s_2s_6_7_1_Mul_DSP_0_U.a ;
wire [1:0] \mul_4s_2s_6_7_1_U8.top_mul_4s_2s_6_7_1_Mul_DSP_0_U.b ;
wire \mul_4s_2s_6_7_1_U8.top_mul_4s_2s_6_7_1_Mul_DSP_0_U.ce ;
wire \mul_4s_2s_6_7_1_U8.top_mul_4s_2s_6_7_1_Mul_DSP_0_U.clk ;
wire [5:0] \mul_4s_2s_6_7_1_U8.top_mul_4s_2s_6_7_1_Mul_DSP_0_U.p ;
wire [5:0] \mul_4s_2s_6_7_1_U8.top_mul_4s_2s_6_7_1_Mul_DSP_0_U.tmp_product ;
wire neg_src_2_fu_1399_p2;
wire neg_src_4_fu_1336_p3;
wire [7:0] op_0;
wire [15:0] op_1;
wire [1:0] op_11;
wire [3:0] op_12_V_fu_606_p2;
wire [21:0] op_13_V_fu_780_p3;
wire [1:0] op_14_V_fu_968_p3;
wire [7:0] op_16_V_fu_1240_p3;
wire [1:0] op_17_V_fu_1409_p3;
wire [1:0] op_18;
wire [3:0] op_19_V_fu_1393_p3;
wire [31:0] op_27;
wire op_27_ap_vld;
wire [7:0] op_2_V_fu_529_p3;
wire [7:0] op_4;
wire [3:0] op_5;
wire [1:0] op_6;
wire [2:0] op_8_V_fu_679_p3;
wire [3:0] or_ln1195_1_fu_643_p1;
wire [3:0] or_ln1195_1_fu_643_p2;
wire [4:0] or_ln1195_fu_629_p2;
wire or_ln384_1_fu_956_p2;
wire or_ln384_fu_506_p2;
wire or_ln410_fu_1291_p2;
wire or_ln412_fu_703_p2;
wire or_ln785_fu_897_p2;
wire or_ln788_1_fu_496_p2;
wire or_ln788_2_fu_940_p2;
wire or_ln788_fu_492_p2;
wire [7:0] or_ln_fu_437_p4;
wire overflow_1_fu_907_p2;
wire overflow_fu_481_p2;
wire [3:0] p_Result_12_fu_1383_p4;
wire p_Result_16_fu_686_p3;
wire p_Result_18_fu_974_p3;
wire p_Result_19_fu_1109_p3;
wire [3:0] p_Result_1_fu_1268_p3;
wire p_Result_20_fu_1416_p3;
wire p_Result_21_fu_1470_p3;
wire p_Result_22_fu_1537_p3;
wire p_Result_25_fu_1281_p3;
wire [3:0] p_Result_29_fu_649_p1;
wire p_Result_2_fu_1060_p3;
wire [3:0] p_Result_30_fu_693_p1;
wire p_Result_30_fu_693_p3;
wire p_Result_31_fu_816_p3;
wire [19:0] p_Result_3_fu_736_p3;
wire p_Result_4_fu_383_p3;
wire [6:0] p_Result_5_fu_456_p3;
wire p_Result_s_fu_286_p3;
wire [2:0] p_Val2_7_fu_1374_p2;
wire [7:0] p_Val2_s_fu_514_p3;
wire r_1_fu_700_p1;
wire [3:0] r_V_2_fu_1086_p1;
wire [3:0] r_V_2_fu_1086_p2;
wire r_fu_1288_p1;
wire [1:0] ret_V_19_fu_1072_p3;
wire [15:0] ret_V_20_fu_324_p2;
wire [3:0] ret_V_21_fu_395_p3;
wire [31:0] ret_V_24_fu_1125_p3;
wire [31:0] ret_V_27_fu_1486_p3;
wire [7:0] ret_V_2_fu_298_p3;
wire [6:0] ret_V_5_fu_581_p2;
wire [1:0] ret_fu_547_p2;
wire [35:0] rhs_10_fu_1251_p3;
wire [32:0] rhs_11_fu_1438_p3;
wire [32:0] rhs_13_fu_1505_p3;
wire rhs_1_fu_281_p2;
wire [8:0] rhs_2_fu_313_p3;
wire [4:0] rhs_5_fu_611_p3;
wire [5:0] rhs_7_fu_719_p3;
wire [24:0] rhs_8_fu_799_p3;
wire [6:0] rhs_fu_574_p3;
wire [1:0] select_ln1118_1_fu_1135_p3;
wire [3:0] select_ln1118_fu_1079_p3;
wire [1:0] select_ln1345_fu_540_p3;
wire [31:0] select_ln1497_fu_402_p3;
wire select_ln340_2_fu_1349_p3;
wire select_ln340_fu_1403_p3;
wire [31:0] select_ln353_2_fu_1428_p3;
wire [6:0] select_ln353_fu_986_p3;
wire [7:0] select_ln384_1_fu_522_p3;
wire [1:0] select_ln384_fu_961_p3;
wire [1:0] select_ln850_1_fu_1067_p3;
wire [3:0] select_ln850_2_fu_390_p3;
wire [31:0] select_ln850_4_fu_1119_p3;
wire [6:0] select_ln850_5_fu_981_p3;
wire [31:0] select_ln850_6_fu_1480_p3;
wire [31:0] select_ln850_7_fu_1547_p3;
wire [31:0] select_ln850_8_fu_1423_p3;
wire [7:0] select_ln850_fu_293_p3;
wire [3:0] sext_ln1193_fu_1173_p0;
wire [3:0] sext_ln1195_fu_625_p0;
wire [4:0] sext_ln1195_fu_625_p1;
wire [3:0] sext_ln367_fu_1379_p1;
wire [12:0] sext_ln727_fu_557_p1;
wire [3:0] sext_ln745_fu_1328_p1;
wire [6:0] sext_ln850_fu_927_p1;
wire \shl_32s_32s_32_7_1_U5.ce ;
wire \shl_32s_32s_32_7_1_U5.clk ;
wire [31:0] \shl_32s_32s_32_7_1_U5.din0 ;
wire [31:0] \shl_32s_32s_32_7_1_U5.din1 ;
wire [31:0] \shl_32s_32s_32_7_1_U5.din1_cast ;
wire [31:0] \shl_32s_32s_32_7_1_U5.din1_mask ;
wire [31:0] \shl_32s_32s_32_7_1_U5.dout ;
wire \shl_32s_32s_32_7_1_U5.reset ;
wire \shl_4s_1ns_4_7_1_U11.ce ;
wire \shl_4s_1ns_4_7_1_U11.clk ;
wire [3:0] \shl_4s_1ns_4_7_1_U11.din0 ;
wire [3:0] \shl_4s_1ns_4_7_1_U11.din1 ;
wire \shl_4s_1ns_4_7_1_U11.din1_cast ;
wire \shl_4s_1ns_4_7_1_U11.din1_mask ;
wire [3:0] \shl_4s_1ns_4_7_1_U11.dout ;
wire \shl_4s_1ns_4_7_1_U11.reset ;
wire [12:0] shl_ln728_1_fu_560_p3;
wire [5:0] shl_ln728_5_fu_586_p3;
wire [7:0] shl_ln_fu_273_p1;
wire [15:0] shl_ln_fu_273_p3;
wire signbit_fu_597_p2;
wire \sub_7s_7ns_7_2_1_U15.ce ;
wire \sub_7s_7ns_7_2_1_U15.clk ;
wire [6:0] \sub_7s_7ns_7_2_1_U15.din0 ;
wire [6:0] \sub_7s_7ns_7_2_1_U15.din1 ;
wire [6:0] \sub_7s_7ns_7_2_1_U15.dout ;
wire \sub_7s_7ns_7_2_1_U15.reset ;
wire [6:0] \sub_7s_7ns_7_2_1_U15.top_sub_7s_7ns_7_2_1_Adder_8_U.a ;
wire [6:0] \sub_7s_7ns_7_2_1_U15.top_sub_7s_7ns_7_2_1_Adder_8_U.ain_s0 ;
wire [6:0] \sub_7s_7ns_7_2_1_U15.top_sub_7s_7ns_7_2_1_Adder_8_U.b ;
wire [6:0] \sub_7s_7ns_7_2_1_U15.top_sub_7s_7ns_7_2_1_Adder_8_U.bin_s0 ;
wire \sub_7s_7ns_7_2_1_U15.top_sub_7s_7ns_7_2_1_Adder_8_U.ce ;
wire \sub_7s_7ns_7_2_1_U15.top_sub_7s_7ns_7_2_1_Adder_8_U.clk ;
wire \sub_7s_7ns_7_2_1_U15.top_sub_7s_7ns_7_2_1_Adder_8_U.facout_s1 ;
wire \sub_7s_7ns_7_2_1_U15.top_sub_7s_7ns_7_2_1_Adder_8_U.facout_s2 ;
wire [2:0] \sub_7s_7ns_7_2_1_U15.top_sub_7s_7ns_7_2_1_Adder_8_U.fas_s1 ;
wire [3:0] \sub_7s_7ns_7_2_1_U15.top_sub_7s_7ns_7_2_1_Adder_8_U.fas_s2 ;
wire \sub_7s_7ns_7_2_1_U15.top_sub_7s_7ns_7_2_1_Adder_8_U.reset ;
wire [6:0] \sub_7s_7ns_7_2_1_U15.top_sub_7s_7ns_7_2_1_Adder_8_U.s ;
wire [2:0] \sub_7s_7ns_7_2_1_U15.top_sub_7s_7ns_7_2_1_Adder_8_U.u1.a ;
wire [2:0] \sub_7s_7ns_7_2_1_U15.top_sub_7s_7ns_7_2_1_Adder_8_U.u1.b ;
wire \sub_7s_7ns_7_2_1_U15.top_sub_7s_7ns_7_2_1_Adder_8_U.u1.cin ;
wire \sub_7s_7ns_7_2_1_U15.top_sub_7s_7ns_7_2_1_Adder_8_U.u1.cout ;
wire [2:0] \sub_7s_7ns_7_2_1_U15.top_sub_7s_7ns_7_2_1_Adder_8_U.u1.s ;
wire [3:0] \sub_7s_7ns_7_2_1_U15.top_sub_7s_7ns_7_2_1_Adder_8_U.u2.a ;
wire [3:0] \sub_7s_7ns_7_2_1_U15.top_sub_7s_7ns_7_2_1_Adder_8_U.u2.b ;
wire \sub_7s_7ns_7_2_1_U15.top_sub_7s_7ns_7_2_1_Adder_8_U.u2.cin ;
wire \sub_7s_7ns_7_2_1_U15.top_sub_7s_7ns_7_2_1_Adder_8_U.u2.cout ;
wire [3:0] \sub_7s_7ns_7_2_1_U15.top_sub_7s_7ns_7_2_1_Adder_8_U.u2.s ;
wire \sub_9ns_9s_9_2_1_U2.ce ;
wire \sub_9ns_9s_9_2_1_U2.clk ;
wire [8:0] \sub_9ns_9s_9_2_1_U2.din0 ;
wire [8:0] \sub_9ns_9s_9_2_1_U2.din1 ;
wire [8:0] \sub_9ns_9s_9_2_1_U2.dout ;
wire \sub_9ns_9s_9_2_1_U2.reset ;
wire [8:0] \sub_9ns_9s_9_2_1_U2.top_sub_9ns_9s_9_2_1_Adder_1_U.a ;
wire [8:0] \sub_9ns_9s_9_2_1_U2.top_sub_9ns_9s_9_2_1_Adder_1_U.ain_s0 ;
wire [8:0] \sub_9ns_9s_9_2_1_U2.top_sub_9ns_9s_9_2_1_Adder_1_U.b ;
wire [8:0] \sub_9ns_9s_9_2_1_U2.top_sub_9ns_9s_9_2_1_Adder_1_U.bin_s0 ;
wire \sub_9ns_9s_9_2_1_U2.top_sub_9ns_9s_9_2_1_Adder_1_U.ce ;
wire \sub_9ns_9s_9_2_1_U2.top_sub_9ns_9s_9_2_1_Adder_1_U.clk ;
wire \sub_9ns_9s_9_2_1_U2.top_sub_9ns_9s_9_2_1_Adder_1_U.facout_s1 ;
wire \sub_9ns_9s_9_2_1_U2.top_sub_9ns_9s_9_2_1_Adder_1_U.facout_s2 ;
wire [3:0] \sub_9ns_9s_9_2_1_U2.top_sub_9ns_9s_9_2_1_Adder_1_U.fas_s1 ;
wire [4:0] \sub_9ns_9s_9_2_1_U2.top_sub_9ns_9s_9_2_1_Adder_1_U.fas_s2 ;
wire \sub_9ns_9s_9_2_1_U2.top_sub_9ns_9s_9_2_1_Adder_1_U.reset ;
wire [8:0] \sub_9ns_9s_9_2_1_U2.top_sub_9ns_9s_9_2_1_Adder_1_U.s ;
wire [3:0] \sub_9ns_9s_9_2_1_U2.top_sub_9ns_9s_9_2_1_Adder_1_U.u1.a ;
wire [3:0] \sub_9ns_9s_9_2_1_U2.top_sub_9ns_9s_9_2_1_Adder_1_U.u1.b ;
wire \sub_9ns_9s_9_2_1_U2.top_sub_9ns_9s_9_2_1_Adder_1_U.u1.cin ;
wire \sub_9ns_9s_9_2_1_U2.top_sub_9ns_9s_9_2_1_Adder_1_U.u1.cout ;
wire [3:0] \sub_9ns_9s_9_2_1_U2.top_sub_9ns_9s_9_2_1_Adder_1_U.u1.s ;
wire [4:0] \sub_9ns_9s_9_2_1_U2.top_sub_9ns_9s_9_2_1_Adder_1_U.u2.a ;
wire [4:0] \sub_9ns_9s_9_2_1_U2.top_sub_9ns_9s_9_2_1_Adder_1_U.u2.b ;
wire \sub_9ns_9s_9_2_1_U2.top_sub_9ns_9s_9_2_1_Adder_1_U.u2.cin ;
wire \sub_9ns_9s_9_2_1_U2.top_sub_9ns_9s_9_2_1_Adder_1_U.u2.cout ;
wire [4:0] \sub_9ns_9s_9_2_1_U2.top_sub_9ns_9s_9_2_1_Adder_1_U.u2.s ;
wire tmp_13_fu_1151_p3;
wire tmp_24_fu_867_p3;
wire [7:0] tmp_26_fu_1004_p3;
wire [1:0] tmp_3_fu_1159_p3;
wire [1:0] tmp_9_fu_834_p3;
wire [3:0] trunc_ln1118_fu_1132_p0;
wire [1:0] trunc_ln1118_fu_1132_p1;
wire [3:0] trunc_ln1195_1_fu_618_p3;
wire trunc_ln1195_fu_553_p1;
wire [3:0] trunc_ln1349_fu_602_p1;
wire trunc_ln718_fu_1142_p1;
wire [2:0] trunc_ln731_fu_511_p1;
wire trunc_ln790_1_fu_913_p1;
wire [1:0] trunc_ln790_fu_433_p1;
wire [2:0] trunc_ln851_1_fu_1031_p1;
wire [7:0] trunc_ln851_2_fu_339_p1;
wire [4:0] trunc_ln851_3_fu_675_p1;
wire trunc_ln851_4_fu_1116_p1;
wire [2:0] trunc_ln851_5_fu_1219_p1;
wire trunc_ln851_6_fu_1477_p1;
wire trunc_ln851_7_fu_1544_p1;
wire [7:0] trunc_ln851_fu_257_p1;
wire [6:0] trunc_ln8_fu_536_p1;
wire underflow_1_fu_951_p2;
wire underflow_fu_501_p2;
wire ush_fu_568_p2;
wire xor_ln410_fu_1223_p2;
wire xor_ln416_fu_823_p2;
wire xor_ln780_fu_874_p2;
wire xor_ln785_1_fu_1344_p2;
wire xor_ln785_2_fu_891_p2;
wire xor_ln785_3_fu_902_p2;
wire xor_ln785_fu_476_p2;
wire xor_ln788_fu_945_p2;
wire [15:0] zext_ln1196_fu_320_p1;
wire [7:0] zext_ln1499_fu_593_p1;


assign _0103_ = icmp_ln851_4_reg_2133 & ap_CS_fsm[35];
assign _0104_ = icmp_ln851_3_reg_1848 & ap_CS_fsm[23];
assign _0105_ = ap_CS_fsm[11] & _0110_;
assign _0106_ = ap_CS_fsm[11] & tmp_reg_1603;
assign _0107_ = ap_CS_fsm[4] & tmp_reg_1603;
assign _0108_ = _0111_ & ap_CS_fsm[0];
assign _0109_ = ap_start & ap_CS_fsm[0];
assign and_ln340_fu_1356_p2 = select_ln340_2_fu_1349_p3 & p_Result_28_reg_2149;
assign and_ln410_fu_1296_p2 = r_V_1_reg_2070[1] & or_ln410_fu_1291_p2;
assign and_ln412_fu_709_p2 = op_5[1] & or_ln412_fu_703_p2;
assign and_ln414_1_fu_1215_p2 = p_Result_27_reg_2034 & icmp_ln414_reg_2050;
assign and_ln414_fu_1145_p2 = op_5[1:0] & select_ln1118_1_fu_1135_p3;
assign and_ln780_fu_880_p2 = xor_ln780_fu_874_p2 & Range2_all_ones_reg_1800;
assign and_ln781_fu_936_p2 = carry_1_reg_1896 & Range1_all_ones_reg_1903;
assign and_ln783_fu_1331_p2 = { p_Val2_6_reg_2143[2], p_Val2_6_reg_2143 } & r_V_2_reg_2028;
assign and_ln788_1_fu_922_p2 = p_Result_32_reg_1879 & and_ln788_fu_916_p2;
assign and_ln788_fu_916_p2 = p_Val2_9_reg_1873[0] & deleted_ones_fu_885_p3;
assign carry_1_fu_828_p2 = xor_ln416_fu_823_p2 & or_ln1195_1_reg_1806[3];
assign neg_src_2_fu_1399_p2 = p_Result_26_reg_2187 & p_Result_24_reg_2076;
assign overflow_1_fu_907_p2 = xor_ln785_3_fu_902_p2 & or_ln785_fu_897_p2;
assign overflow_fu_481_p2 = xor_ln785_fu_476_p2 & icmp_ln785_reg_1705;
assign r_V_2_fu_1086_p2 = select_ln1118_fu_1079_p3 & op_5;
assign ret_V_5_fu_581_p2 = trunc_ln8_reg_1747 & { op_6, 5'h00 };
assign ret_fu_547_p2 = select_ln1345_fu_540_p3 & op_6;
assign underflow_1_fu_951_p2 = xor_ln788_fu_945_p2 & p_Result_29_reg_1812;
assign underflow_fu_501_p2 = p_Result_23_reg_1682 & or_ln788_1_fu_496_p2;
assign xor_ln785_1_fu_1344_p2 = ~ p_Result_27_reg_2034;
assign xor_ln780_fu_874_p2 = ~ or_ln1195_reg_1794[4];
assign xor_ln416_fu_823_p2 = ~ p_Result_32_reg_1879;
assign xor_ln788_fu_945_p2 = ~ or_ln788_2_fu_940_p2;
assign xor_ln785_2_fu_891_p2 = ~ deleted_zeros_fu_862_p3;
assign xor_ln785_3_fu_902_p2 = ~ p_Result_29_reg_1812;
assign xor_ln785_fu_476_p2 = ~ p_Result_23_reg_1682;
assign xor_ln410_fu_1223_p2 = ~ p_Result_24_reg_2076;
assign p_Val2_7_fu_1374_p2 = ~ p_Val2_6_reg_2143;
assign _0110_ = ~ tmp_reg_1603;
assign _0111_ = ~ ap_start;
assign _0112_ = { Range2_all_ones_reg_1800, tmp_23_reg_1823 } == 2'h3;
assign _0113_ = ! { Range2_all_ones_reg_1800, tmp_23_reg_1823 };
assign _0114_ = ! { tmp_4_reg_1688, 7'h00 };
assign _0115_ = ! { trunc_ln790_reg_1700, 5'h00 };
assign _0116_ = ! trunc_ln851_1_reg_1991;
assign _0117_ = ! trunc_ln851_2_reg_1620;
assign _0118_ = ! op_1[7:0];
assign _0119_ = { op_2_V_reg_1741[7], op_2_V_reg_1741[7], op_2_V_reg_1741[7], op_2_V_reg_1741[7], op_2_V_reg_1741[7], op_2_V_reg_1741 } == { op_4, 5'h00 };
always @(posedge \add_26s_26ns_26_2_1_U9.top_add_26s_26ns_26_2_1_Adder_5_U.clk )
\add_26s_26ns_26_2_1_U9.top_add_26s_26ns_26_2_1_Adder_5_U.bin_s1  <= _0121_;
always @(posedge \add_26s_26ns_26_2_1_U9.top_add_26s_26ns_26_2_1_Adder_5_U.clk )
\add_26s_26ns_26_2_1_U9.top_add_26s_26ns_26_2_1_Adder_5_U.ain_s1  <= _0120_;
always @(posedge \add_26s_26ns_26_2_1_U9.top_add_26s_26ns_26_2_1_Adder_5_U.clk )
\add_26s_26ns_26_2_1_U9.top_add_26s_26ns_26_2_1_Adder_5_U.sum_s1  <= _0123_;
always @(posedge \add_26s_26ns_26_2_1_U9.top_add_26s_26ns_26_2_1_Adder_5_U.clk )
\add_26s_26ns_26_2_1_U9.top_add_26s_26ns_26_2_1_Adder_5_U.carry_s1  <= _0122_;
assign _0121_ = \add_26s_26ns_26_2_1_U9.top_add_26s_26ns_26_2_1_Adder_5_U.ce  ? \add_26s_26ns_26_2_1_U9.top_add_26s_26ns_26_2_1_Adder_5_U.b [25:13] : \add_26s_26ns_26_2_1_U9.top_add_26s_26ns_26_2_1_Adder_5_U.bin_s1 ;
assign _0120_ = \add_26s_26ns_26_2_1_U9.top_add_26s_26ns_26_2_1_Adder_5_U.ce  ? \add_26s_26ns_26_2_1_U9.top_add_26s_26ns_26_2_1_Adder_5_U.a [25:13] : \add_26s_26ns_26_2_1_U9.top_add_26s_26ns_26_2_1_Adder_5_U.ain_s1 ;
assign _0122_ = \add_26s_26ns_26_2_1_U9.top_add_26s_26ns_26_2_1_Adder_5_U.ce  ? \add_26s_26ns_26_2_1_U9.top_add_26s_26ns_26_2_1_Adder_5_U.facout_s1  : \add_26s_26ns_26_2_1_U9.top_add_26s_26ns_26_2_1_Adder_5_U.carry_s1 ;
assign _0123_ = \add_26s_26ns_26_2_1_U9.top_add_26s_26ns_26_2_1_Adder_5_U.ce  ? \add_26s_26ns_26_2_1_U9.top_add_26s_26ns_26_2_1_Adder_5_U.fas_s1  : \add_26s_26ns_26_2_1_U9.top_add_26s_26ns_26_2_1_Adder_5_U.sum_s1 ;
assign _0124_ = \add_26s_26ns_26_2_1_U9.top_add_26s_26ns_26_2_1_Adder_5_U.u1.a  + \add_26s_26ns_26_2_1_U9.top_add_26s_26ns_26_2_1_Adder_5_U.u1.b ;
assign { \add_26s_26ns_26_2_1_U9.top_add_26s_26ns_26_2_1_Adder_5_U.u1.cout , \add_26s_26ns_26_2_1_U9.top_add_26s_26ns_26_2_1_Adder_5_U.u1.s  } = _0124_ + \add_26s_26ns_26_2_1_U9.top_add_26s_26ns_26_2_1_Adder_5_U.u1.cin ;
assign _0125_ = \add_26s_26ns_26_2_1_U9.top_add_26s_26ns_26_2_1_Adder_5_U.u2.a  + \add_26s_26ns_26_2_1_U9.top_add_26s_26ns_26_2_1_Adder_5_U.u2.b ;
assign { \add_26s_26ns_26_2_1_U9.top_add_26s_26ns_26_2_1_Adder_5_U.u2.cout , \add_26s_26ns_26_2_1_U9.top_add_26s_26ns_26_2_1_Adder_5_U.u2.s  } = _0125_ + \add_26s_26ns_26_2_1_U9.top_add_26s_26ns_26_2_1_Adder_5_U.u2.cin ;
always @(posedge \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_4_U.clk )
\add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_4_U.bin_s1  <= _0127_;
always @(posedge \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_4_U.clk )
\add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_4_U.ain_s1  <= _0126_;
always @(posedge \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_4_U.clk )
\add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_4_U.sum_s1  <= _0129_;
always @(posedge \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_4_U.clk )
\add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_4_U.carry_s1  <= _0128_;
assign _0127_ = \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_4_U.ce  ? \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_4_U.b [1] : \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_4_U.bin_s1 ;
assign _0126_ = \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_4_U.ce  ? \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_4_U.a [1] : \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_4_U.ain_s1 ;
assign _0128_ = \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_4_U.ce  ? \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_4_U.facout_s1  : \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_4_U.carry_s1 ;
assign _0129_ = \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_4_U.ce  ? \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_4_U.fas_s1  : \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_4_U.sum_s1 ;
assign _0130_ = \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_4_U.u1.a  + \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_4_U.u1.b ;
assign { \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_4_U.u1.cout , \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_4_U.u1.s  } = _0130_ + \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_4_U.u1.cin ;
assign _0131_ = \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_4_U.u2.a  + \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_4_U.u2.b ;
assign { \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_4_U.u2.cout , \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_4_U.u2.s  } = _0131_ + \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_4_U.u2.cin ;
always @(posedge \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_4_U.clk )
\add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_4_U.bin_s1  <= _0133_;
always @(posedge \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_4_U.clk )
\add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_4_U.ain_s1  <= _0132_;
always @(posedge \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_4_U.clk )
\add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_4_U.sum_s1  <= _0135_;
always @(posedge \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_4_U.clk )
\add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_4_U.carry_s1  <= _0134_;
assign _0133_ = \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_4_U.ce  ? \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_4_U.b [1] : \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_4_U.bin_s1 ;
assign _0132_ = \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_4_U.ce  ? \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_4_U.a [1] : \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_4_U.ain_s1 ;
assign _0134_ = \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_4_U.ce  ? \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_4_U.facout_s1  : \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_4_U.carry_s1 ;
assign _0135_ = \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_4_U.ce  ? \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_4_U.fas_s1  : \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_4_U.sum_s1 ;
assign _0136_ = \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_4_U.u1.a  + \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_4_U.u1.b ;
assign { \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_4_U.u1.cout , \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_4_U.u1.s  } = _0136_ + \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_4_U.u1.cin ;
assign _0137_ = \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_4_U.u2.a  + \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_4_U.u2.b ;
assign { \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_4_U.u2.cout , \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_4_U.u2.s  } = _0137_ + \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_4_U.u2.cin ;
always @(posedge \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_4_U.clk )
\add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_4_U.bin_s1  <= _0139_;
always @(posedge \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_4_U.clk )
\add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_4_U.ain_s1  <= _0138_;
always @(posedge \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_4_U.clk )
\add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_4_U.sum_s1  <= _0141_;
always @(posedge \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_4_U.clk )
\add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_4_U.carry_s1  <= _0140_;
assign _0139_ = \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_4_U.ce  ? \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_4_U.b [1] : \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_4_U.bin_s1 ;
assign _0138_ = \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_4_U.ce  ? \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_4_U.a [1] : \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_4_U.ain_s1 ;
assign _0140_ = \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_4_U.ce  ? \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_4_U.facout_s1  : \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_4_U.carry_s1 ;
assign _0141_ = \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_4_U.ce  ? \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_4_U.fas_s1  : \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_4_U.sum_s1 ;
assign _0142_ = \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_4_U.u1.a  + \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_4_U.u1.b ;
assign { \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_4_U.u1.cout , \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_4_U.u1.s  } = _0142_ + \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_4_U.u1.cin ;
assign _0143_ = \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_4_U.u2.a  + \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_4_U.u2.b ;
assign { \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_4_U.u2.cout , \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_4_U.u2.s  } = _0143_ + \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_4_U.u2.cin ;
always @(posedge \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.clk )
\add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s1  <= _0145_;
always @(posedge \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.clk )
\add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s1  <= _0144_;
always @(posedge \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.clk )
\add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.sum_s1  <= _0147_;
always @(posedge \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.clk )
\add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.carry_s1  <= _0146_;
assign _0145_ = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.ce  ? \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.b [31:16] : \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s1 ;
assign _0144_ = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.ce  ? \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.a [31:16] : \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s1 ;
assign _0146_ = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.ce  ? \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.facout_s1  : \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.carry_s1 ;
assign _0147_ = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.ce  ? \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s1  : \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.sum_s1 ;
assign _0148_ = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.a  + \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.b ;
assign { \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cout , \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.s  } = _0148_ + \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cin ;
assign _0149_ = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.a  + \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.b ;
assign { \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cout , \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.s  } = _0149_ + \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cin ;
always @(posedge \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_7_U.clk )
\add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s1  <= _0151_;
always @(posedge \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_7_U.clk )
\add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s1  <= _0150_;
always @(posedge \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_7_U.clk )
\add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_7_U.sum_s1  <= _0153_;
always @(posedge \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_7_U.clk )
\add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_7_U.carry_s1  <= _0152_;
assign _0151_ = \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_7_U.ce  ? \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_7_U.b [31:16] : \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s1 ;
assign _0150_ = \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_7_U.ce  ? \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_7_U.a [31:16] : \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s1 ;
assign _0152_ = \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_7_U.ce  ? \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_7_U.facout_s1  : \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_7_U.carry_s1 ;
assign _0153_ = \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_7_U.ce  ? \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s1  : \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_7_U.sum_s1 ;
assign _0154_ = \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.a  + \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.b ;
assign { \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cout , \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.s  } = _0154_ + \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cin ;
assign _0155_ = \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.a  + \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.b ;
assign { \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cout , \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.s  } = _0155_ + \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cin ;
always @(posedge \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_7_U.clk )
\add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s1  <= _0157_;
always @(posedge \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_7_U.clk )
\add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s1  <= _0156_;
always @(posedge \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_7_U.clk )
\add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_7_U.sum_s1  <= _0159_;
always @(posedge \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_7_U.clk )
\add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_7_U.carry_s1  <= _0158_;
assign _0157_ = \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_7_U.ce  ? \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_7_U.b [31:16] : \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s1 ;
assign _0156_ = \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_7_U.ce  ? \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_7_U.a [31:16] : \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s1 ;
assign _0158_ = \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_7_U.ce  ? \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_7_U.facout_s1  : \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_7_U.carry_s1 ;
assign _0159_ = \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_7_U.ce  ? \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s1  : \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_7_U.sum_s1 ;
assign _0160_ = \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.a  + \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.b ;
assign { \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cout , \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.s  } = _0160_ + \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cin ;
assign _0161_ = \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.a  + \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.b ;
assign { \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cout , \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.s  } = _0161_ + \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cin ;
always @(posedge \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_7_U.clk )
\add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s1  <= _0163_;
always @(posedge \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_7_U.clk )
\add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s1  <= _0162_;
always @(posedge \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_7_U.clk )
\add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_7_U.sum_s1  <= _0165_;
always @(posedge \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_7_U.clk )
\add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_7_U.carry_s1  <= _0164_;
assign _0163_ = \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_7_U.ce  ? \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_7_U.b [31:16] : \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s1 ;
assign _0162_ = \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_7_U.ce  ? \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_7_U.a [31:16] : \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s1 ;
assign _0164_ = \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_7_U.ce  ? \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_7_U.facout_s1  : \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_7_U.carry_s1 ;
assign _0165_ = \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_7_U.ce  ? \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s1  : \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_7_U.sum_s1 ;
assign _0166_ = \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.a  + \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.b ;
assign { \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cout , \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.s  } = _0166_ + \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cin ;
assign _0167_ = \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.a  + \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.b ;
assign { \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cout , \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.s  } = _0167_ + \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cin ;
always @(posedge \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.clk )
\add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.bin_s1  <= _0169_;
always @(posedge \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.clk )
\add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.ain_s1  <= _0168_;
always @(posedge \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.clk )
\add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.sum_s1  <= _0171_;
always @(posedge \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.clk )
\add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.carry_s1  <= _0170_;
assign _0169_ = \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.ce  ? \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.b [31:16] : \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.bin_s1 ;
assign _0168_ = \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.ce  ? \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.a [31:16] : \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.ain_s1 ;
assign _0170_ = \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.ce  ? \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.facout_s1  : \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.carry_s1 ;
assign _0171_ = \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.ce  ? \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.fas_s1  : \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.sum_s1 ;
assign _0172_ = \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.u1.a  + \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.u1.b ;
assign { \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.u1.cout , \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.u1.s  } = _0172_ + \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.u1.cin ;
assign _0173_ = \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.u2.a  + \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.u2.b ;
assign { \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.u2.cout , \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.u2.s  } = _0173_ + \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.u2.cin ;
always @(posedge \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_9_U.clk )
\add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_9_U.bin_s1  <= _0175_;
always @(posedge \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_9_U.clk )
\add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_9_U.ain_s1  <= _0174_;
always @(posedge \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_9_U.clk )
\add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_9_U.sum_s1  <= _0177_;
always @(posedge \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_9_U.clk )
\add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_9_U.carry_s1  <= _0176_;
assign _0175_ = \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_9_U.ce  ? \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_9_U.b [31:16] : \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_9_U.bin_s1 ;
assign _0174_ = \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_9_U.ce  ? \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_9_U.a [31:16] : \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_9_U.ain_s1 ;
assign _0176_ = \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_9_U.ce  ? \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_9_U.facout_s1  : \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_9_U.carry_s1 ;
assign _0177_ = \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_9_U.ce  ? \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_9_U.fas_s1  : \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_9_U.sum_s1 ;
assign _0178_ = \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_9_U.u1.a  + \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_9_U.u1.b ;
assign { \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_9_U.u1.cout , \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_9_U.u1.s  } = _0178_ + \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_9_U.u1.cin ;
assign _0179_ = \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_9_U.u2.a  + \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_9_U.u2.b ;
assign { \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_9_U.u2.cout , \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_9_U.u2.s  } = _0179_ + \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_9_U.u2.cin ;
always @(posedge \add_34s_34s_34_2_1_U12.top_add_34s_34s_34_2_1_Adder_6_U.clk )
\add_34s_34s_34_2_1_U12.top_add_34s_34s_34_2_1_Adder_6_U.bin_s1  <= _0181_;
always @(posedge \add_34s_34s_34_2_1_U12.top_add_34s_34s_34_2_1_Adder_6_U.clk )
\add_34s_34s_34_2_1_U12.top_add_34s_34s_34_2_1_Adder_6_U.ain_s1  <= _0180_;
always @(posedge \add_34s_34s_34_2_1_U12.top_add_34s_34s_34_2_1_Adder_6_U.clk )
\add_34s_34s_34_2_1_U12.top_add_34s_34s_34_2_1_Adder_6_U.sum_s1  <= _0183_;
always @(posedge \add_34s_34s_34_2_1_U12.top_add_34s_34s_34_2_1_Adder_6_U.clk )
\add_34s_34s_34_2_1_U12.top_add_34s_34s_34_2_1_Adder_6_U.carry_s1  <= _0182_;
assign _0181_ = \add_34s_34s_34_2_1_U12.top_add_34s_34s_34_2_1_Adder_6_U.ce  ? \add_34s_34s_34_2_1_U12.top_add_34s_34s_34_2_1_Adder_6_U.b [33:17] : \add_34s_34s_34_2_1_U12.top_add_34s_34s_34_2_1_Adder_6_U.bin_s1 ;
assign _0180_ = \add_34s_34s_34_2_1_U12.top_add_34s_34s_34_2_1_Adder_6_U.ce  ? \add_34s_34s_34_2_1_U12.top_add_34s_34s_34_2_1_Adder_6_U.a [33:17] : \add_34s_34s_34_2_1_U12.top_add_34s_34s_34_2_1_Adder_6_U.ain_s1 ;
assign _0182_ = \add_34s_34s_34_2_1_U12.top_add_34s_34s_34_2_1_Adder_6_U.ce  ? \add_34s_34s_34_2_1_U12.top_add_34s_34s_34_2_1_Adder_6_U.facout_s1  : \add_34s_34s_34_2_1_U12.top_add_34s_34s_34_2_1_Adder_6_U.carry_s1 ;
assign _0183_ = \add_34s_34s_34_2_1_U12.top_add_34s_34s_34_2_1_Adder_6_U.ce  ? \add_34s_34s_34_2_1_U12.top_add_34s_34s_34_2_1_Adder_6_U.fas_s1  : \add_34s_34s_34_2_1_U12.top_add_34s_34s_34_2_1_Adder_6_U.sum_s1 ;
assign _0184_ = \add_34s_34s_34_2_1_U12.top_add_34s_34s_34_2_1_Adder_6_U.u1.a  + \add_34s_34s_34_2_1_U12.top_add_34s_34s_34_2_1_Adder_6_U.u1.b ;
assign { \add_34s_34s_34_2_1_U12.top_add_34s_34s_34_2_1_Adder_6_U.u1.cout , \add_34s_34s_34_2_1_U12.top_add_34s_34s_34_2_1_Adder_6_U.u1.s  } = _0184_ + \add_34s_34s_34_2_1_U12.top_add_34s_34s_34_2_1_Adder_6_U.u1.cin ;
assign _0185_ = \add_34s_34s_34_2_1_U12.top_add_34s_34s_34_2_1_Adder_6_U.u2.a  + \add_34s_34s_34_2_1_U12.top_add_34s_34s_34_2_1_Adder_6_U.u2.b ;
assign { \add_34s_34s_34_2_1_U12.top_add_34s_34s_34_2_1_Adder_6_U.u2.cout , \add_34s_34s_34_2_1_U12.top_add_34s_34s_34_2_1_Adder_6_U.u2.s  } = _0185_ + \add_34s_34s_34_2_1_U12.top_add_34s_34s_34_2_1_Adder_6_U.u2.cin ;
always @(posedge \add_34s_34s_34_2_1_U21.top_add_34s_34s_34_2_1_Adder_6_U.clk )
\add_34s_34s_34_2_1_U21.top_add_34s_34s_34_2_1_Adder_6_U.bin_s1  <= _0187_;
always @(posedge \add_34s_34s_34_2_1_U21.top_add_34s_34s_34_2_1_Adder_6_U.clk )
\add_34s_34s_34_2_1_U21.top_add_34s_34s_34_2_1_Adder_6_U.ain_s1  <= _0186_;
always @(posedge \add_34s_34s_34_2_1_U21.top_add_34s_34s_34_2_1_Adder_6_U.clk )
\add_34s_34s_34_2_1_U21.top_add_34s_34s_34_2_1_Adder_6_U.sum_s1  <= _0189_;
always @(posedge \add_34s_34s_34_2_1_U21.top_add_34s_34s_34_2_1_Adder_6_U.clk )
\add_34s_34s_34_2_1_U21.top_add_34s_34s_34_2_1_Adder_6_U.carry_s1  <= _0188_;
assign _0187_ = \add_34s_34s_34_2_1_U21.top_add_34s_34s_34_2_1_Adder_6_U.ce  ? \add_34s_34s_34_2_1_U21.top_add_34s_34s_34_2_1_Adder_6_U.b [33:17] : \add_34s_34s_34_2_1_U21.top_add_34s_34s_34_2_1_Adder_6_U.bin_s1 ;
assign _0186_ = \add_34s_34s_34_2_1_U21.top_add_34s_34s_34_2_1_Adder_6_U.ce  ? \add_34s_34s_34_2_1_U21.top_add_34s_34s_34_2_1_Adder_6_U.a [33:17] : \add_34s_34s_34_2_1_U21.top_add_34s_34s_34_2_1_Adder_6_U.ain_s1 ;
assign _0188_ = \add_34s_34s_34_2_1_U21.top_add_34s_34s_34_2_1_Adder_6_U.ce  ? \add_34s_34s_34_2_1_U21.top_add_34s_34s_34_2_1_Adder_6_U.facout_s1  : \add_34s_34s_34_2_1_U21.top_add_34s_34s_34_2_1_Adder_6_U.carry_s1 ;
assign _0189_ = \add_34s_34s_34_2_1_U21.top_add_34s_34s_34_2_1_Adder_6_U.ce  ? \add_34s_34s_34_2_1_U21.top_add_34s_34s_34_2_1_Adder_6_U.fas_s1  : \add_34s_34s_34_2_1_U21.top_add_34s_34s_34_2_1_Adder_6_U.sum_s1 ;
assign _0190_ = \add_34s_34s_34_2_1_U21.top_add_34s_34s_34_2_1_Adder_6_U.u1.a  + \add_34s_34s_34_2_1_U21.top_add_34s_34s_34_2_1_Adder_6_U.u1.b ;
assign { \add_34s_34s_34_2_1_U21.top_add_34s_34s_34_2_1_Adder_6_U.u1.cout , \add_34s_34s_34_2_1_U21.top_add_34s_34s_34_2_1_Adder_6_U.u1.s  } = _0190_ + \add_34s_34s_34_2_1_U21.top_add_34s_34s_34_2_1_Adder_6_U.u1.cin ;
assign _0191_ = \add_34s_34s_34_2_1_U21.top_add_34s_34s_34_2_1_Adder_6_U.u2.a  + \add_34s_34s_34_2_1_U21.top_add_34s_34s_34_2_1_Adder_6_U.u2.b ;
assign { \add_34s_34s_34_2_1_U21.top_add_34s_34s_34_2_1_Adder_6_U.u2.cout , \add_34s_34s_34_2_1_U21.top_add_34s_34s_34_2_1_Adder_6_U.u2.s  } = _0191_ + \add_34s_34s_34_2_1_U21.top_add_34s_34s_34_2_1_Adder_6_U.u2.cin ;
always @(posedge \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_6_U.clk )
\add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_6_U.bin_s1  <= _0193_;
always @(posedge \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_6_U.clk )
\add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_6_U.ain_s1  <= _0192_;
always @(posedge \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_6_U.clk )
\add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_6_U.sum_s1  <= _0195_;
always @(posedge \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_6_U.clk )
\add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_6_U.carry_s1  <= _0194_;
assign _0193_ = \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_6_U.ce  ? \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_6_U.b [33:17] : \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_6_U.bin_s1 ;
assign _0192_ = \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_6_U.ce  ? \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_6_U.a [33:17] : \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_6_U.ain_s1 ;
assign _0194_ = \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_6_U.ce  ? \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_6_U.facout_s1  : \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_6_U.carry_s1 ;
assign _0195_ = \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_6_U.ce  ? \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_6_U.fas_s1  : \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_6_U.sum_s1 ;
assign _0196_ = \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_6_U.u1.a  + \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_6_U.u1.b ;
assign { \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_6_U.u1.cout , \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_6_U.u1.s  } = _0196_ + \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_6_U.u1.cin ;
assign _0197_ = \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_6_U.u2.a  + \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_6_U.u2.b ;
assign { \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_6_U.u2.cout , \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_6_U.u2.s  } = _0197_ + \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_6_U.u2.cin ;
always @(posedge \add_37s_37s_37_2_1_U18.top_add_37s_37s_37_2_1_Adder_11_U.clk )
\add_37s_37s_37_2_1_U18.top_add_37s_37s_37_2_1_Adder_11_U.bin_s1  <= _0199_;
always @(posedge \add_37s_37s_37_2_1_U18.top_add_37s_37s_37_2_1_Adder_11_U.clk )
\add_37s_37s_37_2_1_U18.top_add_37s_37s_37_2_1_Adder_11_U.ain_s1  <= _0198_;
always @(posedge \add_37s_37s_37_2_1_U18.top_add_37s_37s_37_2_1_Adder_11_U.clk )
\add_37s_37s_37_2_1_U18.top_add_37s_37s_37_2_1_Adder_11_U.sum_s1  <= _0201_;
always @(posedge \add_37s_37s_37_2_1_U18.top_add_37s_37s_37_2_1_Adder_11_U.clk )
\add_37s_37s_37_2_1_U18.top_add_37s_37s_37_2_1_Adder_11_U.carry_s1  <= _0200_;
assign _0199_ = \add_37s_37s_37_2_1_U18.top_add_37s_37s_37_2_1_Adder_11_U.ce  ? \add_37s_37s_37_2_1_U18.top_add_37s_37s_37_2_1_Adder_11_U.b [36:18] : \add_37s_37s_37_2_1_U18.top_add_37s_37s_37_2_1_Adder_11_U.bin_s1 ;
assign _0198_ = \add_37s_37s_37_2_1_U18.top_add_37s_37s_37_2_1_Adder_11_U.ce  ? \add_37s_37s_37_2_1_U18.top_add_37s_37s_37_2_1_Adder_11_U.a [36:18] : \add_37s_37s_37_2_1_U18.top_add_37s_37s_37_2_1_Adder_11_U.ain_s1 ;
assign _0200_ = \add_37s_37s_37_2_1_U18.top_add_37s_37s_37_2_1_Adder_11_U.ce  ? \add_37s_37s_37_2_1_U18.top_add_37s_37s_37_2_1_Adder_11_U.facout_s1  : \add_37s_37s_37_2_1_U18.top_add_37s_37s_37_2_1_Adder_11_U.carry_s1 ;
assign _0201_ = \add_37s_37s_37_2_1_U18.top_add_37s_37s_37_2_1_Adder_11_U.ce  ? \add_37s_37s_37_2_1_U18.top_add_37s_37s_37_2_1_Adder_11_U.fas_s1  : \add_37s_37s_37_2_1_U18.top_add_37s_37s_37_2_1_Adder_11_U.sum_s1 ;
assign _0202_ = \add_37s_37s_37_2_1_U18.top_add_37s_37s_37_2_1_Adder_11_U.u1.a  + \add_37s_37s_37_2_1_U18.top_add_37s_37s_37_2_1_Adder_11_U.u1.b ;
assign { \add_37s_37s_37_2_1_U18.top_add_37s_37s_37_2_1_Adder_11_U.u1.cout , \add_37s_37s_37_2_1_U18.top_add_37s_37s_37_2_1_Adder_11_U.u1.s  } = _0202_ + \add_37s_37s_37_2_1_U18.top_add_37s_37s_37_2_1_Adder_11_U.u1.cin ;
assign _0203_ = \add_37s_37s_37_2_1_U18.top_add_37s_37s_37_2_1_Adder_11_U.u2.a  + \add_37s_37s_37_2_1_U18.top_add_37s_37s_37_2_1_Adder_11_U.u2.b ;
assign { \add_37s_37s_37_2_1_U18.top_add_37s_37s_37_2_1_Adder_11_U.u2.cout , \add_37s_37s_37_2_1_U18.top_add_37s_37s_37_2_1_Adder_11_U.u2.s  } = _0203_ + \add_37s_37s_37_2_1_U18.top_add_37s_37s_37_2_1_Adder_11_U.u2.cin ;
always @(posedge \add_3s_3ns_3_2_1_U17.top_add_3s_3ns_3_2_1_Adder_10_U.clk )
\add_3s_3ns_3_2_1_U17.top_add_3s_3ns_3_2_1_Adder_10_U.bin_s1  <= _0205_;
always @(posedge \add_3s_3ns_3_2_1_U17.top_add_3s_3ns_3_2_1_Adder_10_U.clk )
\add_3s_3ns_3_2_1_U17.top_add_3s_3ns_3_2_1_Adder_10_U.ain_s1  <= _0204_;
always @(posedge \add_3s_3ns_3_2_1_U17.top_add_3s_3ns_3_2_1_Adder_10_U.clk )
\add_3s_3ns_3_2_1_U17.top_add_3s_3ns_3_2_1_Adder_10_U.sum_s1  <= _0207_;
always @(posedge \add_3s_3ns_3_2_1_U17.top_add_3s_3ns_3_2_1_Adder_10_U.clk )
\add_3s_3ns_3_2_1_U17.top_add_3s_3ns_3_2_1_Adder_10_U.carry_s1  <= _0206_;
assign _0205_ = \add_3s_3ns_3_2_1_U17.top_add_3s_3ns_3_2_1_Adder_10_U.ce  ? \add_3s_3ns_3_2_1_U17.top_add_3s_3ns_3_2_1_Adder_10_U.b [2:1] : \add_3s_3ns_3_2_1_U17.top_add_3s_3ns_3_2_1_Adder_10_U.bin_s1 ;
assign _0204_ = \add_3s_3ns_3_2_1_U17.top_add_3s_3ns_3_2_1_Adder_10_U.ce  ? \add_3s_3ns_3_2_1_U17.top_add_3s_3ns_3_2_1_Adder_10_U.a [2:1] : \add_3s_3ns_3_2_1_U17.top_add_3s_3ns_3_2_1_Adder_10_U.ain_s1 ;
assign _0206_ = \add_3s_3ns_3_2_1_U17.top_add_3s_3ns_3_2_1_Adder_10_U.ce  ? \add_3s_3ns_3_2_1_U17.top_add_3s_3ns_3_2_1_Adder_10_U.facout_s1  : \add_3s_3ns_3_2_1_U17.top_add_3s_3ns_3_2_1_Adder_10_U.carry_s1 ;
assign _0207_ = \add_3s_3ns_3_2_1_U17.top_add_3s_3ns_3_2_1_Adder_10_U.ce  ? \add_3s_3ns_3_2_1_U17.top_add_3s_3ns_3_2_1_Adder_10_U.fas_s1  : \add_3s_3ns_3_2_1_U17.top_add_3s_3ns_3_2_1_Adder_10_U.sum_s1 ;
assign _0208_ = \add_3s_3ns_3_2_1_U17.top_add_3s_3ns_3_2_1_Adder_10_U.u1.a  + \add_3s_3ns_3_2_1_U17.top_add_3s_3ns_3_2_1_Adder_10_U.u1.b ;
assign { \add_3s_3ns_3_2_1_U17.top_add_3s_3ns_3_2_1_Adder_10_U.u1.cout , \add_3s_3ns_3_2_1_U17.top_add_3s_3ns_3_2_1_Adder_10_U.u1.s  } = _0208_ + \add_3s_3ns_3_2_1_U17.top_add_3s_3ns_3_2_1_Adder_10_U.u1.cin ;
assign _0209_ = \add_3s_3ns_3_2_1_U17.top_add_3s_3ns_3_2_1_Adder_10_U.u2.a  + \add_3s_3ns_3_2_1_U17.top_add_3s_3ns_3_2_1_Adder_10_U.u2.b ;
assign { \add_3s_3ns_3_2_1_U17.top_add_3s_3ns_3_2_1_Adder_10_U.u2.cout , \add_3s_3ns_3_2_1_U17.top_add_3s_3ns_3_2_1_Adder_10_U.u2.s  } = _0209_ + \add_3s_3ns_3_2_1_U17.top_add_3s_3ns_3_2_1_Adder_10_U.u2.cin ;
always @(posedge \add_4ns_4ns_4_2_1_U3.top_add_4ns_4ns_4_2_1_Adder_2_U.clk )
\add_4ns_4ns_4_2_1_U3.top_add_4ns_4ns_4_2_1_Adder_2_U.bin_s1  <= _0211_;
always @(posedge \add_4ns_4ns_4_2_1_U3.top_add_4ns_4ns_4_2_1_Adder_2_U.clk )
\add_4ns_4ns_4_2_1_U3.top_add_4ns_4ns_4_2_1_Adder_2_U.ain_s1  <= _0210_;
always @(posedge \add_4ns_4ns_4_2_1_U3.top_add_4ns_4ns_4_2_1_Adder_2_U.clk )
\add_4ns_4ns_4_2_1_U3.top_add_4ns_4ns_4_2_1_Adder_2_U.sum_s1  <= _0213_;
always @(posedge \add_4ns_4ns_4_2_1_U3.top_add_4ns_4ns_4_2_1_Adder_2_U.clk )
\add_4ns_4ns_4_2_1_U3.top_add_4ns_4ns_4_2_1_Adder_2_U.carry_s1  <= _0212_;
assign _0211_ = \add_4ns_4ns_4_2_1_U3.top_add_4ns_4ns_4_2_1_Adder_2_U.ce  ? \add_4ns_4ns_4_2_1_U3.top_add_4ns_4ns_4_2_1_Adder_2_U.b [3:2] : \add_4ns_4ns_4_2_1_U3.top_add_4ns_4ns_4_2_1_Adder_2_U.bin_s1 ;
assign _0210_ = \add_4ns_4ns_4_2_1_U3.top_add_4ns_4ns_4_2_1_Adder_2_U.ce  ? \add_4ns_4ns_4_2_1_U3.top_add_4ns_4ns_4_2_1_Adder_2_U.a [3:2] : \add_4ns_4ns_4_2_1_U3.top_add_4ns_4ns_4_2_1_Adder_2_U.ain_s1 ;
assign _0212_ = \add_4ns_4ns_4_2_1_U3.top_add_4ns_4ns_4_2_1_Adder_2_U.ce  ? \add_4ns_4ns_4_2_1_U3.top_add_4ns_4ns_4_2_1_Adder_2_U.facout_s1  : \add_4ns_4ns_4_2_1_U3.top_add_4ns_4ns_4_2_1_Adder_2_U.carry_s1 ;
assign _0213_ = \add_4ns_4ns_4_2_1_U3.top_add_4ns_4ns_4_2_1_Adder_2_U.ce  ? \add_4ns_4ns_4_2_1_U3.top_add_4ns_4ns_4_2_1_Adder_2_U.fas_s1  : \add_4ns_4ns_4_2_1_U3.top_add_4ns_4ns_4_2_1_Adder_2_U.sum_s1 ;
assign _0214_ = \add_4ns_4ns_4_2_1_U3.top_add_4ns_4ns_4_2_1_Adder_2_U.u1.a  + \add_4ns_4ns_4_2_1_U3.top_add_4ns_4ns_4_2_1_Adder_2_U.u1.b ;
assign { \add_4ns_4ns_4_2_1_U3.top_add_4ns_4ns_4_2_1_Adder_2_U.u1.cout , \add_4ns_4ns_4_2_1_U3.top_add_4ns_4ns_4_2_1_Adder_2_U.u1.s  } = _0214_ + \add_4ns_4ns_4_2_1_U3.top_add_4ns_4ns_4_2_1_Adder_2_U.u1.cin ;
assign _0215_ = \add_4ns_4ns_4_2_1_U3.top_add_4ns_4ns_4_2_1_Adder_2_U.u2.a  + \add_4ns_4ns_4_2_1_U3.top_add_4ns_4ns_4_2_1_Adder_2_U.u2.b ;
assign { \add_4ns_4ns_4_2_1_U3.top_add_4ns_4ns_4_2_1_Adder_2_U.u2.cout , \add_4ns_4ns_4_2_1_U3.top_add_4ns_4ns_4_2_1_Adder_2_U.u2.s  } = _0215_ + \add_4ns_4ns_4_2_1_U3.top_add_4ns_4ns_4_2_1_Adder_2_U.u2.cin ;
always @(posedge \add_7s_7ns_7_2_1_U10.top_add_7s_7ns_7_2_1_Adder_3_U.clk )
\add_7s_7ns_7_2_1_U10.top_add_7s_7ns_7_2_1_Adder_3_U.bin_s1  <= _0217_;
always @(posedge \add_7s_7ns_7_2_1_U10.top_add_7s_7ns_7_2_1_Adder_3_U.clk )
\add_7s_7ns_7_2_1_U10.top_add_7s_7ns_7_2_1_Adder_3_U.ain_s1  <= _0216_;
always @(posedge \add_7s_7ns_7_2_1_U10.top_add_7s_7ns_7_2_1_Adder_3_U.clk )
\add_7s_7ns_7_2_1_U10.top_add_7s_7ns_7_2_1_Adder_3_U.sum_s1  <= _0219_;
always @(posedge \add_7s_7ns_7_2_1_U10.top_add_7s_7ns_7_2_1_Adder_3_U.clk )
\add_7s_7ns_7_2_1_U10.top_add_7s_7ns_7_2_1_Adder_3_U.carry_s1  <= _0218_;
assign _0217_ = \add_7s_7ns_7_2_1_U10.top_add_7s_7ns_7_2_1_Adder_3_U.ce  ? \add_7s_7ns_7_2_1_U10.top_add_7s_7ns_7_2_1_Adder_3_U.b [6:3] : \add_7s_7ns_7_2_1_U10.top_add_7s_7ns_7_2_1_Adder_3_U.bin_s1 ;
assign _0216_ = \add_7s_7ns_7_2_1_U10.top_add_7s_7ns_7_2_1_Adder_3_U.ce  ? \add_7s_7ns_7_2_1_U10.top_add_7s_7ns_7_2_1_Adder_3_U.a [6:3] : \add_7s_7ns_7_2_1_U10.top_add_7s_7ns_7_2_1_Adder_3_U.ain_s1 ;
assign _0218_ = \add_7s_7ns_7_2_1_U10.top_add_7s_7ns_7_2_1_Adder_3_U.ce  ? \add_7s_7ns_7_2_1_U10.top_add_7s_7ns_7_2_1_Adder_3_U.facout_s1  : \add_7s_7ns_7_2_1_U10.top_add_7s_7ns_7_2_1_Adder_3_U.carry_s1 ;
assign _0219_ = \add_7s_7ns_7_2_1_U10.top_add_7s_7ns_7_2_1_Adder_3_U.ce  ? \add_7s_7ns_7_2_1_U10.top_add_7s_7ns_7_2_1_Adder_3_U.fas_s1  : \add_7s_7ns_7_2_1_U10.top_add_7s_7ns_7_2_1_Adder_3_U.sum_s1 ;
assign _0220_ = \add_7s_7ns_7_2_1_U10.top_add_7s_7ns_7_2_1_Adder_3_U.u1.a  + \add_7s_7ns_7_2_1_U10.top_add_7s_7ns_7_2_1_Adder_3_U.u1.b ;
assign { \add_7s_7ns_7_2_1_U10.top_add_7s_7ns_7_2_1_Adder_3_U.u1.cout , \add_7s_7ns_7_2_1_U10.top_add_7s_7ns_7_2_1_Adder_3_U.u1.s  } = _0220_ + \add_7s_7ns_7_2_1_U10.top_add_7s_7ns_7_2_1_Adder_3_U.u1.cin ;
assign _0221_ = \add_7s_7ns_7_2_1_U10.top_add_7s_7ns_7_2_1_Adder_3_U.u2.a  + \add_7s_7ns_7_2_1_U10.top_add_7s_7ns_7_2_1_Adder_3_U.u2.b ;
assign { \add_7s_7ns_7_2_1_U10.top_add_7s_7ns_7_2_1_Adder_3_U.u2.cout , \add_7s_7ns_7_2_1_U10.top_add_7s_7ns_7_2_1_Adder_3_U.u2.s  } = _0221_ + \add_7s_7ns_7_2_1_U10.top_add_7s_7ns_7_2_1_Adder_3_U.u2.cin ;
always @(posedge \add_7s_7ns_7_2_1_U6.top_add_7s_7ns_7_2_1_Adder_3_U.clk )
\add_7s_7ns_7_2_1_U6.top_add_7s_7ns_7_2_1_Adder_3_U.bin_s1  <= _0223_;
always @(posedge \add_7s_7ns_7_2_1_U6.top_add_7s_7ns_7_2_1_Adder_3_U.clk )
\add_7s_7ns_7_2_1_U6.top_add_7s_7ns_7_2_1_Adder_3_U.ain_s1  <= _0222_;
always @(posedge \add_7s_7ns_7_2_1_U6.top_add_7s_7ns_7_2_1_Adder_3_U.clk )
\add_7s_7ns_7_2_1_U6.top_add_7s_7ns_7_2_1_Adder_3_U.sum_s1  <= _0225_;
always @(posedge \add_7s_7ns_7_2_1_U6.top_add_7s_7ns_7_2_1_Adder_3_U.clk )
\add_7s_7ns_7_2_1_U6.top_add_7s_7ns_7_2_1_Adder_3_U.carry_s1  <= _0224_;
assign _0223_ = \add_7s_7ns_7_2_1_U6.top_add_7s_7ns_7_2_1_Adder_3_U.ce  ? \add_7s_7ns_7_2_1_U6.top_add_7s_7ns_7_2_1_Adder_3_U.b [6:3] : \add_7s_7ns_7_2_1_U6.top_add_7s_7ns_7_2_1_Adder_3_U.bin_s1 ;
assign _0222_ = \add_7s_7ns_7_2_1_U6.top_add_7s_7ns_7_2_1_Adder_3_U.ce  ? \add_7s_7ns_7_2_1_U6.top_add_7s_7ns_7_2_1_Adder_3_U.a [6:3] : \add_7s_7ns_7_2_1_U6.top_add_7s_7ns_7_2_1_Adder_3_U.ain_s1 ;
assign _0224_ = \add_7s_7ns_7_2_1_U6.top_add_7s_7ns_7_2_1_Adder_3_U.ce  ? \add_7s_7ns_7_2_1_U6.top_add_7s_7ns_7_2_1_Adder_3_U.facout_s1  : \add_7s_7ns_7_2_1_U6.top_add_7s_7ns_7_2_1_Adder_3_U.carry_s1 ;
assign _0225_ = \add_7s_7ns_7_2_1_U6.top_add_7s_7ns_7_2_1_Adder_3_U.ce  ? \add_7s_7ns_7_2_1_U6.top_add_7s_7ns_7_2_1_Adder_3_U.fas_s1  : \add_7s_7ns_7_2_1_U6.top_add_7s_7ns_7_2_1_Adder_3_U.sum_s1 ;
assign _0226_ = \add_7s_7ns_7_2_1_U6.top_add_7s_7ns_7_2_1_Adder_3_U.u1.a  + \add_7s_7ns_7_2_1_U6.top_add_7s_7ns_7_2_1_Adder_3_U.u1.b ;
assign { \add_7s_7ns_7_2_1_U6.top_add_7s_7ns_7_2_1_Adder_3_U.u1.cout , \add_7s_7ns_7_2_1_U6.top_add_7s_7ns_7_2_1_Adder_3_U.u1.s  } = _0226_ + \add_7s_7ns_7_2_1_U6.top_add_7s_7ns_7_2_1_Adder_3_U.u1.cin ;
assign _0227_ = \add_7s_7ns_7_2_1_U6.top_add_7s_7ns_7_2_1_Adder_3_U.u2.a  + \add_7s_7ns_7_2_1_U6.top_add_7s_7ns_7_2_1_Adder_3_U.u2.b ;
assign { \add_7s_7ns_7_2_1_U6.top_add_7s_7ns_7_2_1_Adder_3_U.u2.cout , \add_7s_7ns_7_2_1_U6.top_add_7s_7ns_7_2_1_Adder_3_U.u2.s  } = _0227_ + \add_7s_7ns_7_2_1_U6.top_add_7s_7ns_7_2_1_Adder_3_U.u2.cin ;
always @(posedge \add_8ns_8ns_8_2_1_U1.top_add_8ns_8ns_8_2_1_Adder_0_U.clk )
\add_8ns_8ns_8_2_1_U1.top_add_8ns_8ns_8_2_1_Adder_0_U.bin_s1  <= _0229_;
always @(posedge \add_8ns_8ns_8_2_1_U1.top_add_8ns_8ns_8_2_1_Adder_0_U.clk )
\add_8ns_8ns_8_2_1_U1.top_add_8ns_8ns_8_2_1_Adder_0_U.ain_s1  <= _0228_;
always @(posedge \add_8ns_8ns_8_2_1_U1.top_add_8ns_8ns_8_2_1_Adder_0_U.clk )
\add_8ns_8ns_8_2_1_U1.top_add_8ns_8ns_8_2_1_Adder_0_U.sum_s1  <= _0231_;
always @(posedge \add_8ns_8ns_8_2_1_U1.top_add_8ns_8ns_8_2_1_Adder_0_U.clk )
\add_8ns_8ns_8_2_1_U1.top_add_8ns_8ns_8_2_1_Adder_0_U.carry_s1  <= _0230_;
assign _0229_ = \add_8ns_8ns_8_2_1_U1.top_add_8ns_8ns_8_2_1_Adder_0_U.ce  ? \add_8ns_8ns_8_2_1_U1.top_add_8ns_8ns_8_2_1_Adder_0_U.b [7:4] : \add_8ns_8ns_8_2_1_U1.top_add_8ns_8ns_8_2_1_Adder_0_U.bin_s1 ;
assign _0228_ = \add_8ns_8ns_8_2_1_U1.top_add_8ns_8ns_8_2_1_Adder_0_U.ce  ? \add_8ns_8ns_8_2_1_U1.top_add_8ns_8ns_8_2_1_Adder_0_U.a [7:4] : \add_8ns_8ns_8_2_1_U1.top_add_8ns_8ns_8_2_1_Adder_0_U.ain_s1 ;
assign _0230_ = \add_8ns_8ns_8_2_1_U1.top_add_8ns_8ns_8_2_1_Adder_0_U.ce  ? \add_8ns_8ns_8_2_1_U1.top_add_8ns_8ns_8_2_1_Adder_0_U.facout_s1  : \add_8ns_8ns_8_2_1_U1.top_add_8ns_8ns_8_2_1_Adder_0_U.carry_s1 ;
assign _0231_ = \add_8ns_8ns_8_2_1_U1.top_add_8ns_8ns_8_2_1_Adder_0_U.ce  ? \add_8ns_8ns_8_2_1_U1.top_add_8ns_8ns_8_2_1_Adder_0_U.fas_s1  : \add_8ns_8ns_8_2_1_U1.top_add_8ns_8ns_8_2_1_Adder_0_U.sum_s1 ;
assign _0232_ = \add_8ns_8ns_8_2_1_U1.top_add_8ns_8ns_8_2_1_Adder_0_U.u1.a  + \add_8ns_8ns_8_2_1_U1.top_add_8ns_8ns_8_2_1_Adder_0_U.u1.b ;
assign { \add_8ns_8ns_8_2_1_U1.top_add_8ns_8ns_8_2_1_Adder_0_U.u1.cout , \add_8ns_8ns_8_2_1_U1.top_add_8ns_8ns_8_2_1_Adder_0_U.u1.s  } = _0232_ + \add_8ns_8ns_8_2_1_U1.top_add_8ns_8ns_8_2_1_Adder_0_U.u1.cin ;
assign _0233_ = \add_8ns_8ns_8_2_1_U1.top_add_8ns_8ns_8_2_1_Adder_0_U.u2.a  + \add_8ns_8ns_8_2_1_U1.top_add_8ns_8ns_8_2_1_Adder_0_U.u2.b ;
assign { \add_8ns_8ns_8_2_1_U1.top_add_8ns_8ns_8_2_1_Adder_0_U.u2.cout , \add_8ns_8ns_8_2_1_U1.top_add_8ns_8ns_8_2_1_Adder_0_U.u2.s  } = _0233_ + \add_8ns_8ns_8_2_1_U1.top_add_8ns_8ns_8_2_1_Adder_0_U.u2.cin ;
always @(posedge \ashr_32s_32s_32_7_1_U4.clk )
\ashr_32s_32s_32_7_1_U4.dout_array[5]  <= _0245_;
always @(posedge \ashr_32s_32s_32_7_1_U4.clk )
\ashr_32s_32s_32_7_1_U4.din1_cast_array[5]  <= _0239_;
always @(posedge \ashr_32s_32s_32_7_1_U4.clk )
\ashr_32s_32s_32_7_1_U4.dout_array[4]  <= _0244_;
always @(posedge \ashr_32s_32s_32_7_1_U4.clk )
\ashr_32s_32s_32_7_1_U4.din1_cast_array[4]  <= _0238_;
always @(posedge \ashr_32s_32s_32_7_1_U4.clk )
\ashr_32s_32s_32_7_1_U4.dout_array[3]  <= _0243_;
always @(posedge \ashr_32s_32s_32_7_1_U4.clk )
\ashr_32s_32s_32_7_1_U4.din1_cast_array[3]  <= _0237_;
always @(posedge \ashr_32s_32s_32_7_1_U4.clk )
\ashr_32s_32s_32_7_1_U4.dout_array[2]  <= _0242_;
always @(posedge \ashr_32s_32s_32_7_1_U4.clk )
\ashr_32s_32s_32_7_1_U4.din1_cast_array[2]  <= _0236_;
always @(posedge \ashr_32s_32s_32_7_1_U4.clk )
\ashr_32s_32s_32_7_1_U4.dout_array[1]  <= _0241_;
always @(posedge \ashr_32s_32s_32_7_1_U4.clk )
\ashr_32s_32s_32_7_1_U4.din1_cast_array[1]  <= _0235_;
always @(posedge \ashr_32s_32s_32_7_1_U4.clk )
\ashr_32s_32s_32_7_1_U4.dout_array[0]  <= _0240_;
always @(posedge \ashr_32s_32s_32_7_1_U4.clk )
\ashr_32s_32s_32_7_1_U4.din1_cast_array[0]  <= _0234_;
assign _0246_ = \ashr_32s_32s_32_7_1_U4.ce  ? \ashr_32s_32s_32_7_1_U4.din1_cast_array[4]  : \ashr_32s_32s_32_7_1_U4.din1_cast_array[5] ;
assign _0239_ = \ashr_32s_32s_32_7_1_U4.reset  ? 32'd0 : _0246_;
assign _0247_ = \ashr_32s_32s_32_7_1_U4.ce  ? _0263_ : \ashr_32s_32s_32_7_1_U4.dout_array[5] ;
assign _0245_ = \ashr_32s_32s_32_7_1_U4.reset  ? 32'd0 : _0247_;
assign _0248_ = \ashr_32s_32s_32_7_1_U4.ce  ? \ashr_32s_32s_32_7_1_U4.din1_cast_array[3]  : \ashr_32s_32s_32_7_1_U4.din1_cast_array[4] ;
assign _0238_ = \ashr_32s_32s_32_7_1_U4.reset  ? 32'd0 : _0248_;
assign _0249_ = \ashr_32s_32s_32_7_1_U4.ce  ? _0262_ : \ashr_32s_32s_32_7_1_U4.dout_array[4] ;
assign _0244_ = \ashr_32s_32s_32_7_1_U4.reset  ? 32'd0 : _0249_;
assign _0250_ = \ashr_32s_32s_32_7_1_U4.ce  ? \ashr_32s_32s_32_7_1_U4.din1_cast_array[2]  : \ashr_32s_32s_32_7_1_U4.din1_cast_array[3] ;
assign _0237_ = \ashr_32s_32s_32_7_1_U4.reset  ? 32'd0 : _0250_;
assign _0251_ = \ashr_32s_32s_32_7_1_U4.ce  ? _0261_ : \ashr_32s_32s_32_7_1_U4.dout_array[3] ;
assign _0243_ = \ashr_32s_32s_32_7_1_U4.reset  ? 32'd0 : _0251_;
assign _0252_ = \ashr_32s_32s_32_7_1_U4.ce  ? \ashr_32s_32s_32_7_1_U4.din1_cast_array[1]  : \ashr_32s_32s_32_7_1_U4.din1_cast_array[2] ;
assign _0236_ = \ashr_32s_32s_32_7_1_U4.reset  ? 32'd0 : _0252_;
assign _0253_ = \ashr_32s_32s_32_7_1_U4.ce  ? _0260_ : \ashr_32s_32s_32_7_1_U4.dout_array[2] ;
assign _0242_ = \ashr_32s_32s_32_7_1_U4.reset  ? 32'd0 : _0253_;
assign _0254_ = \ashr_32s_32s_32_7_1_U4.ce  ? \ashr_32s_32s_32_7_1_U4.din1_cast_array[0]  : \ashr_32s_32s_32_7_1_U4.din1_cast_array[1] ;
assign _0235_ = \ashr_32s_32s_32_7_1_U4.reset  ? 32'd0 : _0254_;
assign _0255_ = \ashr_32s_32s_32_7_1_U4.ce  ? _0259_ : \ashr_32s_32s_32_7_1_U4.dout_array[1] ;
assign _0241_ = \ashr_32s_32s_32_7_1_U4.reset  ? 32'd0 : _0255_;
assign _0256_ = \ashr_32s_32s_32_7_1_U4.ce  ? \ashr_32s_32s_32_7_1_U4.din1  : \ashr_32s_32s_32_7_1_U4.din1_cast_array[0] ;
assign _0234_ = \ashr_32s_32s_32_7_1_U4.reset  ? 32'd0 : _0256_;
assign _0257_ = \ashr_32s_32s_32_7_1_U4.ce  ? _0258_ : \ashr_32s_32s_32_7_1_U4.dout_array[0] ;
assign _0240_ = \ashr_32s_32s_32_7_1_U4.reset  ? 32'd0 : _0257_;
assign _0258_ = $signed(\ashr_32s_32s_32_7_1_U4.din0 ) >>> { \ashr_32s_32s_32_7_1_U4.din1 [31:30], 30'h00000000 };
assign _0259_ = $signed(\ashr_32s_32s_32_7_1_U4.dout_array[0] ) >>> { \ashr_32s_32s_32_7_1_U4.din1_cast_array[0] [29:25], 25'h0000000 };
assign _0260_ = $signed(\ashr_32s_32s_32_7_1_U4.dout_array[1] ) >>> { \ashr_32s_32s_32_7_1_U4.din1_cast_array[1] [24:20], 20'h00000 };
assign _0261_ = $signed(\ashr_32s_32s_32_7_1_U4.dout_array[2] ) >>> { \ashr_32s_32s_32_7_1_U4.din1_cast_array[2] [19:15], 15'h0000 };
assign _0262_ = $signed(\ashr_32s_32s_32_7_1_U4.dout_array[3] ) >>> { \ashr_32s_32s_32_7_1_U4.din1_cast_array[3] [14:10], 10'h000 };
assign _0263_ = $signed(\ashr_32s_32s_32_7_1_U4.dout_array[4] ) >>> { \ashr_32s_32s_32_7_1_U4.din1_cast_array[4] [9:5], 5'h00 };
assign \ashr_32s_32s_32_7_1_U4.dout  = $signed(\ashr_32s_32s_32_7_1_U4.dout_array[5] ) >>> \ashr_32s_32s_32_7_1_U4.din1_cast_array[5] [4:0];
assign \mul_4s_2s_6_7_1_U8.top_mul_4s_2s_6_7_1_Mul_DSP_0_U.tmp_product  = $signed(\mul_4s_2s_6_7_1_U8.top_mul_4s_2s_6_7_1_Mul_DSP_0_U.a_reg0 ) * $signed(\mul_4s_2s_6_7_1_U8.top_mul_4s_2s_6_7_1_Mul_DSP_0_U.b_reg0 );
always @(posedge \mul_4s_2s_6_7_1_U8.top_mul_4s_2s_6_7_1_Mul_DSP_0_U.clk )
\mul_4s_2s_6_7_1_U8.top_mul_4s_2s_6_7_1_Mul_DSP_0_U.a_reg0  <= _0264_;
always @(posedge \mul_4s_2s_6_7_1_U8.top_mul_4s_2s_6_7_1_Mul_DSP_0_U.clk )
\mul_4s_2s_6_7_1_U8.top_mul_4s_2s_6_7_1_Mul_DSP_0_U.b_reg0  <= _0265_;
always @(posedge \mul_4s_2s_6_7_1_U8.top_mul_4s_2s_6_7_1_Mul_DSP_0_U.clk )
\mul_4s_2s_6_7_1_U8.top_mul_4s_2s_6_7_1_Mul_DSP_0_U.buff0  <= _0266_;
always @(posedge \mul_4s_2s_6_7_1_U8.top_mul_4s_2s_6_7_1_Mul_DSP_0_U.clk )
\mul_4s_2s_6_7_1_U8.top_mul_4s_2s_6_7_1_Mul_DSP_0_U.buff1  <= _0267_;
always @(posedge \mul_4s_2s_6_7_1_U8.top_mul_4s_2s_6_7_1_Mul_DSP_0_U.clk )
\mul_4s_2s_6_7_1_U8.top_mul_4s_2s_6_7_1_Mul_DSP_0_U.buff2  <= _0268_;
always @(posedge \mul_4s_2s_6_7_1_U8.top_mul_4s_2s_6_7_1_Mul_DSP_0_U.clk )
\mul_4s_2s_6_7_1_U8.top_mul_4s_2s_6_7_1_Mul_DSP_0_U.buff3  <= _0269_;
always @(posedge \mul_4s_2s_6_7_1_U8.top_mul_4s_2s_6_7_1_Mul_DSP_0_U.clk )
\mul_4s_2s_6_7_1_U8.top_mul_4s_2s_6_7_1_Mul_DSP_0_U.buff4  <= _0270_;
assign _0270_ = \mul_4s_2s_6_7_1_U8.top_mul_4s_2s_6_7_1_Mul_DSP_0_U.ce  ? \mul_4s_2s_6_7_1_U8.top_mul_4s_2s_6_7_1_Mul_DSP_0_U.buff3  : \mul_4s_2s_6_7_1_U8.top_mul_4s_2s_6_7_1_Mul_DSP_0_U.buff4 ;
assign _0269_ = \mul_4s_2s_6_7_1_U8.top_mul_4s_2s_6_7_1_Mul_DSP_0_U.ce  ? \mul_4s_2s_6_7_1_U8.top_mul_4s_2s_6_7_1_Mul_DSP_0_U.buff2  : \mul_4s_2s_6_7_1_U8.top_mul_4s_2s_6_7_1_Mul_DSP_0_U.buff3 ;
assign _0268_ = \mul_4s_2s_6_7_1_U8.top_mul_4s_2s_6_7_1_Mul_DSP_0_U.ce  ? \mul_4s_2s_6_7_1_U8.top_mul_4s_2s_6_7_1_Mul_DSP_0_U.buff1  : \mul_4s_2s_6_7_1_U8.top_mul_4s_2s_6_7_1_Mul_DSP_0_U.buff2 ;
assign _0267_ = \mul_4s_2s_6_7_1_U8.top_mul_4s_2s_6_7_1_Mul_DSP_0_U.ce  ? \mul_4s_2s_6_7_1_U8.top_mul_4s_2s_6_7_1_Mul_DSP_0_U.buff0  : \mul_4s_2s_6_7_1_U8.top_mul_4s_2s_6_7_1_Mul_DSP_0_U.buff1 ;
assign _0266_ = \mul_4s_2s_6_7_1_U8.top_mul_4s_2s_6_7_1_Mul_DSP_0_U.ce  ? \mul_4s_2s_6_7_1_U8.top_mul_4s_2s_6_7_1_Mul_DSP_0_U.tmp_product  : \mul_4s_2s_6_7_1_U8.top_mul_4s_2s_6_7_1_Mul_DSP_0_U.buff0 ;
assign _0265_ = \mul_4s_2s_6_7_1_U8.top_mul_4s_2s_6_7_1_Mul_DSP_0_U.ce  ? \mul_4s_2s_6_7_1_U8.top_mul_4s_2s_6_7_1_Mul_DSP_0_U.b  : \mul_4s_2s_6_7_1_U8.top_mul_4s_2s_6_7_1_Mul_DSP_0_U.b_reg0 ;
assign _0264_ = \mul_4s_2s_6_7_1_U8.top_mul_4s_2s_6_7_1_Mul_DSP_0_U.ce  ? \mul_4s_2s_6_7_1_U8.top_mul_4s_2s_6_7_1_Mul_DSP_0_U.a  : \mul_4s_2s_6_7_1_U8.top_mul_4s_2s_6_7_1_Mul_DSP_0_U.a_reg0 ;
always @(posedge \shl_32s_32s_32_7_1_U5.clk )
\shl_32s_32s_32_7_1_U5.dout_array[5]  <= _0282_;
always @(posedge \shl_32s_32s_32_7_1_U5.clk )
\shl_32s_32s_32_7_1_U5.din1_cast_array[5]  <= _0276_;
always @(posedge \shl_32s_32s_32_7_1_U5.clk )
\shl_32s_32s_32_7_1_U5.dout_array[4]  <= _0281_;
always @(posedge \shl_32s_32s_32_7_1_U5.clk )
\shl_32s_32s_32_7_1_U5.din1_cast_array[4]  <= _0275_;
always @(posedge \shl_32s_32s_32_7_1_U5.clk )
\shl_32s_32s_32_7_1_U5.dout_array[3]  <= _0280_;
always @(posedge \shl_32s_32s_32_7_1_U5.clk )
\shl_32s_32s_32_7_1_U5.din1_cast_array[3]  <= _0274_;
always @(posedge \shl_32s_32s_32_7_1_U5.clk )
\shl_32s_32s_32_7_1_U5.dout_array[2]  <= _0279_;
always @(posedge \shl_32s_32s_32_7_1_U5.clk )
\shl_32s_32s_32_7_1_U5.din1_cast_array[2]  <= _0273_;
always @(posedge \shl_32s_32s_32_7_1_U5.clk )
\shl_32s_32s_32_7_1_U5.dout_array[1]  <= _0278_;
always @(posedge \shl_32s_32s_32_7_1_U5.clk )
\shl_32s_32s_32_7_1_U5.din1_cast_array[1]  <= _0272_;
always @(posedge \shl_32s_32s_32_7_1_U5.clk )
\shl_32s_32s_32_7_1_U5.dout_array[0]  <= _0277_;
always @(posedge \shl_32s_32s_32_7_1_U5.clk )
\shl_32s_32s_32_7_1_U5.din1_cast_array[0]  <= _0271_;
assign _0283_ = \shl_32s_32s_32_7_1_U5.ce  ? \shl_32s_32s_32_7_1_U5.din1_cast_array[4]  : \shl_32s_32s_32_7_1_U5.din1_cast_array[5] ;
assign _0276_ = \shl_32s_32s_32_7_1_U5.reset  ? 32'd0 : _0283_;
assign _0284_ = \shl_32s_32s_32_7_1_U5.ce  ? _0300_ : \shl_32s_32s_32_7_1_U5.dout_array[5] ;
assign _0282_ = \shl_32s_32s_32_7_1_U5.reset  ? 32'd0 : _0284_;
assign _0285_ = \shl_32s_32s_32_7_1_U5.ce  ? \shl_32s_32s_32_7_1_U5.din1_cast_array[3]  : \shl_32s_32s_32_7_1_U5.din1_cast_array[4] ;
assign _0275_ = \shl_32s_32s_32_7_1_U5.reset  ? 32'd0 : _0285_;
assign _0286_ = \shl_32s_32s_32_7_1_U5.ce  ? _0299_ : \shl_32s_32s_32_7_1_U5.dout_array[4] ;
assign _0281_ = \shl_32s_32s_32_7_1_U5.reset  ? 32'd0 : _0286_;
assign _0287_ = \shl_32s_32s_32_7_1_U5.ce  ? \shl_32s_32s_32_7_1_U5.din1_cast_array[2]  : \shl_32s_32s_32_7_1_U5.din1_cast_array[3] ;
assign _0274_ = \shl_32s_32s_32_7_1_U5.reset  ? 32'd0 : _0287_;
assign _0288_ = \shl_32s_32s_32_7_1_U5.ce  ? _0298_ : \shl_32s_32s_32_7_1_U5.dout_array[3] ;
assign _0280_ = \shl_32s_32s_32_7_1_U5.reset  ? 32'd0 : _0288_;
assign _0289_ = \shl_32s_32s_32_7_1_U5.ce  ? \shl_32s_32s_32_7_1_U5.din1_cast_array[1]  : \shl_32s_32s_32_7_1_U5.din1_cast_array[2] ;
assign _0273_ = \shl_32s_32s_32_7_1_U5.reset  ? 32'd0 : _0289_;
assign _0290_ = \shl_32s_32s_32_7_1_U5.ce  ? _0297_ : \shl_32s_32s_32_7_1_U5.dout_array[2] ;
assign _0279_ = \shl_32s_32s_32_7_1_U5.reset  ? 32'd0 : _0290_;
assign _0291_ = \shl_32s_32s_32_7_1_U5.ce  ? \shl_32s_32s_32_7_1_U5.din1_cast_array[0]  : \shl_32s_32s_32_7_1_U5.din1_cast_array[1] ;
assign _0272_ = \shl_32s_32s_32_7_1_U5.reset  ? 32'd0 : _0291_;
assign _0292_ = \shl_32s_32s_32_7_1_U5.ce  ? _0296_ : \shl_32s_32s_32_7_1_U5.dout_array[1] ;
assign _0278_ = \shl_32s_32s_32_7_1_U5.reset  ? 32'd0 : _0292_;
assign _0293_ = \shl_32s_32s_32_7_1_U5.ce  ? \shl_32s_32s_32_7_1_U5.din1  : \shl_32s_32s_32_7_1_U5.din1_cast_array[0] ;
assign _0271_ = \shl_32s_32s_32_7_1_U5.reset  ? 32'd0 : _0293_;
assign _0294_ = \shl_32s_32s_32_7_1_U5.ce  ? _0295_ : \shl_32s_32s_32_7_1_U5.dout_array[0] ;
assign _0277_ = \shl_32s_32s_32_7_1_U5.reset  ? 32'd0 : _0294_;
assign _0295_ = \shl_32s_32s_32_7_1_U5.din0  << { \shl_32s_32s_32_7_1_U5.din1 [31:30], 30'h00000000 };
assign _0296_ = \shl_32s_32s_32_7_1_U5.dout_array[0]  << { \shl_32s_32s_32_7_1_U5.din1_cast_array[0] [29:25], 25'h0000000 };
assign _0297_ = \shl_32s_32s_32_7_1_U5.dout_array[1]  << { \shl_32s_32s_32_7_1_U5.din1_cast_array[1] [24:20], 20'h00000 };
assign _0298_ = \shl_32s_32s_32_7_1_U5.dout_array[2]  << { \shl_32s_32s_32_7_1_U5.din1_cast_array[2] [19:15], 15'h0000 };
assign _0299_ = \shl_32s_32s_32_7_1_U5.dout_array[3]  << { \shl_32s_32s_32_7_1_U5.din1_cast_array[3] [14:10], 10'h000 };
assign _0300_ = \shl_32s_32s_32_7_1_U5.dout_array[4]  << { \shl_32s_32s_32_7_1_U5.din1_cast_array[4] [9:5], 5'h00 };
assign \shl_32s_32s_32_7_1_U5.dout  = \shl_32s_32s_32_7_1_U5.dout_array[5]  << \shl_32s_32s_32_7_1_U5.din1_cast_array[5] [4:0];
always @(posedge \shl_4s_1ns_4_7_1_U11.clk )
\shl_4s_1ns_4_7_1_U11.dout_array[5]  <= _0312_;
always @(posedge \shl_4s_1ns_4_7_1_U11.clk )
\shl_4s_1ns_4_7_1_U11.din1_cast_array[5]  <= _0306_;
always @(posedge \shl_4s_1ns_4_7_1_U11.clk )
\shl_4s_1ns_4_7_1_U11.dout_array[4]  <= _0311_;
always @(posedge \shl_4s_1ns_4_7_1_U11.clk )
\shl_4s_1ns_4_7_1_U11.din1_cast_array[4]  <= _0305_;
always @(posedge \shl_4s_1ns_4_7_1_U11.clk )
\shl_4s_1ns_4_7_1_U11.dout_array[3]  <= _0310_;
always @(posedge \shl_4s_1ns_4_7_1_U11.clk )
\shl_4s_1ns_4_7_1_U11.din1_cast_array[3]  <= _0304_;
always @(posedge \shl_4s_1ns_4_7_1_U11.clk )
\shl_4s_1ns_4_7_1_U11.dout_array[2]  <= _0309_;
always @(posedge \shl_4s_1ns_4_7_1_U11.clk )
\shl_4s_1ns_4_7_1_U11.din1_cast_array[2]  <= _0303_;
always @(posedge \shl_4s_1ns_4_7_1_U11.clk )
\shl_4s_1ns_4_7_1_U11.dout_array[1]  <= _0308_;
always @(posedge \shl_4s_1ns_4_7_1_U11.clk )
\shl_4s_1ns_4_7_1_U11.din1_cast_array[1]  <= _0302_;
always @(posedge \shl_4s_1ns_4_7_1_U11.clk )
\shl_4s_1ns_4_7_1_U11.dout_array[0]  <= _0307_;
always @(posedge \shl_4s_1ns_4_7_1_U11.clk )
\shl_4s_1ns_4_7_1_U11.din1_cast_array[0]  <= _0301_;
assign _0313_ = \shl_4s_1ns_4_7_1_U11.ce  ? \shl_4s_1ns_4_7_1_U11.dout_array[1]  : \shl_4s_1ns_4_7_1_U11.dout_array[2] ;
assign _0309_ = \shl_4s_1ns_4_7_1_U11.reset  ? 4'h0 : _0313_;
assign _0314_ = \shl_4s_1ns_4_7_1_U11.ce  ? \shl_4s_1ns_4_7_1_U11.din1_cast_array[0]  : \shl_4s_1ns_4_7_1_U11.din1_cast_array[1] ;
assign _0302_ = \shl_4s_1ns_4_7_1_U11.reset  ? 1'h0 : _0314_;
assign _0315_ = \shl_4s_1ns_4_7_1_U11.ce  ? \shl_4s_1ns_4_7_1_U11.dout_array[0]  : \shl_4s_1ns_4_7_1_U11.dout_array[1] ;
assign _0308_ = \shl_4s_1ns_4_7_1_U11.reset  ? 4'h0 : _0315_;
assign _0316_ = \shl_4s_1ns_4_7_1_U11.ce  ? \shl_4s_1ns_4_7_1_U11.din1 [0] : \shl_4s_1ns_4_7_1_U11.din1_cast_array[0] ;
assign _0301_ = \shl_4s_1ns_4_7_1_U11.reset  ? 1'h0 : _0316_;
assign _0317_ = \shl_4s_1ns_4_7_1_U11.ce  ? \shl_4s_1ns_4_7_1_U11.din0  : \shl_4s_1ns_4_7_1_U11.dout_array[0] ;
assign _0307_ = \shl_4s_1ns_4_7_1_U11.reset  ? 4'h0 : _0317_;
assign _0318_ = \shl_4s_1ns_4_7_1_U11.ce  ? \shl_4s_1ns_4_7_1_U11.din1_cast_array[4]  : \shl_4s_1ns_4_7_1_U11.din1_cast_array[5] ;
assign _0306_ = \shl_4s_1ns_4_7_1_U11.reset  ? 1'h0 : _0318_;
assign _0319_ = \shl_4s_1ns_4_7_1_U11.ce  ? \shl_4s_1ns_4_7_1_U11.dout_array[4]  : \shl_4s_1ns_4_7_1_U11.dout_array[5] ;
assign _0312_ = \shl_4s_1ns_4_7_1_U11.reset  ? 4'h0 : _0319_;
assign _0320_ = \shl_4s_1ns_4_7_1_U11.ce  ? \shl_4s_1ns_4_7_1_U11.din1_cast_array[3]  : \shl_4s_1ns_4_7_1_U11.din1_cast_array[4] ;
assign _0305_ = \shl_4s_1ns_4_7_1_U11.reset  ? 1'h0 : _0320_;
assign _0321_ = \shl_4s_1ns_4_7_1_U11.ce  ? \shl_4s_1ns_4_7_1_U11.dout_array[3]  : \shl_4s_1ns_4_7_1_U11.dout_array[4] ;
assign _0311_ = \shl_4s_1ns_4_7_1_U11.reset  ? 4'h0 : _0321_;
assign _0322_ = \shl_4s_1ns_4_7_1_U11.ce  ? \shl_4s_1ns_4_7_1_U11.din1_cast_array[2]  : \shl_4s_1ns_4_7_1_U11.din1_cast_array[3] ;
assign _0304_ = \shl_4s_1ns_4_7_1_U11.reset  ? 1'h0 : _0322_;
assign _0323_ = \shl_4s_1ns_4_7_1_U11.ce  ? \shl_4s_1ns_4_7_1_U11.dout_array[2]  : \shl_4s_1ns_4_7_1_U11.dout_array[3] ;
assign _0310_ = \shl_4s_1ns_4_7_1_U11.reset  ? 4'h0 : _0323_;
assign _0324_ = \shl_4s_1ns_4_7_1_U11.ce  ? \shl_4s_1ns_4_7_1_U11.din1_cast_array[1]  : \shl_4s_1ns_4_7_1_U11.din1_cast_array[2] ;
assign _0303_ = \shl_4s_1ns_4_7_1_U11.reset  ? 1'h0 : _0324_;
assign \shl_4s_1ns_4_7_1_U11.dout  = \shl_4s_1ns_4_7_1_U11.dout_array[5]  << \shl_4s_1ns_4_7_1_U11.din1_cast_array[5] ;
assign \sub_7s_7ns_7_2_1_U15.top_sub_7s_7ns_7_2_1_Adder_8_U.bin_s0  = ~ \sub_7s_7ns_7_2_1_U15.top_sub_7s_7ns_7_2_1_Adder_8_U.b ;
always @(posedge \sub_7s_7ns_7_2_1_U15.top_sub_7s_7ns_7_2_1_Adder_8_U.clk )
\sub_7s_7ns_7_2_1_U15.top_sub_7s_7ns_7_2_1_Adder_8_U.bin_s1  <= _0326_;
always @(posedge \sub_7s_7ns_7_2_1_U15.top_sub_7s_7ns_7_2_1_Adder_8_U.clk )
\sub_7s_7ns_7_2_1_U15.top_sub_7s_7ns_7_2_1_Adder_8_U.ain_s1  <= _0325_;
always @(posedge \sub_7s_7ns_7_2_1_U15.top_sub_7s_7ns_7_2_1_Adder_8_U.clk )
\sub_7s_7ns_7_2_1_U15.top_sub_7s_7ns_7_2_1_Adder_8_U.sum_s1  <= _0328_;
always @(posedge \sub_7s_7ns_7_2_1_U15.top_sub_7s_7ns_7_2_1_Adder_8_U.clk )
\sub_7s_7ns_7_2_1_U15.top_sub_7s_7ns_7_2_1_Adder_8_U.carry_s1  <= _0327_;
assign _0326_ = \sub_7s_7ns_7_2_1_U15.top_sub_7s_7ns_7_2_1_Adder_8_U.ce  ? \sub_7s_7ns_7_2_1_U15.top_sub_7s_7ns_7_2_1_Adder_8_U.bin_s0 [6:3] : \sub_7s_7ns_7_2_1_U15.top_sub_7s_7ns_7_2_1_Adder_8_U.bin_s1 ;
assign _0325_ = \sub_7s_7ns_7_2_1_U15.top_sub_7s_7ns_7_2_1_Adder_8_U.ce  ? \sub_7s_7ns_7_2_1_U15.top_sub_7s_7ns_7_2_1_Adder_8_U.a [6:3] : \sub_7s_7ns_7_2_1_U15.top_sub_7s_7ns_7_2_1_Adder_8_U.ain_s1 ;
assign _0327_ = \sub_7s_7ns_7_2_1_U15.top_sub_7s_7ns_7_2_1_Adder_8_U.ce  ? \sub_7s_7ns_7_2_1_U15.top_sub_7s_7ns_7_2_1_Adder_8_U.facout_s1  : \sub_7s_7ns_7_2_1_U15.top_sub_7s_7ns_7_2_1_Adder_8_U.carry_s1 ;
assign _0328_ = \sub_7s_7ns_7_2_1_U15.top_sub_7s_7ns_7_2_1_Adder_8_U.ce  ? \sub_7s_7ns_7_2_1_U15.top_sub_7s_7ns_7_2_1_Adder_8_U.fas_s1  : \sub_7s_7ns_7_2_1_U15.top_sub_7s_7ns_7_2_1_Adder_8_U.sum_s1 ;
assign _0329_ = \sub_7s_7ns_7_2_1_U15.top_sub_7s_7ns_7_2_1_Adder_8_U.u1.a  + \sub_7s_7ns_7_2_1_U15.top_sub_7s_7ns_7_2_1_Adder_8_U.u1.b ;
assign { \sub_7s_7ns_7_2_1_U15.top_sub_7s_7ns_7_2_1_Adder_8_U.u1.cout , \sub_7s_7ns_7_2_1_U15.top_sub_7s_7ns_7_2_1_Adder_8_U.u1.s  } = _0329_ + \sub_7s_7ns_7_2_1_U15.top_sub_7s_7ns_7_2_1_Adder_8_U.u1.cin ;
assign _0330_ = \sub_7s_7ns_7_2_1_U15.top_sub_7s_7ns_7_2_1_Adder_8_U.u2.a  + \sub_7s_7ns_7_2_1_U15.top_sub_7s_7ns_7_2_1_Adder_8_U.u2.b ;
assign { \sub_7s_7ns_7_2_1_U15.top_sub_7s_7ns_7_2_1_Adder_8_U.u2.cout , \sub_7s_7ns_7_2_1_U15.top_sub_7s_7ns_7_2_1_Adder_8_U.u2.s  } = _0330_ + \sub_7s_7ns_7_2_1_U15.top_sub_7s_7ns_7_2_1_Adder_8_U.u2.cin ;
assign \sub_9ns_9s_9_2_1_U2.top_sub_9ns_9s_9_2_1_Adder_1_U.bin_s0  = ~ \sub_9ns_9s_9_2_1_U2.top_sub_9ns_9s_9_2_1_Adder_1_U.b ;
always @(posedge \sub_9ns_9s_9_2_1_U2.top_sub_9ns_9s_9_2_1_Adder_1_U.clk )
\sub_9ns_9s_9_2_1_U2.top_sub_9ns_9s_9_2_1_Adder_1_U.bin_s1  <= _0332_;
always @(posedge \sub_9ns_9s_9_2_1_U2.top_sub_9ns_9s_9_2_1_Adder_1_U.clk )
\sub_9ns_9s_9_2_1_U2.top_sub_9ns_9s_9_2_1_Adder_1_U.ain_s1  <= _0331_;
always @(posedge \sub_9ns_9s_9_2_1_U2.top_sub_9ns_9s_9_2_1_Adder_1_U.clk )
\sub_9ns_9s_9_2_1_U2.top_sub_9ns_9s_9_2_1_Adder_1_U.sum_s1  <= _0334_;
always @(posedge \sub_9ns_9s_9_2_1_U2.top_sub_9ns_9s_9_2_1_Adder_1_U.clk )
\sub_9ns_9s_9_2_1_U2.top_sub_9ns_9s_9_2_1_Adder_1_U.carry_s1  <= _0333_;
assign _0332_ = \sub_9ns_9s_9_2_1_U2.top_sub_9ns_9s_9_2_1_Adder_1_U.ce  ? \sub_9ns_9s_9_2_1_U2.top_sub_9ns_9s_9_2_1_Adder_1_U.bin_s0 [8:4] : \sub_9ns_9s_9_2_1_U2.top_sub_9ns_9s_9_2_1_Adder_1_U.bin_s1 ;
assign _0331_ = \sub_9ns_9s_9_2_1_U2.top_sub_9ns_9s_9_2_1_Adder_1_U.ce  ? \sub_9ns_9s_9_2_1_U2.top_sub_9ns_9s_9_2_1_Adder_1_U.a [8:4] : \sub_9ns_9s_9_2_1_U2.top_sub_9ns_9s_9_2_1_Adder_1_U.ain_s1 ;
assign _0333_ = \sub_9ns_9s_9_2_1_U2.top_sub_9ns_9s_9_2_1_Adder_1_U.ce  ? \sub_9ns_9s_9_2_1_U2.top_sub_9ns_9s_9_2_1_Adder_1_U.facout_s1  : \sub_9ns_9s_9_2_1_U2.top_sub_9ns_9s_9_2_1_Adder_1_U.carry_s1 ;
assign _0334_ = \sub_9ns_9s_9_2_1_U2.top_sub_9ns_9s_9_2_1_Adder_1_U.ce  ? \sub_9ns_9s_9_2_1_U2.top_sub_9ns_9s_9_2_1_Adder_1_U.fas_s1  : \sub_9ns_9s_9_2_1_U2.top_sub_9ns_9s_9_2_1_Adder_1_U.sum_s1 ;
assign _0335_ = \sub_9ns_9s_9_2_1_U2.top_sub_9ns_9s_9_2_1_Adder_1_U.u1.a  + \sub_9ns_9s_9_2_1_U2.top_sub_9ns_9s_9_2_1_Adder_1_U.u1.b ;
assign { \sub_9ns_9s_9_2_1_U2.top_sub_9ns_9s_9_2_1_Adder_1_U.u1.cout , \sub_9ns_9s_9_2_1_U2.top_sub_9ns_9s_9_2_1_Adder_1_U.u1.s  } = _0335_ + \sub_9ns_9s_9_2_1_U2.top_sub_9ns_9s_9_2_1_Adder_1_U.u1.cin ;
assign _0336_ = \sub_9ns_9s_9_2_1_U2.top_sub_9ns_9s_9_2_1_Adder_1_U.u2.a  + \sub_9ns_9s_9_2_1_U2.top_sub_9ns_9s_9_2_1_Adder_1_U.u2.b ;
assign { \sub_9ns_9s_9_2_1_U2.top_sub_9ns_9s_9_2_1_Adder_1_U.u2.cout , \sub_9ns_9s_9_2_1_U2.top_sub_9ns_9s_9_2_1_Adder_1_U.u2.s  } = _0336_ + \sub_9ns_9s_9_2_1_U2.top_sub_9ns_9s_9_2_1_Adder_1_U.u2.cin ;
assign _0337_ = | { and_ln414_fu_1145_p2[1], r_V_2_reg_2028[0] };
assign _0338_ = | { tmp_4_reg_1688, 2'h0, p_Result_s_22_reg_1694 };
assign _0339_ = p_Result_s_22_reg_1694 != 5'h1f;
assign _0340_ = | { trunc_ln851_3_reg_1828, 15'h0000 };
assign _0341_ = | { trunc_ln851_5_reg_2102, 1'h0 };
assign _0342_ = { op_0, 8'h00 } != op_1;
assign _0343_ = op_2_V_reg_1741 != { rhs_1_reg_1590, 5'h00 };
assign op_12_V_fu_606_p2 = op_4[3:0] | ret_V_21_reg_1661;
assign or_ln1195_1_fu_643_p2 = { trunc_ln1195_reg_1757, 3'h0 } | op_5;
assign or_ln1195_fu_629_p2 = { op_5[3], op_5 } | { ret_reg_1752, 3'h0 };
assign or_ln384_1_fu_956_p2 = underflow_1_fu_951_p2 | overflow_1_reg_1925;
assign or_ln384_fu_506_p2 = underflow_fu_501_p2 | overflow_reg_1720;
assign or_ln410_fu_1291_p2 = xor_ln410_reg_2107 | r_V_1_reg_2070[0];
assign or_ln412_fu_703_p2 = or_ln1195_reg_1794[0] | or_ln1195_1_reg_1806[2];
assign or_ln785_fu_897_p2 = xor_ln785_2_fu_891_p2 | p_Result_32_reg_1879;
assign or_ln788_1_fu_496_p2 = or_ln788_fu_492_p2 | icmp_ln786_reg_1726;
assign or_ln788_2_fu_940_p2 = and_ln788_1_reg_1931 | and_ln781_fu_936_p2;
assign or_ln788_fu_492_p2 = icmp_ln790_reg_1715 | icmp_ln786_1_reg_1710;
always @(posedge ap_clk)
ret_V_5_reg_1779[4:0] <= 5'h00;
always @(posedge ap_clk)
trunc_ln851_3_reg_1828 <= 5'h00;
always @(posedge ap_clk)
tmp_1_reg_1858 <= _0087_;
always @(posedge ap_clk)
sub_ln1497_reg_1635 <= _0086_;
always @(posedge ap_clk)
shl_ln1497_reg_1672 <= _0084_;
always @(posedge ap_clk)
ret_V_7_reg_1640 <= _0073_;
always @(posedge ap_clk)
ret_V_28_reg_2267 <= _0068_;
always @(posedge ap_clk)
ret_V_28_cast_reg_2272 <= _0067_;
always @(posedge ap_clk)
ret_V_27_reg_2242 <= _0066_;
always @(posedge ap_clk)
ret_V_26_reg_2225 <= _0065_;
always @(posedge ap_clk)
ret_V_25_cast_reg_2230 <= _0063_;
always @(posedge ap_clk)
ret_V_21_reg_1661 <= _0058_;
always @(posedge ap_clk)
ret_V_2_reg_1597 <= _0069_;
always @(posedge ap_clk)
tmp_reg_1603 <= _0090_;
always @(posedge ap_clk)
ret_V_20_reg_1608 <= _0057_;
always @(posedge ap_clk)
ret_V_8_cast_reg_1613 <= _0074_;
always @(posedge ap_clk)
trunc_ln851_2_reg_1620 <= _0097_;
always @(posedge ap_clk)
ret_V_1_reg_1585 <= _0056_;
always @(posedge ap_clk)
rhs_1_reg_1590 <= _0078_;
always @(posedge ap_clk)
r_V_reg_1979 <= _0053_;
always @(posedge ap_clk)
ret_V_3_cast_reg_1984 <= _0070_;
always @(posedge ap_clk)
trunc_ln851_1_reg_1991 <= _0096_;
always @(posedge ap_clk)
ret_V_23_reg_1996 <= _0061_;
always @(posedge ap_clk)
ret_V_19_cast_reg_2001 <= _0054_;
always @(posedge ap_clk)
p_Val2_9_reg_1873 <= _0050_;
always @(posedge ap_clk)
p_Result_32_reg_1879 <= _0045_;
always @(posedge ap_clk)
ret_V_19_reg_2023 <= _0055_;
always @(posedge ap_clk)
r_V_2_reg_2028 <= _0052_;
always @(posedge ap_clk)
p_Result_27_reg_2034 <= _0042_;
always @(posedge ap_clk)
trunc_ln708_1_reg_2040 <= _0094_;
always @(posedge ap_clk)
ret_V_24_reg_2045 <= _0062_;
always @(posedge ap_clk)
select_ln1497_reg_1677 <= _0079_;
always @(posedge ap_clk)
p_Result_23_reg_1682 <= _0039_;
always @(posedge ap_clk)
tmp_4_reg_1688 <= _0089_;
always @(posedge ap_clk)
p_Result_s_22_reg_1694 <= _0046_;
always @(posedge ap_clk)
trunc_ln790_reg_1700 <= _0095_;
always @(posedge ap_clk)
or_ln384_reg_1731 <= _0036_;
always @(posedge ap_clk)
or_ln384_1_reg_1943 <= _0035_;
always @(posedge ap_clk)
op_2_V_reg_1741 <= _0032_;
always @(posedge ap_clk)
trunc_ln8_reg_1747 <= _0099_;
always @(posedge ap_clk)
ret_reg_1752 <= _0077_;
always @(posedge ap_clk)
trunc_ln1195_reg_1757 <= _0092_;
always @(posedge ap_clk)
op_26_V_reg_2252 <= _0031_;
always @(posedge ap_clk)
p_Val2_4_reg_2182 <= _0047_;
always @(posedge ap_clk)
p_Result_26_reg_2187 <= _0041_;
always @(posedge ap_clk)
op_19_V_reg_2193 <= _0029_;
always @(posedge ap_clk)
op_17_V_reg_2204 <= _0028_;
always @(posedge ap_clk)
select_ln353_2_reg_2210 <= _0080_;
always @(posedge ap_clk)
op_14_V_reg_1953 <= _0027_;
always @(posedge ap_clk)
select_ln353_reg_1959 <= _0081_;
always @(posedge ap_clk)
ret_V_reg_1568 <= _0076_;
always @(posedge ap_clk)
icmp_ln851_reg_1575 <= _0025_;
always @(posedge ap_clk)
xor_ln410_reg_2107 <= _0101_;
always @(posedge ap_clk)
icmp_ln851_4_reg_2133 <= _0024_;
always @(posedge ap_clk)
icmp_ln851_2_reg_1630 <= _0022_;
always @(posedge ap_clk)
icmp_ln851_1_reg_2008 <= _0021_;
always @(posedge ap_clk)
overflow_reg_1720 <= _0038_;
always @(posedge ap_clk)
icmp_ln786_reg_1726 <= _0019_;
always @(posedge ap_clk)
icmp_ln785_reg_1705 <= _0017_;
always @(posedge ap_clk)
icmp_ln786_1_reg_1710 <= _0018_;
always @(posedge ap_clk)
icmp_ln790_reg_1715 <= _0020_;
always @(posedge ap_clk)
icmp_ln414_reg_2050 <= _0016_;
always @(posedge ap_clk)
ashr_ln1497_reg_1667 <= _0014_;
always @(posedge ap_clk)
overflow_1_reg_1925 <= _0037_;
always @(posedge ap_clk)
and_ln788_1_reg_1931 <= _0012_;
always @(posedge ap_clk)
sext_ln850_reg_1936 <= _0083_;
always @(posedge ap_clk)
r_V_1_reg_2070 <= _0051_;
always @(posedge ap_clk)
p_Result_24_reg_2076 <= _0040_;
always @(posedge ap_clk)
trunc_ln1_reg_2082 <= _0093_;
always @(posedge ap_clk)
and_ln414_1_reg_2087 <= _0011_;
always @(posedge ap_clk)
ret_V_9_reg_2092 <= _0075_;
always @(posedge ap_clk)
op_23_V_reg_2097 <= _0030_;
always @(posedge ap_clk)
trunc_ln851_5_reg_2102 <= _0098_;
always @(posedge ap_clk)
and_ln412_reg_1833 <= _0010_;
always @(posedge ap_clk)
icmp_ln851_3_reg_1848 <= _0023_;
always @(posedge ap_clk)
and_ln410_reg_2138 <= _0009_;
always @(posedge ap_clk)
p_Val2_6_reg_2143 <= _0048_;
always @(posedge ap_clk)
p_Result_28_reg_2149 <= _0043_;
always @(posedge ap_clk)
ret_V_25_reg_2155 <= _0064_;
always @(posedge ap_clk)
ret_V_22_cast_reg_2160 <= _0059_;
always @(posedge ap_clk)
sext_ln745_reg_2172 <= _0082_;
always @(posedge ap_clk)
and_ln340_reg_2177 <= _0008_;
always @(posedge ap_clk)
add_ln691_reg_1948 <= _0007_;
always @(posedge ap_clk)
add_ln691_4_reg_2279 <= _0006_;
always @(posedge ap_clk)
add_ln691_3_reg_2237 <= _0005_;
always @(posedge ap_clk)
add_ln691_2_reg_2199 <= _0004_;
always @(posedge ap_clk)
ret_V_3_reg_2013 <= _0071_;
always @(posedge ap_clk)
add_ln691_1_reg_2018 <= _0003_;
always @(posedge ap_clk)
ush_reg_1772 <= _0100_;
always @(posedge ap_clk)
ret_V_5_reg_1779[6:5] <= _0072_;
always @(posedge ap_clk)
signbit_reg_1784 <= _0085_;
always @(posedge ap_clk)
op_12_V_reg_1789 <= _0026_;
always @(posedge ap_clk)
or_ln1195_reg_1794 <= _0034_;
always @(posedge ap_clk)
Range2_all_ones_reg_1800 <= _0002_;
always @(posedge ap_clk)
or_ln1195_1_reg_1806 <= _0033_;
always @(posedge ap_clk)
p_Result_29_reg_1812 <= _0044_;
always @(posedge ap_clk)
p_Val2_8_reg_1818 <= _0049_;
always @(posedge ap_clk)
tmp_23_reg_1823 <= _0088_;
always @(posedge ap_clk)
carry_1_reg_1896 <= _0015_;
always @(posedge ap_clk)
Range1_all_ones_reg_1903 <= _0000_;
always @(posedge ap_clk)
Range1_all_zeros_reg_1910 <= _0001_;
always @(posedge ap_clk)
ret_V_22_reg_1915 <= _0060_;
always @(posedge ap_clk)
tmp_s_reg_1920 <= _0091_;
always @(posedge ap_clk)
ap_CS_fsm <= _0013_;
assign _0102_ = _0109_ ? 2'h2 : 2'h1;
assign _0344_ = ap_CS_fsm == 1'h1;
function [48:0] _0954_;
input [48:0] a;
input [2400:0] b;
input [48:0] s;
case (s)
49'b0000000000000000000000000000000000000000000000001:
_0954_ = b[48:0];
49'b0000000000000000000000000000000000000000000000010:
_0954_ = b[97:49];
49'b0000000000000000000000000000000000000000000000100:
_0954_ = b[146:98];
49'b0000000000000000000000000000000000000000000001000:
_0954_ = b[195:147];
49'b0000000000000000000000000000000000000000000010000:
_0954_ = b[244:196];
49'b0000000000000000000000000000000000000000000100000:
_0954_ = b[293:245];
49'b0000000000000000000000000000000000000000001000000:
_0954_ = b[342:294];
49'b0000000000000000000000000000000000000000010000000:
_0954_ = b[391:343];
49'b0000000000000000000000000000000000000000100000000:
_0954_ = b[440:392];
49'b0000000000000000000000000000000000000001000000000:
_0954_ = b[489:441];
49'b0000000000000000000000000000000000000010000000000:
_0954_ = b[538:490];
49'b0000000000000000000000000000000000000100000000000:
_0954_ = b[587:539];
49'b0000000000000000000000000000000000001000000000000:
_0954_ = b[636:588];
49'b0000000000000000000000000000000000010000000000000:
_0954_ = b[685:637];
49'b0000000000000000000000000000000000100000000000000:
_0954_ = b[734:686];
49'b0000000000000000000000000000000001000000000000000:
_0954_ = b[783:735];
49'b0000000000000000000000000000000010000000000000000:
_0954_ = b[832:784];
49'b0000000000000000000000000000000100000000000000000:
_0954_ = b[881:833];
49'b0000000000000000000000000000001000000000000000000:
_0954_ = b[930:882];
49'b0000000000000000000000000000010000000000000000000:
_0954_ = b[979:931];
49'b0000000000000000000000000000100000000000000000000:
_0954_ = b[1028:980];
49'b0000000000000000000000000001000000000000000000000:
_0954_ = b[1077:1029];
49'b0000000000000000000000000010000000000000000000000:
_0954_ = b[1126:1078];
49'b0000000000000000000000000100000000000000000000000:
_0954_ = b[1175:1127];
49'b0000000000000000000000001000000000000000000000000:
_0954_ = b[1224:1176];
49'b0000000000000000000000010000000000000000000000000:
_0954_ = b[1273:1225];
49'b0000000000000000000000100000000000000000000000000:
_0954_ = b[1322:1274];
49'b0000000000000000000001000000000000000000000000000:
_0954_ = b[1371:1323];
49'b0000000000000000000010000000000000000000000000000:
_0954_ = b[1420:1372];
49'b0000000000000000000100000000000000000000000000000:
_0954_ = b[1469:1421];
49'b0000000000000000001000000000000000000000000000000:
_0954_ = b[1518:1470];
49'b0000000000000000010000000000000000000000000000000:
_0954_ = b[1567:1519];
49'b0000000000000000100000000000000000000000000000000:
_0954_ = b[1616:1568];
49'b0000000000000001000000000000000000000000000000000:
_0954_ = b[1665:1617];
49'b0000000000000010000000000000000000000000000000000:
_0954_ = b[1714:1666];
49'b0000000000000100000000000000000000000000000000000:
_0954_ = b[1763:1715];
49'b0000000000001000000000000000000000000000000000000:
_0954_ = b[1812:1764];
49'b0000000000010000000000000000000000000000000000000:
_0954_ = b[1861:1813];
49'b0000000000100000000000000000000000000000000000000:
_0954_ = b[1910:1862];
49'b0000000001000000000000000000000000000000000000000:
_0954_ = b[1959:1911];
49'b0000000010000000000000000000000000000000000000000:
_0954_ = b[2008:1960];
49'b0000000100000000000000000000000000000000000000000:
_0954_ = b[2057:2009];
49'b0000001000000000000000000000000000000000000000000:
_0954_ = b[2106:2058];
49'b0000010000000000000000000000000000000000000000000:
_0954_ = b[2155:2107];
49'b0000100000000000000000000000000000000000000000000:
_0954_ = b[2204:2156];
49'b0001000000000000000000000000000000000000000000000:
_0954_ = b[2253:2205];
49'b0010000000000000000000000000000000000000000000000:
_0954_ = b[2302:2254];
49'b0100000000000000000000000000000000000000000000000:
_0954_ = b[2351:2303];
49'b1000000000000000000000000000000000000000000000000:
_0954_ = b[2400:2352];
49'b0000000000000000000000000000000000000000000000000:
_0954_ = a;
default:
_0954_ = 49'bx;
endcase
endfunction
assign ap_NS_fsm = _0954_(49'hxxxxxxxxxxxxx, { 47'h000000000000, _0102_, 2352'h000000000002000000000002000000000002000000000002000000000002000000000002000000000002000000000002000000000002000000000002000000000002000000000002000000000002000000000002000000000002000000000002000000000002000000000002000000000002000000000002000000000002000000000002000000000002000000000002000000000002000000000002000000000002000000000002000000000002000000000002000000000002000000000002000000000002000000000002000000000002000000000002000000000002000000000002000000000002000000000002000000000002000000000002000000000002000000000002000000000002000000000002000000000002000000000000000000000001 }, { _0344_, _0392_, _0391_, _0390_, _0389_, _0388_, _0387_, _0386_, _0385_, _0384_, _0383_, _0382_, _0381_, _0380_, _0379_, _0378_, _0377_, _0376_, _0375_, _0374_, _0373_, _0372_, _0371_, _0370_, _0369_, _0368_, _0367_, _0366_, _0365_, _0364_, _0363_, _0362_, _0361_, _0360_, _0359_, _0358_, _0357_, _0356_, _0355_, _0354_, _0353_, _0352_, _0351_, _0350_, _0349_, _0348_, _0347_, _0346_, _0345_ });
assign _0345_ = ap_CS_fsm == 49'h1000000000000;
assign _0346_ = ap_CS_fsm == 48'h800000000000;
assign _0347_ = ap_CS_fsm == 47'h400000000000;
assign _0348_ = ap_CS_fsm == 46'h200000000000;
assign _0349_ = ap_CS_fsm == 45'h100000000000;
assign _0350_ = ap_CS_fsm == 44'h80000000000;
assign _0351_ = ap_CS_fsm == 43'h40000000000;
assign _0352_ = ap_CS_fsm == 42'h20000000000;
assign _0353_ = ap_CS_fsm == 41'h10000000000;
assign _0354_ = ap_CS_fsm == 40'h8000000000;
assign _0355_ = ap_CS_fsm == 39'h4000000000;
assign _0356_ = ap_CS_fsm == 38'h2000000000;
assign _0357_ = ap_CS_fsm == 37'h1000000000;
assign _0358_ = ap_CS_fsm == 36'h800000000;
assign _0359_ = ap_CS_fsm == 35'h400000000;
assign _0360_ = ap_CS_fsm == 34'h200000000;
assign _0361_ = ap_CS_fsm == 33'h100000000;
assign _0362_ = ap_CS_fsm == 32'd2147483648;
assign _0363_ = ap_CS_fsm == 31'h40000000;
assign _0364_ = ap_CS_fsm == 30'h20000000;
assign _0365_ = ap_CS_fsm == 29'h10000000;
assign _0366_ = ap_CS_fsm == 28'h8000000;
assign _0367_ = ap_CS_fsm == 27'h4000000;
assign _0368_ = ap_CS_fsm == 26'h2000000;
assign _0369_ = ap_CS_fsm == 25'h1000000;
assign _0370_ = ap_CS_fsm == 24'h800000;
assign _0371_ = ap_CS_fsm == 23'h400000;
assign _0372_ = ap_CS_fsm == 22'h200000;
assign _0373_ = ap_CS_fsm == 21'h100000;
assign _0374_ = ap_CS_fsm == 20'h80000;
assign _0375_ = ap_CS_fsm == 19'h40000;
assign _0376_ = ap_CS_fsm == 18'h20000;
assign _0377_ = ap_CS_fsm == 17'h10000;
assign _0378_ = ap_CS_fsm == 16'h8000;
assign _0379_ = ap_CS_fsm == 15'h4000;
assign _0380_ = ap_CS_fsm == 14'h2000;
assign _0381_ = ap_CS_fsm == 13'h1000;
assign _0382_ = ap_CS_fsm == 12'h800;
assign _0383_ = ap_CS_fsm == 11'h400;
assign _0384_ = ap_CS_fsm == 10'h200;
assign _0385_ = ap_CS_fsm == 9'h100;
assign _0386_ = ap_CS_fsm == 8'h80;
assign _0387_ = ap_CS_fsm == 7'h40;
assign _0388_ = ap_CS_fsm == 6'h20;
assign _0389_ = ap_CS_fsm == 5'h10;
assign _0390_ = ap_CS_fsm == 4'h8;
assign _0391_ = ap_CS_fsm == 3'h4;
assign _0392_ = ap_CS_fsm == 2'h2;
assign op_27_ap_vld = ap_CS_fsm[48] ? 1'h1 : 1'h0;
assign ap_idle = _0108_ ? 1'h1 : 1'h0;
assign _0087_ = ap_CS_fsm[19] ? grp_fu_730_p2[6:2] : tmp_1_reg_1858;
assign _0086_ = _0107_ ? grp_fu_346_p2 : sub_ln1497_reg_1635;
assign _0084_ = _0106_ ? grp_fu_377_p2 : shl_ln1497_reg_1672;
assign _0073_ = ap_CS_fsm[4] ? grp_fu_357_p2 : ret_V_7_reg_1640;
assign _0067_ = ap_CS_fsm[45] ? grp_fu_1516_p2[32:1] : ret_V_28_cast_reg_2272;
assign _0068_ = ap_CS_fsm[45] ? grp_fu_1516_p2 : ret_V_28_reg_2267;
assign _0066_ = ap_CS_fsm[41] ? ret_V_27_fu_1486_p3 : ret_V_27_reg_2242;
assign _0063_ = ap_CS_fsm[38] ? grp_fu_1449_p2[32:1] : ret_V_25_cast_reg_2230;
assign _0065_ = ap_CS_fsm[38] ? grp_fu_1449_p2 : ret_V_26_reg_2225;
assign _0058_ = ap_CS_fsm[5] ? ret_V_21_fu_395_p3 : ret_V_21_reg_1661;
assign _0097_ = ap_CS_fsm[2] ? ret_V_20_fu_324_p2[7:0] : trunc_ln851_2_reg_1620;
assign _0074_ = ap_CS_fsm[2] ? ret_V_20_fu_324_p2[11:8] : ret_V_8_cast_reg_1613;
assign _0057_ = ap_CS_fsm[2] ? ret_V_20_fu_324_p2 : ret_V_20_reg_1608;
assign _0090_ = ap_CS_fsm[2] ? ret_V_2_fu_298_p3[7] : tmp_reg_1603;
assign _0069_ = ap_CS_fsm[2] ? ret_V_2_fu_298_p3 : ret_V_2_reg_1597;
assign _0078_ = ap_CS_fsm[1] ? rhs_1_fu_281_p2 : rhs_1_reg_1590;
assign _0056_ = ap_CS_fsm[1] ? grp_fu_267_p2 : ret_V_1_reg_1585;
assign _0054_ = ap_CS_fsm[26] ? grp_fu_1015_p2[32:1] : ret_V_19_cast_reg_2001;
assign _0061_ = ap_CS_fsm[26] ? grp_fu_1015_p2 : ret_V_23_reg_1996;
assign _0096_ = ap_CS_fsm[26] ? grp_fu_774_p2[2:0] : trunc_ln851_1_reg_1991;
assign _0070_ = ap_CS_fsm[26] ? grp_fu_774_p2[4:3] : ret_V_3_cast_reg_1984;
assign _0053_ = ap_CS_fsm[26] ? grp_fu_774_p2 : r_V_reg_1979;
assign _0045_ = ap_CS_fsm[20] ? grp_fu_752_p2[1] : p_Result_32_reg_1879;
assign _0050_ = ap_CS_fsm[20] ? grp_fu_752_p2 : p_Val2_9_reg_1873;
assign _0062_ = ap_CS_fsm[29] ? ret_V_24_fu_1125_p3 : ret_V_24_reg_2045;
assign _0094_ = ap_CS_fsm[29] ? r_V_2_fu_1086_p2[3:2] : trunc_ln708_1_reg_2040;
assign _0042_ = ap_CS_fsm[29] ? r_V_2_fu_1086_p2[3] : p_Result_27_reg_2034;
assign _0052_ = ap_CS_fsm[29] ? r_V_2_fu_1086_p2 : r_V_2_reg_2028;
assign _0055_ = ap_CS_fsm[29] ? ret_V_19_fu_1072_p3 : ret_V_19_reg_2023;
assign _0095_ = ap_CS_fsm[12] ? select_ln1497_fu_402_p3[1:0] : trunc_ln790_reg_1700;
assign _0046_ = ap_CS_fsm[12] ? select_ln1497_fu_402_p3[7:3] : p_Result_s_22_reg_1694;
assign _0089_ = ap_CS_fsm[12] ? select_ln1497_fu_402_p3[2] : tmp_4_reg_1688;
assign _0039_ = ap_CS_fsm[12] ? select_ln1497_fu_402_p3[7] : p_Result_23_reg_1682;
assign _0079_ = ap_CS_fsm[12] ? select_ln1497_fu_402_p3 : select_ln1497_reg_1677;
assign _0036_ = ap_CS_fsm[15] ? or_ln384_fu_506_p2 : or_ln384_reg_1731;
assign _0035_ = ap_CS_fsm[23] ? or_ln384_1_fu_956_p2 : or_ln384_1_reg_1943;
assign _0092_ = ap_CS_fsm[16] ? ret_fu_547_p2[0] : trunc_ln1195_reg_1757;
assign _0077_ = ap_CS_fsm[16] ? ret_fu_547_p2 : ret_reg_1752;
assign _0099_ = ap_CS_fsm[16] ? op_2_V_fu_529_p3[6:0] : trunc_ln8_reg_1747;
assign _0032_ = ap_CS_fsm[16] ? op_2_V_fu_529_p3 : op_2_V_reg_1741;
assign _0031_ = ap_CS_fsm[43] ? grp_fu_1497_p2 : op_26_V_reg_2252;
assign _0029_ = ap_CS_fsm[35] ? op_19_V_fu_1393_p3 : op_19_V_reg_2193;
assign _0041_ = ap_CS_fsm[35] ? grp_fu_1323_p2[1] : p_Result_26_reg_2187;
assign _0047_ = ap_CS_fsm[35] ? grp_fu_1323_p2 : p_Val2_4_reg_2182;
assign _0080_ = ap_CS_fsm[36] ? select_ln353_2_fu_1428_p3 : select_ln353_2_reg_2210;
assign _0028_ = ap_CS_fsm[36] ? op_17_V_fu_1409_p3 : op_17_V_reg_2204;
assign _0081_ = ap_CS_fsm[24] ? select_ln353_fu_986_p3 : select_ln353_reg_1959;
assign _0027_ = ap_CS_fsm[24] ? op_14_V_fu_968_p3 : op_14_V_reg_1953;
assign _0025_ = ap_CS_fsm[0] ? icmp_ln851_fu_261_p2 : icmp_ln851_reg_1575;
assign _0076_ = ap_CS_fsm[0] ? op_1[15:8] : ret_V_reg_1568;
assign _0024_ = ap_CS_fsm[32] ? icmp_ln851_4_fu_1275_p2 : icmp_ln851_4_reg_2133;
assign _0101_ = ap_CS_fsm[32] ? xor_ln410_fu_1223_p2 : xor_ln410_reg_2107;
assign _0022_ = ap_CS_fsm[3] ? icmp_ln851_2_fu_352_p2 : icmp_ln851_2_reg_1630;
assign _0021_ = ap_CS_fsm[27] ? icmp_ln851_1_fu_1045_p2 : icmp_ln851_1_reg_2008;
assign _0019_ = ap_CS_fsm[14] ? icmp_ln786_fu_486_p2 : icmp_ln786_reg_1726;
assign _0038_ = ap_CS_fsm[14] ? overflow_fu_481_p2 : overflow_reg_1720;
assign _0020_ = ap_CS_fsm[13] ? icmp_ln790_fu_463_p2 : icmp_ln790_reg_1715;
assign _0018_ = ap_CS_fsm[13] ? icmp_ln786_1_fu_451_p2 : icmp_ln786_1_reg_1710;
assign _0017_ = ap_CS_fsm[13] ? icmp_ln785_fu_445_p2 : icmp_ln785_reg_1705;
assign _0016_ = ap_CS_fsm[30] ? icmp_ln414_fu_1167_p2 : icmp_ln414_reg_2050;
assign _0014_ = _0105_ ? grp_fu_368_p2 : ashr_ln1497_reg_1667;
assign _0083_ = ap_CS_fsm[22] ? { tmp_s_reg_1920[5], tmp_s_reg_1920 } : sext_ln850_reg_1936;
assign _0012_ = ap_CS_fsm[22] ? and_ln788_1_fu_922_p2 : and_ln788_1_reg_1931;
assign _0037_ = ap_CS_fsm[22] ? overflow_1_fu_907_p2 : overflow_1_reg_1925;
assign _0098_ = ap_CS_fsm[31] ? grp_fu_1183_p2[2:0] : trunc_ln851_5_reg_2102;
assign _0030_ = ap_CS_fsm[31] ? grp_fu_1192_p2 : op_23_V_reg_2097;
assign _0075_ = ap_CS_fsm[31] ? grp_fu_1183_p2 : ret_V_9_reg_2092;
assign _0011_ = ap_CS_fsm[31] ? and_ln414_1_fu_1215_p2 : and_ln414_1_reg_2087;
assign _0093_ = ap_CS_fsm[31] ? grp_fu_996_p2[3:2] : trunc_ln1_reg_2082;
assign _0040_ = ap_CS_fsm[31] ? grp_fu_996_p2[3] : p_Result_24_reg_2076;
assign _0051_ = ap_CS_fsm[31] ? grp_fu_996_p2 : r_V_1_reg_2070;
assign _0023_ = ap_CS_fsm[18] ? icmp_ln851_3_fu_743_p2 : icmp_ln851_3_reg_1848;
assign _0010_ = ap_CS_fsm[18] ? and_ln412_fu_709_p2 : and_ln412_reg_1833;
assign _0059_ = ap_CS_fsm[33] ? grp_fu_1262_p2[35:4] : ret_V_22_cast_reg_2160;
assign _0064_ = ap_CS_fsm[33] ? grp_fu_1262_p2 : ret_V_25_reg_2155;
assign _0043_ = ap_CS_fsm[33] ? grp_fu_1234_p2[2] : p_Result_28_reg_2149;
assign _0048_ = ap_CS_fsm[33] ? grp_fu_1234_p2 : p_Val2_6_reg_2143;
assign _0009_ = ap_CS_fsm[33] ? and_ln410_fu_1296_p2 : and_ln410_reg_2138;
assign _0008_ = ap_CS_fsm[34] ? and_ln340_fu_1356_p2 : and_ln340_reg_2177;
assign _0082_ = ap_CS_fsm[34] ? { p_Val2_6_reg_2143[2], p_Val2_6_reg_2143 } : sext_ln745_reg_2172;
assign _0007_ = _0104_ ? grp_fu_930_p2 : add_ln691_reg_1948;
assign _0006_ = ap_CS_fsm[47] ? grp_fu_1532_p2 : add_ln691_4_reg_2279;
assign _0005_ = ap_CS_fsm[40] ? grp_fu_1465_p2 : add_ln691_3_reg_2237;
assign _0004_ = _0103_ ? grp_fu_1361_p2 : add_ln691_2_reg_2199;
assign _0003_ = ap_CS_fsm[28] ? grp_fu_1055_p2 : add_ln691_1_reg_2018;
assign _0071_ = ap_CS_fsm[28] ? grp_fu_1050_p2 : ret_V_3_reg_2013;
assign _0088_ = ap_CS_fsm[17] ? or_ln1195_fu_629_p2[4] : tmp_23_reg_1823;
assign _0049_ = ap_CS_fsm[17] ? or_ln1195_1_fu_643_p2[3:2] : p_Val2_8_reg_1818;
assign _0044_ = ap_CS_fsm[17] ? op_5[3] : p_Result_29_reg_1812;
assign _0033_ = ap_CS_fsm[17] ? or_ln1195_1_fu_643_p2 : or_ln1195_1_reg_1806;
assign _0002_ = ap_CS_fsm[17] ? op_5[3] : Range2_all_ones_reg_1800;
assign _0034_ = ap_CS_fsm[17] ? or_ln1195_fu_629_p2 : or_ln1195_reg_1794;
assign _0026_ = ap_CS_fsm[17] ? op_12_V_fu_606_p2 : op_12_V_reg_1789;
assign _0085_ = ap_CS_fsm[17] ? signbit_fu_597_p2 : signbit_reg_1784;
assign _0072_ = ap_CS_fsm[17] ? ret_V_5_fu_581_p2[6:5] : ret_V_5_reg_1779[6:5];
assign _0100_ = ap_CS_fsm[17] ? ush_fu_568_p2 : ush_reg_1772;
assign _0091_ = ap_CS_fsm[21] ? grp_fu_810_p2[25:20] : tmp_s_reg_1920;
assign _0060_ = ap_CS_fsm[21] ? grp_fu_810_p2 : ret_V_22_reg_1915;
assign _0001_ = ap_CS_fsm[21] ? Range1_all_zeros_fu_846_p2 : Range1_all_zeros_reg_1910;
assign _0000_ = ap_CS_fsm[21] ? Range1_all_ones_fu_840_p2 : Range1_all_ones_reg_1903;
assign _0015_ = ap_CS_fsm[21] ? carry_1_fu_828_p2 : carry_1_reg_1896;
assign _0013_ = ap_rst ? 49'h0000000000001 : ap_NS_fsm;
assign Range1_all_ones_fu_840_p2 = _0112_ ? 1'h1 : 1'h0;
assign Range1_all_zeros_fu_846_p2 = _0113_ ? 1'h1 : 1'h0;
assign deleted_ones_fu_885_p3 = carry_1_reg_1896 ? and_ln780_fu_880_p2 : Range1_all_ones_reg_1903;
assign deleted_zeros_fu_862_p3 = carry_1_reg_1896 ? Range1_all_ones_reg_1903 : Range1_all_zeros_reg_1910;
assign icmp_ln414_fu_1167_p2 = _0337_ ? 1'h1 : 1'h0;
assign icmp_ln785_fu_445_p2 = _0338_ ? 1'h1 : 1'h0;
assign icmp_ln786_1_fu_451_p2 = _0339_ ? 1'h1 : 1'h0;
assign icmp_ln786_fu_486_p2 = _0114_ ? 1'h1 : 1'h0;
assign icmp_ln790_fu_463_p2 = _0115_ ? 1'h1 : 1'h0;
assign icmp_ln851_1_fu_1045_p2 = _0116_ ? 1'h1 : 1'h0;
assign icmp_ln851_2_fu_352_p2 = _0117_ ? 1'h1 : 1'h0;
assign icmp_ln851_3_fu_743_p2 = _0340_ ? 1'h1 : 1'h0;
assign icmp_ln851_4_fu_1275_p2 = _0341_ ? 1'h1 : 1'h0;
assign icmp_ln851_fu_261_p2 = _0118_ ? 1'h1 : 1'h0;
assign op_14_V_fu_968_p3 = or_ln384_1_reg_1943 ? select_ln384_fu_961_p3 : p_Val2_9_reg_1873;
assign op_17_V_fu_1409_p3 = select_ln340_fu_1403_p3 ? 2'h0 : p_Val2_4_reg_2182;
assign op_19_V_fu_1393_p3 = and_ln340_reg_2177 ? { 1'h0, p_Val2_7_fu_1374_p2 } : sext_ln745_reg_2172;
assign op_27 = ret_V_28_reg_2267[33] ? select_ln850_7_fu_1547_p3 : ret_V_28_cast_reg_2272;
assign op_2_V_fu_529_p3 = or_ln384_reg_1731 ? select_ln384_1_fu_522_p3 : { select_ln1497_reg_1677[2:0], 5'h00 };
assign ret_V_19_fu_1072_p3 = r_V_reg_1979[5] ? select_ln850_1_fu_1067_p3 : ret_V_3_cast_reg_1984;
assign ret_V_21_fu_395_p3 = ret_V_20_reg_1608[15] ? select_ln850_2_fu_390_p3 : ret_V_8_cast_reg_1613;
assign ret_V_24_fu_1125_p3 = ret_V_23_reg_1996[33] ? select_ln850_4_fu_1119_p3 : ret_V_19_cast_reg_2001;
assign ret_V_27_fu_1486_p3 = ret_V_26_reg_2225[33] ? select_ln850_6_fu_1480_p3 : ret_V_25_cast_reg_2230;
assign ret_V_2_fu_298_p3 = op_1[15] ? select_ln850_fu_293_p3 : ret_V_reg_1568;
assign rhs_1_fu_281_p2 = _0342_ ? 1'h1 : 1'h0;
assign select_ln1118_1_fu_1135_p3 = ush_reg_1772 ? 2'h3 : 2'h0;
assign select_ln1118_fu_1079_p3 = ush_reg_1772 ? 4'hf : 4'h0;
assign select_ln1345_fu_540_p3 = rhs_1_reg_1590 ? 2'h3 : 2'h0;
assign select_ln1497_fu_402_p3 = tmp_reg_1603 ? shl_ln1497_reg_1672 : ashr_ln1497_reg_1667;
assign select_ln340_2_fu_1349_p3 = p_Result_28_reg_2149 ? xor_ln785_1_fu_1344_p2 : and_ln783_fu_1331_p2[3];
assign select_ln340_fu_1403_p3 = p_Result_26_reg_2187 ? xor_ln410_reg_2107 : neg_src_2_fu_1399_p2;
assign select_ln353_2_fu_1428_p3 = ret_V_25_reg_2155[36] ? select_ln850_8_fu_1423_p3 : ret_V_22_cast_reg_2160;
assign select_ln353_fu_986_p3 = ret_V_22_reg_1915[25] ? select_ln850_5_fu_981_p3 : sext_ln850_reg_1936;
assign select_ln384_1_fu_522_p3 = overflow_reg_1720 ? 8'h7f : 8'h81;
assign select_ln384_fu_961_p3 = overflow_1_reg_1925 ? 2'h1 : 2'h3;
assign select_ln850_1_fu_1067_p3 = icmp_ln851_1_reg_2008 ? ret_V_3_cast_reg_1984 : ret_V_3_reg_2013;
assign select_ln850_2_fu_390_p3 = icmp_ln851_2_reg_1630 ? ret_V_8_cast_reg_1613 : ret_V_7_reg_1640;
assign select_ln850_4_fu_1119_p3 = op_14_V_reg_1953[0] ? add_ln691_1_reg_2018 : ret_V_19_cast_reg_2001;
assign select_ln850_5_fu_981_p3 = icmp_ln851_3_reg_1848 ? add_ln691_reg_1948 : sext_ln850_reg_1936;
assign select_ln850_6_fu_1480_p3 = op_17_V_reg_2204[0] ? add_ln691_3_reg_2237 : ret_V_25_cast_reg_2230;
assign select_ln850_7_fu_1547_p3 = op_19_V_reg_2193[0] ? add_ln691_4_reg_2279 : ret_V_28_cast_reg_2272;
assign select_ln850_8_fu_1423_p3 = icmp_ln851_4_reg_2133 ? add_ln691_2_reg_2199 : ret_V_22_cast_reg_2160;
assign select_ln850_fu_293_p3 = icmp_ln851_reg_1575 ? ret_V_reg_1568 : ret_V_1_reg_1585;
assign signbit_fu_597_p2 = _0343_ ? 1'h1 : 1'h0;
assign ush_fu_568_p2 = _0119_ ? 1'h1 : 1'h0;
assign ret_V_20_fu_324_p2 = { rhs_1_reg_1590, 8'h00 } ^ op_1;
assign Range2_all_ones_fu_635_p1 = op_5;
assign and_ln_fu_469_p3 = { tmp_4_reg_1688, 7'h00 };
assign ap_CS_fsm_state1 = ap_CS_fsm[0];
assign ap_CS_fsm_state12 = ap_CS_fsm[11];
assign ap_CS_fsm_state13 = ap_CS_fsm[12];
assign ap_CS_fsm_state14 = ap_CS_fsm[13];
assign ap_CS_fsm_state15 = ap_CS_fsm[14];
assign ap_CS_fsm_state16 = ap_CS_fsm[15];
assign ap_CS_fsm_state17 = ap_CS_fsm[16];
assign ap_CS_fsm_state18 = ap_CS_fsm[17];
assign ap_CS_fsm_state19 = ap_CS_fsm[18];
assign ap_CS_fsm_state2 = ap_CS_fsm[1];
assign ap_CS_fsm_state20 = ap_CS_fsm[19];
assign ap_CS_fsm_state21 = ap_CS_fsm[20];
assign ap_CS_fsm_state22 = ap_CS_fsm[21];
assign ap_CS_fsm_state23 = ap_CS_fsm[22];
assign ap_CS_fsm_state24 = ap_CS_fsm[23];
assign ap_CS_fsm_state25 = ap_CS_fsm[24];
assign ap_CS_fsm_state26 = ap_CS_fsm[25];
assign ap_CS_fsm_state27 = ap_CS_fsm[26];
assign ap_CS_fsm_state28 = ap_CS_fsm[27];
assign ap_CS_fsm_state29 = ap_CS_fsm[28];
assign ap_CS_fsm_state3 = ap_CS_fsm[2];
assign ap_CS_fsm_state30 = ap_CS_fsm[29];
assign ap_CS_fsm_state31 = ap_CS_fsm[30];
assign ap_CS_fsm_state32 = ap_CS_fsm[31];
assign ap_CS_fsm_state33 = ap_CS_fsm[32];
assign ap_CS_fsm_state34 = ap_CS_fsm[33];
assign ap_CS_fsm_state35 = ap_CS_fsm[34];
assign ap_CS_fsm_state36 = ap_CS_fsm[35];
assign ap_CS_fsm_state37 = ap_CS_fsm[36];
assign ap_CS_fsm_state38 = ap_CS_fsm[37];
assign ap_CS_fsm_state39 = ap_CS_fsm[38];
assign ap_CS_fsm_state4 = ap_CS_fsm[3];
assign ap_CS_fsm_state40 = ap_CS_fsm[39];
assign ap_CS_fsm_state41 = ap_CS_fsm[40];
assign ap_CS_fsm_state42 = ap_CS_fsm[41];
assign ap_CS_fsm_state43 = ap_CS_fsm[42];
assign ap_CS_fsm_state44 = ap_CS_fsm[43];
assign ap_CS_fsm_state45 = ap_CS_fsm[44];
assign ap_CS_fsm_state46 = ap_CS_fsm[45];
assign ap_CS_fsm_state47 = ap_CS_fsm[46];
assign ap_CS_fsm_state48 = ap_CS_fsm[47];
assign ap_CS_fsm_state49 = ap_CS_fsm[48];
assign ap_CS_fsm_state5 = ap_CS_fsm[4];
assign ap_CS_fsm_state6 = ap_CS_fsm[5];
assign ap_done = op_27_ap_vld;
assign ap_ready = op_27_ap_vld;
assign conv_i847_fu_365_p0 = op_0;
assign conv_i847_fu_365_p1 = { op_0[7], op_0[7], op_0[7], op_0[7], op_0[7], op_0[7], op_0[7], op_0[7], op_0[7], op_0[7], op_0[7], op_0[7], op_0[7], op_0[7], op_0[7], op_0[7], op_0[7], op_0[7], op_0[7], op_0[7], op_0[7], op_0[7], op_0[7], op_0[7], op_0 };
assign grp_fu_1015_p0 = { select_ln353_reg_1959[6], select_ln353_reg_1959[6], select_ln353_reg_1959[6], select_ln353_reg_1959[6], select_ln353_reg_1959[6], select_ln353_reg_1959[6], select_ln353_reg_1959[6], select_ln353_reg_1959[6], select_ln353_reg_1959[6], select_ln353_reg_1959[6], select_ln353_reg_1959[6], select_ln353_reg_1959[6], select_ln353_reg_1959[6], select_ln353_reg_1959[6], select_ln353_reg_1959[6], select_ln353_reg_1959[6], select_ln353_reg_1959[6], select_ln353_reg_1959[6], select_ln353_reg_1959[6], select_ln353_reg_1959[6], select_ln353_reg_1959[6], select_ln353_reg_1959[6], select_ln353_reg_1959[6], select_ln353_reg_1959[6], select_ln353_reg_1959[6], select_ln353_reg_1959[6], select_ln353_reg_1959, 1'h0 };
assign grp_fu_1015_p1 = { op_14_V_reg_1953[1], op_14_V_reg_1953[1], op_14_V_reg_1953[1], op_14_V_reg_1953[1], op_14_V_reg_1953[1], op_14_V_reg_1953[1], op_14_V_reg_1953[1], op_14_V_reg_1953[1], op_14_V_reg_1953[1], op_14_V_reg_1953[1], op_14_V_reg_1953[1], op_14_V_reg_1953[1], op_14_V_reg_1953[1], op_14_V_reg_1953[1], op_14_V_reg_1953[1], op_14_V_reg_1953[1], op_14_V_reg_1953[1], op_14_V_reg_1953[1], op_14_V_reg_1953[1], op_14_V_reg_1953[1], op_14_V_reg_1953[1], op_14_V_reg_1953[1], op_14_V_reg_1953[1], op_14_V_reg_1953[1], op_14_V_reg_1953[1], op_14_V_reg_1953[1], op_14_V_reg_1953[1], op_14_V_reg_1953[1], op_14_V_reg_1953[1], op_14_V_reg_1953[1], op_14_V_reg_1953[1], op_14_V_reg_1953[1], op_14_V_reg_1953 };
assign grp_fu_1183_p0 = { op_5[3], op_5[3], op_5[3], op_5 };
assign grp_fu_1183_p1 = { ret_V_21_reg_1661, 3'h0 };
assign grp_fu_1192_p1 = { ret_V_19_reg_2023[1], ret_V_19_reg_2023[1], ret_V_19_reg_2023[1], ret_V_19_reg_2023[1], ret_V_19_reg_2023[1], ret_V_19_reg_2023[1], ret_V_19_reg_2023[1], ret_V_19_reg_2023[1], ret_V_19_reg_2023[1], ret_V_19_reg_2023[1], ret_V_19_reg_2023[1], ret_V_19_reg_2023[1], ret_V_19_reg_2023[1], ret_V_19_reg_2023[1], ret_V_19_reg_2023[1], ret_V_19_reg_2023[1], ret_V_19_reg_2023[1], ret_V_19_reg_2023[1], ret_V_19_reg_2023[1], ret_V_19_reg_2023[1], ret_V_19_reg_2023[1], ret_V_19_reg_2023[1], ret_V_19_reg_2023[1], ret_V_19_reg_2023[1], ret_V_19_reg_2023[1], ret_V_19_reg_2023[1], ret_V_19_reg_2023[1], ret_V_19_reg_2023[1], ret_V_19_reg_2023[1], ret_V_19_reg_2023[1], ret_V_19_reg_2023 };
assign grp_fu_1234_p0 = { trunc_ln708_1_reg_2040[1], trunc_ln708_1_reg_2040 };
assign grp_fu_1234_p1 = { 2'h0, and_ln414_1_reg_2087 };
assign grp_fu_1262_p0 = { op_23_V_reg_2097[31], op_23_V_reg_2097, 4'h0 };
assign grp_fu_1262_p1 = { ret_V_9_reg_2092[6], ret_V_9_reg_2092[6], ret_V_9_reg_2092[6], ret_V_9_reg_2092[6], ret_V_9_reg_2092[6], ret_V_9_reg_2092[6], ret_V_9_reg_2092[6], ret_V_9_reg_2092[6], ret_V_9_reg_2092[6], ret_V_9_reg_2092[6], ret_V_9_reg_2092[6], ret_V_9_reg_2092[6], ret_V_9_reg_2092[6], ret_V_9_reg_2092[6], ret_V_9_reg_2092[6], ret_V_9_reg_2092[6], ret_V_9_reg_2092[6], ret_V_9_reg_2092[6], ret_V_9_reg_2092[6], ret_V_9_reg_2092[6], ret_V_9_reg_2092[6], ret_V_9_reg_2092[6], ret_V_9_reg_2092[6], ret_V_9_reg_2092[6], ret_V_9_reg_2092[6], ret_V_9_reg_2092[6], ret_V_9_reg_2092[6], ret_V_9_reg_2092[6], ret_V_9_reg_2092[6], ret_V_9_reg_2092, 1'h0 };
assign grp_fu_1323_p1 = { 1'h0, and_ln410_reg_2138 };
assign grp_fu_1449_p0 = { select_ln353_2_reg_2210[31], select_ln353_2_reg_2210, 1'h0 };
assign grp_fu_1449_p1 = { op_17_V_reg_2204[1], op_17_V_reg_2204[1], op_17_V_reg_2204[1], op_17_V_reg_2204[1], op_17_V_reg_2204[1], op_17_V_reg_2204[1], op_17_V_reg_2204[1], op_17_V_reg_2204[1], op_17_V_reg_2204[1], op_17_V_reg_2204[1], op_17_V_reg_2204[1], op_17_V_reg_2204[1], op_17_V_reg_2204[1], op_17_V_reg_2204[1], op_17_V_reg_2204[1], op_17_V_reg_2204[1], op_17_V_reg_2204[1], op_17_V_reg_2204[1], op_17_V_reg_2204[1], op_17_V_reg_2204[1], op_17_V_reg_2204[1], op_17_V_reg_2204[1], op_17_V_reg_2204[1], op_17_V_reg_2204[1], op_17_V_reg_2204[1], op_17_V_reg_2204[1], op_17_V_reg_2204[1], op_17_V_reg_2204[1], op_17_V_reg_2204[1], op_17_V_reg_2204[1], op_17_V_reg_2204[1], op_17_V_reg_2204[1], op_17_V_reg_2204 };
assign grp_fu_1497_p1 = { op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18 };
assign grp_fu_1516_p0 = { op_26_V_reg_2252[31], op_26_V_reg_2252, 1'h0 };
assign grp_fu_1516_p1 = { op_19_V_reg_2193[3], op_19_V_reg_2193[3], op_19_V_reg_2193[3], op_19_V_reg_2193[3], op_19_V_reg_2193[3], op_19_V_reg_2193[3], op_19_V_reg_2193[3], op_19_V_reg_2193[3], op_19_V_reg_2193[3], op_19_V_reg_2193[3], op_19_V_reg_2193[3], op_19_V_reg_2193[3], op_19_V_reg_2193[3], op_19_V_reg_2193[3], op_19_V_reg_2193[3], op_19_V_reg_2193[3], op_19_V_reg_2193[3], op_19_V_reg_2193[3], op_19_V_reg_2193[3], op_19_V_reg_2193[3], op_19_V_reg_2193[3], op_19_V_reg_2193[3], op_19_V_reg_2193[3], op_19_V_reg_2193[3], op_19_V_reg_2193[3], op_19_V_reg_2193[3], op_19_V_reg_2193[3], op_19_V_reg_2193[3], op_19_V_reg_2193[3], op_19_V_reg_2193[3], op_19_V_reg_2193 };
assign grp_fu_267_p0 = op_1[15:8];
assign grp_fu_346_p1 = { ret_V_2_reg_1597[7], ret_V_2_reg_1597 };
assign grp_fu_368_p1 = { ret_V_2_reg_1597[7], ret_V_2_reg_1597[7], ret_V_2_reg_1597[7], ret_V_2_reg_1597[7], ret_V_2_reg_1597[7], ret_V_2_reg_1597[7], ret_V_2_reg_1597[7], ret_V_2_reg_1597[7], ret_V_2_reg_1597[7], ret_V_2_reg_1597[7], ret_V_2_reg_1597[7], ret_V_2_reg_1597[7], ret_V_2_reg_1597[7], ret_V_2_reg_1597[7], ret_V_2_reg_1597[7], ret_V_2_reg_1597[7], ret_V_2_reg_1597[7], ret_V_2_reg_1597[7], ret_V_2_reg_1597[7], ret_V_2_reg_1597[7], ret_V_2_reg_1597[7], ret_V_2_reg_1597[7], ret_V_2_reg_1597[7], ret_V_2_reg_1597[7], ret_V_2_reg_1597 };
assign grp_fu_377_p1 = { sub_ln1497_reg_1635[8], sub_ln1497_reg_1635[8], sub_ln1497_reg_1635[8], sub_ln1497_reg_1635[8], sub_ln1497_reg_1635[8], sub_ln1497_reg_1635[8], sub_ln1497_reg_1635[8], sub_ln1497_reg_1635[8], sub_ln1497_reg_1635[8], sub_ln1497_reg_1635[8], sub_ln1497_reg_1635[8], sub_ln1497_reg_1635[8], sub_ln1497_reg_1635[8], sub_ln1497_reg_1635[8], sub_ln1497_reg_1635[8], sub_ln1497_reg_1635[8], sub_ln1497_reg_1635[8], sub_ln1497_reg_1635[8], sub_ln1497_reg_1635[8], sub_ln1497_reg_1635[8], sub_ln1497_reg_1635[8], sub_ln1497_reg_1635[8], sub_ln1497_reg_1635[8], sub_ln1497_reg_1635 };
assign grp_fu_730_p0 = { op_12_V_reg_1789[3], op_12_V_reg_1789, 2'h0 };
assign grp_fu_730_p1 = { 4'h0, signbit_reg_1784, 2'h0 };
assign grp_fu_752_p1 = { 1'h0, and_ln412_reg_1833 };
assign grp_fu_810_p0 = { tmp_1_reg_1858[4], tmp_1_reg_1858, 20'h00000 };
assign grp_fu_810_p1 = { 4'h0, ret_V_5_reg_1779, 15'h0000 };
assign grp_fu_930_p0 = { tmp_s_reg_1920[5], tmp_s_reg_1920 };
assign grp_fu_996_p1 = { 3'h0, ush_reg_1772 };
assign neg_src_4_fu_1336_p3 = and_ln783_fu_1331_p2[3];
assign op_13_V_fu_780_p3 = { ret_V_5_reg_1779, 15'h0000 };
assign op_16_V_fu_1240_p3 = { ret_V_9_reg_2092, 1'h0 };
assign op_8_V_fu_679_p3 = { signbit_reg_1784, 2'h0 };
assign or_ln1195_1_fu_643_p1 = op_5;
assign or_ln_fu_437_p4 = { tmp_4_reg_1688, 2'h0, p_Result_s_22_reg_1694 };
assign p_Result_12_fu_1383_p4 = { 1'h0, p_Val2_7_fu_1374_p2 };
assign p_Result_16_fu_686_p3 = or_ln1195_1_reg_1806[2];
assign p_Result_18_fu_974_p3 = ret_V_22_reg_1915[25];
assign p_Result_19_fu_1109_p3 = ret_V_23_reg_1996[33];
assign p_Result_1_fu_1268_p3 = { trunc_ln851_5_reg_2102, 1'h0 };
assign p_Result_20_fu_1416_p3 = ret_V_25_reg_2155[36];
assign p_Result_21_fu_1470_p3 = ret_V_26_reg_2225[33];
assign p_Result_22_fu_1537_p3 = ret_V_28_reg_2267[33];
assign p_Result_25_fu_1281_p3 = r_V_1_reg_2070[1];
assign p_Result_29_fu_649_p1 = op_5;
assign p_Result_2_fu_1060_p3 = r_V_reg_1979[5];
assign p_Result_30_fu_693_p1 = op_5;
assign p_Result_30_fu_693_p3 = op_5[1];
assign p_Result_31_fu_816_p3 = or_ln1195_1_reg_1806[3];
assign p_Result_3_fu_736_p3 = { trunc_ln851_3_reg_1828, 15'h0000 };
assign p_Result_4_fu_383_p3 = ret_V_20_reg_1608[15];
assign p_Result_5_fu_456_p3 = { trunc_ln790_reg_1700, 5'h00 };
assign p_Result_s_fu_286_p3 = op_1[15];
assign p_Val2_s_fu_514_p3 = { select_ln1497_reg_1677[2:0], 5'h00 };
assign r_1_fu_700_p1 = or_ln1195_reg_1794[0];
assign r_V_2_fu_1086_p1 = op_5;
assign r_fu_1288_p1 = r_V_1_reg_2070[0];
assign rhs_10_fu_1251_p3 = { op_23_V_reg_2097, 4'h0 };
assign rhs_11_fu_1438_p3 = { select_ln353_2_reg_2210, 1'h0 };
assign rhs_13_fu_1505_p3 = { op_26_V_reg_2252, 1'h0 };
assign rhs_2_fu_313_p3 = { rhs_1_reg_1590, 8'h00 };
assign rhs_5_fu_611_p3 = { ret_reg_1752, 3'h0 };
assign rhs_7_fu_719_p3 = { op_12_V_reg_1789, 2'h0 };
assign rhs_8_fu_799_p3 = { tmp_1_reg_1858, 20'h00000 };
assign rhs_fu_574_p3 = { op_6, 5'h00 };
assign sext_ln1193_fu_1173_p0 = op_5;
assign sext_ln1195_fu_625_p0 = op_5;
assign sext_ln1195_fu_625_p1 = { op_5[3], op_5 };
assign sext_ln367_fu_1379_p1 = { p_Val2_7_fu_1374_p2[2], p_Val2_7_fu_1374_p2 };
assign sext_ln727_fu_557_p1 = { op_2_V_reg_1741[7], op_2_V_reg_1741[7], op_2_V_reg_1741[7], op_2_V_reg_1741[7], op_2_V_reg_1741[7], op_2_V_reg_1741 };
assign sext_ln745_fu_1328_p1 = { p_Val2_6_reg_2143[2], p_Val2_6_reg_2143 };
assign sext_ln850_fu_927_p1 = { tmp_s_reg_1920[5], tmp_s_reg_1920 };
assign shl_ln728_1_fu_560_p3 = { op_4, 5'h00 };
assign shl_ln728_5_fu_586_p3 = { rhs_1_reg_1590, 5'h00 };
assign shl_ln_fu_273_p1 = op_0;
assign shl_ln_fu_273_p3 = { op_0, 8'h00 };
assign tmp_13_fu_1151_p3 = and_ln414_fu_1145_p2[1];
assign tmp_24_fu_867_p3 = or_ln1195_reg_1794[4];
assign tmp_26_fu_1004_p3 = { select_ln353_reg_1959, 1'h0 };
assign tmp_3_fu_1159_p3 = { and_ln414_fu_1145_p2[1], r_V_2_reg_2028[0] };
assign tmp_9_fu_834_p3 = { Range2_all_ones_reg_1800, tmp_23_reg_1823 };
assign trunc_ln1118_fu_1132_p0 = op_5;
assign trunc_ln1118_fu_1132_p1 = op_5[1:0];
assign trunc_ln1195_1_fu_618_p3 = { trunc_ln1195_reg_1757, 3'h0 };
assign trunc_ln1195_fu_553_p1 = ret_fu_547_p2[0];
assign trunc_ln1349_fu_602_p1 = op_4[3:0];
assign trunc_ln718_fu_1142_p1 = r_V_2_reg_2028[0];
assign trunc_ln731_fu_511_p1 = select_ln1497_reg_1677[2:0];
assign trunc_ln790_1_fu_913_p1 = p_Val2_9_reg_1873[0];
assign trunc_ln790_fu_433_p1 = select_ln1497_fu_402_p3[1:0];
assign trunc_ln851_1_fu_1031_p1 = grp_fu_774_p2[2:0];
assign trunc_ln851_2_fu_339_p1 = ret_V_20_fu_324_p2[7:0];
assign trunc_ln851_3_fu_675_p1 = ret_V_5_fu_581_p2[4:0];
assign trunc_ln851_4_fu_1116_p1 = op_14_V_reg_1953[0];
assign trunc_ln851_5_fu_1219_p1 = grp_fu_1183_p2[2:0];
assign trunc_ln851_6_fu_1477_p1 = op_17_V_reg_2204[0];
assign trunc_ln851_7_fu_1544_p1 = op_19_V_reg_2193[0];
assign trunc_ln851_fu_257_p1 = op_1[7:0];
assign trunc_ln8_fu_536_p1 = op_2_V_fu_529_p3[6:0];
assign zext_ln1196_fu_320_p1 = { 7'h00, rhs_1_reg_1590, 8'h00 };
assign zext_ln1499_fu_593_p1 = { 2'h0, rhs_1_reg_1590, 5'h00 };
assign \sub_9ns_9s_9_2_1_U2.top_sub_9ns_9s_9_2_1_Adder_1_U.ain_s0  = \sub_9ns_9s_9_2_1_U2.top_sub_9ns_9s_9_2_1_Adder_1_U.a ;
assign \sub_9ns_9s_9_2_1_U2.top_sub_9ns_9s_9_2_1_Adder_1_U.s  = { \sub_9ns_9s_9_2_1_U2.top_sub_9ns_9s_9_2_1_Adder_1_U.fas_s2 , \sub_9ns_9s_9_2_1_U2.top_sub_9ns_9s_9_2_1_Adder_1_U.sum_s1  };
assign \sub_9ns_9s_9_2_1_U2.top_sub_9ns_9s_9_2_1_Adder_1_U.u2.a  = \sub_9ns_9s_9_2_1_U2.top_sub_9ns_9s_9_2_1_Adder_1_U.ain_s1 ;
assign \sub_9ns_9s_9_2_1_U2.top_sub_9ns_9s_9_2_1_Adder_1_U.u2.b  = \sub_9ns_9s_9_2_1_U2.top_sub_9ns_9s_9_2_1_Adder_1_U.bin_s1 ;
assign \sub_9ns_9s_9_2_1_U2.top_sub_9ns_9s_9_2_1_Adder_1_U.u2.cin  = \sub_9ns_9s_9_2_1_U2.top_sub_9ns_9s_9_2_1_Adder_1_U.carry_s1 ;
assign \sub_9ns_9s_9_2_1_U2.top_sub_9ns_9s_9_2_1_Adder_1_U.facout_s2  = \sub_9ns_9s_9_2_1_U2.top_sub_9ns_9s_9_2_1_Adder_1_U.u2.cout ;
assign \sub_9ns_9s_9_2_1_U2.top_sub_9ns_9s_9_2_1_Adder_1_U.fas_s2  = \sub_9ns_9s_9_2_1_U2.top_sub_9ns_9s_9_2_1_Adder_1_U.u2.s ;
assign \sub_9ns_9s_9_2_1_U2.top_sub_9ns_9s_9_2_1_Adder_1_U.u1.a  = \sub_9ns_9s_9_2_1_U2.top_sub_9ns_9s_9_2_1_Adder_1_U.a [3:0];
assign \sub_9ns_9s_9_2_1_U2.top_sub_9ns_9s_9_2_1_Adder_1_U.u1.b  = \sub_9ns_9s_9_2_1_U2.top_sub_9ns_9s_9_2_1_Adder_1_U.bin_s0 [3:0];
assign \sub_9ns_9s_9_2_1_U2.top_sub_9ns_9s_9_2_1_Adder_1_U.u1.cin  = 1'h1;
assign \sub_9ns_9s_9_2_1_U2.top_sub_9ns_9s_9_2_1_Adder_1_U.facout_s1  = \sub_9ns_9s_9_2_1_U2.top_sub_9ns_9s_9_2_1_Adder_1_U.u1.cout ;
assign \sub_9ns_9s_9_2_1_U2.top_sub_9ns_9s_9_2_1_Adder_1_U.fas_s1  = \sub_9ns_9s_9_2_1_U2.top_sub_9ns_9s_9_2_1_Adder_1_U.u1.s ;
assign \sub_9ns_9s_9_2_1_U2.top_sub_9ns_9s_9_2_1_Adder_1_U.a  = \sub_9ns_9s_9_2_1_U2.din0 ;
assign \sub_9ns_9s_9_2_1_U2.top_sub_9ns_9s_9_2_1_Adder_1_U.b  = \sub_9ns_9s_9_2_1_U2.din1 ;
assign \sub_9ns_9s_9_2_1_U2.top_sub_9ns_9s_9_2_1_Adder_1_U.ce  = \sub_9ns_9s_9_2_1_U2.ce ;
assign \sub_9ns_9s_9_2_1_U2.top_sub_9ns_9s_9_2_1_Adder_1_U.clk  = \sub_9ns_9s_9_2_1_U2.clk ;
assign \sub_9ns_9s_9_2_1_U2.top_sub_9ns_9s_9_2_1_Adder_1_U.reset  = \sub_9ns_9s_9_2_1_U2.reset ;
assign \sub_9ns_9s_9_2_1_U2.dout  = \sub_9ns_9s_9_2_1_U2.top_sub_9ns_9s_9_2_1_Adder_1_U.s ;
assign \sub_9ns_9s_9_2_1_U2.ce  = 1'h1;
assign \sub_9ns_9s_9_2_1_U2.clk  = ap_clk;
assign \sub_9ns_9s_9_2_1_U2.din0  = 9'h000;
assign \sub_9ns_9s_9_2_1_U2.din1  = { ret_V_2_reg_1597[7], ret_V_2_reg_1597 };
assign grp_fu_346_p2 = \sub_9ns_9s_9_2_1_U2.dout ;
assign \sub_9ns_9s_9_2_1_U2.reset  = ap_rst;
assign \sub_7s_7ns_7_2_1_U15.top_sub_7s_7ns_7_2_1_Adder_8_U.ain_s0  = \sub_7s_7ns_7_2_1_U15.top_sub_7s_7ns_7_2_1_Adder_8_U.a ;
assign \sub_7s_7ns_7_2_1_U15.top_sub_7s_7ns_7_2_1_Adder_8_U.s  = { \sub_7s_7ns_7_2_1_U15.top_sub_7s_7ns_7_2_1_Adder_8_U.fas_s2 , \sub_7s_7ns_7_2_1_U15.top_sub_7s_7ns_7_2_1_Adder_8_U.sum_s1  };
assign \sub_7s_7ns_7_2_1_U15.top_sub_7s_7ns_7_2_1_Adder_8_U.u2.a  = \sub_7s_7ns_7_2_1_U15.top_sub_7s_7ns_7_2_1_Adder_8_U.ain_s1 ;
assign \sub_7s_7ns_7_2_1_U15.top_sub_7s_7ns_7_2_1_Adder_8_U.u2.b  = \sub_7s_7ns_7_2_1_U15.top_sub_7s_7ns_7_2_1_Adder_8_U.bin_s1 ;
assign \sub_7s_7ns_7_2_1_U15.top_sub_7s_7ns_7_2_1_Adder_8_U.u2.cin  = \sub_7s_7ns_7_2_1_U15.top_sub_7s_7ns_7_2_1_Adder_8_U.carry_s1 ;
assign \sub_7s_7ns_7_2_1_U15.top_sub_7s_7ns_7_2_1_Adder_8_U.facout_s2  = \sub_7s_7ns_7_2_1_U15.top_sub_7s_7ns_7_2_1_Adder_8_U.u2.cout ;
assign \sub_7s_7ns_7_2_1_U15.top_sub_7s_7ns_7_2_1_Adder_8_U.fas_s2  = \sub_7s_7ns_7_2_1_U15.top_sub_7s_7ns_7_2_1_Adder_8_U.u2.s ;
assign \sub_7s_7ns_7_2_1_U15.top_sub_7s_7ns_7_2_1_Adder_8_U.u1.a  = \sub_7s_7ns_7_2_1_U15.top_sub_7s_7ns_7_2_1_Adder_8_U.a [2:0];
assign \sub_7s_7ns_7_2_1_U15.top_sub_7s_7ns_7_2_1_Adder_8_U.u1.b  = \sub_7s_7ns_7_2_1_U15.top_sub_7s_7ns_7_2_1_Adder_8_U.bin_s0 [2:0];
assign \sub_7s_7ns_7_2_1_U15.top_sub_7s_7ns_7_2_1_Adder_8_U.u1.cin  = 1'h1;
assign \sub_7s_7ns_7_2_1_U15.top_sub_7s_7ns_7_2_1_Adder_8_U.facout_s1  = \sub_7s_7ns_7_2_1_U15.top_sub_7s_7ns_7_2_1_Adder_8_U.u1.cout ;
assign \sub_7s_7ns_7_2_1_U15.top_sub_7s_7ns_7_2_1_Adder_8_U.fas_s1  = \sub_7s_7ns_7_2_1_U15.top_sub_7s_7ns_7_2_1_Adder_8_U.u1.s ;
assign \sub_7s_7ns_7_2_1_U15.top_sub_7s_7ns_7_2_1_Adder_8_U.a  = \sub_7s_7ns_7_2_1_U15.din0 ;
assign \sub_7s_7ns_7_2_1_U15.top_sub_7s_7ns_7_2_1_Adder_8_U.b  = \sub_7s_7ns_7_2_1_U15.din1 ;
assign \sub_7s_7ns_7_2_1_U15.top_sub_7s_7ns_7_2_1_Adder_8_U.ce  = \sub_7s_7ns_7_2_1_U15.ce ;
assign \sub_7s_7ns_7_2_1_U15.top_sub_7s_7ns_7_2_1_Adder_8_U.clk  = \sub_7s_7ns_7_2_1_U15.clk ;
assign \sub_7s_7ns_7_2_1_U15.top_sub_7s_7ns_7_2_1_Adder_8_U.reset  = \sub_7s_7ns_7_2_1_U15.reset ;
assign \sub_7s_7ns_7_2_1_U15.dout  = \sub_7s_7ns_7_2_1_U15.top_sub_7s_7ns_7_2_1_Adder_8_U.s ;
assign \sub_7s_7ns_7_2_1_U15.ce  = 1'h1;
assign \sub_7s_7ns_7_2_1_U15.clk  = ap_clk;
assign \sub_7s_7ns_7_2_1_U15.din0  = { op_5[3], op_5[3], op_5[3], op_5 };
assign \sub_7s_7ns_7_2_1_U15.din1  = { ret_V_21_reg_1661, 3'h0 };
assign grp_fu_1183_p2 = \sub_7s_7ns_7_2_1_U15.dout ;
assign \sub_7s_7ns_7_2_1_U15.reset  = ap_rst;
assign \shl_4s_1ns_4_7_1_U11.din1_cast  = \shl_4s_1ns_4_7_1_U11.din1 [0];
assign \shl_4s_1ns_4_7_1_U11.din1_mask  = 1'h1;
assign \shl_4s_1ns_4_7_1_U11.ce  = 1'h1;
assign \shl_4s_1ns_4_7_1_U11.clk  = ap_clk;
assign \shl_4s_1ns_4_7_1_U11.din0  = op_5;
assign \shl_4s_1ns_4_7_1_U11.din1  = { 3'h0, ush_reg_1772 };
assign grp_fu_996_p2 = \shl_4s_1ns_4_7_1_U11.dout ;
assign \shl_4s_1ns_4_7_1_U11.reset  = ap_rst;
assign \shl_32s_32s_32_7_1_U5.din1_cast  = \shl_32s_32s_32_7_1_U5.din1 ;
assign \shl_32s_32s_32_7_1_U5.din1_mask  = 32'd31;
assign \shl_32s_32s_32_7_1_U5.ce  = 1'h1;
assign \shl_32s_32s_32_7_1_U5.clk  = ap_clk;
assign \shl_32s_32s_32_7_1_U5.din0  = { op_0[7], op_0[7], op_0[7], op_0[7], op_0[7], op_0[7], op_0[7], op_0[7], op_0[7], op_0[7], op_0[7], op_0[7], op_0[7], op_0[7], op_0[7], op_0[7], op_0[7], op_0[7], op_0[7], op_0[7], op_0[7], op_0[7], op_0[7], op_0[7], op_0 };
assign \shl_32s_32s_32_7_1_U5.din1  = { sub_ln1497_reg_1635[8], sub_ln1497_reg_1635[8], sub_ln1497_reg_1635[8], sub_ln1497_reg_1635[8], sub_ln1497_reg_1635[8], sub_ln1497_reg_1635[8], sub_ln1497_reg_1635[8], sub_ln1497_reg_1635[8], sub_ln1497_reg_1635[8], sub_ln1497_reg_1635[8], sub_ln1497_reg_1635[8], sub_ln1497_reg_1635[8], sub_ln1497_reg_1635[8], sub_ln1497_reg_1635[8], sub_ln1497_reg_1635[8], sub_ln1497_reg_1635[8], sub_ln1497_reg_1635[8], sub_ln1497_reg_1635[8], sub_ln1497_reg_1635[8], sub_ln1497_reg_1635[8], sub_ln1497_reg_1635[8], sub_ln1497_reg_1635[8], sub_ln1497_reg_1635[8], sub_ln1497_reg_1635 };
assign grp_fu_377_p2 = \shl_32s_32s_32_7_1_U5.dout ;
assign \shl_32s_32s_32_7_1_U5.reset  = ap_rst;
assign \mul_4s_2s_6_7_1_U8.top_mul_4s_2s_6_7_1_Mul_DSP_0_U.p  = \mul_4s_2s_6_7_1_U8.top_mul_4s_2s_6_7_1_Mul_DSP_0_U.buff4 ;
assign \mul_4s_2s_6_7_1_U8.top_mul_4s_2s_6_7_1_Mul_DSP_0_U.a  = \mul_4s_2s_6_7_1_U8.din0 ;
assign \mul_4s_2s_6_7_1_U8.top_mul_4s_2s_6_7_1_Mul_DSP_0_U.b  = \mul_4s_2s_6_7_1_U8.din1 ;
assign \mul_4s_2s_6_7_1_U8.top_mul_4s_2s_6_7_1_Mul_DSP_0_U.ce  = \mul_4s_2s_6_7_1_U8.ce ;
assign \mul_4s_2s_6_7_1_U8.top_mul_4s_2s_6_7_1_Mul_DSP_0_U.clk  = \mul_4s_2s_6_7_1_U8.clk ;
assign \mul_4s_2s_6_7_1_U8.dout  = \mul_4s_2s_6_7_1_U8.top_mul_4s_2s_6_7_1_Mul_DSP_0_U.p ;
assign \mul_4s_2s_6_7_1_U8.ce  = 1'h1;
assign \mul_4s_2s_6_7_1_U8.clk  = ap_clk;
assign \mul_4s_2s_6_7_1_U8.din0  = op_5;
assign \mul_4s_2s_6_7_1_U8.din1  = op_11;
assign grp_fu_774_p2 = \mul_4s_2s_6_7_1_U8.dout ;
assign \mul_4s_2s_6_7_1_U8.reset  = ap_rst;
assign \ashr_32s_32s_32_7_1_U4.din1_cast  = \ashr_32s_32s_32_7_1_U4.din1 ;
assign \ashr_32s_32s_32_7_1_U4.din1_mask  = 32'd31;
assign \ashr_32s_32s_32_7_1_U4.ce  = 1'h1;
assign \ashr_32s_32s_32_7_1_U4.clk  = ap_clk;
assign \ashr_32s_32s_32_7_1_U4.din0  = { op_0[7], op_0[7], op_0[7], op_0[7], op_0[7], op_0[7], op_0[7], op_0[7], op_0[7], op_0[7], op_0[7], op_0[7], op_0[7], op_0[7], op_0[7], op_0[7], op_0[7], op_0[7], op_0[7], op_0[7], op_0[7], op_0[7], op_0[7], op_0[7], op_0 };
assign \ashr_32s_32s_32_7_1_U4.din1  = { ret_V_2_reg_1597[7], ret_V_2_reg_1597[7], ret_V_2_reg_1597[7], ret_V_2_reg_1597[7], ret_V_2_reg_1597[7], ret_V_2_reg_1597[7], ret_V_2_reg_1597[7], ret_V_2_reg_1597[7], ret_V_2_reg_1597[7], ret_V_2_reg_1597[7], ret_V_2_reg_1597[7], ret_V_2_reg_1597[7], ret_V_2_reg_1597[7], ret_V_2_reg_1597[7], ret_V_2_reg_1597[7], ret_V_2_reg_1597[7], ret_V_2_reg_1597[7], ret_V_2_reg_1597[7], ret_V_2_reg_1597[7], ret_V_2_reg_1597[7], ret_V_2_reg_1597[7], ret_V_2_reg_1597[7], ret_V_2_reg_1597[7], ret_V_2_reg_1597[7], ret_V_2_reg_1597 };
assign grp_fu_368_p2 = \ashr_32s_32s_32_7_1_U4.dout ;
assign \ashr_32s_32s_32_7_1_U4.reset  = ap_rst;
assign \add_8ns_8ns_8_2_1_U1.top_add_8ns_8ns_8_2_1_Adder_0_U.ain_s0  = \add_8ns_8ns_8_2_1_U1.top_add_8ns_8ns_8_2_1_Adder_0_U.a ;
assign \add_8ns_8ns_8_2_1_U1.top_add_8ns_8ns_8_2_1_Adder_0_U.bin_s0  = \add_8ns_8ns_8_2_1_U1.top_add_8ns_8ns_8_2_1_Adder_0_U.b ;
assign \add_8ns_8ns_8_2_1_U1.top_add_8ns_8ns_8_2_1_Adder_0_U.s  = { \add_8ns_8ns_8_2_1_U1.top_add_8ns_8ns_8_2_1_Adder_0_U.fas_s2 , \add_8ns_8ns_8_2_1_U1.top_add_8ns_8ns_8_2_1_Adder_0_U.sum_s1  };
assign \add_8ns_8ns_8_2_1_U1.top_add_8ns_8ns_8_2_1_Adder_0_U.u2.a  = \add_8ns_8ns_8_2_1_U1.top_add_8ns_8ns_8_2_1_Adder_0_U.ain_s1 ;
assign \add_8ns_8ns_8_2_1_U1.top_add_8ns_8ns_8_2_1_Adder_0_U.u2.b  = \add_8ns_8ns_8_2_1_U1.top_add_8ns_8ns_8_2_1_Adder_0_U.bin_s1 ;
assign \add_8ns_8ns_8_2_1_U1.top_add_8ns_8ns_8_2_1_Adder_0_U.u2.cin  = \add_8ns_8ns_8_2_1_U1.top_add_8ns_8ns_8_2_1_Adder_0_U.carry_s1 ;
assign \add_8ns_8ns_8_2_1_U1.top_add_8ns_8ns_8_2_1_Adder_0_U.facout_s2  = \add_8ns_8ns_8_2_1_U1.top_add_8ns_8ns_8_2_1_Adder_0_U.u2.cout ;
assign \add_8ns_8ns_8_2_1_U1.top_add_8ns_8ns_8_2_1_Adder_0_U.fas_s2  = \add_8ns_8ns_8_2_1_U1.top_add_8ns_8ns_8_2_1_Adder_0_U.u2.s ;
assign \add_8ns_8ns_8_2_1_U1.top_add_8ns_8ns_8_2_1_Adder_0_U.u1.a  = \add_8ns_8ns_8_2_1_U1.top_add_8ns_8ns_8_2_1_Adder_0_U.a [3:0];
assign \add_8ns_8ns_8_2_1_U1.top_add_8ns_8ns_8_2_1_Adder_0_U.u1.b  = \add_8ns_8ns_8_2_1_U1.top_add_8ns_8ns_8_2_1_Adder_0_U.b [3:0];
assign \add_8ns_8ns_8_2_1_U1.top_add_8ns_8ns_8_2_1_Adder_0_U.u1.cin  = 1'h0;
assign \add_8ns_8ns_8_2_1_U1.top_add_8ns_8ns_8_2_1_Adder_0_U.facout_s1  = \add_8ns_8ns_8_2_1_U1.top_add_8ns_8ns_8_2_1_Adder_0_U.u1.cout ;
assign \add_8ns_8ns_8_2_1_U1.top_add_8ns_8ns_8_2_1_Adder_0_U.fas_s1  = \add_8ns_8ns_8_2_1_U1.top_add_8ns_8ns_8_2_1_Adder_0_U.u1.s ;
assign \add_8ns_8ns_8_2_1_U1.top_add_8ns_8ns_8_2_1_Adder_0_U.a  = \add_8ns_8ns_8_2_1_U1.din0 ;
assign \add_8ns_8ns_8_2_1_U1.top_add_8ns_8ns_8_2_1_Adder_0_U.b  = \add_8ns_8ns_8_2_1_U1.din1 ;
assign \add_8ns_8ns_8_2_1_U1.top_add_8ns_8ns_8_2_1_Adder_0_U.ce  = \add_8ns_8ns_8_2_1_U1.ce ;
assign \add_8ns_8ns_8_2_1_U1.top_add_8ns_8ns_8_2_1_Adder_0_U.clk  = \add_8ns_8ns_8_2_1_U1.clk ;
assign \add_8ns_8ns_8_2_1_U1.top_add_8ns_8ns_8_2_1_Adder_0_U.reset  = \add_8ns_8ns_8_2_1_U1.reset ;
assign \add_8ns_8ns_8_2_1_U1.dout  = \add_8ns_8ns_8_2_1_U1.top_add_8ns_8ns_8_2_1_Adder_0_U.s ;
assign \add_8ns_8ns_8_2_1_U1.ce  = 1'h1;
assign \add_8ns_8ns_8_2_1_U1.clk  = ap_clk;
assign \add_8ns_8ns_8_2_1_U1.din0  = op_1[15:8];
assign \add_8ns_8ns_8_2_1_U1.din1  = 8'h01;
assign grp_fu_267_p2 = \add_8ns_8ns_8_2_1_U1.dout ;
assign \add_8ns_8ns_8_2_1_U1.reset  = ap_rst;
assign \add_7s_7ns_7_2_1_U6.top_add_7s_7ns_7_2_1_Adder_3_U.ain_s0  = \add_7s_7ns_7_2_1_U6.top_add_7s_7ns_7_2_1_Adder_3_U.a ;
assign \add_7s_7ns_7_2_1_U6.top_add_7s_7ns_7_2_1_Adder_3_U.bin_s0  = \add_7s_7ns_7_2_1_U6.top_add_7s_7ns_7_2_1_Adder_3_U.b ;
assign \add_7s_7ns_7_2_1_U6.top_add_7s_7ns_7_2_1_Adder_3_U.s  = { \add_7s_7ns_7_2_1_U6.top_add_7s_7ns_7_2_1_Adder_3_U.fas_s2 , \add_7s_7ns_7_2_1_U6.top_add_7s_7ns_7_2_1_Adder_3_U.sum_s1  };
assign \add_7s_7ns_7_2_1_U6.top_add_7s_7ns_7_2_1_Adder_3_U.u2.a  = \add_7s_7ns_7_2_1_U6.top_add_7s_7ns_7_2_1_Adder_3_U.ain_s1 ;
assign \add_7s_7ns_7_2_1_U6.top_add_7s_7ns_7_2_1_Adder_3_U.u2.b  = \add_7s_7ns_7_2_1_U6.top_add_7s_7ns_7_2_1_Adder_3_U.bin_s1 ;
assign \add_7s_7ns_7_2_1_U6.top_add_7s_7ns_7_2_1_Adder_3_U.u2.cin  = \add_7s_7ns_7_2_1_U6.top_add_7s_7ns_7_2_1_Adder_3_U.carry_s1 ;
assign \add_7s_7ns_7_2_1_U6.top_add_7s_7ns_7_2_1_Adder_3_U.facout_s2  = \add_7s_7ns_7_2_1_U6.top_add_7s_7ns_7_2_1_Adder_3_U.u2.cout ;
assign \add_7s_7ns_7_2_1_U6.top_add_7s_7ns_7_2_1_Adder_3_U.fas_s2  = \add_7s_7ns_7_2_1_U6.top_add_7s_7ns_7_2_1_Adder_3_U.u2.s ;
assign \add_7s_7ns_7_2_1_U6.top_add_7s_7ns_7_2_1_Adder_3_U.u1.a  = \add_7s_7ns_7_2_1_U6.top_add_7s_7ns_7_2_1_Adder_3_U.a [2:0];
assign \add_7s_7ns_7_2_1_U6.top_add_7s_7ns_7_2_1_Adder_3_U.u1.b  = \add_7s_7ns_7_2_1_U6.top_add_7s_7ns_7_2_1_Adder_3_U.b [2:0];
assign \add_7s_7ns_7_2_1_U6.top_add_7s_7ns_7_2_1_Adder_3_U.u1.cin  = 1'h0;
assign \add_7s_7ns_7_2_1_U6.top_add_7s_7ns_7_2_1_Adder_3_U.facout_s1  = \add_7s_7ns_7_2_1_U6.top_add_7s_7ns_7_2_1_Adder_3_U.u1.cout ;
assign \add_7s_7ns_7_2_1_U6.top_add_7s_7ns_7_2_1_Adder_3_U.fas_s1  = \add_7s_7ns_7_2_1_U6.top_add_7s_7ns_7_2_1_Adder_3_U.u1.s ;
assign \add_7s_7ns_7_2_1_U6.top_add_7s_7ns_7_2_1_Adder_3_U.a  = \add_7s_7ns_7_2_1_U6.din0 ;
assign \add_7s_7ns_7_2_1_U6.top_add_7s_7ns_7_2_1_Adder_3_U.b  = \add_7s_7ns_7_2_1_U6.din1 ;
assign \add_7s_7ns_7_2_1_U6.top_add_7s_7ns_7_2_1_Adder_3_U.ce  = \add_7s_7ns_7_2_1_U6.ce ;
assign \add_7s_7ns_7_2_1_U6.top_add_7s_7ns_7_2_1_Adder_3_U.clk  = \add_7s_7ns_7_2_1_U6.clk ;
assign \add_7s_7ns_7_2_1_U6.top_add_7s_7ns_7_2_1_Adder_3_U.reset  = \add_7s_7ns_7_2_1_U6.reset ;
assign \add_7s_7ns_7_2_1_U6.dout  = \add_7s_7ns_7_2_1_U6.top_add_7s_7ns_7_2_1_Adder_3_U.s ;
assign \add_7s_7ns_7_2_1_U6.ce  = 1'h1;
assign \add_7s_7ns_7_2_1_U6.clk  = ap_clk;
assign \add_7s_7ns_7_2_1_U6.din0  = { op_12_V_reg_1789[3], op_12_V_reg_1789, 2'h0 };
assign \add_7s_7ns_7_2_1_U6.din1  = { 4'h0, signbit_reg_1784, 2'h0 };
assign grp_fu_730_p2 = \add_7s_7ns_7_2_1_U6.dout ;
assign \add_7s_7ns_7_2_1_U6.reset  = ap_rst;
assign \add_7s_7ns_7_2_1_U10.top_add_7s_7ns_7_2_1_Adder_3_U.ain_s0  = \add_7s_7ns_7_2_1_U10.top_add_7s_7ns_7_2_1_Adder_3_U.a ;
assign \add_7s_7ns_7_2_1_U10.top_add_7s_7ns_7_2_1_Adder_3_U.bin_s0  = \add_7s_7ns_7_2_1_U10.top_add_7s_7ns_7_2_1_Adder_3_U.b ;
assign \add_7s_7ns_7_2_1_U10.top_add_7s_7ns_7_2_1_Adder_3_U.s  = { \add_7s_7ns_7_2_1_U10.top_add_7s_7ns_7_2_1_Adder_3_U.fas_s2 , \add_7s_7ns_7_2_1_U10.top_add_7s_7ns_7_2_1_Adder_3_U.sum_s1  };
assign \add_7s_7ns_7_2_1_U10.top_add_7s_7ns_7_2_1_Adder_3_U.u2.a  = \add_7s_7ns_7_2_1_U10.top_add_7s_7ns_7_2_1_Adder_3_U.ain_s1 ;
assign \add_7s_7ns_7_2_1_U10.top_add_7s_7ns_7_2_1_Adder_3_U.u2.b  = \add_7s_7ns_7_2_1_U10.top_add_7s_7ns_7_2_1_Adder_3_U.bin_s1 ;
assign \add_7s_7ns_7_2_1_U10.top_add_7s_7ns_7_2_1_Adder_3_U.u2.cin  = \add_7s_7ns_7_2_1_U10.top_add_7s_7ns_7_2_1_Adder_3_U.carry_s1 ;
assign \add_7s_7ns_7_2_1_U10.top_add_7s_7ns_7_2_1_Adder_3_U.facout_s2  = \add_7s_7ns_7_2_1_U10.top_add_7s_7ns_7_2_1_Adder_3_U.u2.cout ;
assign \add_7s_7ns_7_2_1_U10.top_add_7s_7ns_7_2_1_Adder_3_U.fas_s2  = \add_7s_7ns_7_2_1_U10.top_add_7s_7ns_7_2_1_Adder_3_U.u2.s ;
assign \add_7s_7ns_7_2_1_U10.top_add_7s_7ns_7_2_1_Adder_3_U.u1.a  = \add_7s_7ns_7_2_1_U10.top_add_7s_7ns_7_2_1_Adder_3_U.a [2:0];
assign \add_7s_7ns_7_2_1_U10.top_add_7s_7ns_7_2_1_Adder_3_U.u1.b  = \add_7s_7ns_7_2_1_U10.top_add_7s_7ns_7_2_1_Adder_3_U.b [2:0];
assign \add_7s_7ns_7_2_1_U10.top_add_7s_7ns_7_2_1_Adder_3_U.u1.cin  = 1'h0;
assign \add_7s_7ns_7_2_1_U10.top_add_7s_7ns_7_2_1_Adder_3_U.facout_s1  = \add_7s_7ns_7_2_1_U10.top_add_7s_7ns_7_2_1_Adder_3_U.u1.cout ;
assign \add_7s_7ns_7_2_1_U10.top_add_7s_7ns_7_2_1_Adder_3_U.fas_s1  = \add_7s_7ns_7_2_1_U10.top_add_7s_7ns_7_2_1_Adder_3_U.u1.s ;
assign \add_7s_7ns_7_2_1_U10.top_add_7s_7ns_7_2_1_Adder_3_U.a  = \add_7s_7ns_7_2_1_U10.din0 ;
assign \add_7s_7ns_7_2_1_U10.top_add_7s_7ns_7_2_1_Adder_3_U.b  = \add_7s_7ns_7_2_1_U10.din1 ;
assign \add_7s_7ns_7_2_1_U10.top_add_7s_7ns_7_2_1_Adder_3_U.ce  = \add_7s_7ns_7_2_1_U10.ce ;
assign \add_7s_7ns_7_2_1_U10.top_add_7s_7ns_7_2_1_Adder_3_U.clk  = \add_7s_7ns_7_2_1_U10.clk ;
assign \add_7s_7ns_7_2_1_U10.top_add_7s_7ns_7_2_1_Adder_3_U.reset  = \add_7s_7ns_7_2_1_U10.reset ;
assign \add_7s_7ns_7_2_1_U10.dout  = \add_7s_7ns_7_2_1_U10.top_add_7s_7ns_7_2_1_Adder_3_U.s ;
assign \add_7s_7ns_7_2_1_U10.ce  = 1'h1;
assign \add_7s_7ns_7_2_1_U10.clk  = ap_clk;
assign \add_7s_7ns_7_2_1_U10.din0  = { tmp_s_reg_1920[5], tmp_s_reg_1920 };
assign \add_7s_7ns_7_2_1_U10.din1  = 7'h01;
assign grp_fu_930_p2 = \add_7s_7ns_7_2_1_U10.dout ;
assign \add_7s_7ns_7_2_1_U10.reset  = ap_rst;
assign \add_4ns_4ns_4_2_1_U3.top_add_4ns_4ns_4_2_1_Adder_2_U.ain_s0  = \add_4ns_4ns_4_2_1_U3.top_add_4ns_4ns_4_2_1_Adder_2_U.a ;
assign \add_4ns_4ns_4_2_1_U3.top_add_4ns_4ns_4_2_1_Adder_2_U.bin_s0  = \add_4ns_4ns_4_2_1_U3.top_add_4ns_4ns_4_2_1_Adder_2_U.b ;
assign \add_4ns_4ns_4_2_1_U3.top_add_4ns_4ns_4_2_1_Adder_2_U.s  = { \add_4ns_4ns_4_2_1_U3.top_add_4ns_4ns_4_2_1_Adder_2_U.fas_s2 , \add_4ns_4ns_4_2_1_U3.top_add_4ns_4ns_4_2_1_Adder_2_U.sum_s1  };
assign \add_4ns_4ns_4_2_1_U3.top_add_4ns_4ns_4_2_1_Adder_2_U.u2.a  = \add_4ns_4ns_4_2_1_U3.top_add_4ns_4ns_4_2_1_Adder_2_U.ain_s1 ;
assign \add_4ns_4ns_4_2_1_U3.top_add_4ns_4ns_4_2_1_Adder_2_U.u2.b  = \add_4ns_4ns_4_2_1_U3.top_add_4ns_4ns_4_2_1_Adder_2_U.bin_s1 ;
assign \add_4ns_4ns_4_2_1_U3.top_add_4ns_4ns_4_2_1_Adder_2_U.u2.cin  = \add_4ns_4ns_4_2_1_U3.top_add_4ns_4ns_4_2_1_Adder_2_U.carry_s1 ;
assign \add_4ns_4ns_4_2_1_U3.top_add_4ns_4ns_4_2_1_Adder_2_U.facout_s2  = \add_4ns_4ns_4_2_1_U3.top_add_4ns_4ns_4_2_1_Adder_2_U.u2.cout ;
assign \add_4ns_4ns_4_2_1_U3.top_add_4ns_4ns_4_2_1_Adder_2_U.fas_s2  = \add_4ns_4ns_4_2_1_U3.top_add_4ns_4ns_4_2_1_Adder_2_U.u2.s ;
assign \add_4ns_4ns_4_2_1_U3.top_add_4ns_4ns_4_2_1_Adder_2_U.u1.a  = \add_4ns_4ns_4_2_1_U3.top_add_4ns_4ns_4_2_1_Adder_2_U.a [1:0];
assign \add_4ns_4ns_4_2_1_U3.top_add_4ns_4ns_4_2_1_Adder_2_U.u1.b  = \add_4ns_4ns_4_2_1_U3.top_add_4ns_4ns_4_2_1_Adder_2_U.b [1:0];
assign \add_4ns_4ns_4_2_1_U3.top_add_4ns_4ns_4_2_1_Adder_2_U.u1.cin  = 1'h0;
assign \add_4ns_4ns_4_2_1_U3.top_add_4ns_4ns_4_2_1_Adder_2_U.facout_s1  = \add_4ns_4ns_4_2_1_U3.top_add_4ns_4ns_4_2_1_Adder_2_U.u1.cout ;
assign \add_4ns_4ns_4_2_1_U3.top_add_4ns_4ns_4_2_1_Adder_2_U.fas_s1  = \add_4ns_4ns_4_2_1_U3.top_add_4ns_4ns_4_2_1_Adder_2_U.u1.s ;
assign \add_4ns_4ns_4_2_1_U3.top_add_4ns_4ns_4_2_1_Adder_2_U.a  = \add_4ns_4ns_4_2_1_U3.din0 ;
assign \add_4ns_4ns_4_2_1_U3.top_add_4ns_4ns_4_2_1_Adder_2_U.b  = \add_4ns_4ns_4_2_1_U3.din1 ;
assign \add_4ns_4ns_4_2_1_U3.top_add_4ns_4ns_4_2_1_Adder_2_U.ce  = \add_4ns_4ns_4_2_1_U3.ce ;
assign \add_4ns_4ns_4_2_1_U3.top_add_4ns_4ns_4_2_1_Adder_2_U.clk  = \add_4ns_4ns_4_2_1_U3.clk ;
assign \add_4ns_4ns_4_2_1_U3.top_add_4ns_4ns_4_2_1_Adder_2_U.reset  = \add_4ns_4ns_4_2_1_U3.reset ;
assign \add_4ns_4ns_4_2_1_U3.dout  = \add_4ns_4ns_4_2_1_U3.top_add_4ns_4ns_4_2_1_Adder_2_U.s ;
assign \add_4ns_4ns_4_2_1_U3.ce  = 1'h1;
assign \add_4ns_4ns_4_2_1_U3.clk  = ap_clk;
assign \add_4ns_4ns_4_2_1_U3.din0  = ret_V_8_cast_reg_1613;
assign \add_4ns_4ns_4_2_1_U3.din1  = 4'h1;
assign grp_fu_357_p2 = \add_4ns_4ns_4_2_1_U3.dout ;
assign \add_4ns_4ns_4_2_1_U3.reset  = ap_rst;
assign \add_3s_3ns_3_2_1_U17.top_add_3s_3ns_3_2_1_Adder_10_U.ain_s0  = \add_3s_3ns_3_2_1_U17.top_add_3s_3ns_3_2_1_Adder_10_U.a ;
assign \add_3s_3ns_3_2_1_U17.top_add_3s_3ns_3_2_1_Adder_10_U.bin_s0  = \add_3s_3ns_3_2_1_U17.top_add_3s_3ns_3_2_1_Adder_10_U.b ;
assign \add_3s_3ns_3_2_1_U17.top_add_3s_3ns_3_2_1_Adder_10_U.s  = { \add_3s_3ns_3_2_1_U17.top_add_3s_3ns_3_2_1_Adder_10_U.fas_s2 , \add_3s_3ns_3_2_1_U17.top_add_3s_3ns_3_2_1_Adder_10_U.sum_s1  };
assign \add_3s_3ns_3_2_1_U17.top_add_3s_3ns_3_2_1_Adder_10_U.u2.a  = \add_3s_3ns_3_2_1_U17.top_add_3s_3ns_3_2_1_Adder_10_U.ain_s1 ;
assign \add_3s_3ns_3_2_1_U17.top_add_3s_3ns_3_2_1_Adder_10_U.u2.b  = \add_3s_3ns_3_2_1_U17.top_add_3s_3ns_3_2_1_Adder_10_U.bin_s1 ;
assign \add_3s_3ns_3_2_1_U17.top_add_3s_3ns_3_2_1_Adder_10_U.u2.cin  = \add_3s_3ns_3_2_1_U17.top_add_3s_3ns_3_2_1_Adder_10_U.carry_s1 ;
assign \add_3s_3ns_3_2_1_U17.top_add_3s_3ns_3_2_1_Adder_10_U.facout_s2  = \add_3s_3ns_3_2_1_U17.top_add_3s_3ns_3_2_1_Adder_10_U.u2.cout ;
assign \add_3s_3ns_3_2_1_U17.top_add_3s_3ns_3_2_1_Adder_10_U.fas_s2  = \add_3s_3ns_3_2_1_U17.top_add_3s_3ns_3_2_1_Adder_10_U.u2.s ;
assign \add_3s_3ns_3_2_1_U17.top_add_3s_3ns_3_2_1_Adder_10_U.u1.a  = \add_3s_3ns_3_2_1_U17.top_add_3s_3ns_3_2_1_Adder_10_U.a [0];
assign \add_3s_3ns_3_2_1_U17.top_add_3s_3ns_3_2_1_Adder_10_U.u1.b  = \add_3s_3ns_3_2_1_U17.top_add_3s_3ns_3_2_1_Adder_10_U.b [0];
assign \add_3s_3ns_3_2_1_U17.top_add_3s_3ns_3_2_1_Adder_10_U.u1.cin  = 1'h0;
assign \add_3s_3ns_3_2_1_U17.top_add_3s_3ns_3_2_1_Adder_10_U.facout_s1  = \add_3s_3ns_3_2_1_U17.top_add_3s_3ns_3_2_1_Adder_10_U.u1.cout ;
assign \add_3s_3ns_3_2_1_U17.top_add_3s_3ns_3_2_1_Adder_10_U.fas_s1  = \add_3s_3ns_3_2_1_U17.top_add_3s_3ns_3_2_1_Adder_10_U.u1.s ;
assign \add_3s_3ns_3_2_1_U17.top_add_3s_3ns_3_2_1_Adder_10_U.a  = \add_3s_3ns_3_2_1_U17.din0 ;
assign \add_3s_3ns_3_2_1_U17.top_add_3s_3ns_3_2_1_Adder_10_U.b  = \add_3s_3ns_3_2_1_U17.din1 ;
assign \add_3s_3ns_3_2_1_U17.top_add_3s_3ns_3_2_1_Adder_10_U.ce  = \add_3s_3ns_3_2_1_U17.ce ;
assign \add_3s_3ns_3_2_1_U17.top_add_3s_3ns_3_2_1_Adder_10_U.clk  = \add_3s_3ns_3_2_1_U17.clk ;
assign \add_3s_3ns_3_2_1_U17.top_add_3s_3ns_3_2_1_Adder_10_U.reset  = \add_3s_3ns_3_2_1_U17.reset ;
assign \add_3s_3ns_3_2_1_U17.dout  = \add_3s_3ns_3_2_1_U17.top_add_3s_3ns_3_2_1_Adder_10_U.s ;
assign \add_3s_3ns_3_2_1_U17.ce  = 1'h1;
assign \add_3s_3ns_3_2_1_U17.clk  = ap_clk;
assign \add_3s_3ns_3_2_1_U17.din0  = { trunc_ln708_1_reg_2040[1], trunc_ln708_1_reg_2040 };
assign \add_3s_3ns_3_2_1_U17.din1  = { 2'h0, and_ln414_1_reg_2087 };
assign grp_fu_1234_p2 = \add_3s_3ns_3_2_1_U17.dout ;
assign \add_3s_3ns_3_2_1_U17.reset  = ap_rst;
assign \add_37s_37s_37_2_1_U18.top_add_37s_37s_37_2_1_Adder_11_U.ain_s0  = \add_37s_37s_37_2_1_U18.top_add_37s_37s_37_2_1_Adder_11_U.a ;
assign \add_37s_37s_37_2_1_U18.top_add_37s_37s_37_2_1_Adder_11_U.bin_s0  = \add_37s_37s_37_2_1_U18.top_add_37s_37s_37_2_1_Adder_11_U.b ;
assign \add_37s_37s_37_2_1_U18.top_add_37s_37s_37_2_1_Adder_11_U.s  = { \add_37s_37s_37_2_1_U18.top_add_37s_37s_37_2_1_Adder_11_U.fas_s2 , \add_37s_37s_37_2_1_U18.top_add_37s_37s_37_2_1_Adder_11_U.sum_s1  };
assign \add_37s_37s_37_2_1_U18.top_add_37s_37s_37_2_1_Adder_11_U.u2.a  = \add_37s_37s_37_2_1_U18.top_add_37s_37s_37_2_1_Adder_11_U.ain_s1 ;
assign \add_37s_37s_37_2_1_U18.top_add_37s_37s_37_2_1_Adder_11_U.u2.b  = \add_37s_37s_37_2_1_U18.top_add_37s_37s_37_2_1_Adder_11_U.bin_s1 ;
assign \add_37s_37s_37_2_1_U18.top_add_37s_37s_37_2_1_Adder_11_U.u2.cin  = \add_37s_37s_37_2_1_U18.top_add_37s_37s_37_2_1_Adder_11_U.carry_s1 ;
assign \add_37s_37s_37_2_1_U18.top_add_37s_37s_37_2_1_Adder_11_U.facout_s2  = \add_37s_37s_37_2_1_U18.top_add_37s_37s_37_2_1_Adder_11_U.u2.cout ;
assign \add_37s_37s_37_2_1_U18.top_add_37s_37s_37_2_1_Adder_11_U.fas_s2  = \add_37s_37s_37_2_1_U18.top_add_37s_37s_37_2_1_Adder_11_U.u2.s ;
assign \add_37s_37s_37_2_1_U18.top_add_37s_37s_37_2_1_Adder_11_U.u1.a  = \add_37s_37s_37_2_1_U18.top_add_37s_37s_37_2_1_Adder_11_U.a [17:0];
assign \add_37s_37s_37_2_1_U18.top_add_37s_37s_37_2_1_Adder_11_U.u1.b  = \add_37s_37s_37_2_1_U18.top_add_37s_37s_37_2_1_Adder_11_U.b [17:0];
assign \add_37s_37s_37_2_1_U18.top_add_37s_37s_37_2_1_Adder_11_U.u1.cin  = 1'h0;
assign \add_37s_37s_37_2_1_U18.top_add_37s_37s_37_2_1_Adder_11_U.facout_s1  = \add_37s_37s_37_2_1_U18.top_add_37s_37s_37_2_1_Adder_11_U.u1.cout ;
assign \add_37s_37s_37_2_1_U18.top_add_37s_37s_37_2_1_Adder_11_U.fas_s1  = \add_37s_37s_37_2_1_U18.top_add_37s_37s_37_2_1_Adder_11_U.u1.s ;
assign \add_37s_37s_37_2_1_U18.top_add_37s_37s_37_2_1_Adder_11_U.a  = \add_37s_37s_37_2_1_U18.din0 ;
assign \add_37s_37s_37_2_1_U18.top_add_37s_37s_37_2_1_Adder_11_U.b  = \add_37s_37s_37_2_1_U18.din1 ;
assign \add_37s_37s_37_2_1_U18.top_add_37s_37s_37_2_1_Adder_11_U.ce  = \add_37s_37s_37_2_1_U18.ce ;
assign \add_37s_37s_37_2_1_U18.top_add_37s_37s_37_2_1_Adder_11_U.clk  = \add_37s_37s_37_2_1_U18.clk ;
assign \add_37s_37s_37_2_1_U18.top_add_37s_37s_37_2_1_Adder_11_U.reset  = \add_37s_37s_37_2_1_U18.reset ;
assign \add_37s_37s_37_2_1_U18.dout  = \add_37s_37s_37_2_1_U18.top_add_37s_37s_37_2_1_Adder_11_U.s ;
assign \add_37s_37s_37_2_1_U18.ce  = 1'h1;
assign \add_37s_37s_37_2_1_U18.clk  = ap_clk;
assign \add_37s_37s_37_2_1_U18.din0  = { op_23_V_reg_2097[31], op_23_V_reg_2097, 4'h0 };
assign \add_37s_37s_37_2_1_U18.din1  = { ret_V_9_reg_2092[6], ret_V_9_reg_2092[6], ret_V_9_reg_2092[6], ret_V_9_reg_2092[6], ret_V_9_reg_2092[6], ret_V_9_reg_2092[6], ret_V_9_reg_2092[6], ret_V_9_reg_2092[6], ret_V_9_reg_2092[6], ret_V_9_reg_2092[6], ret_V_9_reg_2092[6], ret_V_9_reg_2092[6], ret_V_9_reg_2092[6], ret_V_9_reg_2092[6], ret_V_9_reg_2092[6], ret_V_9_reg_2092[6], ret_V_9_reg_2092[6], ret_V_9_reg_2092[6], ret_V_9_reg_2092[6], ret_V_9_reg_2092[6], ret_V_9_reg_2092[6], ret_V_9_reg_2092[6], ret_V_9_reg_2092[6], ret_V_9_reg_2092[6], ret_V_9_reg_2092[6], ret_V_9_reg_2092[6], ret_V_9_reg_2092[6], ret_V_9_reg_2092[6], ret_V_9_reg_2092[6], ret_V_9_reg_2092, 1'h0 };
assign grp_fu_1262_p2 = \add_37s_37s_37_2_1_U18.dout ;
assign \add_37s_37s_37_2_1_U18.reset  = ap_rst;
assign \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_6_U.ain_s0  = \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_6_U.a ;
assign \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_6_U.bin_s0  = \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_6_U.b ;
assign \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_6_U.s  = { \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_6_U.fas_s2 , \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_6_U.sum_s1  };
assign \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_6_U.u2.a  = \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_6_U.ain_s1 ;
assign \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_6_U.u2.b  = \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_6_U.bin_s1 ;
assign \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_6_U.u2.cin  = \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_6_U.carry_s1 ;
assign \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_6_U.facout_s2  = \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_6_U.u2.cout ;
assign \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_6_U.fas_s2  = \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_6_U.u2.s ;
assign \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_6_U.u1.a  = \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_6_U.a [16:0];
assign \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_6_U.u1.b  = \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_6_U.b [16:0];
assign \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_6_U.u1.cin  = 1'h0;
assign \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_6_U.facout_s1  = \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_6_U.u1.cout ;
assign \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_6_U.fas_s1  = \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_6_U.u1.s ;
assign \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_6_U.a  = \add_34s_34s_34_2_1_U24.din0 ;
assign \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_6_U.b  = \add_34s_34s_34_2_1_U24.din1 ;
assign \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_6_U.ce  = \add_34s_34s_34_2_1_U24.ce ;
assign \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_6_U.clk  = \add_34s_34s_34_2_1_U24.clk ;
assign \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_6_U.reset  = \add_34s_34s_34_2_1_U24.reset ;
assign \add_34s_34s_34_2_1_U24.dout  = \add_34s_34s_34_2_1_U24.top_add_34s_34s_34_2_1_Adder_6_U.s ;
assign \add_34s_34s_34_2_1_U24.ce  = 1'h1;
assign \add_34s_34s_34_2_1_U24.clk  = ap_clk;
assign \add_34s_34s_34_2_1_U24.din0  = { op_26_V_reg_2252[31], op_26_V_reg_2252, 1'h0 };
assign \add_34s_34s_34_2_1_U24.din1  = { op_19_V_reg_2193[3], op_19_V_reg_2193[3], op_19_V_reg_2193[3], op_19_V_reg_2193[3], op_19_V_reg_2193[3], op_19_V_reg_2193[3], op_19_V_reg_2193[3], op_19_V_reg_2193[3], op_19_V_reg_2193[3], op_19_V_reg_2193[3], op_19_V_reg_2193[3], op_19_V_reg_2193[3], op_19_V_reg_2193[3], op_19_V_reg_2193[3], op_19_V_reg_2193[3], op_19_V_reg_2193[3], op_19_V_reg_2193[3], op_19_V_reg_2193[3], op_19_V_reg_2193[3], op_19_V_reg_2193[3], op_19_V_reg_2193[3], op_19_V_reg_2193[3], op_19_V_reg_2193[3], op_19_V_reg_2193[3], op_19_V_reg_2193[3], op_19_V_reg_2193[3], op_19_V_reg_2193[3], op_19_V_reg_2193[3], op_19_V_reg_2193[3], op_19_V_reg_2193[3], op_19_V_reg_2193 };
assign grp_fu_1516_p2 = \add_34s_34s_34_2_1_U24.dout ;
assign \add_34s_34s_34_2_1_U24.reset  = ap_rst;
assign \add_34s_34s_34_2_1_U21.top_add_34s_34s_34_2_1_Adder_6_U.ain_s0  = \add_34s_34s_34_2_1_U21.top_add_34s_34s_34_2_1_Adder_6_U.a ;
assign \add_34s_34s_34_2_1_U21.top_add_34s_34s_34_2_1_Adder_6_U.bin_s0  = \add_34s_34s_34_2_1_U21.top_add_34s_34s_34_2_1_Adder_6_U.b ;
assign \add_34s_34s_34_2_1_U21.top_add_34s_34s_34_2_1_Adder_6_U.s  = { \add_34s_34s_34_2_1_U21.top_add_34s_34s_34_2_1_Adder_6_U.fas_s2 , \add_34s_34s_34_2_1_U21.top_add_34s_34s_34_2_1_Adder_6_U.sum_s1  };
assign \add_34s_34s_34_2_1_U21.top_add_34s_34s_34_2_1_Adder_6_U.u2.a  = \add_34s_34s_34_2_1_U21.top_add_34s_34s_34_2_1_Adder_6_U.ain_s1 ;
assign \add_34s_34s_34_2_1_U21.top_add_34s_34s_34_2_1_Adder_6_U.u2.b  = \add_34s_34s_34_2_1_U21.top_add_34s_34s_34_2_1_Adder_6_U.bin_s1 ;
assign \add_34s_34s_34_2_1_U21.top_add_34s_34s_34_2_1_Adder_6_U.u2.cin  = \add_34s_34s_34_2_1_U21.top_add_34s_34s_34_2_1_Adder_6_U.carry_s1 ;
assign \add_34s_34s_34_2_1_U21.top_add_34s_34s_34_2_1_Adder_6_U.facout_s2  = \add_34s_34s_34_2_1_U21.top_add_34s_34s_34_2_1_Adder_6_U.u2.cout ;
assign \add_34s_34s_34_2_1_U21.top_add_34s_34s_34_2_1_Adder_6_U.fas_s2  = \add_34s_34s_34_2_1_U21.top_add_34s_34s_34_2_1_Adder_6_U.u2.s ;
assign \add_34s_34s_34_2_1_U21.top_add_34s_34s_34_2_1_Adder_6_U.u1.a  = \add_34s_34s_34_2_1_U21.top_add_34s_34s_34_2_1_Adder_6_U.a [16:0];
assign \add_34s_34s_34_2_1_U21.top_add_34s_34s_34_2_1_Adder_6_U.u1.b  = \add_34s_34s_34_2_1_U21.top_add_34s_34s_34_2_1_Adder_6_U.b [16:0];
assign \add_34s_34s_34_2_1_U21.top_add_34s_34s_34_2_1_Adder_6_U.u1.cin  = 1'h0;
assign \add_34s_34s_34_2_1_U21.top_add_34s_34s_34_2_1_Adder_6_U.facout_s1  = \add_34s_34s_34_2_1_U21.top_add_34s_34s_34_2_1_Adder_6_U.u1.cout ;
assign \add_34s_34s_34_2_1_U21.top_add_34s_34s_34_2_1_Adder_6_U.fas_s1  = \add_34s_34s_34_2_1_U21.top_add_34s_34s_34_2_1_Adder_6_U.u1.s ;
assign \add_34s_34s_34_2_1_U21.top_add_34s_34s_34_2_1_Adder_6_U.a  = \add_34s_34s_34_2_1_U21.din0 ;
assign \add_34s_34s_34_2_1_U21.top_add_34s_34s_34_2_1_Adder_6_U.b  = \add_34s_34s_34_2_1_U21.din1 ;
assign \add_34s_34s_34_2_1_U21.top_add_34s_34s_34_2_1_Adder_6_U.ce  = \add_34s_34s_34_2_1_U21.ce ;
assign \add_34s_34s_34_2_1_U21.top_add_34s_34s_34_2_1_Adder_6_U.clk  = \add_34s_34s_34_2_1_U21.clk ;
assign \add_34s_34s_34_2_1_U21.top_add_34s_34s_34_2_1_Adder_6_U.reset  = \add_34s_34s_34_2_1_U21.reset ;
assign \add_34s_34s_34_2_1_U21.dout  = \add_34s_34s_34_2_1_U21.top_add_34s_34s_34_2_1_Adder_6_U.s ;
assign \add_34s_34s_34_2_1_U21.ce  = 1'h1;
assign \add_34s_34s_34_2_1_U21.clk  = ap_clk;
assign \add_34s_34s_34_2_1_U21.din0  = { select_ln353_2_reg_2210[31], select_ln353_2_reg_2210, 1'h0 };
assign \add_34s_34s_34_2_1_U21.din1  = { op_17_V_reg_2204[1], op_17_V_reg_2204[1], op_17_V_reg_2204[1], op_17_V_reg_2204[1], op_17_V_reg_2204[1], op_17_V_reg_2204[1], op_17_V_reg_2204[1], op_17_V_reg_2204[1], op_17_V_reg_2204[1], op_17_V_reg_2204[1], op_17_V_reg_2204[1], op_17_V_reg_2204[1], op_17_V_reg_2204[1], op_17_V_reg_2204[1], op_17_V_reg_2204[1], op_17_V_reg_2204[1], op_17_V_reg_2204[1], op_17_V_reg_2204[1], op_17_V_reg_2204[1], op_17_V_reg_2204[1], op_17_V_reg_2204[1], op_17_V_reg_2204[1], op_17_V_reg_2204[1], op_17_V_reg_2204[1], op_17_V_reg_2204[1], op_17_V_reg_2204[1], op_17_V_reg_2204[1], op_17_V_reg_2204[1], op_17_V_reg_2204[1], op_17_V_reg_2204[1], op_17_V_reg_2204[1], op_17_V_reg_2204[1], op_17_V_reg_2204 };
assign grp_fu_1449_p2 = \add_34s_34s_34_2_1_U21.dout ;
assign \add_34s_34s_34_2_1_U21.reset  = ap_rst;
assign \add_34s_34s_34_2_1_U12.top_add_34s_34s_34_2_1_Adder_6_U.ain_s0  = \add_34s_34s_34_2_1_U12.top_add_34s_34s_34_2_1_Adder_6_U.a ;
assign \add_34s_34s_34_2_1_U12.top_add_34s_34s_34_2_1_Adder_6_U.bin_s0  = \add_34s_34s_34_2_1_U12.top_add_34s_34s_34_2_1_Adder_6_U.b ;
assign \add_34s_34s_34_2_1_U12.top_add_34s_34s_34_2_1_Adder_6_U.s  = { \add_34s_34s_34_2_1_U12.top_add_34s_34s_34_2_1_Adder_6_U.fas_s2 , \add_34s_34s_34_2_1_U12.top_add_34s_34s_34_2_1_Adder_6_U.sum_s1  };
assign \add_34s_34s_34_2_1_U12.top_add_34s_34s_34_2_1_Adder_6_U.u2.a  = \add_34s_34s_34_2_1_U12.top_add_34s_34s_34_2_1_Adder_6_U.ain_s1 ;
assign \add_34s_34s_34_2_1_U12.top_add_34s_34s_34_2_1_Adder_6_U.u2.b  = \add_34s_34s_34_2_1_U12.top_add_34s_34s_34_2_1_Adder_6_U.bin_s1 ;
assign \add_34s_34s_34_2_1_U12.top_add_34s_34s_34_2_1_Adder_6_U.u2.cin  = \add_34s_34s_34_2_1_U12.top_add_34s_34s_34_2_1_Adder_6_U.carry_s1 ;
assign \add_34s_34s_34_2_1_U12.top_add_34s_34s_34_2_1_Adder_6_U.facout_s2  = \add_34s_34s_34_2_1_U12.top_add_34s_34s_34_2_1_Adder_6_U.u2.cout ;
assign \add_34s_34s_34_2_1_U12.top_add_34s_34s_34_2_1_Adder_6_U.fas_s2  = \add_34s_34s_34_2_1_U12.top_add_34s_34s_34_2_1_Adder_6_U.u2.s ;
assign \add_34s_34s_34_2_1_U12.top_add_34s_34s_34_2_1_Adder_6_U.u1.a  = \add_34s_34s_34_2_1_U12.top_add_34s_34s_34_2_1_Adder_6_U.a [16:0];
assign \add_34s_34s_34_2_1_U12.top_add_34s_34s_34_2_1_Adder_6_U.u1.b  = \add_34s_34s_34_2_1_U12.top_add_34s_34s_34_2_1_Adder_6_U.b [16:0];
assign \add_34s_34s_34_2_1_U12.top_add_34s_34s_34_2_1_Adder_6_U.u1.cin  = 1'h0;
assign \add_34s_34s_34_2_1_U12.top_add_34s_34s_34_2_1_Adder_6_U.facout_s1  = \add_34s_34s_34_2_1_U12.top_add_34s_34s_34_2_1_Adder_6_U.u1.cout ;
assign \add_34s_34s_34_2_1_U12.top_add_34s_34s_34_2_1_Adder_6_U.fas_s1  = \add_34s_34s_34_2_1_U12.top_add_34s_34s_34_2_1_Adder_6_U.u1.s ;
assign \add_34s_34s_34_2_1_U12.top_add_34s_34s_34_2_1_Adder_6_U.a  = \add_34s_34s_34_2_1_U12.din0 ;
assign \add_34s_34s_34_2_1_U12.top_add_34s_34s_34_2_1_Adder_6_U.b  = \add_34s_34s_34_2_1_U12.din1 ;
assign \add_34s_34s_34_2_1_U12.top_add_34s_34s_34_2_1_Adder_6_U.ce  = \add_34s_34s_34_2_1_U12.ce ;
assign \add_34s_34s_34_2_1_U12.top_add_34s_34s_34_2_1_Adder_6_U.clk  = \add_34s_34s_34_2_1_U12.clk ;
assign \add_34s_34s_34_2_1_U12.top_add_34s_34s_34_2_1_Adder_6_U.reset  = \add_34s_34s_34_2_1_U12.reset ;
assign \add_34s_34s_34_2_1_U12.dout  = \add_34s_34s_34_2_1_U12.top_add_34s_34s_34_2_1_Adder_6_U.s ;
assign \add_34s_34s_34_2_1_U12.ce  = 1'h1;
assign \add_34s_34s_34_2_1_U12.clk  = ap_clk;
assign \add_34s_34s_34_2_1_U12.din0  = { select_ln353_reg_1959[6], select_ln353_reg_1959[6], select_ln353_reg_1959[6], select_ln353_reg_1959[6], select_ln353_reg_1959[6], select_ln353_reg_1959[6], select_ln353_reg_1959[6], select_ln353_reg_1959[6], select_ln353_reg_1959[6], select_ln353_reg_1959[6], select_ln353_reg_1959[6], select_ln353_reg_1959[6], select_ln353_reg_1959[6], select_ln353_reg_1959[6], select_ln353_reg_1959[6], select_ln353_reg_1959[6], select_ln353_reg_1959[6], select_ln353_reg_1959[6], select_ln353_reg_1959[6], select_ln353_reg_1959[6], select_ln353_reg_1959[6], select_ln353_reg_1959[6], select_ln353_reg_1959[6], select_ln353_reg_1959[6], select_ln353_reg_1959[6], select_ln353_reg_1959[6], select_ln353_reg_1959, 1'h0 };
assign \add_34s_34s_34_2_1_U12.din1  = { op_14_V_reg_1953[1], op_14_V_reg_1953[1], op_14_V_reg_1953[1], op_14_V_reg_1953[1], op_14_V_reg_1953[1], op_14_V_reg_1953[1], op_14_V_reg_1953[1], op_14_V_reg_1953[1], op_14_V_reg_1953[1], op_14_V_reg_1953[1], op_14_V_reg_1953[1], op_14_V_reg_1953[1], op_14_V_reg_1953[1], op_14_V_reg_1953[1], op_14_V_reg_1953[1], op_14_V_reg_1953[1], op_14_V_reg_1953[1], op_14_V_reg_1953[1], op_14_V_reg_1953[1], op_14_V_reg_1953[1], op_14_V_reg_1953[1], op_14_V_reg_1953[1], op_14_V_reg_1953[1], op_14_V_reg_1953[1], op_14_V_reg_1953[1], op_14_V_reg_1953[1], op_14_V_reg_1953[1], op_14_V_reg_1953[1], op_14_V_reg_1953[1], op_14_V_reg_1953[1], op_14_V_reg_1953[1], op_14_V_reg_1953[1], op_14_V_reg_1953 };
assign grp_fu_1015_p2 = \add_34s_34s_34_2_1_U12.dout ;
assign \add_34s_34s_34_2_1_U12.reset  = ap_rst;
assign \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_9_U.ain_s0  = \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_9_U.a ;
assign \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_9_U.bin_s0  = \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_9_U.b ;
assign \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_9_U.s  = { \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_9_U.fas_s2 , \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_9_U.sum_s1  };
assign \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_9_U.u2.a  = \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_9_U.ain_s1 ;
assign \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_9_U.u2.b  = \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_9_U.bin_s1 ;
assign \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_9_U.u2.cin  = \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_9_U.carry_s1 ;
assign \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_9_U.facout_s2  = \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_9_U.u2.cout ;
assign \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_9_U.fas_s2  = \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_9_U.u2.s ;
assign \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_9_U.u1.a  = \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_9_U.a [15:0];
assign \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_9_U.u1.b  = \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_9_U.b [15:0];
assign \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_9_U.u1.cin  = 1'h0;
assign \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_9_U.facout_s1  = \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_9_U.u1.cout ;
assign \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_9_U.fas_s1  = \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_9_U.u1.s ;
assign \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_9_U.a  = \add_32ns_32s_32_2_1_U23.din0 ;
assign \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_9_U.b  = \add_32ns_32s_32_2_1_U23.din1 ;
assign \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_9_U.ce  = \add_32ns_32s_32_2_1_U23.ce ;
assign \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_9_U.clk  = \add_32ns_32s_32_2_1_U23.clk ;
assign \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_9_U.reset  = \add_32ns_32s_32_2_1_U23.reset ;
assign \add_32ns_32s_32_2_1_U23.dout  = \add_32ns_32s_32_2_1_U23.top_add_32ns_32s_32_2_1_Adder_9_U.s ;
assign \add_32ns_32s_32_2_1_U23.ce  = 1'h1;
assign \add_32ns_32s_32_2_1_U23.clk  = ap_clk;
assign \add_32ns_32s_32_2_1_U23.din0  = ret_V_27_reg_2242;
assign \add_32ns_32s_32_2_1_U23.din1  = { op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18 };
assign grp_fu_1497_p2 = \add_32ns_32s_32_2_1_U23.dout ;
assign \add_32ns_32s_32_2_1_U23.reset  = ap_rst;
assign \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.ain_s0  = \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.a ;
assign \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.bin_s0  = \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.b ;
assign \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.s  = { \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.fas_s2 , \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.sum_s1  };
assign \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.u2.a  = \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.ain_s1 ;
assign \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.u2.b  = \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.bin_s1 ;
assign \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.u2.cin  = \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.carry_s1 ;
assign \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.facout_s2  = \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.u2.cout ;
assign \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.fas_s2  = \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.u2.s ;
assign \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.u1.a  = \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.a [15:0];
assign \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.u1.b  = \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.b [15:0];
assign \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.u1.cin  = 1'h0;
assign \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.facout_s1  = \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.u1.cout ;
assign \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.fas_s1  = \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.u1.s ;
assign \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.a  = \add_32ns_32s_32_2_1_U16.din0 ;
assign \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.b  = \add_32ns_32s_32_2_1_U16.din1 ;
assign \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.ce  = \add_32ns_32s_32_2_1_U16.ce ;
assign \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.clk  = \add_32ns_32s_32_2_1_U16.clk ;
assign \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.reset  = \add_32ns_32s_32_2_1_U16.reset ;
assign \add_32ns_32s_32_2_1_U16.dout  = \add_32ns_32s_32_2_1_U16.top_add_32ns_32s_32_2_1_Adder_9_U.s ;
assign \add_32ns_32s_32_2_1_U16.ce  = 1'h1;
assign \add_32ns_32s_32_2_1_U16.clk  = ap_clk;
assign \add_32ns_32s_32_2_1_U16.din0  = ret_V_24_reg_2045;
assign \add_32ns_32s_32_2_1_U16.din1  = { ret_V_19_reg_2023[1], ret_V_19_reg_2023[1], ret_V_19_reg_2023[1], ret_V_19_reg_2023[1], ret_V_19_reg_2023[1], ret_V_19_reg_2023[1], ret_V_19_reg_2023[1], ret_V_19_reg_2023[1], ret_V_19_reg_2023[1], ret_V_19_reg_2023[1], ret_V_19_reg_2023[1], ret_V_19_reg_2023[1], ret_V_19_reg_2023[1], ret_V_19_reg_2023[1], ret_V_19_reg_2023[1], ret_V_19_reg_2023[1], ret_V_19_reg_2023[1], ret_V_19_reg_2023[1], ret_V_19_reg_2023[1], ret_V_19_reg_2023[1], ret_V_19_reg_2023[1], ret_V_19_reg_2023[1], ret_V_19_reg_2023[1], ret_V_19_reg_2023[1], ret_V_19_reg_2023[1], ret_V_19_reg_2023[1], ret_V_19_reg_2023[1], ret_V_19_reg_2023[1], ret_V_19_reg_2023[1], ret_V_19_reg_2023[1], ret_V_19_reg_2023 };
assign grp_fu_1192_p2 = \add_32ns_32s_32_2_1_U16.dout ;
assign \add_32ns_32s_32_2_1_U16.reset  = ap_rst;
assign \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s0  = \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_7_U.a ;
assign \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s0  = \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_7_U.b ;
assign \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_7_U.s  = { \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s2 , \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_7_U.sum_s1  };
assign \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.a  = \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s1 ;
assign \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.b  = \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s1 ;
assign \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cin  = \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_7_U.carry_s1 ;
assign \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_7_U.facout_s2  = \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cout ;
assign \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s2  = \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.s ;
assign \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.a  = \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_7_U.a [15:0];
assign \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.b  = \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_7_U.b [15:0];
assign \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cin  = 1'h0;
assign \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_7_U.facout_s1  = \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cout ;
assign \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s1  = \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.s ;
assign \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_7_U.a  = \add_32ns_32ns_32_2_1_U25.din0 ;
assign \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_7_U.b  = \add_32ns_32ns_32_2_1_U25.din1 ;
assign \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_7_U.ce  = \add_32ns_32ns_32_2_1_U25.ce ;
assign \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_7_U.clk  = \add_32ns_32ns_32_2_1_U25.clk ;
assign \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_7_U.reset  = \add_32ns_32ns_32_2_1_U25.reset ;
assign \add_32ns_32ns_32_2_1_U25.dout  = \add_32ns_32ns_32_2_1_U25.top_add_32ns_32ns_32_2_1_Adder_7_U.s ;
assign \add_32ns_32ns_32_2_1_U25.ce  = 1'h1;
assign \add_32ns_32ns_32_2_1_U25.clk  = ap_clk;
assign \add_32ns_32ns_32_2_1_U25.din0  = ret_V_28_cast_reg_2272;
assign \add_32ns_32ns_32_2_1_U25.din1  = 32'd1;
assign grp_fu_1532_p2 = \add_32ns_32ns_32_2_1_U25.dout ;
assign \add_32ns_32ns_32_2_1_U25.reset  = ap_rst;
assign \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s0  = \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_7_U.a ;
assign \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s0  = \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_7_U.b ;
assign \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_7_U.s  = { \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s2 , \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_7_U.sum_s1  };
assign \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.a  = \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s1 ;
assign \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.b  = \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s1 ;
assign \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cin  = \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_7_U.carry_s1 ;
assign \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_7_U.facout_s2  = \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cout ;
assign \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s2  = \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.s ;
assign \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.a  = \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_7_U.a [15:0];
assign \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.b  = \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_7_U.b [15:0];
assign \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cin  = 1'h0;
assign \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_7_U.facout_s1  = \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cout ;
assign \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s1  = \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.s ;
assign \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_7_U.a  = \add_32ns_32ns_32_2_1_U22.din0 ;
assign \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_7_U.b  = \add_32ns_32ns_32_2_1_U22.din1 ;
assign \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_7_U.ce  = \add_32ns_32ns_32_2_1_U22.ce ;
assign \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_7_U.clk  = \add_32ns_32ns_32_2_1_U22.clk ;
assign \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_7_U.reset  = \add_32ns_32ns_32_2_1_U22.reset ;
assign \add_32ns_32ns_32_2_1_U22.dout  = \add_32ns_32ns_32_2_1_U22.top_add_32ns_32ns_32_2_1_Adder_7_U.s ;
assign \add_32ns_32ns_32_2_1_U22.ce  = 1'h1;
assign \add_32ns_32ns_32_2_1_U22.clk  = ap_clk;
assign \add_32ns_32ns_32_2_1_U22.din0  = ret_V_25_cast_reg_2230;
assign \add_32ns_32ns_32_2_1_U22.din1  = 32'd1;
assign grp_fu_1465_p2 = \add_32ns_32ns_32_2_1_U22.dout ;
assign \add_32ns_32ns_32_2_1_U22.reset  = ap_rst;
assign \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s0  = \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_7_U.a ;
assign \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s0  = \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_7_U.b ;
assign \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_7_U.s  = { \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s2 , \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_7_U.sum_s1  };
assign \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.a  = \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s1 ;
assign \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.b  = \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s1 ;
assign \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cin  = \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_7_U.carry_s1 ;
assign \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_7_U.facout_s2  = \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cout ;
assign \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s2  = \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.s ;
assign \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.a  = \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_7_U.a [15:0];
assign \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.b  = \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_7_U.b [15:0];
assign \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cin  = 1'h0;
assign \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_7_U.facout_s1  = \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cout ;
assign \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s1  = \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.s ;
assign \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_7_U.a  = \add_32ns_32ns_32_2_1_U20.din0 ;
assign \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_7_U.b  = \add_32ns_32ns_32_2_1_U20.din1 ;
assign \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_7_U.ce  = \add_32ns_32ns_32_2_1_U20.ce ;
assign \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_7_U.clk  = \add_32ns_32ns_32_2_1_U20.clk ;
assign \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_7_U.reset  = \add_32ns_32ns_32_2_1_U20.reset ;
assign \add_32ns_32ns_32_2_1_U20.dout  = \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_7_U.s ;
assign \add_32ns_32ns_32_2_1_U20.ce  = 1'h1;
assign \add_32ns_32ns_32_2_1_U20.clk  = ap_clk;
assign \add_32ns_32ns_32_2_1_U20.din0  = ret_V_22_cast_reg_2160;
assign \add_32ns_32ns_32_2_1_U20.din1  = 32'd1;
assign grp_fu_1361_p2 = \add_32ns_32ns_32_2_1_U20.dout ;
assign \add_32ns_32ns_32_2_1_U20.reset  = ap_rst;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s0  = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.a ;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s0  = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.b ;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.s  = { \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s2 , \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.sum_s1  };
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.a  = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s1 ;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.b  = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s1 ;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cin  = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.carry_s1 ;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.facout_s2  = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cout ;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s2  = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.s ;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.a  = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.a [15:0];
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.b  = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.b [15:0];
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cin  = 1'h0;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.facout_s1  = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cout ;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s1  = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.s ;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.a  = \add_32ns_32ns_32_2_1_U14.din0 ;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.b  = \add_32ns_32ns_32_2_1_U14.din1 ;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.ce  = \add_32ns_32ns_32_2_1_U14.ce ;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.clk  = \add_32ns_32ns_32_2_1_U14.clk ;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.reset  = \add_32ns_32ns_32_2_1_U14.reset ;
assign \add_32ns_32ns_32_2_1_U14.dout  = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.s ;
assign \add_32ns_32ns_32_2_1_U14.ce  = 1'h1;
assign \add_32ns_32ns_32_2_1_U14.clk  = ap_clk;
assign \add_32ns_32ns_32_2_1_U14.din0  = ret_V_19_cast_reg_2001;
assign \add_32ns_32ns_32_2_1_U14.din1  = 32'd1;
assign grp_fu_1055_p2 = \add_32ns_32ns_32_2_1_U14.dout ;
assign \add_32ns_32ns_32_2_1_U14.reset  = ap_rst;
assign \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_4_U.ain_s0  = \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_4_U.a ;
assign \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_4_U.bin_s0  = \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_4_U.b ;
assign \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_4_U.s  = { \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_4_U.fas_s2 , \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_4_U.sum_s1  };
assign \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_4_U.u2.a  = \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_4_U.ain_s1 ;
assign \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_4_U.u2.b  = \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_4_U.bin_s1 ;
assign \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_4_U.u2.cin  = \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_4_U.carry_s1 ;
assign \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_4_U.facout_s2  = \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_4_U.u2.cout ;
assign \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_4_U.fas_s2  = \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_4_U.u2.s ;
assign \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_4_U.u1.a  = \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_4_U.a [0];
assign \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_4_U.u1.b  = \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_4_U.b [0];
assign \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_4_U.u1.cin  = 1'h0;
assign \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_4_U.facout_s1  = \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_4_U.u1.cout ;
assign \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_4_U.fas_s1  = \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_4_U.u1.s ;
assign \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_4_U.a  = \add_2ns_2ns_2_2_1_U7.din0 ;
assign \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_4_U.b  = \add_2ns_2ns_2_2_1_U7.din1 ;
assign \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_4_U.ce  = \add_2ns_2ns_2_2_1_U7.ce ;
assign \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_4_U.clk  = \add_2ns_2ns_2_2_1_U7.clk ;
assign \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_4_U.reset  = \add_2ns_2ns_2_2_1_U7.reset ;
assign \add_2ns_2ns_2_2_1_U7.dout  = \add_2ns_2ns_2_2_1_U7.top_add_2ns_2ns_2_2_1_Adder_4_U.s ;
assign \add_2ns_2ns_2_2_1_U7.ce  = 1'h1;
assign \add_2ns_2ns_2_2_1_U7.clk  = ap_clk;
assign \add_2ns_2ns_2_2_1_U7.din0  = p_Val2_8_reg_1818;
assign \add_2ns_2ns_2_2_1_U7.din1  = { 1'h0, and_ln412_reg_1833 };
assign grp_fu_752_p2 = \add_2ns_2ns_2_2_1_U7.dout ;
assign \add_2ns_2ns_2_2_1_U7.reset  = ap_rst;
assign \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_4_U.ain_s0  = \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_4_U.a ;
assign \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_4_U.bin_s0  = \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_4_U.b ;
assign \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_4_U.s  = { \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_4_U.fas_s2 , \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_4_U.sum_s1  };
assign \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_4_U.u2.a  = \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_4_U.ain_s1 ;
assign \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_4_U.u2.b  = \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_4_U.bin_s1 ;
assign \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_4_U.u2.cin  = \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_4_U.carry_s1 ;
assign \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_4_U.facout_s2  = \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_4_U.u2.cout ;
assign \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_4_U.fas_s2  = \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_4_U.u2.s ;
assign \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_4_U.u1.a  = \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_4_U.a [0];
assign \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_4_U.u1.b  = \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_4_U.b [0];
assign \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_4_U.u1.cin  = 1'h0;
assign \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_4_U.facout_s1  = \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_4_U.u1.cout ;
assign \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_4_U.fas_s1  = \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_4_U.u1.s ;
assign \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_4_U.a  = \add_2ns_2ns_2_2_1_U19.din0 ;
assign \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_4_U.b  = \add_2ns_2ns_2_2_1_U19.din1 ;
assign \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_4_U.ce  = \add_2ns_2ns_2_2_1_U19.ce ;
assign \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_4_U.clk  = \add_2ns_2ns_2_2_1_U19.clk ;
assign \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_4_U.reset  = \add_2ns_2ns_2_2_1_U19.reset ;
assign \add_2ns_2ns_2_2_1_U19.dout  = \add_2ns_2ns_2_2_1_U19.top_add_2ns_2ns_2_2_1_Adder_4_U.s ;
assign \add_2ns_2ns_2_2_1_U19.ce  = 1'h1;
assign \add_2ns_2ns_2_2_1_U19.clk  = ap_clk;
assign \add_2ns_2ns_2_2_1_U19.din0  = trunc_ln1_reg_2082;
assign \add_2ns_2ns_2_2_1_U19.din1  = { 1'h0, and_ln410_reg_2138 };
assign grp_fu_1323_p2 = \add_2ns_2ns_2_2_1_U19.dout ;
assign \add_2ns_2ns_2_2_1_U19.reset  = ap_rst;
assign \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_4_U.ain_s0  = \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_4_U.a ;
assign \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_4_U.bin_s0  = \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_4_U.b ;
assign \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_4_U.s  = { \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_4_U.fas_s2 , \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_4_U.sum_s1  };
assign \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_4_U.u2.a  = \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_4_U.ain_s1 ;
assign \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_4_U.u2.b  = \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_4_U.bin_s1 ;
assign \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_4_U.u2.cin  = \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_4_U.carry_s1 ;
assign \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_4_U.facout_s2  = \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_4_U.u2.cout ;
assign \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_4_U.fas_s2  = \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_4_U.u2.s ;
assign \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_4_U.u1.a  = \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_4_U.a [0];
assign \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_4_U.u1.b  = \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_4_U.b [0];
assign \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_4_U.u1.cin  = 1'h0;
assign \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_4_U.facout_s1  = \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_4_U.u1.cout ;
assign \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_4_U.fas_s1  = \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_4_U.u1.s ;
assign \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_4_U.a  = \add_2ns_2ns_2_2_1_U13.din0 ;
assign \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_4_U.b  = \add_2ns_2ns_2_2_1_U13.din1 ;
assign \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_4_U.ce  = \add_2ns_2ns_2_2_1_U13.ce ;
assign \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_4_U.clk  = \add_2ns_2ns_2_2_1_U13.clk ;
assign \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_4_U.reset  = \add_2ns_2ns_2_2_1_U13.reset ;
assign \add_2ns_2ns_2_2_1_U13.dout  = \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_4_U.s ;
assign \add_2ns_2ns_2_2_1_U13.ce  = 1'h1;
assign \add_2ns_2ns_2_2_1_U13.clk  = ap_clk;
assign \add_2ns_2ns_2_2_1_U13.din0  = ret_V_3_cast_reg_1984;
assign \add_2ns_2ns_2_2_1_U13.din1  = 2'h1;
assign grp_fu_1050_p2 = \add_2ns_2ns_2_2_1_U13.dout ;
assign \add_2ns_2ns_2_2_1_U13.reset  = ap_rst;
assign \add_26s_26ns_26_2_1_U9.top_add_26s_26ns_26_2_1_Adder_5_U.ain_s0  = \add_26s_26ns_26_2_1_U9.top_add_26s_26ns_26_2_1_Adder_5_U.a ;
assign \add_26s_26ns_26_2_1_U9.top_add_26s_26ns_26_2_1_Adder_5_U.bin_s0  = \add_26s_26ns_26_2_1_U9.top_add_26s_26ns_26_2_1_Adder_5_U.b ;
assign \add_26s_26ns_26_2_1_U9.top_add_26s_26ns_26_2_1_Adder_5_U.s  = { \add_26s_26ns_26_2_1_U9.top_add_26s_26ns_26_2_1_Adder_5_U.fas_s2 , \add_26s_26ns_26_2_1_U9.top_add_26s_26ns_26_2_1_Adder_5_U.sum_s1  };
assign \add_26s_26ns_26_2_1_U9.top_add_26s_26ns_26_2_1_Adder_5_U.u2.a  = \add_26s_26ns_26_2_1_U9.top_add_26s_26ns_26_2_1_Adder_5_U.ain_s1 ;
assign \add_26s_26ns_26_2_1_U9.top_add_26s_26ns_26_2_1_Adder_5_U.u2.b  = \add_26s_26ns_26_2_1_U9.top_add_26s_26ns_26_2_1_Adder_5_U.bin_s1 ;
assign \add_26s_26ns_26_2_1_U9.top_add_26s_26ns_26_2_1_Adder_5_U.u2.cin  = \add_26s_26ns_26_2_1_U9.top_add_26s_26ns_26_2_1_Adder_5_U.carry_s1 ;
assign \add_26s_26ns_26_2_1_U9.top_add_26s_26ns_26_2_1_Adder_5_U.facout_s2  = \add_26s_26ns_26_2_1_U9.top_add_26s_26ns_26_2_1_Adder_5_U.u2.cout ;
assign \add_26s_26ns_26_2_1_U9.top_add_26s_26ns_26_2_1_Adder_5_U.fas_s2  = \add_26s_26ns_26_2_1_U9.top_add_26s_26ns_26_2_1_Adder_5_U.u2.s ;
assign \add_26s_26ns_26_2_1_U9.top_add_26s_26ns_26_2_1_Adder_5_U.u1.a  = \add_26s_26ns_26_2_1_U9.top_add_26s_26ns_26_2_1_Adder_5_U.a [12:0];
assign \add_26s_26ns_26_2_1_U9.top_add_26s_26ns_26_2_1_Adder_5_U.u1.b  = \add_26s_26ns_26_2_1_U9.top_add_26s_26ns_26_2_1_Adder_5_U.b [12:0];
assign \add_26s_26ns_26_2_1_U9.top_add_26s_26ns_26_2_1_Adder_5_U.u1.cin  = 1'h0;
assign \add_26s_26ns_26_2_1_U9.top_add_26s_26ns_26_2_1_Adder_5_U.facout_s1  = \add_26s_26ns_26_2_1_U9.top_add_26s_26ns_26_2_1_Adder_5_U.u1.cout ;
assign \add_26s_26ns_26_2_1_U9.top_add_26s_26ns_26_2_1_Adder_5_U.fas_s1  = \add_26s_26ns_26_2_1_U9.top_add_26s_26ns_26_2_1_Adder_5_U.u1.s ;
assign \add_26s_26ns_26_2_1_U9.top_add_26s_26ns_26_2_1_Adder_5_U.a  = \add_26s_26ns_26_2_1_U9.din0 ;
assign \add_26s_26ns_26_2_1_U9.top_add_26s_26ns_26_2_1_Adder_5_U.b  = \add_26s_26ns_26_2_1_U9.din1 ;
assign \add_26s_26ns_26_2_1_U9.top_add_26s_26ns_26_2_1_Adder_5_U.ce  = \add_26s_26ns_26_2_1_U9.ce ;
assign \add_26s_26ns_26_2_1_U9.top_add_26s_26ns_26_2_1_Adder_5_U.clk  = \add_26s_26ns_26_2_1_U9.clk ;
assign \add_26s_26ns_26_2_1_U9.top_add_26s_26ns_26_2_1_Adder_5_U.reset  = \add_26s_26ns_26_2_1_U9.reset ;
assign \add_26s_26ns_26_2_1_U9.dout  = \add_26s_26ns_26_2_1_U9.top_add_26s_26ns_26_2_1_Adder_5_U.s ;
assign \add_26s_26ns_26_2_1_U9.ce  = 1'h1;
assign \add_26s_26ns_26_2_1_U9.clk  = ap_clk;
assign \add_26s_26ns_26_2_1_U9.din0  = { tmp_1_reg_1858[4], tmp_1_reg_1858, 20'h00000 };
assign \add_26s_26ns_26_2_1_U9.din1  = { 4'h0, ret_V_5_reg_1779, 15'h0000 };
assign grp_fu_810_p2 = \add_26s_26ns_26_2_1_U9.dout ;
assign \add_26s_26ns_26_2_1_U9.reset  = ap_rst;
endmodule


// Machine B:
// Processed by function `add_clk_enable_signal` in `verilog_tricks.py`.
// Processed by function `remove_reset_signal` in `verilog_tricks.py`.
module top_B (
  ap_clk,
  ap_start,
  ap_done,
  ap_idle,
  ap_ready,
  op_0,
  op_1,
  op_4,
  op_5,
  op_6,
  op_11,
  op_18,
  op_27,
  op_27_ap_vld,
clk_enable
);
input clk_enable;


input ap_clk;
wire ap_rst;
assign ap_rst = op_27_ap_vld;
input ap_start;
input [7:0] op_0;
input [15:0] op_1;
input [1:0] op_11;
input [1:0] op_18;
input [7:0] op_4;
input [3:0] op_5;
input [1:0] op_6;
output ap_done;
output ap_idle;
output ap_ready;
output [31:0] op_27;
output op_27_ap_vld;


reg [31:0] add_ln691_1_reg_1821;
reg [6:0] add_ln691_reg_1795;
reg [9:0] ap_CS_fsm = 10'h001;
reg icmp_ln786_1_reg_1708;
reg icmp_ln786_reg_1703;
reg icmp_ln790_reg_1713;
reg icmp_ln851_3_reg_1751;
reg icmp_ln851_4_reg_1859;
reg [1:0] op_14_V_reg_1805;
reg [1:0] op_17_V_reg_1864;
reg [3:0] op_19_V_reg_1763;
reg [31:0] op_26_V_reg_1881;
reg or_ln384_1_reg_1779;
reg overflow_1_reg_1774;
reg overflow_reg_1697;
reg p_Result_23_reg_1692;
reg p_Result_24_reg_1826;
reg p_Result_26_reg_1841;
reg [1:0] p_Val2_4_reg_1836;
reg [1:0] p_Val2_9_reg_1769;
reg [31:0] ret_V_19_cast_reg_1815;
reg [1:0] ret_V_19_reg_1800;
reg [3:0] ret_V_21_reg_1718;
reg [31:0] ret_V_22_cast_reg_1852;
reg [33:0] ret_V_23_reg_1810;
reg [31:0] ret_V_25_cast_reg_1874;
reg [33:0] ret_V_26_reg_1869;
reg [31:0] ret_V_28_cast_reg_1891;
reg [33:0] ret_V_28_reg_1886;
reg [7:0] ret_V_2_reg_1669;
reg [6:0] ret_V_5_reg_1731;
reg [1:0] ret_reg_1736;
reg rhs_1_reg_1680;
reg [31:0] select_ln1497_reg_1687;
reg [6:0] sext_ln850_reg_1789;
reg [8:0] sub_ln1497_reg_1675;
reg [4:0] tmp_1_reg_1746;
reg trunc_ln1195_reg_1741;
reg ush_reg_1724;
reg xor_ln410_reg_1831;
reg [5:0] _161_;
reg [35:0] _170_;
wire [31:0] _000_;
wire [6:0] _001_;
wire [9:0] _002_;
wire _003_;
wire _004_;
wire _005_;
wire _006_;
wire _007_;
wire [1:0] _008_;
wire [1:0] _009_;
wire [3:0] _010_;
wire [31:0] _011_;
wire _012_;
wire _013_;
wire _014_;
wire _015_;
wire _016_;
wire _017_;
wire [1:0] _018_;
wire [1:0] _019_;
wire [31:0] _020_;
wire [1:0] _021_;
wire [3:0] _022_;
wire [31:0] _023_;
wire [5:0] _024_;
wire [33:0] _025_;
wire [31:0] _026_;
wire [35:0] _027_;
wire [33:0] _028_;
wire [31:0] _029_;
wire [33:0] _030_;
wire [7:0] _031_;
wire [1:0] _032_;
wire [1:0] _033_;
wire _034_;
wire [31:0] _035_;
wire [6:0] _036_;
wire [8:0] _037_;
wire [4:0] _038_;
wire _039_;
wire _040_;
wire _041_;
wire [1:0] _042_;
wire _043_;
wire _044_;
wire _045_;
wire _046_;
wire _047_;
wire _048_;
wire _049_;
wire _050_;
wire _051_;
wire _052_;
wire _053_;
wire _054_;
wire _055_;
wire _056_;
wire _057_;
wire _058_;
wire _059_;
wire _060_;
wire _061_;
wire _062_;
wire _063_;
wire _064_;
wire _065_;
wire _066_;
wire _067_;
wire _068_;
wire _069_;
wire _070_;
wire _071_;
wire Range1_all_ones_fu_1014_p2;
wire Range1_all_zeros_fu_1020_p2;
wire [3:0] Range2_all_ones_fu_896_p1;
wire Range2_all_ones_fu_896_p3;
wire [31:0] add_ln691_1_fu_1300_p2;
wire [31:0] add_ln691_2_fu_1510_p2;
wire [31:0] add_ln691_3_fu_1570_p2;
wire [31:0] add_ln691_4_fu_1639_p2;
wire [6:0] add_ln691_fu_1167_p2;
wire and_ln340_fu_838_p2;
wire and_ln410_fu_1356_p2;
wire and_ln412_fu_962_p2;
wire and_ln414_1_fu_782_p2;
wire [1:0] and_ln414_fu_754_p2;
wire and_ln780_fu_1048_p2;
wire and_ln781_fu_1062_p2;
wire [3:0] and_ln783_fu_810_p2;
wire and_ln788_1_fu_1102_p2;
wire and_ln788_fu_1096_p2;
wire [7:0] and_ln_fu_373_p3;
wire ap_CS_fsm_state1;
wire ap_CS_fsm_state10;
wire ap_CS_fsm_state2;
wire ap_CS_fsm_state3;
wire ap_CS_fsm_state4;
wire ap_CS_fsm_state5;
wire ap_CS_fsm_state6;
wire ap_CS_fsm_state7;
wire ap_CS_fsm_state8;
wire ap_CS_fsm_state9;
wire [9:0] ap_NS_fsm;
wire ap_clk;
wire ap_done;
wire ap_idle;
wire ap_ready;
wire ap_rst;
wire ap_start;
wire [31:0] ashr_ln1497_fu_334_p2;
wire carry_1_fu_992_p2;
wire [7:0] conv_i847_fu_331_p0;
wire [31:0] conv_i847_fu_331_p1;
wire deleted_ones_fu_1054_p3;
wire deleted_zeros_fu_1026_p3;
wire icmp_ln414_fu_776_p2;
wire icmp_ln785_fu_401_p2;
wire icmp_ln786_1_fu_425_p2;
wire icmp_ln786_fu_419_p2;
wire icmp_ln790_fu_443_p2;
wire icmp_ln851_1_fu_1208_p2;
wire icmp_ln851_2_fu_487_p2;
wire icmp_ln851_3_fu_691_p2;
wire icmp_ln851_4_fu_1480_p2;
wire icmp_ln851_fu_269_p2;
wire [3:0] \mul_4s_2s_6_1_1_U1.din0 ;
wire [1:0] \mul_4s_2s_6_1_1_U1.din1 ;
wire [5:0] \mul_4s_2s_6_1_1_U1.dout ;
wire [3:0] \mul_4s_2s_6_1_1_U1.top_mul_4s_2s_6_1_1_Multiplier_0_U.a ;
wire [1:0] \mul_4s_2s_6_1_1_U1.top_mul_4s_2s_6_1_1_Multiplier_0_U.b ;
wire [5:0] \mul_4s_2s_6_1_1_U1.top_mul_4s_2s_6_1_1_Multiplier_0_U.p ;
wire neg_src_2_fu_1486_p2;
wire neg_src_4_fu_816_p3;
wire [7:0] op_0;
wire [15:0] op_1;
wire [1:0] op_11;
wire [3:0] op_12_V_fu_638_p2;
wire [21:0] op_13_V_fu_697_p3;
wire [1:0] op_14_V_fu_1243_p3;
wire [7:0] op_16_V_fu_1396_p3;
wire [1:0] op_17_V_fu_1496_p3;
wire [1:0] op_18;
wire [3:0] op_19_V_fu_864_p3;
wire [31:0] op_23_V_fu_1430_p2;
wire [31:0] op_26_V_fu_1593_p2;
wire [31:0] op_27;
wire op_27_ap_vld;
wire [7:0] op_2_V_fu_552_p3;
wire [7:0] op_4;
wire [3:0] op_5;
wire [1:0] op_6;
wire [2:0] op_8_V_fu_613_p3;
wire [3:0] or_ln1195_1_fu_904_p1;
wire [3:0] or_ln1195_1_fu_904_p2;
wire [4:0] or_ln1195_fu_890_p2;
wire or_ln384_1_fu_1126_p2;
wire or_ln384_fu_547_p2;
wire or_ln410_fu_1350_p2;
wire or_ln412_fu_956_p2;
wire or_ln785_fu_1074_p2;
wire or_ln788_1_fu_530_p2;
wire or_ln788_2_fu_1108_p2;
wire or_ln788_fu_526_p2;
wire [7:0] or_ln_fu_391_p4;
wire overflow_1_fu_1086_p2;
wire overflow_fu_413_p2;
wire [3:0] p_Result_12_fu_854_p4;
wire p_Result_16_fu_928_p3;
wire p_Result_18_fu_1249_p3;
wire p_Result_19_fu_1404_p3;
wire [3:0] p_Result_1_fu_1472_p3;
wire p_Result_20_fu_1503_p3;
wire p_Result_21_fu_1560_p3;
wire p_Result_22_fu_1629_p3;
wire p_Result_23_fu_357_p3;
wire p_Result_24_fu_1314_p3;
wire p_Result_25_fu_1332_p3;
wire p_Result_27_fu_728_p3;
wire p_Result_28_fu_802_p3;
wire [3:0] p_Result_29_fu_910_p1;
wire p_Result_29_fu_910_p3;
wire p_Result_2_fu_1196_p3;
wire [3:0] p_Result_30_fu_936_p1;
wire p_Result_30_fu_936_p3;
wire p_Result_31_fu_948_p3;
wire p_Result_32_fu_978_p3;
wire [19:0] p_Result_3_fu_683_p3;
wire p_Result_4_fu_475_p3;
wire [6:0] p_Result_5_fu_435_p3;
wire [4:0] p_Result_s_22_fu_381_p4;
wire p_Result_s_fu_257_p3;
wire [6:0] p_Val2_11_fu_663_p2;
wire [1:0] p_Val2_4_fu_1366_p2;
wire [2:0] p_Val2_6_fu_792_p2;
wire [2:0] p_Val2_7_fu_844_p2;
wire [1:0] p_Val2_8_fu_918_p4;
wire [1:0] p_Val2_9_fu_972_p2;
wire [7:0] p_Val2_s_fu_518_p3;
wire r_1_fu_944_p1;
wire [3:0] r_V_1_fu_1309_p0;
wire [3:0] r_V_1_fu_1309_p2;
wire [3:0] r_V_2_fu_722_p1;
wire [3:0] r_V_2_fu_722_p2;
wire [5:0] r_V_fu_1180_p2;
wire r_fu_1340_p1;
wire [31:0] ret_V_19_cast_fu_1290_p4;
wire [1:0] ret_V_19_fu_1228_p3;
wire [7:0] ret_V_1_fu_275_p2;
wire [15:0] ret_V_20_fu_460_p2;
wire [3:0] ret_V_21_fu_507_p3;
wire [25:0] ret_V_22_fu_1147_p2;
wire [25:0] ret_V_22_reg_1784;
wire [33:0] ret_V_23_fu_1284_p2;
wire [31:0] ret_V_24_fu_1420_p3;
wire [36:0] ret_V_25_fu_1452_p2;
wire [36:0] ret_V_25_reg_1847;
wire [33:0] ret_V_26_fu_1544_p2;
wire [31:0] ret_V_27_fu_1582_p3;
wire [33:0] ret_V_28_fu_1613_p2;
wire [7:0] ret_V_2_fu_289_p3;
wire [1:0] ret_V_3_cast_fu_1186_p4;
wire [1:0] ret_V_3_fu_1214_p2;
wire [6:0] ret_V_5_fu_590_p2;
wire [3:0] ret_V_7_fu_493_p2;
wire [3:0] ret_V_8_cast_fu_465_p4;
wire [6:0] ret_V_9_fu_1390_p2;
wire [7:0] ret_V_fu_247_p4;
wire [1:0] ret_fu_628_p2;
wire [35:0] rhs_10_fu_1440_p3;
wire [32:0] rhs_11_fu_1532_p3;
wire [32:0] rhs_13_fu_1602_p3;
wire rhs_1_fu_315_p2;
wire [8:0] rhs_2_fu_449_p3;
wire [6:0] rhs_4_fu_1383_p3;
wire [4:0] rhs_5_fu_872_p3;
wire [5:0] rhs_7_fu_651_p3;
wire [24:0] rhs_8_fu_1136_p3;
wire [6:0] rhs_fu_582_p3;
wire [1:0] select_ln1118_1_fu_715_p3;
wire [3:0] select_ln1118_fu_704_p3;
wire [1:0] select_ln1345_fu_621_p3;
wire [31:0] select_ln1497_fu_349_p3;
wire select_ln340_2_fu_830_p3;
wire select_ln340_fu_1490_p3;
wire [31:0] select_ln353_2_fu_1525_p3;
wire [6:0] select_ln353_fu_1265_p3;
wire [7:0] select_ln384_1_fu_540_p3;
wire [1:0] select_ln384_fu_1236_p3;
wire [1:0] select_ln850_1_fu_1220_p3;
wire [3:0] select_ln850_2_fu_499_p3;
wire [31:0] select_ln850_4_fu_1414_p3;
wire [6:0] select_ln850_5_fu_1260_p3;
wire [31:0] select_ln850_6_fu_1575_p3;
wire [31:0] select_ln850_7_fu_1644_p3;
wire [31:0] select_ln850_8_fu_1519_p3;
wire [7:0] select_ln850_fu_281_p3;
wire [25:0] sext_ln1192_1_fu_1143_p1;
wire [33:0] sext_ln1192_2_fu_1280_p1;
wire [36:0] sext_ln1192_3_fu_1448_p1;
wire [33:0] sext_ln1192_4_fu_1540_p1;
wire [33:0] sext_ln1192_5_fu_1609_p1;
wire [6:0] sext_ln1192_fu_659_p1;
wire [3:0] sext_ln1193_fu_1380_p0;
wire [6:0] sext_ln1193_fu_1380_p1;
wire [3:0] sext_ln1195_fu_886_p0;
wire [4:0] sext_ln1195_fu_886_p1;
wire [31:0] sext_ln1497_1_fu_340_p1;
wire [8:0] sext_ln1497_fu_297_p1;
wire [3:0] sext_ln367_fu_850_p1;
wire [31:0] sext_ln545_fu_321_p1;
wire [31:0] sext_ln69_1_fu_1589_p1;
wire [31:0] sext_ln69_fu_1427_p1;
wire [36:0] sext_ln703_1_fu_1436_p1;
wire [33:0] sext_ln703_2_fu_1515_p1;
wire [33:0] sext_ln703_3_fu_1599_p1;
wire [33:0] sext_ln703_fu_1256_p1;
wire [2:0] sext_ln713_fu_746_p1;
wire [12:0] sext_ln727_fu_564_p1;
wire [3:0] sext_ln745_fu_798_p1;
wire [6:0] sext_ln850_fu_1163_p1;
wire [31:0] shl_ln1497_fu_343_p2;
wire [12:0] shl_ln728_1_fu_568_p3;
wire [5:0] shl_ln728_5_fu_596_p3;
wire [7:0] shl_ln_fu_307_p1;
wire [15:0] shl_ln_fu_307_p3;
wire signbit_fu_607_p2;
wire [8:0] sub_ln1497_fu_301_p2;
wire tmp_13_fu_760_p3;
wire tmp_23_fu_998_p3;
wire tmp_24_fu_1034_p3;
wire [7:0] tmp_26_fu_1272_p3;
wire [1:0] tmp_3_fu_768_p3;
wire tmp_4_fu_365_p3;
wire [1:0] tmp_9_fu_1006_p3;
wire tmp_fu_324_p3;
wire [5:0] tmp_s_fu_1153_p4;
wire [3:0] trunc_ln1118_fu_711_p0;
wire [1:0] trunc_ln1118_fu_711_p1;
wire [3:0] trunc_ln1195_1_fu_879_p3;
wire trunc_ln1195_fu_643_p1;
wire [3:0] trunc_ln1349_fu_634_p1;
wire [1:0] trunc_ln1_fu_1322_p4;
wire [1:0] trunc_ln708_1_fu_736_p4;
wire trunc_ln718_fu_750_p1;
wire [2:0] trunc_ln731_fu_515_p1;
wire trunc_ln790_1_fu_1092_p1;
wire [1:0] trunc_ln790_fu_431_p1;
wire [2:0] trunc_ln851_1_fu_1204_p1;
wire [7:0] trunc_ln851_2_fu_483_p1;
wire [4:0] trunc_ln851_3_fu_679_p1;
wire trunc_ln851_4_fu_1411_p1;
wire [2:0] trunc_ln851_5_fu_1468_p1;
wire trunc_ln851_6_fu_1567_p1;
wire trunc_ln851_7_fu_1636_p1;
wire [7:0] trunc_ln851_fu_265_p1;
wire [6:0] trunc_ln8_fu_560_p1;
wire underflow_1_fu_1120_p2;
wire underflow_fu_535_p2;
wire ush_fu_576_p2;
wire xor_ln410_fu_1344_p2;
wire xor_ln416_fu_986_p2;
wire xor_ln780_fu_1042_p2;
wire xor_ln785_1_fu_824_p2;
wire xor_ln785_2_fu_1068_p2;
wire xor_ln785_3_fu_1080_p2;
wire xor_ln785_fu_407_p2;
wire xor_ln788_fu_1114_p2;
wire [25:0] zext_ln1192_fu_1132_p1;
wire [15:0] zext_ln1196_fu_456_p1;
wire [3:0] zext_ln1380_fu_1306_p1;
wire [7:0] zext_ln1499_fu_603_p1;
wire [2:0] zext_ln415_1_fu_788_p1;
wire [1:0] zext_ln415_2_fu_968_p1;
wire [1:0] zext_ln415_fu_1362_p1;
wire [6:0] zext_ln703_fu_647_p1;


assign add_ln691_1_fu_1300_p2 = { ret_V_23_fu_1284_p2[33], ret_V_23_fu_1284_p2[33], ret_V_23_fu_1284_p2[33], ret_V_23_fu_1284_p2[33], ret_V_23_fu_1284_p2[33], ret_V_23_fu_1284_p2[33], ret_V_23_fu_1284_p2[33], ret_V_23_fu_1284_p2[33], ret_V_23_fu_1284_p2[33], ret_V_23_fu_1284_p2[33], ret_V_23_fu_1284_p2[33], ret_V_23_fu_1284_p2[33], ret_V_23_fu_1284_p2[33], ret_V_23_fu_1284_p2[33], ret_V_23_fu_1284_p2[33], ret_V_23_fu_1284_p2[33], ret_V_23_fu_1284_p2[33], ret_V_23_fu_1284_p2[33], ret_V_23_fu_1284_p2[33], ret_V_23_fu_1284_p2[33], ret_V_23_fu_1284_p2[33], ret_V_23_fu_1284_p2[33], ret_V_23_fu_1284_p2[33], ret_V_23_fu_1284_p2[33], ret_V_23_fu_1284_p2[33], ret_V_23_fu_1284_p2[7:1] } + 1'h1;
assign add_ln691_2_fu_1510_p2 = ret_V_22_cast_reg_1852 + 1'h1;
assign add_ln691_3_fu_1570_p2 = ret_V_25_cast_reg_1874 + 1'h1;
assign add_ln691_4_fu_1639_p2 = ret_V_28_cast_reg_1891 + 1'h1;
assign add_ln691_fu_1167_p2 = $signed(ret_V_22_fu_1147_p2[25:20]) + $signed(2'h1);
assign op_23_V_fu_1430_p2 = $signed(ret_V_24_fu_1420_p3) + $signed(ret_V_19_reg_1800);
assign op_26_V_fu_1593_p2 = $signed(ret_V_27_fu_1582_p3) + $signed(op_18);
assign p_Val2_11_fu_663_p2 = $signed({ op_12_V_fu_638_p2, 2'h0 }) + $signed({ 1'h0, signbit_fu_607_p2, 2'h0 });
assign p_Val2_4_fu_1366_p2 = r_V_1_fu_1309_p2[3:2] + and_ln410_fu_1356_p2;
assign p_Val2_6_fu_792_p2 = $signed(r_V_2_fu_722_p2[3:2]) + $signed({ 1'h0, and_ln414_1_fu_782_p2 });
assign p_Val2_9_fu_972_p2 = or_ln1195_1_fu_904_p2[3:2] + and_ln412_fu_962_p2;
assign ret_V_1_fu_275_p2 = op_1[15:8] + 1'h1;
assign ret_V_22_fu_1147_p2 = $signed({ tmp_1_reg_1746, 20'h00000 }) + $signed({ 1'h0, ret_V_5_reg_1731, 15'h0000 });
assign { ret_V_23_fu_1284_p2[33], ret_V_23_fu_1284_p2[7:0] } = $signed({ select_ln353_fu_1265_p3, 1'h0 }) + $signed(op_14_V_fu_1243_p3);
assign ret_V_25_fu_1452_p2 = $signed({ op_23_V_fu_1430_p2, 4'h0 }) + $signed({ ret_V_9_fu_1390_p2, 1'h0 });
assign ret_V_26_fu_1544_p2 = $signed({ select_ln353_2_fu_1525_p3, 1'h0 }) + $signed(op_17_V_fu_1496_p3);
assign ret_V_28_fu_1613_p2 = $signed({ op_26_V_reg_1881, 1'h0 }) + $signed(op_19_V_reg_1763);
assign ret_V_3_fu_1214_p2 = r_V_fu_1180_p2[4:3] + 1'h1;
assign ret_V_7_fu_493_p2 = ret_V_20_fu_460_p2[11:8] + 1'h1;
assign underflow_1_fu_1120_p2 = xor_ln788_fu_1114_p2 & op_5[3];
assign underflow_fu_535_p2 = p_Result_23_reg_1692 & or_ln788_1_fu_530_p2;
assign _043_ = icmp_ln851_3_reg_1751 & ap_CS_fsm[3];
assign _044_ = ap_CS_fsm[0] & _047_;
assign _045_ = ap_CS_fsm[0] & ap_start;
assign and_ln340_fu_838_p2 = select_ln340_2_fu_830_p3 & p_Val2_6_fu_792_p2[2];
assign and_ln410_fu_1356_p2 = r_V_1_fu_1309_p2[1] & or_ln410_fu_1350_p2;
assign and_ln412_fu_962_p2 = op_5[1] & or_ln412_fu_956_p2;
assign and_ln414_1_fu_782_p2 = r_V_2_fu_722_p2[3] & icmp_ln414_fu_776_p2;
assign and_ln414_fu_754_p2 = op_5[1:0] & select_ln1118_1_fu_715_p3;
assign and_ln780_fu_1048_p2 = xor_ln780_fu_1042_p2 & op_5[3];
assign and_ln781_fu_1062_p2 = carry_1_fu_992_p2 & Range1_all_ones_fu_1014_p2;
assign and_ln783_fu_810_p2 = { p_Val2_6_fu_792_p2[2], p_Val2_6_fu_792_p2 } & r_V_2_fu_722_p2;
assign and_ln788_1_fu_1102_p2 = p_Val2_9_fu_972_p2[1] & and_ln788_fu_1096_p2;
assign and_ln788_fu_1096_p2 = p_Val2_9_fu_972_p2[0] & deleted_ones_fu_1054_p3;
assign carry_1_fu_992_p2 = xor_ln416_fu_986_p2 & or_ln1195_1_fu_904_p2[3];
assign neg_src_2_fu_1486_p2 = p_Result_26_reg_1841 & p_Result_24_reg_1826;
assign overflow_1_fu_1086_p2 = xor_ln785_3_fu_1080_p2 & or_ln785_fu_1074_p2;
assign overflow_fu_413_p2 = xor_ln785_fu_407_p2 & icmp_ln785_fu_401_p2;
assign r_V_2_fu_722_p2 = select_ln1118_fu_704_p3 & op_5;
assign ret_V_5_fu_590_p2 = op_2_V_fu_552_p3[6:0] & { op_6, 5'h00 };
assign ret_fu_628_p2 = select_ln1345_fu_621_p3 & op_6;
assign xor_ln785_1_fu_824_p2 = ~ r_V_2_fu_722_p2[3];
assign xor_ln410_fu_1344_p2 = ~ r_V_1_fu_1309_p2[3];
assign xor_ln780_fu_1042_p2 = ~ or_ln1195_fu_890_p2[4];
assign xor_ln416_fu_986_p2 = ~ p_Val2_9_fu_972_p2[1];
assign xor_ln785_2_fu_1068_p2 = ~ deleted_zeros_fu_1026_p3;
assign xor_ln785_3_fu_1080_p2 = ~ op_5[3];
assign xor_ln788_fu_1114_p2 = ~ or_ln788_2_fu_1108_p2;
assign xor_ln785_fu_407_p2 = ~ select_ln1497_fu_349_p3[7];
assign p_Val2_7_fu_844_p2 = ~ p_Val2_6_fu_792_p2;
assign _046_ = { op_2_V_fu_552_p3[7], op_2_V_fu_552_p3[7], op_2_V_fu_552_p3[7], op_2_V_fu_552_p3[7], op_2_V_fu_552_p3[7], op_2_V_fu_552_p3 } == { op_4, 5'h00 };
assign _047_ = ~ ap_start;
assign _048_ = { op_5[3], or_ln1195_fu_890_p2[4] } == 2'h3;
assign _049_ = ! { op_5[3], or_ln1195_fu_890_p2[4] };
assign _050_ = ! { select_ln1497_fu_349_p3[2], 7'h00 };
assign _051_ = ! { select_ln1497_fu_349_p3[1:0], 5'h00 };
assign _052_ = ! r_V_fu_1180_p2[2:0];
assign _053_ = ! ret_V_20_fu_460_p2[7:0];
assign _054_ = ! op_1[7:0];
assign \mul_4s_2s_6_1_1_U1.top_mul_4s_2s_6_1_1_Multiplier_0_U.p  = $signed(\mul_4s_2s_6_1_1_U1.top_mul_4s_2s_6_1_1_Multiplier_0_U.a ) * $signed(\mul_4s_2s_6_1_1_U1.top_mul_4s_2s_6_1_1_Multiplier_0_U.b );
assign _055_ = | { and_ln414_fu_754_p2[1], r_V_2_fu_722_p2[0] };
assign _056_ = | { select_ln1497_fu_349_p3[2], 2'h0, select_ln1497_fu_349_p3[7:3] };
assign _057_ = select_ln1497_fu_349_p3[7:3] != 5'h1f;
assign _058_ = | { ret_V_5_fu_590_p2[4:0], 15'h0000 };
assign _059_ = | { ret_V_9_fu_1390_p2[2:0], 1'h0 };
assign _060_ = { op_0, 8'h00 } != op_1;
assign _061_ = op_2_V_fu_552_p3 != { rhs_1_reg_1680, 5'h00 };
assign op_12_V_fu_638_p2 = op_4[3:0] | ret_V_21_reg_1718;
assign or_ln1195_1_fu_904_p2 = { trunc_ln1195_reg_1741, 3'h0 } | op_5;
assign or_ln1195_fu_890_p2 = { op_5[3], op_5 } | { ret_reg_1736, 3'h0 };
assign or_ln384_1_fu_1126_p2 = underflow_1_fu_1120_p2 | overflow_1_fu_1086_p2;
assign or_ln384_fu_547_p2 = underflow_fu_535_p2 | overflow_reg_1697;
assign or_ln410_fu_1350_p2 = xor_ln410_fu_1344_p2 | r_V_1_fu_1309_p2[0];
assign or_ln412_fu_956_p2 = or_ln1195_fu_890_p2[0] | or_ln1195_1_fu_904_p2[2];
assign or_ln785_fu_1074_p2 = xor_ln785_2_fu_1068_p2 | p_Val2_9_fu_972_p2[1];
assign or_ln788_1_fu_530_p2 = or_ln788_fu_526_p2 | icmp_ln786_reg_1703;
assign or_ln788_2_fu_1108_p2 = and_ln788_1_fu_1102_p2 | and_ln781_fu_1062_p2;
assign or_ln788_fu_526_p2 = icmp_ln790_reg_1713 | icmp_ln786_1_reg_1708;
always @(posedge ap_clk)
ret_V_5_reg_1731[4:0] <= 5'h00;
always @(posedge ap_clk)
ret_V_2_reg_1669 <= _031_;
always @(posedge ap_clk)
sub_ln1497_reg_1675 <= _037_;
always @(posedge ap_clk)
rhs_1_reg_1680 <= _034_;
always @(posedge ap_clk)
ret_V_28_reg_1886 <= _030_;
always @(posedge ap_clk)
ret_V_28_cast_reg_1891 <= _029_;
always @(posedge ap_clk)
op_26_V_reg_1881 <= _011_;
always @(posedge ap_clk)
op_19_V_reg_1763 <= _010_;
always @(posedge ap_clk)
p_Val2_9_reg_1769 <= _019_;
always @(posedge ap_clk)
overflow_1_reg_1774 <= _013_;
always @(posedge ap_clk)
or_ln384_1_reg_1779 <= _012_;
always @(posedge ap_clk)
_161_ <= _024_;
assign ret_V_22_reg_1784[25:20] = _161_;
always @(posedge ap_clk)
sext_ln850_reg_1789 <= _036_;
always @(posedge ap_clk)
op_17_V_reg_1864 <= _009_;
always @(posedge ap_clk)
ret_V_26_reg_1869 <= _028_;
always @(posedge ap_clk)
ret_V_25_cast_reg_1874 <= _026_;
always @(posedge ap_clk)
p_Result_24_reg_1826 <= _016_;
always @(posedge ap_clk)
xor_ln410_reg_1831 <= _041_;
always @(posedge ap_clk)
p_Val2_4_reg_1836 <= _018_;
always @(posedge ap_clk)
p_Result_26_reg_1841 <= _017_;
always @(posedge ap_clk)
_170_ <= _027_;
assign ret_V_25_reg_1847[36:1] = _170_;
always @(posedge ap_clk)
ret_V_22_cast_reg_1852 <= _023_;
always @(posedge ap_clk)
icmp_ln851_4_reg_1859 <= _007_;
always @(posedge ap_clk)
ush_reg_1724 <= _040_;
always @(posedge ap_clk)
ret_V_5_reg_1731[6:5] <= _032_;
always @(posedge ap_clk)
ret_reg_1736 <= _033_;
always @(posedge ap_clk)
trunc_ln1195_reg_1741 <= _039_;
always @(posedge ap_clk)
tmp_1_reg_1746 <= _038_;
always @(posedge ap_clk)
icmp_ln851_3_reg_1751 <= _006_;
always @(posedge ap_clk)
select_ln1497_reg_1687 <= _035_;
always @(posedge ap_clk)
p_Result_23_reg_1692 <= _015_;
always @(posedge ap_clk)
overflow_reg_1697 <= _014_;
always @(posedge ap_clk)
icmp_ln786_reg_1703 <= _004_;
always @(posedge ap_clk)
icmp_ln786_1_reg_1708 <= _003_;
always @(posedge ap_clk)
icmp_ln790_reg_1713 <= _005_;
always @(posedge ap_clk)
ret_V_21_reg_1718 <= _022_;
always @(posedge ap_clk)
add_ln691_reg_1795 <= _001_;
always @(posedge ap_clk)
ret_V_19_reg_1800 <= _021_;
always @(posedge ap_clk)
op_14_V_reg_1805 <= _008_;
always @(posedge ap_clk)
ret_V_23_reg_1810 <= _025_;
always @(posedge ap_clk)
ret_V_19_cast_reg_1815 <= _020_;
always @(posedge ap_clk)
add_ln691_1_reg_1821 <= _000_;
always @(posedge ap_clk)
ap_CS_fsm <= _002_;
assign _042_ = _045_ ? 2'h2 : 2'h1;
assign _062_ = ap_CS_fsm == 1'h1;
function [9:0] _195_;
input [9:0] a;
input [99:0] b;
input [9:0] s;
case (s)
10'b0000000001:
_195_ = b[9:0];
10'b0000000010:
_195_ = b[19:10];
10'b0000000100:
_195_ = b[29:20];
10'b0000001000:
_195_ = b[39:30];
10'b0000010000:
_195_ = b[49:40];
10'b0000100000:
_195_ = b[59:50];
10'b0001000000:
_195_ = b[69:60];
10'b0010000000:
_195_ = b[79:70];
10'b0100000000:
_195_ = b[89:80];
10'b1000000000:
_195_ = b[99:90];
10'b0000000000:
_195_ = a;
default:
_195_ = 10'bx;
endcase
endfunction
assign ap_NS_fsm = _195_(10'hxxx, { 8'h00, _042_, 90'h00402010080402010080001 }, { _062_, _071_, _070_, _069_, _068_, _067_, _066_, _065_, _064_, _063_ });
assign _063_ = ap_CS_fsm == 10'h200;
assign _064_ = ap_CS_fsm == 9'h100;
assign _065_ = ap_CS_fsm == 8'h80;
assign _066_ = ap_CS_fsm == 7'h40;
assign _067_ = ap_CS_fsm == 6'h20;
assign _068_ = ap_CS_fsm == 5'h10;
assign _069_ = ap_CS_fsm == 4'h8;
assign _070_ = ap_CS_fsm == 3'h4;
assign _071_ = ap_CS_fsm == 2'h2;
assign op_27_ap_vld = ap_CS_fsm[9] ? 1'h1 : 1'h0;
assign ap_idle = _044_ ? 1'h1 : 1'h0;
assign _034_ = ap_CS_fsm[0] ? rhs_1_fu_315_p2 : rhs_1_reg_1680;
assign _037_ = ap_CS_fsm[0] ? sub_ln1497_fu_301_p2 : sub_ln1497_reg_1675;
assign _031_ = ap_CS_fsm[0] ? ret_V_2_fu_289_p3 : ret_V_2_reg_1669;
assign _029_ = ap_CS_fsm[8] ? ret_V_28_fu_1613_p2[32:1] : ret_V_28_cast_reg_1891;
assign _030_ = ap_CS_fsm[8] ? ret_V_28_fu_1613_p2 : ret_V_28_reg_1886;
assign _011_ = ap_CS_fsm[7] ? op_26_V_fu_1593_p2 : op_26_V_reg_1881;
assign _036_ = ap_CS_fsm[3] ? { ret_V_22_fu_1147_p2[25], ret_V_22_fu_1147_p2[25:20] } : sext_ln850_reg_1789;
assign _024_ = ap_CS_fsm[3] ? ret_V_22_fu_1147_p2[25:20] : ret_V_22_reg_1784[25:20];
assign _012_ = ap_CS_fsm[3] ? or_ln384_1_fu_1126_p2 : or_ln384_1_reg_1779;
assign _013_ = ap_CS_fsm[3] ? overflow_1_fu_1086_p2 : overflow_1_reg_1774;
assign _019_ = ap_CS_fsm[3] ? p_Val2_9_fu_972_p2 : p_Val2_9_reg_1769;
assign _010_ = ap_CS_fsm[3] ? op_19_V_fu_864_p3 : op_19_V_reg_1763;
assign _026_ = ap_CS_fsm[6] ? ret_V_26_fu_1544_p2[32:1] : ret_V_25_cast_reg_1874;
assign _028_ = ap_CS_fsm[6] ? ret_V_26_fu_1544_p2 : ret_V_26_reg_1869;
assign _009_ = ap_CS_fsm[6] ? op_17_V_fu_1496_p3 : op_17_V_reg_1864;
assign _007_ = ap_CS_fsm[5] ? icmp_ln851_4_fu_1480_p2 : icmp_ln851_4_reg_1859;
assign _023_ = ap_CS_fsm[5] ? ret_V_25_fu_1452_p2[35:4] : ret_V_22_cast_reg_1852;
assign _027_ = ap_CS_fsm[5] ? ret_V_25_fu_1452_p2[36:1] : ret_V_25_reg_1847[36:1];
assign _017_ = ap_CS_fsm[5] ? p_Val2_4_fu_1366_p2[1] : p_Result_26_reg_1841;
assign _018_ = ap_CS_fsm[5] ? p_Val2_4_fu_1366_p2 : p_Val2_4_reg_1836;
assign _041_ = ap_CS_fsm[5] ? xor_ln410_fu_1344_p2 : xor_ln410_reg_1831;
assign _016_ = ap_CS_fsm[5] ? r_V_1_fu_1309_p2[3] : p_Result_24_reg_1826;
assign _006_ = ap_CS_fsm[2] ? icmp_ln851_3_fu_691_p2 : icmp_ln851_3_reg_1751;
assign _038_ = ap_CS_fsm[2] ? p_Val2_11_fu_663_p2[6:2] : tmp_1_reg_1746;
assign _039_ = ap_CS_fsm[2] ? ret_fu_628_p2[0] : trunc_ln1195_reg_1741;
assign _033_ = ap_CS_fsm[2] ? ret_fu_628_p2 : ret_reg_1736;
assign _032_ = ap_CS_fsm[2] ? ret_V_5_fu_590_p2[6:5] : ret_V_5_reg_1731[6:5];
assign _040_ = ap_CS_fsm[2] ? ush_fu_576_p2 : ush_reg_1724;
assign _022_ = ap_CS_fsm[1] ? ret_V_21_fu_507_p3 : ret_V_21_reg_1718;
assign _005_ = ap_CS_fsm[1] ? icmp_ln790_fu_443_p2 : icmp_ln790_reg_1713;
assign _003_ = ap_CS_fsm[1] ? icmp_ln786_1_fu_425_p2 : icmp_ln786_1_reg_1708;
assign _004_ = ap_CS_fsm[1] ? icmp_ln786_fu_419_p2 : icmp_ln786_reg_1703;
assign _014_ = ap_CS_fsm[1] ? overflow_fu_413_p2 : overflow_reg_1697;
assign _015_ = ap_CS_fsm[1] ? select_ln1497_fu_349_p3[7] : p_Result_23_reg_1692;
assign _035_ = ap_CS_fsm[1] ? select_ln1497_fu_349_p3 : select_ln1497_reg_1687;
assign _001_ = _043_ ? add_ln691_fu_1167_p2 : add_ln691_reg_1795;
assign _000_ = ap_CS_fsm[4] ? add_ln691_1_fu_1300_p2 : add_ln691_1_reg_1821;
assign _020_ = ap_CS_fsm[4] ? { ret_V_23_fu_1284_p2[33], ret_V_23_fu_1284_p2[33], ret_V_23_fu_1284_p2[33], ret_V_23_fu_1284_p2[33], ret_V_23_fu_1284_p2[33], ret_V_23_fu_1284_p2[33], ret_V_23_fu_1284_p2[33], ret_V_23_fu_1284_p2[33], ret_V_23_fu_1284_p2[33], ret_V_23_fu_1284_p2[33], ret_V_23_fu_1284_p2[33], ret_V_23_fu_1284_p2[33], ret_V_23_fu_1284_p2[33], ret_V_23_fu_1284_p2[33], ret_V_23_fu_1284_p2[33], ret_V_23_fu_1284_p2[33], ret_V_23_fu_1284_p2[33], ret_V_23_fu_1284_p2[33], ret_V_23_fu_1284_p2[33], ret_V_23_fu_1284_p2[33], ret_V_23_fu_1284_p2[33], ret_V_23_fu_1284_p2[33], ret_V_23_fu_1284_p2[33], ret_V_23_fu_1284_p2[33], ret_V_23_fu_1284_p2[33], ret_V_23_fu_1284_p2[7:1] } : ret_V_19_cast_reg_1815;
assign _025_ = ap_CS_fsm[4] ? { ret_V_23_fu_1284_p2[33], ret_V_23_fu_1284_p2[33], ret_V_23_fu_1284_p2[33], ret_V_23_fu_1284_p2[33], ret_V_23_fu_1284_p2[33], ret_V_23_fu_1284_p2[33], ret_V_23_fu_1284_p2[33], ret_V_23_fu_1284_p2[33], ret_V_23_fu_1284_p2[33], ret_V_23_fu_1284_p2[33], ret_V_23_fu_1284_p2[33], ret_V_23_fu_1284_p2[33], ret_V_23_fu_1284_p2[33], ret_V_23_fu_1284_p2[33], ret_V_23_fu_1284_p2[33], ret_V_23_fu_1284_p2[33], ret_V_23_fu_1284_p2[33], ret_V_23_fu_1284_p2[33], ret_V_23_fu_1284_p2[33], ret_V_23_fu_1284_p2[33], ret_V_23_fu_1284_p2[33], ret_V_23_fu_1284_p2[33], ret_V_23_fu_1284_p2[33], ret_V_23_fu_1284_p2[33], ret_V_23_fu_1284_p2[33], ret_V_23_fu_1284_p2[33], ret_V_23_fu_1284_p2[7:0] } : ret_V_23_reg_1810;
assign _008_ = ap_CS_fsm[4] ? op_14_V_fu_1243_p3 : op_14_V_reg_1805;
assign _021_ = ap_CS_fsm[4] ? ret_V_19_fu_1228_p3 : ret_V_19_reg_1800;
assign _002_ = ap_rst ? 10'h001 : ap_NS_fsm;
assign r_V_1_fu_1309_p2 = $signed(op_5) << ush_reg_1724;
assign shl_ln1497_fu_343_p2 = $signed(op_0) << { sub_ln1497_reg_1675[8], sub_ln1497_reg_1675[8], sub_ln1497_reg_1675[8], sub_ln1497_reg_1675[8], sub_ln1497_reg_1675[8], sub_ln1497_reg_1675[8], sub_ln1497_reg_1675[8], sub_ln1497_reg_1675[8], sub_ln1497_reg_1675[8], sub_ln1497_reg_1675[8], sub_ln1497_reg_1675[8], sub_ln1497_reg_1675[8], sub_ln1497_reg_1675[8], sub_ln1497_reg_1675[8], sub_ln1497_reg_1675[8], sub_ln1497_reg_1675[8], sub_ln1497_reg_1675[8], sub_ln1497_reg_1675[8], sub_ln1497_reg_1675[8], sub_ln1497_reg_1675[8], sub_ln1497_reg_1675[8], sub_ln1497_reg_1675[8], sub_ln1497_reg_1675[8], sub_ln1497_reg_1675 };
assign ashr_ln1497_fu_334_p2 = $signed(op_0) >>> { ret_V_2_reg_1669[7], ret_V_2_reg_1669[7], ret_V_2_reg_1669[7], ret_V_2_reg_1669[7], ret_V_2_reg_1669[7], ret_V_2_reg_1669[7], ret_V_2_reg_1669[7], ret_V_2_reg_1669[7], ret_V_2_reg_1669[7], ret_V_2_reg_1669[7], ret_V_2_reg_1669[7], ret_V_2_reg_1669[7], ret_V_2_reg_1669[7], ret_V_2_reg_1669[7], ret_V_2_reg_1669[7], ret_V_2_reg_1669[7], ret_V_2_reg_1669[7], ret_V_2_reg_1669[7], ret_V_2_reg_1669[7], ret_V_2_reg_1669[7], ret_V_2_reg_1669[7], ret_V_2_reg_1669[7], ret_V_2_reg_1669[7], ret_V_2_reg_1669[7], ret_V_2_reg_1669 };
assign ret_V_9_fu_1390_p2 = $signed(op_5) - $signed({ ret_V_21_reg_1718, 3'h0 });
assign sub_ln1497_fu_301_p2 = $signed(1'h0) - $signed(ret_V_2_fu_289_p3);
assign ush_fu_576_p2 = _046_ ? 1'h1 : 1'h0;
assign Range1_all_ones_fu_1014_p2 = _048_ ? 1'h1 : 1'h0;
assign Range1_all_zeros_fu_1020_p2 = _049_ ? 1'h1 : 1'h0;
assign deleted_ones_fu_1054_p3 = carry_1_fu_992_p2 ? and_ln780_fu_1048_p2 : Range1_all_ones_fu_1014_p2;
assign deleted_zeros_fu_1026_p3 = carry_1_fu_992_p2 ? Range1_all_ones_fu_1014_p2 : Range1_all_zeros_fu_1020_p2;
assign icmp_ln414_fu_776_p2 = _055_ ? 1'h1 : 1'h0;
assign icmp_ln785_fu_401_p2 = _056_ ? 1'h1 : 1'h0;
assign icmp_ln786_1_fu_425_p2 = _057_ ? 1'h1 : 1'h0;
assign icmp_ln786_fu_419_p2 = _050_ ? 1'h1 : 1'h0;
assign icmp_ln790_fu_443_p2 = _051_ ? 1'h1 : 1'h0;
assign icmp_ln851_1_fu_1208_p2 = _052_ ? 1'h1 : 1'h0;
assign icmp_ln851_2_fu_487_p2 = _053_ ? 1'h1 : 1'h0;
assign icmp_ln851_3_fu_691_p2 = _058_ ? 1'h1 : 1'h0;
assign icmp_ln851_4_fu_1480_p2 = _059_ ? 1'h1 : 1'h0;
assign icmp_ln851_fu_269_p2 = _054_ ? 1'h1 : 1'h0;
assign op_14_V_fu_1243_p3 = or_ln384_1_reg_1779 ? select_ln384_fu_1236_p3 : p_Val2_9_reg_1769;
assign op_17_V_fu_1496_p3 = select_ln340_fu_1490_p3 ? 2'h0 : p_Val2_4_reg_1836;
assign op_19_V_fu_864_p3 = and_ln340_fu_838_p2 ? { 1'h0, p_Val2_7_fu_844_p2 } : { p_Val2_6_fu_792_p2[2], p_Val2_6_fu_792_p2 };
assign op_27 = ret_V_28_reg_1886[33] ? select_ln850_7_fu_1644_p3 : ret_V_28_cast_reg_1891;
assign op_2_V_fu_552_p3 = or_ln384_fu_547_p2 ? select_ln384_1_fu_540_p3 : { select_ln1497_reg_1687[2:0], 5'h00 };
assign ret_V_19_fu_1228_p3 = r_V_fu_1180_p2[5] ? select_ln850_1_fu_1220_p3 : r_V_fu_1180_p2[4:3];
assign ret_V_21_fu_507_p3 = ret_V_20_fu_460_p2[15] ? select_ln850_2_fu_499_p3 : ret_V_20_fu_460_p2[11:8];
assign ret_V_24_fu_1420_p3 = ret_V_23_reg_1810[33] ? select_ln850_4_fu_1414_p3 : ret_V_19_cast_reg_1815;
assign ret_V_27_fu_1582_p3 = ret_V_26_reg_1869[33] ? select_ln850_6_fu_1575_p3 : ret_V_25_cast_reg_1874;
assign ret_V_2_fu_289_p3 = op_1[15] ? select_ln850_fu_281_p3 : { 1'h0, op_1[14:8] };
assign rhs_1_fu_315_p2 = _060_ ? 1'h1 : 1'h0;
assign select_ln1118_1_fu_715_p3 = ush_reg_1724 ? 2'h3 : 2'h0;
assign select_ln1118_fu_704_p3 = ush_reg_1724 ? 4'hf : 4'h0;
assign select_ln1345_fu_621_p3 = rhs_1_reg_1680 ? 2'h3 : 2'h0;
assign select_ln1497_fu_349_p3 = ret_V_2_reg_1669[7] ? shl_ln1497_fu_343_p2 : ashr_ln1497_fu_334_p2;
assign select_ln340_2_fu_830_p3 = p_Val2_6_fu_792_p2[2] ? xor_ln785_1_fu_824_p2 : and_ln783_fu_810_p2[3];
assign select_ln340_fu_1490_p3 = p_Result_26_reg_1841 ? xor_ln410_reg_1831 : neg_src_2_fu_1486_p2;
assign select_ln353_2_fu_1525_p3 = ret_V_25_reg_1847[36] ? select_ln850_8_fu_1519_p3 : ret_V_22_cast_reg_1852;
assign select_ln353_fu_1265_p3 = ret_V_22_reg_1784[25] ? select_ln850_5_fu_1260_p3 : sext_ln850_reg_1789;
assign select_ln384_1_fu_540_p3 = overflow_reg_1697 ? 8'h7f : 8'h81;
assign select_ln384_fu_1236_p3 = overflow_1_reg_1774 ? 2'h1 : 2'h3;
assign select_ln850_1_fu_1220_p3 = icmp_ln851_1_fu_1208_p2 ? r_V_fu_1180_p2[4:3] : ret_V_3_fu_1214_p2;
assign select_ln850_2_fu_499_p3 = icmp_ln851_2_fu_487_p2 ? ret_V_20_fu_460_p2[11:8] : ret_V_7_fu_493_p2;
assign select_ln850_4_fu_1414_p3 = op_14_V_reg_1805[0] ? add_ln691_1_reg_1821 : ret_V_19_cast_reg_1815;
assign select_ln850_5_fu_1260_p3 = icmp_ln851_3_reg_1751 ? add_ln691_reg_1795 : sext_ln850_reg_1789;
assign select_ln850_6_fu_1575_p3 = op_17_V_reg_1864[0] ? add_ln691_3_fu_1570_p2 : ret_V_25_cast_reg_1874;
assign select_ln850_7_fu_1644_p3 = op_19_V_reg_1763[0] ? add_ln691_4_fu_1639_p2 : ret_V_28_cast_reg_1891;
assign select_ln850_8_fu_1519_p3 = icmp_ln851_4_reg_1859 ? add_ln691_2_fu_1510_p2 : ret_V_22_cast_reg_1852;
assign select_ln850_fu_281_p3 = icmp_ln851_fu_269_p2 ? { 1'h1, op_1[14:8] } : ret_V_1_fu_275_p2;
assign signbit_fu_607_p2 = _061_ ? 1'h1 : 1'h0;
assign ret_V_20_fu_460_p2 = { rhs_1_reg_1680, 8'h00 } ^ op_1;
assign Range2_all_ones_fu_896_p1 = op_5;
assign Range2_all_ones_fu_896_p3 = op_5[3];
assign and_ln_fu_373_p3 = { select_ln1497_fu_349_p3[2], 7'h00 };
assign ap_CS_fsm_state1 = ap_CS_fsm[0];
assign ap_CS_fsm_state10 = ap_CS_fsm[9];
assign ap_CS_fsm_state2 = ap_CS_fsm[1];
assign ap_CS_fsm_state3 = ap_CS_fsm[2];
assign ap_CS_fsm_state4 = ap_CS_fsm[3];
assign ap_CS_fsm_state5 = ap_CS_fsm[4];
assign ap_CS_fsm_state6 = ap_CS_fsm[5];
assign ap_CS_fsm_state7 = ap_CS_fsm[6];
assign ap_CS_fsm_state8 = ap_CS_fsm[7];
assign ap_CS_fsm_state9 = ap_CS_fsm[8];
assign ap_done = op_27_ap_vld;
assign ap_ready = op_27_ap_vld;
assign conv_i847_fu_331_p0 = op_0;
assign conv_i847_fu_331_p1 = { op_0[7], op_0[7], op_0[7], op_0[7], op_0[7], op_0[7], op_0[7], op_0[7], op_0[7], op_0[7], op_0[7], op_0[7], op_0[7], op_0[7], op_0[7], op_0[7], op_0[7], op_0[7], op_0[7], op_0[7], op_0[7], op_0[7], op_0[7], op_0[7], op_0 };
assign neg_src_4_fu_816_p3 = and_ln783_fu_810_p2[3];
assign op_13_V_fu_697_p3 = { ret_V_5_reg_1731, 15'h0000 };
assign op_16_V_fu_1396_p3 = { ret_V_9_fu_1390_p2, 1'h0 };
assign op_8_V_fu_613_p3 = { signbit_fu_607_p2, 2'h0 };
assign or_ln1195_1_fu_904_p1 = op_5;
assign or_ln_fu_391_p4 = { select_ln1497_fu_349_p3[2], 2'h0, select_ln1497_fu_349_p3[7:3] };
assign p_Result_12_fu_854_p4 = { 1'h0, p_Val2_7_fu_844_p2 };
assign p_Result_16_fu_928_p3 = or_ln1195_1_fu_904_p2[2];
assign p_Result_18_fu_1249_p3 = ret_V_22_reg_1784[25];
assign p_Result_19_fu_1404_p3 = ret_V_23_reg_1810[33];
assign p_Result_1_fu_1472_p3 = { ret_V_9_fu_1390_p2[2:0], 1'h0 };
assign p_Result_20_fu_1503_p3 = ret_V_25_reg_1847[36];
assign p_Result_21_fu_1560_p3 = ret_V_26_reg_1869[33];
assign p_Result_22_fu_1629_p3 = ret_V_28_reg_1886[33];
assign p_Result_23_fu_357_p3 = select_ln1497_fu_349_p3[7];
assign p_Result_24_fu_1314_p3 = r_V_1_fu_1309_p2[3];
assign p_Result_25_fu_1332_p3 = r_V_1_fu_1309_p2[1];
assign p_Result_27_fu_728_p3 = r_V_2_fu_722_p2[3];
assign p_Result_28_fu_802_p3 = p_Val2_6_fu_792_p2[2];
assign p_Result_29_fu_910_p1 = op_5;
assign p_Result_29_fu_910_p3 = op_5[3];
assign p_Result_2_fu_1196_p3 = r_V_fu_1180_p2[5];
assign p_Result_30_fu_936_p1 = op_5;
assign p_Result_30_fu_936_p3 = op_5[1];
assign p_Result_31_fu_948_p3 = or_ln1195_1_fu_904_p2[3];
assign p_Result_32_fu_978_p3 = p_Val2_9_fu_972_p2[1];
assign p_Result_3_fu_683_p3 = { ret_V_5_fu_590_p2[4:0], 15'h0000 };
assign p_Result_4_fu_475_p3 = ret_V_20_fu_460_p2[15];
assign p_Result_5_fu_435_p3 = { select_ln1497_fu_349_p3[1:0], 5'h00 };
assign p_Result_s_22_fu_381_p4 = select_ln1497_fu_349_p3[7:3];
assign p_Result_s_fu_257_p3 = op_1[15];
assign p_Val2_8_fu_918_p4 = or_ln1195_1_fu_904_p2[3:2];
assign p_Val2_s_fu_518_p3 = { select_ln1497_reg_1687[2:0], 5'h00 };
assign r_1_fu_944_p1 = or_ln1195_fu_890_p2[0];
assign r_V_1_fu_1309_p0 = op_5;
assign r_V_2_fu_722_p1 = op_5;
assign r_fu_1340_p1 = r_V_1_fu_1309_p2[0];
assign ret_V_19_cast_fu_1290_p4 = { ret_V_23_fu_1284_p2[33], ret_V_23_fu_1284_p2[33], ret_V_23_fu_1284_p2[33], ret_V_23_fu_1284_p2[33], ret_V_23_fu_1284_p2[33], ret_V_23_fu_1284_p2[33], ret_V_23_fu_1284_p2[33], ret_V_23_fu_1284_p2[33], ret_V_23_fu_1284_p2[33], ret_V_23_fu_1284_p2[33], ret_V_23_fu_1284_p2[33], ret_V_23_fu_1284_p2[33], ret_V_23_fu_1284_p2[33], ret_V_23_fu_1284_p2[33], ret_V_23_fu_1284_p2[33], ret_V_23_fu_1284_p2[33], ret_V_23_fu_1284_p2[33], ret_V_23_fu_1284_p2[33], ret_V_23_fu_1284_p2[33], ret_V_23_fu_1284_p2[33], ret_V_23_fu_1284_p2[33], ret_V_23_fu_1284_p2[33], ret_V_23_fu_1284_p2[33], ret_V_23_fu_1284_p2[33], ret_V_23_fu_1284_p2[33], ret_V_23_fu_1284_p2[7:1] };
assign ret_V_23_fu_1284_p2[32:8] = { ret_V_23_fu_1284_p2[33], ret_V_23_fu_1284_p2[33], ret_V_23_fu_1284_p2[33], ret_V_23_fu_1284_p2[33], ret_V_23_fu_1284_p2[33], ret_V_23_fu_1284_p2[33], ret_V_23_fu_1284_p2[33], ret_V_23_fu_1284_p2[33], ret_V_23_fu_1284_p2[33], ret_V_23_fu_1284_p2[33], ret_V_23_fu_1284_p2[33], ret_V_23_fu_1284_p2[33], ret_V_23_fu_1284_p2[33], ret_V_23_fu_1284_p2[33], ret_V_23_fu_1284_p2[33], ret_V_23_fu_1284_p2[33], ret_V_23_fu_1284_p2[33], ret_V_23_fu_1284_p2[33], ret_V_23_fu_1284_p2[33], ret_V_23_fu_1284_p2[33], ret_V_23_fu_1284_p2[33], ret_V_23_fu_1284_p2[33], ret_V_23_fu_1284_p2[33], ret_V_23_fu_1284_p2[33], ret_V_23_fu_1284_p2[33] };
assign ret_V_3_cast_fu_1186_p4 = r_V_fu_1180_p2[4:3];
assign ret_V_8_cast_fu_465_p4 = ret_V_20_fu_460_p2[11:8];
assign ret_V_fu_247_p4 = op_1[15:8];
assign rhs_10_fu_1440_p3 = { op_23_V_fu_1430_p2, 4'h0 };
assign rhs_11_fu_1532_p3 = { select_ln353_2_fu_1525_p3, 1'h0 };
assign rhs_13_fu_1602_p3 = { op_26_V_reg_1881, 1'h0 };
assign rhs_2_fu_449_p3 = { rhs_1_reg_1680, 8'h00 };
assign rhs_4_fu_1383_p3 = { ret_V_21_reg_1718, 3'h0 };
assign rhs_5_fu_872_p3 = { ret_reg_1736, 3'h0 };
assign rhs_7_fu_651_p3 = { op_12_V_fu_638_p2, 2'h0 };
assign rhs_8_fu_1136_p3 = { tmp_1_reg_1746, 20'h00000 };
assign rhs_fu_582_p3 = { op_6, 5'h00 };
assign sext_ln1192_1_fu_1143_p1 = { tmp_1_reg_1746[4], tmp_1_reg_1746, 20'h00000 };
assign sext_ln1192_2_fu_1280_p1 = { select_ln353_fu_1265_p3[6], select_ln353_fu_1265_p3[6], select_ln353_fu_1265_p3[6], select_ln353_fu_1265_p3[6], select_ln353_fu_1265_p3[6], select_ln353_fu_1265_p3[6], select_ln353_fu_1265_p3[6], select_ln353_fu_1265_p3[6], select_ln353_fu_1265_p3[6], select_ln353_fu_1265_p3[6], select_ln353_fu_1265_p3[6], select_ln353_fu_1265_p3[6], select_ln353_fu_1265_p3[6], select_ln353_fu_1265_p3[6], select_ln353_fu_1265_p3[6], select_ln353_fu_1265_p3[6], select_ln353_fu_1265_p3[6], select_ln353_fu_1265_p3[6], select_ln353_fu_1265_p3[6], select_ln353_fu_1265_p3[6], select_ln353_fu_1265_p3[6], select_ln353_fu_1265_p3[6], select_ln353_fu_1265_p3[6], select_ln353_fu_1265_p3[6], select_ln353_fu_1265_p3[6], select_ln353_fu_1265_p3[6], select_ln353_fu_1265_p3, 1'h0 };
assign sext_ln1192_3_fu_1448_p1 = { op_23_V_fu_1430_p2[31], op_23_V_fu_1430_p2, 4'h0 };
assign sext_ln1192_4_fu_1540_p1 = { select_ln353_2_fu_1525_p3[31], select_ln353_2_fu_1525_p3, 1'h0 };
assign sext_ln1192_5_fu_1609_p1 = { op_26_V_reg_1881[31], op_26_V_reg_1881, 1'h0 };
assign sext_ln1192_fu_659_p1 = { op_12_V_fu_638_p2[3], op_12_V_fu_638_p2, 2'h0 };
assign sext_ln1193_fu_1380_p0 = op_5;
assign sext_ln1193_fu_1380_p1 = { op_5[3], op_5[3], op_5[3], op_5 };
assign sext_ln1195_fu_886_p0 = op_5;
assign sext_ln1195_fu_886_p1 = { op_5[3], op_5 };
assign sext_ln1497_1_fu_340_p1 = { sub_ln1497_reg_1675[8], sub_ln1497_reg_1675[8], sub_ln1497_reg_1675[8], sub_ln1497_reg_1675[8], sub_ln1497_reg_1675[8], sub_ln1497_reg_1675[8], sub_ln1497_reg_1675[8], sub_ln1497_reg_1675[8], sub_ln1497_reg_1675[8], sub_ln1497_reg_1675[8], sub_ln1497_reg_1675[8], sub_ln1497_reg_1675[8], sub_ln1497_reg_1675[8], sub_ln1497_reg_1675[8], sub_ln1497_reg_1675[8], sub_ln1497_reg_1675[8], sub_ln1497_reg_1675[8], sub_ln1497_reg_1675[8], sub_ln1497_reg_1675[8], sub_ln1497_reg_1675[8], sub_ln1497_reg_1675[8], sub_ln1497_reg_1675[8], sub_ln1497_reg_1675[8], sub_ln1497_reg_1675 };
assign sext_ln1497_fu_297_p1 = { ret_V_2_fu_289_p3[7], ret_V_2_fu_289_p3 };
assign sext_ln367_fu_850_p1 = { p_Val2_7_fu_844_p2[2], p_Val2_7_fu_844_p2 };
assign sext_ln545_fu_321_p1 = { ret_V_2_reg_1669[7], ret_V_2_reg_1669[7], ret_V_2_reg_1669[7], ret_V_2_reg_1669[7], ret_V_2_reg_1669[7], ret_V_2_reg_1669[7], ret_V_2_reg_1669[7], ret_V_2_reg_1669[7], ret_V_2_reg_1669[7], ret_V_2_reg_1669[7], ret_V_2_reg_1669[7], ret_V_2_reg_1669[7], ret_V_2_reg_1669[7], ret_V_2_reg_1669[7], ret_V_2_reg_1669[7], ret_V_2_reg_1669[7], ret_V_2_reg_1669[7], ret_V_2_reg_1669[7], ret_V_2_reg_1669[7], ret_V_2_reg_1669[7], ret_V_2_reg_1669[7], ret_V_2_reg_1669[7], ret_V_2_reg_1669[7], ret_V_2_reg_1669[7], ret_V_2_reg_1669 };
assign sext_ln69_1_fu_1589_p1 = { op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18 };
assign sext_ln69_fu_1427_p1 = { ret_V_19_reg_1800[1], ret_V_19_reg_1800[1], ret_V_19_reg_1800[1], ret_V_19_reg_1800[1], ret_V_19_reg_1800[1], ret_V_19_reg_1800[1], ret_V_19_reg_1800[1], ret_V_19_reg_1800[1], ret_V_19_reg_1800[1], ret_V_19_reg_1800[1], ret_V_19_reg_1800[1], ret_V_19_reg_1800[1], ret_V_19_reg_1800[1], ret_V_19_reg_1800[1], ret_V_19_reg_1800[1], ret_V_19_reg_1800[1], ret_V_19_reg_1800[1], ret_V_19_reg_1800[1], ret_V_19_reg_1800[1], ret_V_19_reg_1800[1], ret_V_19_reg_1800[1], ret_V_19_reg_1800[1], ret_V_19_reg_1800[1], ret_V_19_reg_1800[1], ret_V_19_reg_1800[1], ret_V_19_reg_1800[1], ret_V_19_reg_1800[1], ret_V_19_reg_1800[1], ret_V_19_reg_1800[1], ret_V_19_reg_1800[1], ret_V_19_reg_1800 };
assign sext_ln703_1_fu_1436_p1 = { ret_V_9_fu_1390_p2[6], ret_V_9_fu_1390_p2[6], ret_V_9_fu_1390_p2[6], ret_V_9_fu_1390_p2[6], ret_V_9_fu_1390_p2[6], ret_V_9_fu_1390_p2[6], ret_V_9_fu_1390_p2[6], ret_V_9_fu_1390_p2[6], ret_V_9_fu_1390_p2[6], ret_V_9_fu_1390_p2[6], ret_V_9_fu_1390_p2[6], ret_V_9_fu_1390_p2[6], ret_V_9_fu_1390_p2[6], ret_V_9_fu_1390_p2[6], ret_V_9_fu_1390_p2[6], ret_V_9_fu_1390_p2[6], ret_V_9_fu_1390_p2[6], ret_V_9_fu_1390_p2[6], ret_V_9_fu_1390_p2[6], ret_V_9_fu_1390_p2[6], ret_V_9_fu_1390_p2[6], ret_V_9_fu_1390_p2[6], ret_V_9_fu_1390_p2[6], ret_V_9_fu_1390_p2[6], ret_V_9_fu_1390_p2[6], ret_V_9_fu_1390_p2[6], ret_V_9_fu_1390_p2[6], ret_V_9_fu_1390_p2[6], ret_V_9_fu_1390_p2[6], ret_V_9_fu_1390_p2, 1'h0 };
assign sext_ln703_2_fu_1515_p1 = { op_17_V_fu_1496_p3[1], op_17_V_fu_1496_p3[1], op_17_V_fu_1496_p3[1], op_17_V_fu_1496_p3[1], op_17_V_fu_1496_p3[1], op_17_V_fu_1496_p3[1], op_17_V_fu_1496_p3[1], op_17_V_fu_1496_p3[1], op_17_V_fu_1496_p3[1], op_17_V_fu_1496_p3[1], op_17_V_fu_1496_p3[1], op_17_V_fu_1496_p3[1], op_17_V_fu_1496_p3[1], op_17_V_fu_1496_p3[1], op_17_V_fu_1496_p3[1], op_17_V_fu_1496_p3[1], op_17_V_fu_1496_p3[1], op_17_V_fu_1496_p3[1], op_17_V_fu_1496_p3[1], op_17_V_fu_1496_p3[1], op_17_V_fu_1496_p3[1], op_17_V_fu_1496_p3[1], op_17_V_fu_1496_p3[1], op_17_V_fu_1496_p3[1], op_17_V_fu_1496_p3[1], op_17_V_fu_1496_p3[1], op_17_V_fu_1496_p3[1], op_17_V_fu_1496_p3[1], op_17_V_fu_1496_p3[1], op_17_V_fu_1496_p3[1], op_17_V_fu_1496_p3[1], op_17_V_fu_1496_p3[1], op_17_V_fu_1496_p3 };
assign sext_ln703_3_fu_1599_p1 = { op_19_V_reg_1763[3], op_19_V_reg_1763[3], op_19_V_reg_1763[3], op_19_V_reg_1763[3], op_19_V_reg_1763[3], op_19_V_reg_1763[3], op_19_V_reg_1763[3], op_19_V_reg_1763[3], op_19_V_reg_1763[3], op_19_V_reg_1763[3], op_19_V_reg_1763[3], op_19_V_reg_1763[3], op_19_V_reg_1763[3], op_19_V_reg_1763[3], op_19_V_reg_1763[3], op_19_V_reg_1763[3], op_19_V_reg_1763[3], op_19_V_reg_1763[3], op_19_V_reg_1763[3], op_19_V_reg_1763[3], op_19_V_reg_1763[3], op_19_V_reg_1763[3], op_19_V_reg_1763[3], op_19_V_reg_1763[3], op_19_V_reg_1763[3], op_19_V_reg_1763[3], op_19_V_reg_1763[3], op_19_V_reg_1763[3], op_19_V_reg_1763[3], op_19_V_reg_1763[3], op_19_V_reg_1763 };
assign sext_ln703_fu_1256_p1 = { op_14_V_fu_1243_p3[1], op_14_V_fu_1243_p3[1], op_14_V_fu_1243_p3[1], op_14_V_fu_1243_p3[1], op_14_V_fu_1243_p3[1], op_14_V_fu_1243_p3[1], op_14_V_fu_1243_p3[1], op_14_V_fu_1243_p3[1], op_14_V_fu_1243_p3[1], op_14_V_fu_1243_p3[1], op_14_V_fu_1243_p3[1], op_14_V_fu_1243_p3[1], op_14_V_fu_1243_p3[1], op_14_V_fu_1243_p3[1], op_14_V_fu_1243_p3[1], op_14_V_fu_1243_p3[1], op_14_V_fu_1243_p3[1], op_14_V_fu_1243_p3[1], op_14_V_fu_1243_p3[1], op_14_V_fu_1243_p3[1], op_14_V_fu_1243_p3[1], op_14_V_fu_1243_p3[1], op_14_V_fu_1243_p3[1], op_14_V_fu_1243_p3[1], op_14_V_fu_1243_p3[1], op_14_V_fu_1243_p3[1], op_14_V_fu_1243_p3[1], op_14_V_fu_1243_p3[1], op_14_V_fu_1243_p3[1], op_14_V_fu_1243_p3[1], op_14_V_fu_1243_p3[1], op_14_V_fu_1243_p3[1], op_14_V_fu_1243_p3 };
assign sext_ln713_fu_746_p1 = { r_V_2_fu_722_p2[3], r_V_2_fu_722_p2[3:2] };
assign sext_ln727_fu_564_p1 = { op_2_V_fu_552_p3[7], op_2_V_fu_552_p3[7], op_2_V_fu_552_p3[7], op_2_V_fu_552_p3[7], op_2_V_fu_552_p3[7], op_2_V_fu_552_p3 };
assign sext_ln745_fu_798_p1 = { p_Val2_6_fu_792_p2[2], p_Val2_6_fu_792_p2 };
assign sext_ln850_fu_1163_p1 = { ret_V_22_fu_1147_p2[25], ret_V_22_fu_1147_p2[25:20] };
assign shl_ln728_1_fu_568_p3 = { op_4, 5'h00 };
assign shl_ln728_5_fu_596_p3 = { rhs_1_reg_1680, 5'h00 };
assign shl_ln_fu_307_p1 = op_0;
assign shl_ln_fu_307_p3 = { op_0, 8'h00 };
assign tmp_13_fu_760_p3 = and_ln414_fu_754_p2[1];
assign tmp_23_fu_998_p3 = or_ln1195_fu_890_p2[4];
assign tmp_24_fu_1034_p3 = or_ln1195_fu_890_p2[4];
assign tmp_26_fu_1272_p3 = { select_ln353_fu_1265_p3, 1'h0 };
assign tmp_3_fu_768_p3 = { and_ln414_fu_754_p2[1], r_V_2_fu_722_p2[0] };
assign tmp_4_fu_365_p3 = select_ln1497_fu_349_p3[2];
assign tmp_9_fu_1006_p3 = { op_5[3], or_ln1195_fu_890_p2[4] };
assign tmp_fu_324_p3 = ret_V_2_reg_1669[7];
assign tmp_s_fu_1153_p4 = ret_V_22_fu_1147_p2[25:20];
assign trunc_ln1118_fu_711_p0 = op_5;
assign trunc_ln1118_fu_711_p1 = op_5[1:0];
assign trunc_ln1195_1_fu_879_p3 = { trunc_ln1195_reg_1741, 3'h0 };
assign trunc_ln1195_fu_643_p1 = ret_fu_628_p2[0];
assign trunc_ln1349_fu_634_p1 = op_4[3:0];
assign trunc_ln1_fu_1322_p4 = r_V_1_fu_1309_p2[3:2];
assign trunc_ln708_1_fu_736_p4 = r_V_2_fu_722_p2[3:2];
assign trunc_ln718_fu_750_p1 = r_V_2_fu_722_p2[0];
assign trunc_ln731_fu_515_p1 = select_ln1497_reg_1687[2:0];
assign trunc_ln790_1_fu_1092_p1 = p_Val2_9_fu_972_p2[0];
assign trunc_ln790_fu_431_p1 = select_ln1497_fu_349_p3[1:0];
assign trunc_ln851_1_fu_1204_p1 = r_V_fu_1180_p2[2:0];
assign trunc_ln851_2_fu_483_p1 = ret_V_20_fu_460_p2[7:0];
assign trunc_ln851_3_fu_679_p1 = ret_V_5_fu_590_p2[4:0];
assign trunc_ln851_4_fu_1411_p1 = op_14_V_reg_1805[0];
assign trunc_ln851_5_fu_1468_p1 = ret_V_9_fu_1390_p2[2:0];
assign trunc_ln851_6_fu_1567_p1 = op_17_V_reg_1864[0];
assign trunc_ln851_7_fu_1636_p1 = op_19_V_reg_1763[0];
assign trunc_ln851_fu_265_p1 = op_1[7:0];
assign trunc_ln8_fu_560_p1 = op_2_V_fu_552_p3[6:0];
assign zext_ln1192_fu_1132_p1 = { 4'h0, ret_V_5_reg_1731, 15'h0000 };
assign zext_ln1196_fu_456_p1 = { 7'h00, rhs_1_reg_1680, 8'h00 };
assign zext_ln1380_fu_1306_p1 = { 3'h0, ush_reg_1724 };
assign zext_ln1499_fu_603_p1 = { 2'h0, rhs_1_reg_1680, 5'h00 };
assign zext_ln415_1_fu_788_p1 = { 2'h0, and_ln414_1_fu_782_p2 };
assign zext_ln415_2_fu_968_p1 = { 1'h0, and_ln412_fu_962_p2 };
assign zext_ln415_fu_1362_p1 = { 1'h0, and_ln410_fu_1356_p2 };
assign zext_ln703_fu_647_p1 = { 4'h0, signbit_fu_607_p2, 2'h0 };
assign \mul_4s_2s_6_1_1_U1.top_mul_4s_2s_6_1_1_Multiplier_0_U.a  = \mul_4s_2s_6_1_1_U1.din0 ;
assign \mul_4s_2s_6_1_1_U1.top_mul_4s_2s_6_1_1_Multiplier_0_U.b  = \mul_4s_2s_6_1_1_U1.din1 ;
assign \mul_4s_2s_6_1_1_U1.dout  = \mul_4s_2s_6_1_1_U1.top_mul_4s_2s_6_1_1_Multiplier_0_U.p ;
assign \mul_4s_2s_6_1_1_U1.din0  = op_5;
assign \mul_4s_2s_6_1_1_U1.din1  = op_11;
assign r_V_fu_1180_p2 = \mul_4s_2s_6_1_1_U1.dout ;
endmodule


// Product machine:
module top_A_times_top_B (ap_start, op_0, op_1, op_11, op_18, op_4, op_5, op_6, ap_clk, unsafe_signal);
input ap_start;
input [7:0] op_0;
input [15:0] op_1;
input [1:0] op_11;
input [1:0] op_18;
input [7:0] op_4;
input [3:0] op_5;
input [1:0] op_6;
input ap_clk;
output unsafe_signal;
reg _setup;
initial _setup = 1'b0;
always @ (posedge ap_clk) _setup <= 1'b1;
reg ap_start_internal;
always @ (posedge ap_clk) if (!_setup) ap_start_internal <= ap_start;
reg [7:0] op_0_internal;
always @ (posedge ap_clk) if (!_setup) op_0_internal <= op_0;
reg [15:0] op_1_internal;
always @ (posedge ap_clk) if (!_setup) op_1_internal <= op_1;
reg [1:0] op_11_internal;
always @ (posedge ap_clk) if (!_setup) op_11_internal <= op_11;
reg [1:0] op_18_internal;
always @ (posedge ap_clk) if (!_setup) op_18_internal <= op_18;
reg [7:0] op_4_internal;
always @ (posedge ap_clk) if (!_setup) op_4_internal <= op_4;
reg [3:0] op_5_internal;
always @ (posedge ap_clk) if (!_setup) op_5_internal <= op_5;
reg [1:0] op_6_internal;
always @ (posedge ap_clk) if (!_setup) op_6_internal <= op_6;
wire ap_done_A;
wire ap_done_B;
wire ap_done_eq;
assign ap_done_eq = ap_done_A == ap_done_B;
wire ap_idle_A;
wire ap_idle_B;
wire ap_idle_eq;
assign ap_idle_eq = ap_idle_A == ap_idle_B;
wire ap_ready_A;
wire ap_ready_B;
wire ap_ready_eq;
assign ap_ready_eq = ap_ready_A == ap_ready_B;
wire [31:0] op_27_A;
wire [31:0] op_27_B;
wire op_27_eq;
assign op_27_eq = op_27_A == op_27_B;
wire op_27_ap_vld_A;
wire op_27_ap_vld_B;
wire clk_enable_A;
wire clk_enable_B;
assign clk_enable_A = _setup & (~op_27_ap_vld_A | op_27_ap_vld_B);
assign clk_enable_B = _setup;
wire divergent;
assign divergent = ~(ap_done_eq & ap_idle_eq & ap_ready_eq & op_27_eq);
assign unsafe_signal = op_27_ap_vld_A & op_27_ap_vld_B & divergent;
top_A instance_A (
    .ap_clk(ap_clk),
    .clk_enable(clk_enable_A),
    .ap_start(ap_start_internal),
    .op_0(op_0_internal),
    .op_1(op_1_internal),
    .op_11(op_11_internal),
    .op_18(op_18_internal),
    .op_4(op_4_internal),
    .op_5(op_5_internal),
    .op_6(op_6_internal),
    .ap_done(ap_done_A),
    .ap_idle(ap_idle_A),
    .ap_ready(ap_ready_A),
    .op_27(op_27_A),
    .op_27_ap_vld(op_27_ap_vld_A)
);
top_B instance_B (
    .ap_clk(ap_clk),
    .clk_enable(clk_enable_B),
    .ap_start(ap_start_internal),
    .op_0(op_0_internal),
    .op_1(op_1_internal),
    .op_11(op_11_internal),
    .op_18(op_18_internal),
    .op_4(op_4_internal),
    .op_5(op_5_internal),
    .op_6(op_6_internal),
    .ap_done(ap_done_B),
    .ap_idle(ap_idle_B),
    .ap_ready(ap_ready_B),
    .op_27(op_27_B),
    .op_27_ap_vld(op_27_ap_vld_B)
);
endmodule
