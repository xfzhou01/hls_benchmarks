// Processed by function `construct_kairos` in `verilog_tricks.py`.
// Machine A:
// Processed by function `add_clk_enable_signal` in `verilog_tricks.py`.
// Processed by function `remove_reset_signal` in `verilog_tricks.py`.
module top_A (
  ap_clk,
  ap_start,
  ap_done,
  ap_idle,
  ap_ready,
  op_0,
  op_2,
  op_4,
  op_6,
  op_7,
  op_8,
  op_10,
  op_12,
  op_14,
  op_15,
  op_16,
  op_18,
  op_31,
  op_31_ap_vld,
clk_enable
);
input clk_enable;


input ap_clk;
wire ap_rst;
assign ap_rst = op_31_ap_vld;
input ap_start;
input [7:0] op_0;
input [7:0] op_10;
input [1:0] op_12;
input [7:0] op_14;
input [7:0] op_15;
input op_16;
input [3:0] op_18;
input [3:0] op_2;
input [7:0] op_4;
input [7:0] op_6;
input [7:0] op_7;
input [3:0] op_8;
output ap_done;
output ap_idle;
output ap_ready;
output [31:0] op_31;
output op_31_ap_vld;


reg [31:0] add_ln691_reg_642;
reg [4:0] add_ln69_5_reg_679;
reg [8:0] add_ln69_reg_620;
reg [7:0] ap_CS_fsm = 8'h01;
reg icmp_ln851_1_reg_669;
reg icmp_ln886_reg_610;
reg op_17_V_reg_652;
reg [10:0] op_21_V_reg_615;
reg [31:0] op_25_V_reg_647;
reg [5:0] ret_V_11_reg_594;
reg [33:0] ret_V_12_reg_630;
reg [36:0] ret_V_14_reg_657;
reg [31:0] ret_V_15_reg_674;
reg [31:0] ret_V_19_cast_reg_662;
reg [4:0] ret_V_2_reg_605;
reg [31:0] ret_V_8_cast_reg_635;
reg [4:0] ret_V_reg_599;
reg [9:0] ret_reg_589;
wire [31:0] _000_;
wire [4:0] _001_;
wire [8:0] _002_;
wire [7:0] _003_;
wire _004_;
wire _005_;
wire _006_;
wire [10:0] _007_;
wire [31:0] _008_;
wire [5:0] _009_;
wire [33:0] _010_;
wire [36:0] _011_;
wire [31:0] _012_;
wire [31:0] _013_;
wire [4:0] _014_;
wire [31:0] _015_;
wire [4:0] _016_;
wire [9:0] _017_;
wire [1:0] _018_;
wire _019_;
wire _020_;
wire _021_;
wire _022_;
wire _023_;
wire _024_;
wire _025_;
wire _026_;
wire _027_;
wire _028_;
wire _029_;
wire _030_;
wire _031_;
wire _032_;
wire _033_;
wire [31:0] add_ln691_1_fu_523_p2;
wire [31:0] add_ln691_fu_367_p2;
wire [31:0] add_ln69_3_fu_569_p2;
wire [1:0] add_ln69_4_fu_549_p2;
wire [4:0] add_ln69_5_fu_559_p2;
wire [8:0] add_ln69_fu_317_p2;
wire ap_CS_fsm_state1;
wire ap_CS_fsm_state2;
wire ap_CS_fsm_state3;
wire ap_CS_fsm_state4;
wire ap_CS_fsm_state5;
wire ap_CS_fsm_state6;
wire ap_CS_fsm_state7;
wire ap_CS_fsm_state8;
wire [7:0] ap_NS_fsm;
wire ap_clk;
wire ap_done;
wire ap_idle;
wire ap_ready;
wire ap_rst;
wire ap_start;
wire icmp_ln851_1_fu_507_p2;
wire icmp_ln851_fu_430_p2;
wire [7:0] icmp_ln886_fu_245_p0;
wire icmp_ln886_fu_245_p2;
wire [7:0] op_0;
wire [7:0] op_10;
wire [1:0] op_12;
wire [7:0] op_14;
wire [7:0] op_15;
wire op_16;
wire op_17_V_fu_466_p2;
wire [3:0] op_18;
wire [3:0] op_2;
wire [11:0] op_23_V_fu_329_p2;
wire [31:0] op_25_V_fu_398_p2;
wire [31:0] op_31;
wire op_31_ap_vld;
wire [7:0] op_4;
wire [7:0] op_6;
wire [7:0] op_7;
wire [3:0] op_8;
wire [15:0] op_9_V_fu_251_p3;
wire p_Result_1_fu_418_p3;
wire p_Result_2_fu_372_p3;
wire p_Result_3_fu_516_p3;
wire p_Result_s_fu_258_p3;
wire [16:0] p_Val2_2_fu_297_p2;
wire [5:0] ret_V_11_fu_223_p2;
wire [33:0] ret_V_12_fu_351_p2;
wire [31:0] ret_V_13_fu_388_p3;
wire [36:0] ret_V_14_fu_487_p2;
wire [31:0] ret_V_15_fu_534_p3;
wire [4:0] ret_V_2_fu_239_p2;
wire [2:0] ret_V_3_fu_404_p4;
wire [3:0] ret_V_4_fu_436_p2;
wire [3:0] ret_V_5_fu_450_p3;
wire [4:0] ret_V_fu_229_p4;
wire [9:0] ret_fu_201_p2;
wire [10:0] rhs_1_fu_285_p3;
wire [35:0] rhs_4_fu_476_p3;
wire [4:0] rhs_fu_211_p3;
wire [31:0] select_ln850_2_fu_382_p3;
wire [31:0] select_ln850_3_fu_528_p3;
wire [4:0] select_ln850_4_fu_272_p3;
wire [4:0] select_ln850_5_fu_278_p3;
wire [3:0] select_ln850_fu_442_p3;
wire [16:0] sext_ln1192_1_fu_268_p1;
wire [16:0] sext_ln1192_2_fu_293_p1;
wire [33:0] sext_ln1192_3_fu_347_p1;
wire [36:0] sext_ln1192_4_fu_483_p1;
wire [5:0] sext_ln1192_fu_219_p1;
wire [11:0] sext_ln20_fu_323_p1;
wire [7:0] sext_ln215_fu_193_p0;
wire [9:0] sext_ln215_fu_193_p1;
wire [1:0] sext_ln703_1_fu_335_p0;
wire [33:0] sext_ln703_1_fu_335_p1;
wire [7:0] sext_ln703_2_fu_472_p0;
wire [36:0] sext_ln703_2_fu_472_p1;
wire [3:0] sext_ln703_fu_207_p0;
wire [5:0] sext_ln703_fu_207_p1;
wire [3:0] sext_ln835_fu_414_p1;
wire [8:0] sext_ln886_fu_458_p1;
wire [12:0] tmp_3_fu_339_p3;
wire [4:0] trunc_ln851_1_fu_426_p1;
wire [1:0] trunc_ln851_2_fu_379_p0;
wire trunc_ln851_2_fu_379_p1;
wire [7:0] trunc_ln851_3_fu_503_p0;
wire [3:0] trunc_ln851_3_fu_503_p1;
wire [3:0] trunc_ln851_fu_265_p0;
wire trunc_ln851_fu_265_p1;
wire [1:0] zext_ln17_fu_513_p1;
wire [9:0] zext_ln215_fu_197_p1;
wire [31:0] zext_ln69_1_fu_395_p1;
wire [31:0] zext_ln69_2_fu_565_p1;
wire [11:0] zext_ln69_3_fu_326_p1;
wire [1:0] zext_ln69_4_fu_541_p1;
wire [4:0] zext_ln69_5_fu_545_p1;
wire [4:0] zext_ln69_6_fu_555_p1;
wire [31:0] zext_ln69_7_fu_574_p1;
wire [8:0] zext_ln69_fu_313_p1;
wire [8:0] zext_ln886_fu_462_p1;


assign add_ln691_1_fu_523_p2 = ret_V_19_cast_reg_662 + 1'h1;
assign add_ln691_fu_367_p2 = ret_V_8_cast_reg_635 + 1'h1;
assign add_ln69_3_fu_569_p2 = ret_V_15_reg_674 + op_15;
assign add_ln69_4_fu_549_p2 = op_16 + op_17_V_reg_652;
assign add_ln69_5_fu_559_p2 = add_ln69_4_fu_549_p2 + op_18;
assign add_ln69_fu_317_p2 = op_10 + 1'h1;
assign op_23_V_fu_329_p2 = $signed({ 1'h0, add_ln69_reg_620 }) + $signed(op_21_V_reg_615);
assign op_25_V_fu_398_p2 = ret_V_13_fu_388_p3 + icmp_ln886_reg_610;
assign op_31 = add_ln69_5_reg_679 + add_ln69_3_fu_569_p2;
assign p_Val2_2_fu_297_p2 = $signed({ select_ln850_5_fu_278_p3, 6'h00 }) + $signed({ ret_reg_589, 6'h00 });
assign ret_V_11_fu_223_p2 = $signed({ op_8, 1'h0 }) + $signed(op_2);
assign { ret_V_12_fu_351_p2[33], ret_V_12_fu_351_p2[12:0] } = $signed({ op_23_V_fu_329_p2, 1'h0 }) + $signed(op_12);
assign ret_V_14_fu_487_p2 = $signed({ op_25_V_reg_647, 4'h0 }) + $signed(op_14);
assign ret_V_2_fu_239_p2 = ret_V_11_fu_223_p2[5:1] + 1'h1;
assign ret_V_4_fu_436_p2 = $signed(op_0[7:5]) + $signed(2'h1);
assign _019_ = ap_CS_fsm[0] & _021_;
assign _020_ = ap_CS_fsm[0] & ap_start;
assign _021_ = ~ ap_start;
assign _022_ = ! op_0[4:0];
assign _023_ = $signed(op_4) > $signed(1'h0);
assign _024_ = $signed(ret_V_5_fu_450_p3) > $signed({ 1'h0, op_7 });
assign _025_ = | op_14[3:0];
always @(posedge ap_clk)
ret_V_12_reg_630 <= _010_;
always @(posedge ap_clk)
ret_V_8_cast_reg_635 <= _015_;
always @(posedge ap_clk)
op_25_V_reg_647 <= _008_;
always @(posedge ap_clk)
ret_reg_589 <= _017_;
always @(posedge ap_clk)
ret_V_11_reg_594 <= _009_;
always @(posedge ap_clk)
ret_V_reg_599 <= _016_;
always @(posedge ap_clk)
ret_V_2_reg_605 <= _014_;
always @(posedge ap_clk)
icmp_ln886_reg_610 <= _005_;
always @(posedge ap_clk)
op_17_V_reg_652 <= _006_;
always @(posedge ap_clk)
ret_V_14_reg_657 <= _011_;
always @(posedge ap_clk)
ret_V_19_cast_reg_662 <= _013_;
always @(posedge ap_clk)
icmp_ln851_1_reg_669 <= _004_;
always @(posedge ap_clk)
op_21_V_reg_615 <= _007_;
always @(posedge ap_clk)
add_ln69_reg_620 <= _002_;
always @(posedge ap_clk)
ret_V_15_reg_674 <= _012_;
always @(posedge ap_clk)
add_ln69_5_reg_679 <= _001_;
always @(posedge ap_clk)
add_ln691_reg_642 <= _000_;
always @(posedge ap_clk)
ap_CS_fsm <= _003_;
assign ap_idle = _019_ ? 1'h1 : 1'h0;
assign ap_done = ap_CS_fsm[7] ? 1'h1 : 1'h0;
assign _015_ = ap_CS_fsm[2] ? { ret_V_12_fu_351_p2[33], ret_V_12_fu_351_p2[33], ret_V_12_fu_351_p2[33], ret_V_12_fu_351_p2[33], ret_V_12_fu_351_p2[33], ret_V_12_fu_351_p2[33], ret_V_12_fu_351_p2[33], ret_V_12_fu_351_p2[33], ret_V_12_fu_351_p2[33], ret_V_12_fu_351_p2[33], ret_V_12_fu_351_p2[33], ret_V_12_fu_351_p2[33], ret_V_12_fu_351_p2[33], ret_V_12_fu_351_p2[33], ret_V_12_fu_351_p2[33], ret_V_12_fu_351_p2[33], ret_V_12_fu_351_p2[33], ret_V_12_fu_351_p2[33], ret_V_12_fu_351_p2[33], ret_V_12_fu_351_p2[33], ret_V_12_fu_351_p2[12:1] } : ret_V_8_cast_reg_635;
assign _010_ = ap_CS_fsm[2] ? { ret_V_12_fu_351_p2[33], ret_V_12_fu_351_p2[33], ret_V_12_fu_351_p2[33], ret_V_12_fu_351_p2[33], ret_V_12_fu_351_p2[33], ret_V_12_fu_351_p2[33], ret_V_12_fu_351_p2[33], ret_V_12_fu_351_p2[33], ret_V_12_fu_351_p2[33], ret_V_12_fu_351_p2[33], ret_V_12_fu_351_p2[33], ret_V_12_fu_351_p2[33], ret_V_12_fu_351_p2[33], ret_V_12_fu_351_p2[33], ret_V_12_fu_351_p2[33], ret_V_12_fu_351_p2[33], ret_V_12_fu_351_p2[33], ret_V_12_fu_351_p2[33], ret_V_12_fu_351_p2[33], ret_V_12_fu_351_p2[33], ret_V_12_fu_351_p2[33], ret_V_12_fu_351_p2[12:0] } : ret_V_12_reg_630;
assign _008_ = ap_CS_fsm[4] ? op_25_V_fu_398_p2 : op_25_V_reg_647;
assign _005_ = ap_CS_fsm[0] ? icmp_ln886_fu_245_p2 : icmp_ln886_reg_610;
assign _014_ = ap_CS_fsm[0] ? ret_V_2_fu_239_p2 : ret_V_2_reg_605;
assign _016_ = ap_CS_fsm[0] ? ret_V_11_fu_223_p2[5:1] : ret_V_reg_599;
assign _009_ = ap_CS_fsm[0] ? ret_V_11_fu_223_p2 : ret_V_11_reg_594;
assign _017_ = ap_CS_fsm[0] ? ret_fu_201_p2 : ret_reg_589;
assign _004_ = ap_CS_fsm[5] ? icmp_ln851_1_fu_507_p2 : icmp_ln851_1_reg_669;
assign _013_ = ap_CS_fsm[5] ? ret_V_14_fu_487_p2[35:4] : ret_V_19_cast_reg_662;
assign _011_ = ap_CS_fsm[5] ? ret_V_14_fu_487_p2 : ret_V_14_reg_657;
assign _006_ = ap_CS_fsm[5] ? op_17_V_fu_466_p2 : op_17_V_reg_652;
assign _002_ = ap_CS_fsm[1] ? add_ln69_fu_317_p2 : add_ln69_reg_620;
assign _007_ = ap_CS_fsm[1] ? p_Val2_2_fu_297_p2[16:6] : op_21_V_reg_615;
assign _001_ = ap_CS_fsm[6] ? add_ln69_5_fu_559_p2 : add_ln69_5_reg_679;
assign _012_ = ap_CS_fsm[6] ? ret_V_15_fu_534_p3 : ret_V_15_reg_674;
assign _000_ = ap_CS_fsm[3] ? add_ln691_fu_367_p2 : add_ln691_reg_642;
assign _003_ = ap_rst ? 8'h01 : ap_NS_fsm;
assign _018_ = _020_ ? 2'h2 : 2'h1;
assign _026_ = ap_CS_fsm == 1'h1;
function [7:0] _096_;
input [7:0] a;
input [63:0] b;
input [7:0] s;
case (s)
8'b00000001:
_096_ = b[7:0];
8'b00000010:
_096_ = b[15:8];
8'b00000100:
_096_ = b[23:16];
8'b00001000:
_096_ = b[31:24];
8'b00010000:
_096_ = b[39:32];
8'b00100000:
_096_ = b[47:40];
8'b01000000:
_096_ = b[55:48];
8'b10000000:
_096_ = b[63:56];
8'b00000000:
_096_ = a;
default:
_096_ = 8'bx;
endcase
endfunction
assign ap_NS_fsm = _096_(8'hxx, { 6'h00, _018_, 56'h04081020408001 }, { _026_, _033_, _032_, _031_, _030_, _029_, _028_, _027_ });
assign _027_ = ap_CS_fsm == 8'h80;
assign _028_ = ap_CS_fsm == 7'h40;
assign _029_ = ap_CS_fsm == 6'h20;
assign _030_ = ap_CS_fsm == 5'h10;
assign _031_ = ap_CS_fsm == 4'h8;
assign _032_ = ap_CS_fsm == 3'h4;
assign _033_ = ap_CS_fsm == 2'h2;
assign ret_fu_201_p2 = $signed(op_4) - $signed({ 1'h0, op_6 });
assign icmp_ln851_1_fu_507_p2 = _025_ ? 1'h1 : 1'h0;
assign icmp_ln851_fu_430_p2 = _022_ ? 1'h1 : 1'h0;
assign icmp_ln886_fu_245_p2 = _023_ ? 1'h1 : 1'h0;
assign op_17_V_fu_466_p2 = _024_ ? 1'h1 : 1'h0;
assign ret_V_13_fu_388_p3 = ret_V_12_reg_630[33] ? select_ln850_2_fu_382_p3 : ret_V_8_cast_reg_635;
assign ret_V_15_fu_534_p3 = ret_V_14_reg_657[36] ? select_ln850_3_fu_528_p3 : ret_V_19_cast_reg_662;
assign ret_V_5_fu_450_p3 = op_0[7] ? select_ln850_fu_442_p3 : { 2'h0, op_0[6:5] };
assign select_ln850_2_fu_382_p3 = op_12[0] ? add_ln691_reg_642 : ret_V_8_cast_reg_635;
assign select_ln850_3_fu_528_p3 = icmp_ln851_1_reg_669 ? add_ln691_1_fu_523_p2 : ret_V_19_cast_reg_662;
assign select_ln850_4_fu_272_p3 = op_2[0] ? ret_V_2_reg_605 : ret_V_reg_599;
assign select_ln850_5_fu_278_p3 = ret_V_11_reg_594[5] ? select_ln850_4_fu_272_p3 : ret_V_reg_599;
assign select_ln850_fu_442_p3 = icmp_ln851_fu_430_p2 ? { 2'h3, op_0[6:5] } : ret_V_4_fu_436_p2;
assign ap_CS_fsm_state1 = ap_CS_fsm[0];
assign ap_CS_fsm_state2 = ap_CS_fsm[1];
assign ap_CS_fsm_state3 = ap_CS_fsm[2];
assign ap_CS_fsm_state4 = ap_CS_fsm[3];
assign ap_CS_fsm_state5 = ap_CS_fsm[4];
assign ap_CS_fsm_state6 = ap_CS_fsm[5];
assign ap_CS_fsm_state7 = ap_CS_fsm[6];
assign ap_CS_fsm_state8 = ap_CS_fsm[7];
assign ap_ready = ap_done;
assign icmp_ln886_fu_245_p0 = op_4;
assign op_31_ap_vld = ap_done;
assign op_9_V_fu_251_p3 = { ret_reg_589, 6'h00 };
assign p_Result_1_fu_418_p3 = op_0[7];
assign p_Result_2_fu_372_p3 = ret_V_12_reg_630[33];
assign p_Result_3_fu_516_p3 = ret_V_14_reg_657[36];
assign p_Result_s_fu_258_p3 = ret_V_11_reg_594[5];
assign ret_V_12_fu_351_p2[32:13] = { ret_V_12_fu_351_p2[33], ret_V_12_fu_351_p2[33], ret_V_12_fu_351_p2[33], ret_V_12_fu_351_p2[33], ret_V_12_fu_351_p2[33], ret_V_12_fu_351_p2[33], ret_V_12_fu_351_p2[33], ret_V_12_fu_351_p2[33], ret_V_12_fu_351_p2[33], ret_V_12_fu_351_p2[33], ret_V_12_fu_351_p2[33], ret_V_12_fu_351_p2[33], ret_V_12_fu_351_p2[33], ret_V_12_fu_351_p2[33], ret_V_12_fu_351_p2[33], ret_V_12_fu_351_p2[33], ret_V_12_fu_351_p2[33], ret_V_12_fu_351_p2[33], ret_V_12_fu_351_p2[33], ret_V_12_fu_351_p2[33] };
assign ret_V_3_fu_404_p4 = op_0[7:5];
assign ret_V_fu_229_p4 = ret_V_11_fu_223_p2[5:1];
assign rhs_1_fu_285_p3 = { select_ln850_5_fu_278_p3, 6'h00 };
assign rhs_4_fu_476_p3 = { op_25_V_reg_647, 4'h0 };
assign rhs_fu_211_p3 = { op_8, 1'h0 };
assign sext_ln1192_1_fu_268_p1 = { ret_reg_589[9], ret_reg_589, 6'h00 };
assign sext_ln1192_2_fu_293_p1 = { select_ln850_5_fu_278_p3[4], select_ln850_5_fu_278_p3[4], select_ln850_5_fu_278_p3[4], select_ln850_5_fu_278_p3[4], select_ln850_5_fu_278_p3[4], select_ln850_5_fu_278_p3[4], select_ln850_5_fu_278_p3, 6'h00 };
assign sext_ln1192_3_fu_347_p1 = { op_23_V_fu_329_p2[11], op_23_V_fu_329_p2[11], op_23_V_fu_329_p2[11], op_23_V_fu_329_p2[11], op_23_V_fu_329_p2[11], op_23_V_fu_329_p2[11], op_23_V_fu_329_p2[11], op_23_V_fu_329_p2[11], op_23_V_fu_329_p2[11], op_23_V_fu_329_p2[11], op_23_V_fu_329_p2[11], op_23_V_fu_329_p2[11], op_23_V_fu_329_p2[11], op_23_V_fu_329_p2[11], op_23_V_fu_329_p2[11], op_23_V_fu_329_p2[11], op_23_V_fu_329_p2[11], op_23_V_fu_329_p2[11], op_23_V_fu_329_p2[11], op_23_V_fu_329_p2[11], op_23_V_fu_329_p2[11], op_23_V_fu_329_p2, 1'h0 };
assign sext_ln1192_4_fu_483_p1 = { op_25_V_reg_647[31], op_25_V_reg_647, 4'h0 };
assign sext_ln1192_fu_219_p1 = { op_8[3], op_8, 1'h0 };
assign sext_ln20_fu_323_p1 = { op_21_V_reg_615[10], op_21_V_reg_615 };
assign sext_ln215_fu_193_p0 = op_4;
assign sext_ln215_fu_193_p1 = { op_4[7], op_4[7], op_4 };
assign sext_ln703_1_fu_335_p0 = op_12;
assign sext_ln703_1_fu_335_p1 = { op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12 };
assign sext_ln703_2_fu_472_p0 = op_14;
assign sext_ln703_2_fu_472_p1 = { op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14 };
assign sext_ln703_fu_207_p0 = op_2;
assign sext_ln703_fu_207_p1 = { op_2[3], op_2[3], op_2 };
assign sext_ln835_fu_414_p1 = { op_0[7], op_0[7:5] };
assign sext_ln886_fu_458_p1 = { ret_V_5_fu_450_p3[3], ret_V_5_fu_450_p3[3], ret_V_5_fu_450_p3[3], ret_V_5_fu_450_p3[3], ret_V_5_fu_450_p3[3], ret_V_5_fu_450_p3 };
assign tmp_3_fu_339_p3 = { op_23_V_fu_329_p2, 1'h0 };
assign trunc_ln851_1_fu_426_p1 = op_0[4:0];
assign trunc_ln851_2_fu_379_p0 = op_12;
assign trunc_ln851_2_fu_379_p1 = op_12[0];
assign trunc_ln851_3_fu_503_p0 = op_14;
assign trunc_ln851_3_fu_503_p1 = op_14[3:0];
assign trunc_ln851_fu_265_p0 = op_2;
assign trunc_ln851_fu_265_p1 = op_2[0];
assign zext_ln17_fu_513_p1 = { 1'h0, op_17_V_reg_652 };
assign zext_ln215_fu_197_p1 = { 2'h0, op_6 };
assign zext_ln69_1_fu_395_p1 = { 31'h00000000, icmp_ln886_reg_610 };
assign zext_ln69_2_fu_565_p1 = { 24'h000000, op_15 };
assign zext_ln69_3_fu_326_p1 = { 3'h0, add_ln69_reg_620 };
assign zext_ln69_4_fu_541_p1 = { 1'h0, op_16 };
assign zext_ln69_5_fu_545_p1 = { 1'h0, op_18 };
assign zext_ln69_6_fu_555_p1 = { 3'h0, add_ln69_4_fu_549_p2 };
assign zext_ln69_7_fu_574_p1 = { 27'h0000000, add_ln69_5_reg_679 };
assign zext_ln69_fu_313_p1 = { 1'h0, op_10 };
assign zext_ln886_fu_462_p1 = { 1'h0, op_7 };
endmodule


// Machine B:
// Processed by function `add_clk_enable_signal` in `verilog_tricks.py`.
// Processed by function `remove_reset_signal` in `verilog_tricks.py`.
module top_B (
  ap_clk,
  ap_start,
  ap_done,
  ap_idle,
  ap_ready,
  op_0,
  op_2,
  op_4,
  op_6,
  op_7,
  op_8,
  op_10,
  op_12,
  op_14,
  op_15,
  op_16,
  op_18,
  op_31,
  op_31_ap_vld,
clk_enable
);
input clk_enable;


input ap_clk;
wire ap_rst;
assign ap_rst = op_31_ap_vld;
input ap_start;
input [7:0] op_0;
input [7:0] op_10;
input [1:0] op_12;
input [7:0] op_14;
input [7:0] op_15;
input op_16;
input [3:0] op_18;
input [3:0] op_2;
input [7:0] op_4;
input [7:0] op_6;
input [7:0] op_7;
input [3:0] op_8;
output ap_done;
output ap_idle;
output ap_ready;
output [31:0] op_31;
output op_31_ap_vld;


reg [5:0] \add_12ns_12s_12_2_1_U6.top_add_12ns_12s_12_2_1_Adder_5_U.ain_s1 ;
reg [5:0] \add_12ns_12s_12_2_1_U6.top_add_12ns_12s_12_2_1_Adder_5_U.bin_s1 ;
reg \add_12ns_12s_12_2_1_U6.top_add_12ns_12s_12_2_1_Adder_5_U.carry_s1 ;
reg [5:0] \add_12ns_12s_12_2_1_U6.top_add_12ns_12s_12_2_1_Adder_5_U.sum_s1 ;
reg [8:0] \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.ain_s1 ;
reg [8:0] \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.bin_s1 ;
reg \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.carry_s1 ;
reg [7:0] \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.sum_s1 ;
reg \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_10_U.ain_s1 ;
reg \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_10_U.bin_s1 ;
reg \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_10_U.carry_s1 ;
reg \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_10_U.sum_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s1 ;
reg \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.carry_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.sum_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s1 ;
reg \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.carry_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.sum_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s1 ;
reg \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.carry_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.sum_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s1 ;
reg \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_7_U.carry_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_7_U.sum_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s1 ;
reg \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.carry_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.sum_s1 ;
reg [16:0] \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_6_U.ain_s1 ;
reg [16:0] \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_6_U.bin_s1 ;
reg \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_6_U.carry_s1 ;
reg [16:0] \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_6_U.sum_s1 ;
reg [18:0] \add_37s_37s_37_2_1_U11.top_add_37s_37s_37_2_1_Adder_9_U.ain_s1 ;
reg [18:0] \add_37s_37s_37_2_1_U11.top_add_37s_37s_37_2_1_Adder_9_U.bin_s1 ;
reg \add_37s_37s_37_2_1_U11.top_add_37s_37s_37_2_1_Adder_9_U.carry_s1 ;
reg [17:0] \add_37s_37s_37_2_1_U11.top_add_37s_37s_37_2_1_Adder_9_U.sum_s1 ;
reg [1:0] \add_4s_4ns_4_2_1_U10.top_add_4s_4ns_4_2_1_Adder_8_U.ain_s1 ;
reg [1:0] \add_4s_4ns_4_2_1_U10.top_add_4s_4ns_4_2_1_Adder_8_U.bin_s1 ;
reg \add_4s_4ns_4_2_1_U10.top_add_4s_4ns_4_2_1_Adder_8_U.carry_s1 ;
reg [1:0] \add_4s_4ns_4_2_1_U10.top_add_4s_4ns_4_2_1_Adder_8_U.sum_s1 ;
reg [2:0] \add_5ns_5ns_5_2_1_U15.top_add_5ns_5ns_5_2_1_Adder_1_U.ain_s1 ;
reg [2:0] \add_5ns_5ns_5_2_1_U15.top_add_5ns_5ns_5_2_1_Adder_1_U.bin_s1 ;
reg \add_5ns_5ns_5_2_1_U15.top_add_5ns_5ns_5_2_1_Adder_1_U.carry_s1 ;
reg [1:0] \add_5ns_5ns_5_2_1_U15.top_add_5ns_5ns_5_2_1_Adder_1_U.sum_s1 ;
reg [2:0] \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.ain_s1 ;
reg [2:0] \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.bin_s1 ;
reg \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.carry_s1 ;
reg [1:0] \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.sum_s1 ;
reg [2:0] \add_6s_6s_6_2_1_U1.top_add_6s_6s_6_2_1_Adder_0_U.ain_s1 ;
reg [2:0] \add_6s_6s_6_2_1_U1.top_add_6s_6s_6_2_1_Adder_0_U.bin_s1 ;
reg \add_6s_6s_6_2_1_U1.top_add_6s_6s_6_2_1_Adder_0_U.carry_s1 ;
reg [2:0] \add_6s_6s_6_2_1_U1.top_add_6s_6s_6_2_1_Adder_0_U.sum_s1 ;
reg [4:0] \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.ain_s1 ;
reg [4:0] \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.bin_s1 ;
reg \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.carry_s1 ;
reg [3:0] \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.sum_s1 ;
reg [31:0] add_ln691_1_reg_775;
reg [31:0] add_ln691_reg_696;
reg [31:0] add_ln69_3_reg_810;
reg [1:0] add_ln69_4_reg_790;
reg [4:0] add_ln69_5_reg_815;
reg [8:0] add_ln69_reg_649;
reg [24:0] ap_CS_fsm = 25'h0000001;
reg icmp_ln851_1_reg_743;
reg icmp_ln851_reg_728;
reg icmp_ln886_reg_614;
reg op_17_V_reg_765;
reg [10:0] op_21_V_reg_644;
reg [11:0] op_23_V_reg_664;
reg [31:0] op_25_V_reg_711;
reg [5:0] ret_V_11_reg_587;
reg [33:0] ret_V_12_reg_684;
reg [31:0] ret_V_13_reg_701;
reg [36:0] ret_V_14_reg_753;
reg [31:0] ret_V_15_reg_785;
reg [31:0] ret_V_19_cast_reg_758;
reg [4:0] ret_V_2_reg_609;
reg [3:0] ret_V_4_reg_748;
reg [31:0] ret_V_8_cast_reg_689;
reg [4:0] ret_V_reg_592;
reg [9:0] ret_reg_619;
reg [4:0] select_ln850_5_reg_624;
reg [3:0] sext_ln835_reg_721;
reg [4:0] \sub_10s_10ns_10_2_1_U3.top_sub_10s_10ns_10_2_1_Adder_2_U.ain_s1 ;
reg [4:0] \sub_10s_10ns_10_2_1_U3.top_sub_10s_10ns_10_2_1_Adder_2_U.bin_s1 ;
reg \sub_10s_10ns_10_2_1_U3.top_sub_10s_10ns_10_2_1_Adder_2_U.carry_s1 ;
reg [4:0] \sub_10s_10ns_10_2_1_U3.top_sub_10s_10ns_10_2_1_Adder_2_U.sum_s1 ;
wire [31:0] _000_;
wire [31:0] _001_;
wire [31:0] _002_;
wire [1:0] _003_;
wire [4:0] _004_;
wire [8:0] _005_;
wire [24:0] _006_;
wire _007_;
wire _008_;
wire _009_;
wire _010_;
wire [10:0] _011_;
wire [11:0] _012_;
wire [31:0] _013_;
wire [5:0] _014_;
wire [33:0] _015_;
wire [31:0] _016_;
wire [36:0] _017_;
wire [31:0] _018_;
wire [31:0] _019_;
wire [4:0] _020_;
wire [3:0] _021_;
wire [31:0] _022_;
wire [4:0] _023_;
wire [9:0] _024_;
wire [4:0] _025_;
wire [3:0] _026_;
wire [1:0] _027_;
wire _028_;
wire _029_;
wire _030_;
wire _031_;
wire _032_;
wire [5:0] _033_;
wire [5:0] _034_;
wire _035_;
wire [5:0] _036_;
wire [6:0] _037_;
wire [6:0] _038_;
wire [8:0] _039_;
wire [8:0] _040_;
wire _041_;
wire [7:0] _042_;
wire [8:0] _043_;
wire [9:0] _044_;
wire _045_;
wire _046_;
wire _047_;
wire _048_;
wire [1:0] _049_;
wire [1:0] _050_;
wire [15:0] _051_;
wire [15:0] _052_;
wire _053_;
wire [15:0] _054_;
wire [16:0] _055_;
wire [16:0] _056_;
wire [15:0] _057_;
wire [15:0] _058_;
wire _059_;
wire [15:0] _060_;
wire [16:0] _061_;
wire [16:0] _062_;
wire [15:0] _063_;
wire [15:0] _064_;
wire _065_;
wire [15:0] _066_;
wire [16:0] _067_;
wire [16:0] _068_;
wire [15:0] _069_;
wire [15:0] _070_;
wire _071_;
wire [15:0] _072_;
wire [16:0] _073_;
wire [16:0] _074_;
wire [15:0] _075_;
wire [15:0] _076_;
wire _077_;
wire [15:0] _078_;
wire [16:0] _079_;
wire [16:0] _080_;
wire [16:0] _081_;
wire [16:0] _082_;
wire _083_;
wire [16:0] _084_;
wire [17:0] _085_;
wire [17:0] _086_;
wire [18:0] _087_;
wire [18:0] _088_;
wire _089_;
wire [17:0] _090_;
wire [18:0] _091_;
wire [19:0] _092_;
wire [1:0] _093_;
wire [1:0] _094_;
wire _095_;
wire [1:0] _096_;
wire [2:0] _097_;
wire [2:0] _098_;
wire [2:0] _099_;
wire [2:0] _100_;
wire _101_;
wire [1:0] _102_;
wire [2:0] _103_;
wire [3:0] _104_;
wire [2:0] _105_;
wire [2:0] _106_;
wire _107_;
wire [1:0] _108_;
wire [2:0] _109_;
wire [3:0] _110_;
wire [2:0] _111_;
wire [2:0] _112_;
wire _113_;
wire [2:0] _114_;
wire [3:0] _115_;
wire [3:0] _116_;
wire [4:0] _117_;
wire [4:0] _118_;
wire _119_;
wire [3:0] _120_;
wire [4:0] _121_;
wire [5:0] _122_;
wire [4:0] _123_;
wire [4:0] _124_;
wire _125_;
wire [4:0] _126_;
wire [5:0] _127_;
wire [5:0] _128_;
wire _129_;
wire _130_;
wire _131_;
wire _132_;
wire _133_;
wire _134_;
wire _135_;
wire _136_;
wire _137_;
wire _138_;
wire _139_;
wire _140_;
wire _141_;
wire _142_;
wire _143_;
wire _144_;
wire _145_;
wire _146_;
wire _147_;
wire _148_;
wire _149_;
wire _150_;
wire _151_;
wire _152_;
wire _153_;
wire _154_;
wire _155_;
wire _156_;
wire \add_12ns_12s_12_2_1_U6.ce ;
wire \add_12ns_12s_12_2_1_U6.clk ;
wire [11:0] \add_12ns_12s_12_2_1_U6.din0 ;
wire [11:0] \add_12ns_12s_12_2_1_U6.din1 ;
wire [11:0] \add_12ns_12s_12_2_1_U6.dout ;
wire \add_12ns_12s_12_2_1_U6.reset ;
wire [11:0] \add_12ns_12s_12_2_1_U6.top_add_12ns_12s_12_2_1_Adder_5_U.a ;
wire [11:0] \add_12ns_12s_12_2_1_U6.top_add_12ns_12s_12_2_1_Adder_5_U.ain_s0 ;
wire [11:0] \add_12ns_12s_12_2_1_U6.top_add_12ns_12s_12_2_1_Adder_5_U.b ;
wire [11:0] \add_12ns_12s_12_2_1_U6.top_add_12ns_12s_12_2_1_Adder_5_U.bin_s0 ;
wire \add_12ns_12s_12_2_1_U6.top_add_12ns_12s_12_2_1_Adder_5_U.ce ;
wire \add_12ns_12s_12_2_1_U6.top_add_12ns_12s_12_2_1_Adder_5_U.clk ;
wire \add_12ns_12s_12_2_1_U6.top_add_12ns_12s_12_2_1_Adder_5_U.facout_s1 ;
wire \add_12ns_12s_12_2_1_U6.top_add_12ns_12s_12_2_1_Adder_5_U.facout_s2 ;
wire [5:0] \add_12ns_12s_12_2_1_U6.top_add_12ns_12s_12_2_1_Adder_5_U.fas_s1 ;
wire [5:0] \add_12ns_12s_12_2_1_U6.top_add_12ns_12s_12_2_1_Adder_5_U.fas_s2 ;
wire \add_12ns_12s_12_2_1_U6.top_add_12ns_12s_12_2_1_Adder_5_U.reset ;
wire [11:0] \add_12ns_12s_12_2_1_U6.top_add_12ns_12s_12_2_1_Adder_5_U.s ;
wire [5:0] \add_12ns_12s_12_2_1_U6.top_add_12ns_12s_12_2_1_Adder_5_U.u1.a ;
wire [5:0] \add_12ns_12s_12_2_1_U6.top_add_12ns_12s_12_2_1_Adder_5_U.u1.b ;
wire \add_12ns_12s_12_2_1_U6.top_add_12ns_12s_12_2_1_Adder_5_U.u1.cin ;
wire \add_12ns_12s_12_2_1_U6.top_add_12ns_12s_12_2_1_Adder_5_U.u1.cout ;
wire [5:0] \add_12ns_12s_12_2_1_U6.top_add_12ns_12s_12_2_1_Adder_5_U.u1.s ;
wire [5:0] \add_12ns_12s_12_2_1_U6.top_add_12ns_12s_12_2_1_Adder_5_U.u2.a ;
wire [5:0] \add_12ns_12s_12_2_1_U6.top_add_12ns_12s_12_2_1_Adder_5_U.u2.b ;
wire \add_12ns_12s_12_2_1_U6.top_add_12ns_12s_12_2_1_Adder_5_U.u2.cin ;
wire \add_12ns_12s_12_2_1_U6.top_add_12ns_12s_12_2_1_Adder_5_U.u2.cout ;
wire [5:0] \add_12ns_12s_12_2_1_U6.top_add_12ns_12s_12_2_1_Adder_5_U.u2.s ;
wire \add_17s_17s_17_2_1_U4.ce ;
wire \add_17s_17s_17_2_1_U4.clk ;
wire [16:0] \add_17s_17s_17_2_1_U4.din0 ;
wire [16:0] \add_17s_17s_17_2_1_U4.din1 ;
wire [16:0] \add_17s_17s_17_2_1_U4.dout ;
wire \add_17s_17s_17_2_1_U4.reset ;
wire [16:0] \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.a ;
wire [16:0] \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.ain_s0 ;
wire [16:0] \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.b ;
wire [16:0] \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.bin_s0 ;
wire \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.ce ;
wire \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.clk ;
wire \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.facout_s1 ;
wire \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.facout_s2 ;
wire [7:0] \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.fas_s1 ;
wire [8:0] \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.fas_s2 ;
wire \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.reset ;
wire [16:0] \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.s ;
wire [7:0] \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.u1.a ;
wire [7:0] \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.u1.b ;
wire \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.u1.cin ;
wire \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.u1.cout ;
wire [7:0] \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.u1.s ;
wire [8:0] \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.u2.a ;
wire [8:0] \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.u2.b ;
wire \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.u2.cin ;
wire \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.u2.cout ;
wire [8:0] \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.u2.s ;
wire \add_2ns_2ns_2_2_1_U13.ce ;
wire \add_2ns_2ns_2_2_1_U13.clk ;
wire [1:0] \add_2ns_2ns_2_2_1_U13.din0 ;
wire [1:0] \add_2ns_2ns_2_2_1_U13.din1 ;
wire [1:0] \add_2ns_2ns_2_2_1_U13.dout ;
wire \add_2ns_2ns_2_2_1_U13.reset ;
wire [1:0] \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_10_U.a ;
wire [1:0] \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_10_U.ain_s0 ;
wire [1:0] \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_10_U.b ;
wire [1:0] \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_10_U.bin_s0 ;
wire \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_10_U.ce ;
wire \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_10_U.clk ;
wire \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_10_U.facout_s1 ;
wire \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_10_U.facout_s2 ;
wire \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_10_U.fas_s1 ;
wire \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_10_U.fas_s2 ;
wire \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_10_U.reset ;
wire [1:0] \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_10_U.s ;
wire \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_10_U.u1.a ;
wire \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_10_U.u1.b ;
wire \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_10_U.u1.cin ;
wire \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_10_U.u1.cout ;
wire \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_10_U.u1.s ;
wire \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_10_U.u2.a ;
wire \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_10_U.u2.b ;
wire \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_10_U.u2.cin ;
wire \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_10_U.u2.cout ;
wire \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_10_U.u2.s ;
wire \add_32ns_32ns_32_2_1_U12.ce ;
wire \add_32ns_32ns_32_2_1_U12.clk ;
wire [31:0] \add_32ns_32ns_32_2_1_U12.din0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U12.din1 ;
wire [31:0] \add_32ns_32ns_32_2_1_U12.dout ;
wire \add_32ns_32ns_32_2_1_U12.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.a ;
wire [31:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.b ;
wire [31:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s0 ;
wire \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.ce ;
wire \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.clk ;
wire \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.facout_s1 ;
wire \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.facout_s2 ;
wire [15:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s1 ;
wire [15:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s2 ;
wire \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.b ;
wire \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cin ;
wire \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.b ;
wire \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cin ;
wire \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.s ;
wire \add_32ns_32ns_32_2_1_U14.ce ;
wire \add_32ns_32ns_32_2_1_U14.clk ;
wire [31:0] \add_32ns_32ns_32_2_1_U14.din0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U14.din1 ;
wire [31:0] \add_32ns_32ns_32_2_1_U14.dout ;
wire \add_32ns_32ns_32_2_1_U14.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.a ;
wire [31:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.b ;
wire [31:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s0 ;
wire \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.ce ;
wire \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.clk ;
wire \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.facout_s1 ;
wire \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.facout_s2 ;
wire [15:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s1 ;
wire [15:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s2 ;
wire \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.b ;
wire \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cin ;
wire \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.b ;
wire \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cin ;
wire \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.s ;
wire \add_32ns_32ns_32_2_1_U16.ce ;
wire \add_32ns_32ns_32_2_1_U16.clk ;
wire [31:0] \add_32ns_32ns_32_2_1_U16.din0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U16.din1 ;
wire [31:0] \add_32ns_32ns_32_2_1_U16.dout ;
wire \add_32ns_32ns_32_2_1_U16.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.a ;
wire [31:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.b ;
wire [31:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s0 ;
wire \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.ce ;
wire \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.clk ;
wire \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.facout_s1 ;
wire \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.facout_s2 ;
wire [15:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s1 ;
wire [15:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s2 ;
wire \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.b ;
wire \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cin ;
wire \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.b ;
wire \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cin ;
wire \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.s ;
wire \add_32ns_32ns_32_2_1_U8.ce ;
wire \add_32ns_32ns_32_2_1_U8.clk ;
wire [31:0] \add_32ns_32ns_32_2_1_U8.din0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U8.din1 ;
wire [31:0] \add_32ns_32ns_32_2_1_U8.dout ;
wire \add_32ns_32ns_32_2_1_U8.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_7_U.a ;
wire [31:0] \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_7_U.b ;
wire [31:0] \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s0 ;
wire \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_7_U.ce ;
wire \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_7_U.clk ;
wire \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_7_U.facout_s1 ;
wire \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_7_U.facout_s2 ;
wire [15:0] \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s1 ;
wire [15:0] \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s2 ;
wire \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_7_U.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_7_U.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.b ;
wire \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cin ;
wire \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.b ;
wire \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cin ;
wire \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.s ;
wire \add_32ns_32ns_32_2_1_U9.ce ;
wire \add_32ns_32ns_32_2_1_U9.clk ;
wire [31:0] \add_32ns_32ns_32_2_1_U9.din0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U9.din1 ;
wire [31:0] \add_32ns_32ns_32_2_1_U9.dout ;
wire \add_32ns_32ns_32_2_1_U9.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.a ;
wire [31:0] \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.b ;
wire [31:0] \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s0 ;
wire \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.ce ;
wire \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.clk ;
wire \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.facout_s1 ;
wire \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.facout_s2 ;
wire [15:0] \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s1 ;
wire [15:0] \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s2 ;
wire \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.b ;
wire \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cin ;
wire \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.b ;
wire \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cin ;
wire \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.s ;
wire \add_34s_34s_34_2_1_U7.ce ;
wire \add_34s_34s_34_2_1_U7.clk ;
wire [33:0] \add_34s_34s_34_2_1_U7.din0 ;
wire [33:0] \add_34s_34s_34_2_1_U7.din1 ;
wire [33:0] \add_34s_34s_34_2_1_U7.dout ;
wire \add_34s_34s_34_2_1_U7.reset ;
wire [33:0] \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_6_U.a ;
wire [33:0] \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_6_U.ain_s0 ;
wire [33:0] \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_6_U.b ;
wire [33:0] \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_6_U.bin_s0 ;
wire \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_6_U.ce ;
wire \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_6_U.clk ;
wire \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_6_U.facout_s1 ;
wire \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_6_U.facout_s2 ;
wire [16:0] \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_6_U.fas_s1 ;
wire [16:0] \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_6_U.fas_s2 ;
wire \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_6_U.reset ;
wire [33:0] \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_6_U.s ;
wire [16:0] \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_6_U.u1.a ;
wire [16:0] \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_6_U.u1.b ;
wire \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_6_U.u1.cin ;
wire \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_6_U.u1.cout ;
wire [16:0] \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_6_U.u1.s ;
wire [16:0] \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_6_U.u2.a ;
wire [16:0] \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_6_U.u2.b ;
wire \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_6_U.u2.cin ;
wire \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_6_U.u2.cout ;
wire [16:0] \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_6_U.u2.s ;
wire \add_37s_37s_37_2_1_U11.ce ;
wire \add_37s_37s_37_2_1_U11.clk ;
wire [36:0] \add_37s_37s_37_2_1_U11.din0 ;
wire [36:0] \add_37s_37s_37_2_1_U11.din1 ;
wire [36:0] \add_37s_37s_37_2_1_U11.dout ;
wire \add_37s_37s_37_2_1_U11.reset ;
wire [36:0] \add_37s_37s_37_2_1_U11.top_add_37s_37s_37_2_1_Adder_9_U.a ;
wire [36:0] \add_37s_37s_37_2_1_U11.top_add_37s_37s_37_2_1_Adder_9_U.ain_s0 ;
wire [36:0] \add_37s_37s_37_2_1_U11.top_add_37s_37s_37_2_1_Adder_9_U.b ;
wire [36:0] \add_37s_37s_37_2_1_U11.top_add_37s_37s_37_2_1_Adder_9_U.bin_s0 ;
wire \add_37s_37s_37_2_1_U11.top_add_37s_37s_37_2_1_Adder_9_U.ce ;
wire \add_37s_37s_37_2_1_U11.top_add_37s_37s_37_2_1_Adder_9_U.clk ;
wire \add_37s_37s_37_2_1_U11.top_add_37s_37s_37_2_1_Adder_9_U.facout_s1 ;
wire \add_37s_37s_37_2_1_U11.top_add_37s_37s_37_2_1_Adder_9_U.facout_s2 ;
wire [17:0] \add_37s_37s_37_2_1_U11.top_add_37s_37s_37_2_1_Adder_9_U.fas_s1 ;
wire [18:0] \add_37s_37s_37_2_1_U11.top_add_37s_37s_37_2_1_Adder_9_U.fas_s2 ;
wire \add_37s_37s_37_2_1_U11.top_add_37s_37s_37_2_1_Adder_9_U.reset ;
wire [36:0] \add_37s_37s_37_2_1_U11.top_add_37s_37s_37_2_1_Adder_9_U.s ;
wire [17:0] \add_37s_37s_37_2_1_U11.top_add_37s_37s_37_2_1_Adder_9_U.u1.a ;
wire [17:0] \add_37s_37s_37_2_1_U11.top_add_37s_37s_37_2_1_Adder_9_U.u1.b ;
wire \add_37s_37s_37_2_1_U11.top_add_37s_37s_37_2_1_Adder_9_U.u1.cin ;
wire \add_37s_37s_37_2_1_U11.top_add_37s_37s_37_2_1_Adder_9_U.u1.cout ;
wire [17:0] \add_37s_37s_37_2_1_U11.top_add_37s_37s_37_2_1_Adder_9_U.u1.s ;
wire [18:0] \add_37s_37s_37_2_1_U11.top_add_37s_37s_37_2_1_Adder_9_U.u2.a ;
wire [18:0] \add_37s_37s_37_2_1_U11.top_add_37s_37s_37_2_1_Adder_9_U.u2.b ;
wire \add_37s_37s_37_2_1_U11.top_add_37s_37s_37_2_1_Adder_9_U.u2.cin ;
wire \add_37s_37s_37_2_1_U11.top_add_37s_37s_37_2_1_Adder_9_U.u2.cout ;
wire [18:0] \add_37s_37s_37_2_1_U11.top_add_37s_37s_37_2_1_Adder_9_U.u2.s ;
wire \add_4s_4ns_4_2_1_U10.ce ;
wire \add_4s_4ns_4_2_1_U10.clk ;
wire [3:0] \add_4s_4ns_4_2_1_U10.din0 ;
wire [3:0] \add_4s_4ns_4_2_1_U10.din1 ;
wire [3:0] \add_4s_4ns_4_2_1_U10.dout ;
wire \add_4s_4ns_4_2_1_U10.reset ;
wire [3:0] \add_4s_4ns_4_2_1_U10.top_add_4s_4ns_4_2_1_Adder_8_U.a ;
wire [3:0] \add_4s_4ns_4_2_1_U10.top_add_4s_4ns_4_2_1_Adder_8_U.ain_s0 ;
wire [3:0] \add_4s_4ns_4_2_1_U10.top_add_4s_4ns_4_2_1_Adder_8_U.b ;
wire [3:0] \add_4s_4ns_4_2_1_U10.top_add_4s_4ns_4_2_1_Adder_8_U.bin_s0 ;
wire \add_4s_4ns_4_2_1_U10.top_add_4s_4ns_4_2_1_Adder_8_U.ce ;
wire \add_4s_4ns_4_2_1_U10.top_add_4s_4ns_4_2_1_Adder_8_U.clk ;
wire \add_4s_4ns_4_2_1_U10.top_add_4s_4ns_4_2_1_Adder_8_U.facout_s1 ;
wire \add_4s_4ns_4_2_1_U10.top_add_4s_4ns_4_2_1_Adder_8_U.facout_s2 ;
wire [1:0] \add_4s_4ns_4_2_1_U10.top_add_4s_4ns_4_2_1_Adder_8_U.fas_s1 ;
wire [1:0] \add_4s_4ns_4_2_1_U10.top_add_4s_4ns_4_2_1_Adder_8_U.fas_s2 ;
wire \add_4s_4ns_4_2_1_U10.top_add_4s_4ns_4_2_1_Adder_8_U.reset ;
wire [3:0] \add_4s_4ns_4_2_1_U10.top_add_4s_4ns_4_2_1_Adder_8_U.s ;
wire [1:0] \add_4s_4ns_4_2_1_U10.top_add_4s_4ns_4_2_1_Adder_8_U.u1.a ;
wire [1:0] \add_4s_4ns_4_2_1_U10.top_add_4s_4ns_4_2_1_Adder_8_U.u1.b ;
wire \add_4s_4ns_4_2_1_U10.top_add_4s_4ns_4_2_1_Adder_8_U.u1.cin ;
wire \add_4s_4ns_4_2_1_U10.top_add_4s_4ns_4_2_1_Adder_8_U.u1.cout ;
wire [1:0] \add_4s_4ns_4_2_1_U10.top_add_4s_4ns_4_2_1_Adder_8_U.u1.s ;
wire [1:0] \add_4s_4ns_4_2_1_U10.top_add_4s_4ns_4_2_1_Adder_8_U.u2.a ;
wire [1:0] \add_4s_4ns_4_2_1_U10.top_add_4s_4ns_4_2_1_Adder_8_U.u2.b ;
wire \add_4s_4ns_4_2_1_U10.top_add_4s_4ns_4_2_1_Adder_8_U.u2.cin ;
wire \add_4s_4ns_4_2_1_U10.top_add_4s_4ns_4_2_1_Adder_8_U.u2.cout ;
wire [1:0] \add_4s_4ns_4_2_1_U10.top_add_4s_4ns_4_2_1_Adder_8_U.u2.s ;
wire \add_5ns_5ns_5_2_1_U15.ce ;
wire \add_5ns_5ns_5_2_1_U15.clk ;
wire [4:0] \add_5ns_5ns_5_2_1_U15.din0 ;
wire [4:0] \add_5ns_5ns_5_2_1_U15.din1 ;
wire [4:0] \add_5ns_5ns_5_2_1_U15.dout ;
wire \add_5ns_5ns_5_2_1_U15.reset ;
wire [4:0] \add_5ns_5ns_5_2_1_U15.top_add_5ns_5ns_5_2_1_Adder_1_U.a ;
wire [4:0] \add_5ns_5ns_5_2_1_U15.top_add_5ns_5ns_5_2_1_Adder_1_U.ain_s0 ;
wire [4:0] \add_5ns_5ns_5_2_1_U15.top_add_5ns_5ns_5_2_1_Adder_1_U.b ;
wire [4:0] \add_5ns_5ns_5_2_1_U15.top_add_5ns_5ns_5_2_1_Adder_1_U.bin_s0 ;
wire \add_5ns_5ns_5_2_1_U15.top_add_5ns_5ns_5_2_1_Adder_1_U.ce ;
wire \add_5ns_5ns_5_2_1_U15.top_add_5ns_5ns_5_2_1_Adder_1_U.clk ;
wire \add_5ns_5ns_5_2_1_U15.top_add_5ns_5ns_5_2_1_Adder_1_U.facout_s1 ;
wire \add_5ns_5ns_5_2_1_U15.top_add_5ns_5ns_5_2_1_Adder_1_U.facout_s2 ;
wire [1:0] \add_5ns_5ns_5_2_1_U15.top_add_5ns_5ns_5_2_1_Adder_1_U.fas_s1 ;
wire [2:0] \add_5ns_5ns_5_2_1_U15.top_add_5ns_5ns_5_2_1_Adder_1_U.fas_s2 ;
wire \add_5ns_5ns_5_2_1_U15.top_add_5ns_5ns_5_2_1_Adder_1_U.reset ;
wire [4:0] \add_5ns_5ns_5_2_1_U15.top_add_5ns_5ns_5_2_1_Adder_1_U.s ;
wire [1:0] \add_5ns_5ns_5_2_1_U15.top_add_5ns_5ns_5_2_1_Adder_1_U.u1.a ;
wire [1:0] \add_5ns_5ns_5_2_1_U15.top_add_5ns_5ns_5_2_1_Adder_1_U.u1.b ;
wire \add_5ns_5ns_5_2_1_U15.top_add_5ns_5ns_5_2_1_Adder_1_U.u1.cin ;
wire \add_5ns_5ns_5_2_1_U15.top_add_5ns_5ns_5_2_1_Adder_1_U.u1.cout ;
wire [1:0] \add_5ns_5ns_5_2_1_U15.top_add_5ns_5ns_5_2_1_Adder_1_U.u1.s ;
wire [2:0] \add_5ns_5ns_5_2_1_U15.top_add_5ns_5ns_5_2_1_Adder_1_U.u2.a ;
wire [2:0] \add_5ns_5ns_5_2_1_U15.top_add_5ns_5ns_5_2_1_Adder_1_U.u2.b ;
wire \add_5ns_5ns_5_2_1_U15.top_add_5ns_5ns_5_2_1_Adder_1_U.u2.cin ;
wire \add_5ns_5ns_5_2_1_U15.top_add_5ns_5ns_5_2_1_Adder_1_U.u2.cout ;
wire [2:0] \add_5ns_5ns_5_2_1_U15.top_add_5ns_5ns_5_2_1_Adder_1_U.u2.s ;
wire \add_5ns_5ns_5_2_1_U2.ce ;
wire \add_5ns_5ns_5_2_1_U2.clk ;
wire [4:0] \add_5ns_5ns_5_2_1_U2.din0 ;
wire [4:0] \add_5ns_5ns_5_2_1_U2.din1 ;
wire [4:0] \add_5ns_5ns_5_2_1_U2.dout ;
wire \add_5ns_5ns_5_2_1_U2.reset ;
wire [4:0] \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.a ;
wire [4:0] \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.ain_s0 ;
wire [4:0] \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.b ;
wire [4:0] \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.bin_s0 ;
wire \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.ce ;
wire \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.clk ;
wire \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.facout_s1 ;
wire \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.facout_s2 ;
wire [1:0] \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.fas_s1 ;
wire [2:0] \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.fas_s2 ;
wire \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.reset ;
wire [4:0] \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.s ;
wire [1:0] \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.u1.a ;
wire [1:0] \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.u1.b ;
wire \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.u1.cin ;
wire \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.u1.cout ;
wire [1:0] \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.u1.s ;
wire [2:0] \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.u2.a ;
wire [2:0] \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.u2.b ;
wire \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.u2.cin ;
wire \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.u2.cout ;
wire [2:0] \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.u2.s ;
wire \add_6s_6s_6_2_1_U1.ce ;
wire \add_6s_6s_6_2_1_U1.clk ;
wire [5:0] \add_6s_6s_6_2_1_U1.din0 ;
wire [5:0] \add_6s_6s_6_2_1_U1.din1 ;
wire [5:0] \add_6s_6s_6_2_1_U1.dout ;
wire \add_6s_6s_6_2_1_U1.reset ;
wire [5:0] \add_6s_6s_6_2_1_U1.top_add_6s_6s_6_2_1_Adder_0_U.a ;
wire [5:0] \add_6s_6s_6_2_1_U1.top_add_6s_6s_6_2_1_Adder_0_U.ain_s0 ;
wire [5:0] \add_6s_6s_6_2_1_U1.top_add_6s_6s_6_2_1_Adder_0_U.b ;
wire [5:0] \add_6s_6s_6_2_1_U1.top_add_6s_6s_6_2_1_Adder_0_U.bin_s0 ;
wire \add_6s_6s_6_2_1_U1.top_add_6s_6s_6_2_1_Adder_0_U.ce ;
wire \add_6s_6s_6_2_1_U1.top_add_6s_6s_6_2_1_Adder_0_U.clk ;
wire \add_6s_6s_6_2_1_U1.top_add_6s_6s_6_2_1_Adder_0_U.facout_s1 ;
wire \add_6s_6s_6_2_1_U1.top_add_6s_6s_6_2_1_Adder_0_U.facout_s2 ;
wire [2:0] \add_6s_6s_6_2_1_U1.top_add_6s_6s_6_2_1_Adder_0_U.fas_s1 ;
wire [2:0] \add_6s_6s_6_2_1_U1.top_add_6s_6s_6_2_1_Adder_0_U.fas_s2 ;
wire \add_6s_6s_6_2_1_U1.top_add_6s_6s_6_2_1_Adder_0_U.reset ;
wire [5:0] \add_6s_6s_6_2_1_U1.top_add_6s_6s_6_2_1_Adder_0_U.s ;
wire [2:0] \add_6s_6s_6_2_1_U1.top_add_6s_6s_6_2_1_Adder_0_U.u1.a ;
wire [2:0] \add_6s_6s_6_2_1_U1.top_add_6s_6s_6_2_1_Adder_0_U.u1.b ;
wire \add_6s_6s_6_2_1_U1.top_add_6s_6s_6_2_1_Adder_0_U.u1.cin ;
wire \add_6s_6s_6_2_1_U1.top_add_6s_6s_6_2_1_Adder_0_U.u1.cout ;
wire [2:0] \add_6s_6s_6_2_1_U1.top_add_6s_6s_6_2_1_Adder_0_U.u1.s ;
wire [2:0] \add_6s_6s_6_2_1_U1.top_add_6s_6s_6_2_1_Adder_0_U.u2.a ;
wire [2:0] \add_6s_6s_6_2_1_U1.top_add_6s_6s_6_2_1_Adder_0_U.u2.b ;
wire \add_6s_6s_6_2_1_U1.top_add_6s_6s_6_2_1_Adder_0_U.u2.cin ;
wire \add_6s_6s_6_2_1_U1.top_add_6s_6s_6_2_1_Adder_0_U.u2.cout ;
wire [2:0] \add_6s_6s_6_2_1_U1.top_add_6s_6s_6_2_1_Adder_0_U.u2.s ;
wire \add_9ns_9ns_9_2_1_U5.ce ;
wire \add_9ns_9ns_9_2_1_U5.clk ;
wire [8:0] \add_9ns_9ns_9_2_1_U5.din0 ;
wire [8:0] \add_9ns_9ns_9_2_1_U5.din1 ;
wire [8:0] \add_9ns_9ns_9_2_1_U5.dout ;
wire \add_9ns_9ns_9_2_1_U5.reset ;
wire [8:0] \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.a ;
wire [8:0] \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.ain_s0 ;
wire [8:0] \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.b ;
wire [8:0] \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.bin_s0 ;
wire \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.ce ;
wire \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.clk ;
wire \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.facout_s1 ;
wire \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.facout_s2 ;
wire [3:0] \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.fas_s1 ;
wire [4:0] \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.fas_s2 ;
wire \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.reset ;
wire [8:0] \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.s ;
wire [3:0] \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.u1.a ;
wire [3:0] \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.u1.b ;
wire \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.u1.cin ;
wire \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.u1.cout ;
wire [3:0] \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.u1.s ;
wire [4:0] \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.u2.a ;
wire [4:0] \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.u2.b ;
wire \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.u2.cin ;
wire \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.u2.cout ;
wire [4:0] \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.u2.s ;
wire ap_CS_fsm_state1;
wire ap_CS_fsm_state10;
wire ap_CS_fsm_state11;
wire ap_CS_fsm_state12;
wire ap_CS_fsm_state13;
wire ap_CS_fsm_state14;
wire ap_CS_fsm_state15;
wire ap_CS_fsm_state16;
wire ap_CS_fsm_state17;
wire ap_CS_fsm_state18;
wire ap_CS_fsm_state19;
wire ap_CS_fsm_state2;
wire ap_CS_fsm_state20;
wire ap_CS_fsm_state21;
wire ap_CS_fsm_state22;
wire ap_CS_fsm_state23;
wire ap_CS_fsm_state24;
wire ap_CS_fsm_state25;
wire ap_CS_fsm_state3;
wire ap_CS_fsm_state4;
wire ap_CS_fsm_state5;
wire ap_CS_fsm_state6;
wire ap_CS_fsm_state7;
wire ap_CS_fsm_state8;
wire ap_CS_fsm_state9;
wire [24:0] ap_NS_fsm;
wire ap_clk;
wire ap_done;
wire ap_idle;
wire ap_ready;
wire ap_rst;
wire ap_start;
wire [5:0] grp_fu_209_p0;
wire [5:0] grp_fu_209_p1;
wire [5:0] grp_fu_209_p2;
wire [4:0] grp_fu_225_p2;
wire [9:0] grp_fu_238_p0;
wire [9:0] grp_fu_238_p1;
wire [9:0] grp_fu_238_p2;
wire [16:0] grp_fu_295_p0;
wire [16:0] grp_fu_295_p1;
wire [16:0] grp_fu_295_p2;
wire [8:0] grp_fu_305_p0;
wire [8:0] grp_fu_305_p2;
wire [11:0] grp_fu_327_p0;
wire [11:0] grp_fu_327_p1;
wire [11:0] grp_fu_327_p2;
wire [33:0] grp_fu_348_p0;
wire [33:0] grp_fu_348_p1;
wire [33:0] grp_fu_348_p2;
wire [31:0] grp_fu_364_p2;
wire [31:0] grp_fu_395_p1;
wire [31:0] grp_fu_395_p2;
wire [3:0] grp_fu_424_p0;
wire [3:0] grp_fu_424_p2;
wire [36:0] grp_fu_445_p0;
wire [36:0] grp_fu_445_p1;
wire [36:0] grp_fu_445_p2;
wire [31:0] grp_fu_504_p2;
wire [1:0] grp_fu_516_p0;
wire [1:0] grp_fu_516_p1;
wire [1:0] grp_fu_516_p2;
wire [31:0] grp_fu_549_p1;
wire [31:0] grp_fu_549_p2;
wire [4:0] grp_fu_557_p0;
wire [4:0] grp_fu_557_p1;
wire [4:0] grp_fu_557_p2;
wire [31:0] grp_fu_566_p0;
wire [31:0] grp_fu_566_p2;
wire icmp_ln851_1_fu_455_p2;
wire icmp_ln851_fu_418_p2;
wire [7:0] icmp_ln886_fu_244_p0;
wire icmp_ln886_fu_244_p2;
wire [7:0] op_0;
wire [7:0] op_10;
wire [1:0] op_12;
wire [7:0] op_14;
wire [7:0] op_15;
wire op_16;
wire op_17_V_fu_498_p2;
wire [3:0] op_18;
wire [3:0] op_2;
wire [31:0] op_31;
wire op_31_ap_vld;
wire [7:0] op_4;
wire [7:0] op_6;
wire [7:0] op_7;
wire [3:0] op_8;
wire [15:0] op_9_V_fu_273_p3;
wire p_Result_1_fu_471_p3;
wire p_Result_2_fu_369_p3;
wire p_Result_3_fu_522_p3;
wire p_Result_s_fu_250_p3;
wire [31:0] ret_V_13_fu_385_p3;
wire [31:0] ret_V_15_fu_534_p3;
wire [2:0] ret_V_3_fu_400_p4;
wire [3:0] ret_V_5_fu_483_p3;
wire [10:0] rhs_1_fu_284_p3;
wire [35:0] rhs_4_fu_434_p3;
wire [4:0] rhs_fu_197_p3;
wire [31:0] select_ln850_2_fu_379_p3;
wire [31:0] select_ln850_3_fu_529_p3;
wire [4:0] select_ln850_4_fu_260_p3;
wire [4:0] select_ln850_5_fu_266_p3;
wire [3:0] select_ln850_fu_478_p3;
wire [7:0] sext_ln215_fu_230_p0;
wire [1:0] sext_ln703_1_fu_333_p0;
wire [7:0] sext_ln703_2_fu_430_p0;
wire [3:0] sext_ln703_fu_193_p0;
wire [3:0] sext_ln835_fu_410_p1;
wire [8:0] sext_ln886_fu_490_p1;
wire \sub_10s_10ns_10_2_1_U3.ce ;
wire \sub_10s_10ns_10_2_1_U3.clk ;
wire [9:0] \sub_10s_10ns_10_2_1_U3.din0 ;
wire [9:0] \sub_10s_10ns_10_2_1_U3.din1 ;
wire [9:0] \sub_10s_10ns_10_2_1_U3.dout ;
wire \sub_10s_10ns_10_2_1_U3.reset ;
wire [9:0] \sub_10s_10ns_10_2_1_U3.top_sub_10s_10ns_10_2_1_Adder_2_U.a ;
wire [9:0] \sub_10s_10ns_10_2_1_U3.top_sub_10s_10ns_10_2_1_Adder_2_U.ain_s0 ;
wire [9:0] \sub_10s_10ns_10_2_1_U3.top_sub_10s_10ns_10_2_1_Adder_2_U.b ;
wire [9:0] \sub_10s_10ns_10_2_1_U3.top_sub_10s_10ns_10_2_1_Adder_2_U.bin_s0 ;
wire \sub_10s_10ns_10_2_1_U3.top_sub_10s_10ns_10_2_1_Adder_2_U.ce ;
wire \sub_10s_10ns_10_2_1_U3.top_sub_10s_10ns_10_2_1_Adder_2_U.clk ;
wire \sub_10s_10ns_10_2_1_U3.top_sub_10s_10ns_10_2_1_Adder_2_U.facout_s1 ;
wire \sub_10s_10ns_10_2_1_U3.top_sub_10s_10ns_10_2_1_Adder_2_U.facout_s2 ;
wire [4:0] \sub_10s_10ns_10_2_1_U3.top_sub_10s_10ns_10_2_1_Adder_2_U.fas_s1 ;
wire [4:0] \sub_10s_10ns_10_2_1_U3.top_sub_10s_10ns_10_2_1_Adder_2_U.fas_s2 ;
wire \sub_10s_10ns_10_2_1_U3.top_sub_10s_10ns_10_2_1_Adder_2_U.reset ;
wire [9:0] \sub_10s_10ns_10_2_1_U3.top_sub_10s_10ns_10_2_1_Adder_2_U.s ;
wire [4:0] \sub_10s_10ns_10_2_1_U3.top_sub_10s_10ns_10_2_1_Adder_2_U.u1.a ;
wire [4:0] \sub_10s_10ns_10_2_1_U3.top_sub_10s_10ns_10_2_1_Adder_2_U.u1.b ;
wire \sub_10s_10ns_10_2_1_U3.top_sub_10s_10ns_10_2_1_Adder_2_U.u1.cin ;
wire \sub_10s_10ns_10_2_1_U3.top_sub_10s_10ns_10_2_1_Adder_2_U.u1.cout ;
wire [4:0] \sub_10s_10ns_10_2_1_U3.top_sub_10s_10ns_10_2_1_Adder_2_U.u1.s ;
wire [4:0] \sub_10s_10ns_10_2_1_U3.top_sub_10s_10ns_10_2_1_Adder_2_U.u2.a ;
wire [4:0] \sub_10s_10ns_10_2_1_U3.top_sub_10s_10ns_10_2_1_Adder_2_U.u2.b ;
wire \sub_10s_10ns_10_2_1_U3.top_sub_10s_10ns_10_2_1_Adder_2_U.u2.cin ;
wire \sub_10s_10ns_10_2_1_U3.top_sub_10s_10ns_10_2_1_Adder_2_U.u2.cout ;
wire [4:0] \sub_10s_10ns_10_2_1_U3.top_sub_10s_10ns_10_2_1_Adder_2_U.u2.s ;
wire [12:0] tmp_3_fu_337_p3;
wire [4:0] trunc_ln851_1_fu_414_p1;
wire [1:0] trunc_ln851_2_fu_376_p0;
wire trunc_ln851_2_fu_376_p1;
wire [7:0] trunc_ln851_3_fu_451_p0;
wire [3:0] trunc_ln851_3_fu_451_p1;
wire [3:0] trunc_ln851_fu_257_p0;
wire trunc_ln851_fu_257_p1;
wire [8:0] zext_ln886_fu_494_p1;


assign _028_ = ap_CS_fsm[19] & icmp_ln851_1_reg_743;
assign _029_ = _031_ & ap_CS_fsm[0];
assign _030_ = ap_start & ap_CS_fsm[0];
assign _031_ = ~ ap_start;
assign _032_ = ! op_0[4:0];
always @(posedge \add_12ns_12s_12_2_1_U6.top_add_12ns_12s_12_2_1_Adder_5_U.clk )
\add_12ns_12s_12_2_1_U6.top_add_12ns_12s_12_2_1_Adder_5_U.bin_s1  <= _034_;
always @(posedge \add_12ns_12s_12_2_1_U6.top_add_12ns_12s_12_2_1_Adder_5_U.clk )
\add_12ns_12s_12_2_1_U6.top_add_12ns_12s_12_2_1_Adder_5_U.ain_s1  <= _033_;
always @(posedge \add_12ns_12s_12_2_1_U6.top_add_12ns_12s_12_2_1_Adder_5_U.clk )
\add_12ns_12s_12_2_1_U6.top_add_12ns_12s_12_2_1_Adder_5_U.sum_s1  <= _036_;
always @(posedge \add_12ns_12s_12_2_1_U6.top_add_12ns_12s_12_2_1_Adder_5_U.clk )
\add_12ns_12s_12_2_1_U6.top_add_12ns_12s_12_2_1_Adder_5_U.carry_s1  <= _035_;
assign _034_ = \add_12ns_12s_12_2_1_U6.top_add_12ns_12s_12_2_1_Adder_5_U.ce  ? \add_12ns_12s_12_2_1_U6.top_add_12ns_12s_12_2_1_Adder_5_U.b [11:6] : \add_12ns_12s_12_2_1_U6.top_add_12ns_12s_12_2_1_Adder_5_U.bin_s1 ;
assign _033_ = \add_12ns_12s_12_2_1_U6.top_add_12ns_12s_12_2_1_Adder_5_U.ce  ? \add_12ns_12s_12_2_1_U6.top_add_12ns_12s_12_2_1_Adder_5_U.a [11:6] : \add_12ns_12s_12_2_1_U6.top_add_12ns_12s_12_2_1_Adder_5_U.ain_s1 ;
assign _035_ = \add_12ns_12s_12_2_1_U6.top_add_12ns_12s_12_2_1_Adder_5_U.ce  ? \add_12ns_12s_12_2_1_U6.top_add_12ns_12s_12_2_1_Adder_5_U.facout_s1  : \add_12ns_12s_12_2_1_U6.top_add_12ns_12s_12_2_1_Adder_5_U.carry_s1 ;
assign _036_ = \add_12ns_12s_12_2_1_U6.top_add_12ns_12s_12_2_1_Adder_5_U.ce  ? \add_12ns_12s_12_2_1_U6.top_add_12ns_12s_12_2_1_Adder_5_U.fas_s1  : \add_12ns_12s_12_2_1_U6.top_add_12ns_12s_12_2_1_Adder_5_U.sum_s1 ;
assign _037_ = \add_12ns_12s_12_2_1_U6.top_add_12ns_12s_12_2_1_Adder_5_U.u1.a  + \add_12ns_12s_12_2_1_U6.top_add_12ns_12s_12_2_1_Adder_5_U.u1.b ;
assign { \add_12ns_12s_12_2_1_U6.top_add_12ns_12s_12_2_1_Adder_5_U.u1.cout , \add_12ns_12s_12_2_1_U6.top_add_12ns_12s_12_2_1_Adder_5_U.u1.s  } = _037_ + \add_12ns_12s_12_2_1_U6.top_add_12ns_12s_12_2_1_Adder_5_U.u1.cin ;
assign _038_ = \add_12ns_12s_12_2_1_U6.top_add_12ns_12s_12_2_1_Adder_5_U.u2.a  + \add_12ns_12s_12_2_1_U6.top_add_12ns_12s_12_2_1_Adder_5_U.u2.b ;
assign { \add_12ns_12s_12_2_1_U6.top_add_12ns_12s_12_2_1_Adder_5_U.u2.cout , \add_12ns_12s_12_2_1_U6.top_add_12ns_12s_12_2_1_Adder_5_U.u2.s  } = _038_ + \add_12ns_12s_12_2_1_U6.top_add_12ns_12s_12_2_1_Adder_5_U.u2.cin ;
always @(posedge \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.clk )
\add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.bin_s1  <= _040_;
always @(posedge \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.clk )
\add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.ain_s1  <= _039_;
always @(posedge \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.clk )
\add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.sum_s1  <= _042_;
always @(posedge \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.clk )
\add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.carry_s1  <= _041_;
assign _040_ = \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.ce  ? \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.b [16:8] : \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.bin_s1 ;
assign _039_ = \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.ce  ? \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.a [16:8] : \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.ain_s1 ;
assign _041_ = \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.ce  ? \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.facout_s1  : \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.carry_s1 ;
assign _042_ = \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.ce  ? \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.fas_s1  : \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.sum_s1 ;
assign _043_ = \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.u1.a  + \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.u1.b ;
assign { \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.u1.cout , \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.u1.s  } = _043_ + \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.u1.cin ;
assign _044_ = \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.u2.a  + \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.u2.b ;
assign { \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.u2.cout , \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.u2.s  } = _044_ + \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.u2.cin ;
always @(posedge \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_10_U.clk )
\add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_10_U.bin_s1  <= _046_;
always @(posedge \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_10_U.clk )
\add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_10_U.ain_s1  <= _045_;
always @(posedge \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_10_U.clk )
\add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_10_U.sum_s1  <= _048_;
always @(posedge \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_10_U.clk )
\add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_10_U.carry_s1  <= _047_;
assign _046_ = \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_10_U.ce  ? \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_10_U.b [1] : \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_10_U.bin_s1 ;
assign _045_ = \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_10_U.ce  ? \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_10_U.a [1] : \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_10_U.ain_s1 ;
assign _047_ = \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_10_U.ce  ? \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_10_U.facout_s1  : \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_10_U.carry_s1 ;
assign _048_ = \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_10_U.ce  ? \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_10_U.fas_s1  : \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_10_U.sum_s1 ;
assign _049_ = \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_10_U.u1.a  + \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_10_U.u1.b ;
assign { \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_10_U.u1.cout , \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_10_U.u1.s  } = _049_ + \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_10_U.u1.cin ;
assign _050_ = \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_10_U.u2.a  + \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_10_U.u2.b ;
assign { \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_10_U.u2.cout , \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_10_U.u2.s  } = _050_ + \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_10_U.u2.cin ;
always @(posedge \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.clk )
\add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s1  <= _052_;
always @(posedge \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.clk )
\add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s1  <= _051_;
always @(posedge \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.clk )
\add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.sum_s1  <= _054_;
always @(posedge \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.clk )
\add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.carry_s1  <= _053_;
assign _052_ = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.ce  ? \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.b [31:16] : \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s1 ;
assign _051_ = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.ce  ? \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.a [31:16] : \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s1 ;
assign _053_ = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.ce  ? \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.facout_s1  : \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.carry_s1 ;
assign _054_ = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.ce  ? \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s1  : \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.sum_s1 ;
assign _055_ = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.a  + \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.b ;
assign { \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cout , \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.s  } = _055_ + \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cin ;
assign _056_ = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.a  + \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.b ;
assign { \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cout , \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.s  } = _056_ + \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cin ;
always @(posedge \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.clk )
\add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s1  <= _058_;
always @(posedge \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.clk )
\add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s1  <= _057_;
always @(posedge \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.clk )
\add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.sum_s1  <= _060_;
always @(posedge \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.clk )
\add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.carry_s1  <= _059_;
assign _058_ = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.ce  ? \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.b [31:16] : \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s1 ;
assign _057_ = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.ce  ? \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.a [31:16] : \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s1 ;
assign _059_ = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.ce  ? \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.facout_s1  : \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.carry_s1 ;
assign _060_ = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.ce  ? \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s1  : \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.sum_s1 ;
assign _061_ = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.a  + \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.b ;
assign { \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cout , \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.s  } = _061_ + \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cin ;
assign _062_ = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.a  + \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.b ;
assign { \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cout , \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.s  } = _062_ + \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cin ;
always @(posedge \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.clk )
\add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s1  <= _064_;
always @(posedge \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.clk )
\add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s1  <= _063_;
always @(posedge \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.clk )
\add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.sum_s1  <= _066_;
always @(posedge \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.clk )
\add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.carry_s1  <= _065_;
assign _064_ = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.ce  ? \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.b [31:16] : \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s1 ;
assign _063_ = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.ce  ? \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.a [31:16] : \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s1 ;
assign _065_ = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.ce  ? \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.facout_s1  : \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.carry_s1 ;
assign _066_ = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.ce  ? \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s1  : \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.sum_s1 ;
assign _067_ = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.a  + \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.b ;
assign { \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cout , \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.s  } = _067_ + \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cin ;
assign _068_ = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.a  + \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.b ;
assign { \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cout , \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.s  } = _068_ + \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cin ;
always @(posedge \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_7_U.clk )
\add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s1  <= _070_;
always @(posedge \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_7_U.clk )
\add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s1  <= _069_;
always @(posedge \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_7_U.clk )
\add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_7_U.sum_s1  <= _072_;
always @(posedge \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_7_U.clk )
\add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_7_U.carry_s1  <= _071_;
assign _070_ = \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_7_U.ce  ? \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_7_U.b [31:16] : \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s1 ;
assign _069_ = \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_7_U.ce  ? \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_7_U.a [31:16] : \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s1 ;
assign _071_ = \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_7_U.ce  ? \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_7_U.facout_s1  : \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_7_U.carry_s1 ;
assign _072_ = \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_7_U.ce  ? \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s1  : \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_7_U.sum_s1 ;
assign _073_ = \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.a  + \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.b ;
assign { \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cout , \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.s  } = _073_ + \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cin ;
assign _074_ = \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.a  + \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.b ;
assign { \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cout , \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.s  } = _074_ + \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cin ;
always @(posedge \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.clk )
\add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s1  <= _076_;
always @(posedge \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.clk )
\add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s1  <= _075_;
always @(posedge \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.clk )
\add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.sum_s1  <= _078_;
always @(posedge \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.clk )
\add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.carry_s1  <= _077_;
assign _076_ = \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.ce  ? \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.b [31:16] : \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s1 ;
assign _075_ = \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.ce  ? \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.a [31:16] : \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s1 ;
assign _077_ = \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.ce  ? \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.facout_s1  : \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.carry_s1 ;
assign _078_ = \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.ce  ? \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s1  : \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.sum_s1 ;
assign _079_ = \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.a  + \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.b ;
assign { \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cout , \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.s  } = _079_ + \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cin ;
assign _080_ = \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.a  + \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.b ;
assign { \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cout , \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.s  } = _080_ + \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cin ;
always @(posedge \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_6_U.clk )
\add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_6_U.bin_s1  <= _082_;
always @(posedge \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_6_U.clk )
\add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_6_U.ain_s1  <= _081_;
always @(posedge \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_6_U.clk )
\add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_6_U.sum_s1  <= _084_;
always @(posedge \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_6_U.clk )
\add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_6_U.carry_s1  <= _083_;
assign _082_ = \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_6_U.ce  ? \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_6_U.b [33:17] : \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_6_U.bin_s1 ;
assign _081_ = \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_6_U.ce  ? \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_6_U.a [33:17] : \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_6_U.ain_s1 ;
assign _083_ = \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_6_U.ce  ? \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_6_U.facout_s1  : \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_6_U.carry_s1 ;
assign _084_ = \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_6_U.ce  ? \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_6_U.fas_s1  : \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_6_U.sum_s1 ;
assign _085_ = \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_6_U.u1.a  + \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_6_U.u1.b ;
assign { \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_6_U.u1.cout , \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_6_U.u1.s  } = _085_ + \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_6_U.u1.cin ;
assign _086_ = \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_6_U.u2.a  + \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_6_U.u2.b ;
assign { \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_6_U.u2.cout , \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_6_U.u2.s  } = _086_ + \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_6_U.u2.cin ;
always @(posedge \add_37s_37s_37_2_1_U11.top_add_37s_37s_37_2_1_Adder_9_U.clk )
\add_37s_37s_37_2_1_U11.top_add_37s_37s_37_2_1_Adder_9_U.bin_s1  <= _088_;
always @(posedge \add_37s_37s_37_2_1_U11.top_add_37s_37s_37_2_1_Adder_9_U.clk )
\add_37s_37s_37_2_1_U11.top_add_37s_37s_37_2_1_Adder_9_U.ain_s1  <= _087_;
always @(posedge \add_37s_37s_37_2_1_U11.top_add_37s_37s_37_2_1_Adder_9_U.clk )
\add_37s_37s_37_2_1_U11.top_add_37s_37s_37_2_1_Adder_9_U.sum_s1  <= _090_;
always @(posedge \add_37s_37s_37_2_1_U11.top_add_37s_37s_37_2_1_Adder_9_U.clk )
\add_37s_37s_37_2_1_U11.top_add_37s_37s_37_2_1_Adder_9_U.carry_s1  <= _089_;
assign _088_ = \add_37s_37s_37_2_1_U11.top_add_37s_37s_37_2_1_Adder_9_U.ce  ? \add_37s_37s_37_2_1_U11.top_add_37s_37s_37_2_1_Adder_9_U.b [36:18] : \add_37s_37s_37_2_1_U11.top_add_37s_37s_37_2_1_Adder_9_U.bin_s1 ;
assign _087_ = \add_37s_37s_37_2_1_U11.top_add_37s_37s_37_2_1_Adder_9_U.ce  ? \add_37s_37s_37_2_1_U11.top_add_37s_37s_37_2_1_Adder_9_U.a [36:18] : \add_37s_37s_37_2_1_U11.top_add_37s_37s_37_2_1_Adder_9_U.ain_s1 ;
assign _089_ = \add_37s_37s_37_2_1_U11.top_add_37s_37s_37_2_1_Adder_9_U.ce  ? \add_37s_37s_37_2_1_U11.top_add_37s_37s_37_2_1_Adder_9_U.facout_s1  : \add_37s_37s_37_2_1_U11.top_add_37s_37s_37_2_1_Adder_9_U.carry_s1 ;
assign _090_ = \add_37s_37s_37_2_1_U11.top_add_37s_37s_37_2_1_Adder_9_U.ce  ? \add_37s_37s_37_2_1_U11.top_add_37s_37s_37_2_1_Adder_9_U.fas_s1  : \add_37s_37s_37_2_1_U11.top_add_37s_37s_37_2_1_Adder_9_U.sum_s1 ;
assign _091_ = \add_37s_37s_37_2_1_U11.top_add_37s_37s_37_2_1_Adder_9_U.u1.a  + \add_37s_37s_37_2_1_U11.top_add_37s_37s_37_2_1_Adder_9_U.u1.b ;
assign { \add_37s_37s_37_2_1_U11.top_add_37s_37s_37_2_1_Adder_9_U.u1.cout , \add_37s_37s_37_2_1_U11.top_add_37s_37s_37_2_1_Adder_9_U.u1.s  } = _091_ + \add_37s_37s_37_2_1_U11.top_add_37s_37s_37_2_1_Adder_9_U.u1.cin ;
assign _092_ = \add_37s_37s_37_2_1_U11.top_add_37s_37s_37_2_1_Adder_9_U.u2.a  + \add_37s_37s_37_2_1_U11.top_add_37s_37s_37_2_1_Adder_9_U.u2.b ;
assign { \add_37s_37s_37_2_1_U11.top_add_37s_37s_37_2_1_Adder_9_U.u2.cout , \add_37s_37s_37_2_1_U11.top_add_37s_37s_37_2_1_Adder_9_U.u2.s  } = _092_ + \add_37s_37s_37_2_1_U11.top_add_37s_37s_37_2_1_Adder_9_U.u2.cin ;
always @(posedge \add_4s_4ns_4_2_1_U10.top_add_4s_4ns_4_2_1_Adder_8_U.clk )
\add_4s_4ns_4_2_1_U10.top_add_4s_4ns_4_2_1_Adder_8_U.bin_s1  <= _094_;
always @(posedge \add_4s_4ns_4_2_1_U10.top_add_4s_4ns_4_2_1_Adder_8_U.clk )
\add_4s_4ns_4_2_1_U10.top_add_4s_4ns_4_2_1_Adder_8_U.ain_s1  <= _093_;
always @(posedge \add_4s_4ns_4_2_1_U10.top_add_4s_4ns_4_2_1_Adder_8_U.clk )
\add_4s_4ns_4_2_1_U10.top_add_4s_4ns_4_2_1_Adder_8_U.sum_s1  <= _096_;
always @(posedge \add_4s_4ns_4_2_1_U10.top_add_4s_4ns_4_2_1_Adder_8_U.clk )
\add_4s_4ns_4_2_1_U10.top_add_4s_4ns_4_2_1_Adder_8_U.carry_s1  <= _095_;
assign _094_ = \add_4s_4ns_4_2_1_U10.top_add_4s_4ns_4_2_1_Adder_8_U.ce  ? \add_4s_4ns_4_2_1_U10.top_add_4s_4ns_4_2_1_Adder_8_U.b [3:2] : \add_4s_4ns_4_2_1_U10.top_add_4s_4ns_4_2_1_Adder_8_U.bin_s1 ;
assign _093_ = \add_4s_4ns_4_2_1_U10.top_add_4s_4ns_4_2_1_Adder_8_U.ce  ? \add_4s_4ns_4_2_1_U10.top_add_4s_4ns_4_2_1_Adder_8_U.a [3:2] : \add_4s_4ns_4_2_1_U10.top_add_4s_4ns_4_2_1_Adder_8_U.ain_s1 ;
assign _095_ = \add_4s_4ns_4_2_1_U10.top_add_4s_4ns_4_2_1_Adder_8_U.ce  ? \add_4s_4ns_4_2_1_U10.top_add_4s_4ns_4_2_1_Adder_8_U.facout_s1  : \add_4s_4ns_4_2_1_U10.top_add_4s_4ns_4_2_1_Adder_8_U.carry_s1 ;
assign _096_ = \add_4s_4ns_4_2_1_U10.top_add_4s_4ns_4_2_1_Adder_8_U.ce  ? \add_4s_4ns_4_2_1_U10.top_add_4s_4ns_4_2_1_Adder_8_U.fas_s1  : \add_4s_4ns_4_2_1_U10.top_add_4s_4ns_4_2_1_Adder_8_U.sum_s1 ;
assign _097_ = \add_4s_4ns_4_2_1_U10.top_add_4s_4ns_4_2_1_Adder_8_U.u1.a  + \add_4s_4ns_4_2_1_U10.top_add_4s_4ns_4_2_1_Adder_8_U.u1.b ;
assign { \add_4s_4ns_4_2_1_U10.top_add_4s_4ns_4_2_1_Adder_8_U.u1.cout , \add_4s_4ns_4_2_1_U10.top_add_4s_4ns_4_2_1_Adder_8_U.u1.s  } = _097_ + \add_4s_4ns_4_2_1_U10.top_add_4s_4ns_4_2_1_Adder_8_U.u1.cin ;
assign _098_ = \add_4s_4ns_4_2_1_U10.top_add_4s_4ns_4_2_1_Adder_8_U.u2.a  + \add_4s_4ns_4_2_1_U10.top_add_4s_4ns_4_2_1_Adder_8_U.u2.b ;
assign { \add_4s_4ns_4_2_1_U10.top_add_4s_4ns_4_2_1_Adder_8_U.u2.cout , \add_4s_4ns_4_2_1_U10.top_add_4s_4ns_4_2_1_Adder_8_U.u2.s  } = _098_ + \add_4s_4ns_4_2_1_U10.top_add_4s_4ns_4_2_1_Adder_8_U.u2.cin ;
always @(posedge \add_5ns_5ns_5_2_1_U15.top_add_5ns_5ns_5_2_1_Adder_1_U.clk )
\add_5ns_5ns_5_2_1_U15.top_add_5ns_5ns_5_2_1_Adder_1_U.bin_s1  <= _100_;
always @(posedge \add_5ns_5ns_5_2_1_U15.top_add_5ns_5ns_5_2_1_Adder_1_U.clk )
\add_5ns_5ns_5_2_1_U15.top_add_5ns_5ns_5_2_1_Adder_1_U.ain_s1  <= _099_;
always @(posedge \add_5ns_5ns_5_2_1_U15.top_add_5ns_5ns_5_2_1_Adder_1_U.clk )
\add_5ns_5ns_5_2_1_U15.top_add_5ns_5ns_5_2_1_Adder_1_U.sum_s1  <= _102_;
always @(posedge \add_5ns_5ns_5_2_1_U15.top_add_5ns_5ns_5_2_1_Adder_1_U.clk )
\add_5ns_5ns_5_2_1_U15.top_add_5ns_5ns_5_2_1_Adder_1_U.carry_s1  <= _101_;
assign _100_ = \add_5ns_5ns_5_2_1_U15.top_add_5ns_5ns_5_2_1_Adder_1_U.ce  ? \add_5ns_5ns_5_2_1_U15.top_add_5ns_5ns_5_2_1_Adder_1_U.b [4:2] : \add_5ns_5ns_5_2_1_U15.top_add_5ns_5ns_5_2_1_Adder_1_U.bin_s1 ;
assign _099_ = \add_5ns_5ns_5_2_1_U15.top_add_5ns_5ns_5_2_1_Adder_1_U.ce  ? \add_5ns_5ns_5_2_1_U15.top_add_5ns_5ns_5_2_1_Adder_1_U.a [4:2] : \add_5ns_5ns_5_2_1_U15.top_add_5ns_5ns_5_2_1_Adder_1_U.ain_s1 ;
assign _101_ = \add_5ns_5ns_5_2_1_U15.top_add_5ns_5ns_5_2_1_Adder_1_U.ce  ? \add_5ns_5ns_5_2_1_U15.top_add_5ns_5ns_5_2_1_Adder_1_U.facout_s1  : \add_5ns_5ns_5_2_1_U15.top_add_5ns_5ns_5_2_1_Adder_1_U.carry_s1 ;
assign _102_ = \add_5ns_5ns_5_2_1_U15.top_add_5ns_5ns_5_2_1_Adder_1_U.ce  ? \add_5ns_5ns_5_2_1_U15.top_add_5ns_5ns_5_2_1_Adder_1_U.fas_s1  : \add_5ns_5ns_5_2_1_U15.top_add_5ns_5ns_5_2_1_Adder_1_U.sum_s1 ;
assign _103_ = \add_5ns_5ns_5_2_1_U15.top_add_5ns_5ns_5_2_1_Adder_1_U.u1.a  + \add_5ns_5ns_5_2_1_U15.top_add_5ns_5ns_5_2_1_Adder_1_U.u1.b ;
assign { \add_5ns_5ns_5_2_1_U15.top_add_5ns_5ns_5_2_1_Adder_1_U.u1.cout , \add_5ns_5ns_5_2_1_U15.top_add_5ns_5ns_5_2_1_Adder_1_U.u1.s  } = _103_ + \add_5ns_5ns_5_2_1_U15.top_add_5ns_5ns_5_2_1_Adder_1_U.u1.cin ;
assign _104_ = \add_5ns_5ns_5_2_1_U15.top_add_5ns_5ns_5_2_1_Adder_1_U.u2.a  + \add_5ns_5ns_5_2_1_U15.top_add_5ns_5ns_5_2_1_Adder_1_U.u2.b ;
assign { \add_5ns_5ns_5_2_1_U15.top_add_5ns_5ns_5_2_1_Adder_1_U.u2.cout , \add_5ns_5ns_5_2_1_U15.top_add_5ns_5ns_5_2_1_Adder_1_U.u2.s  } = _104_ + \add_5ns_5ns_5_2_1_U15.top_add_5ns_5ns_5_2_1_Adder_1_U.u2.cin ;
always @(posedge \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.clk )
\add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.bin_s1  <= _106_;
always @(posedge \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.clk )
\add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.ain_s1  <= _105_;
always @(posedge \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.clk )
\add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.sum_s1  <= _108_;
always @(posedge \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.clk )
\add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.carry_s1  <= _107_;
assign _106_ = \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.ce  ? \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.b [4:2] : \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.bin_s1 ;
assign _105_ = \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.ce  ? \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.a [4:2] : \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.ain_s1 ;
assign _107_ = \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.ce  ? \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.facout_s1  : \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.carry_s1 ;
assign _108_ = \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.ce  ? \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.fas_s1  : \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.sum_s1 ;
assign _109_ = \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.u1.a  + \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.u1.b ;
assign { \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.u1.cout , \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.u1.s  } = _109_ + \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.u1.cin ;
assign _110_ = \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.u2.a  + \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.u2.b ;
assign { \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.u2.cout , \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.u2.s  } = _110_ + \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.u2.cin ;
always @(posedge \add_6s_6s_6_2_1_U1.top_add_6s_6s_6_2_1_Adder_0_U.clk )
\add_6s_6s_6_2_1_U1.top_add_6s_6s_6_2_1_Adder_0_U.bin_s1  <= _112_;
always @(posedge \add_6s_6s_6_2_1_U1.top_add_6s_6s_6_2_1_Adder_0_U.clk )
\add_6s_6s_6_2_1_U1.top_add_6s_6s_6_2_1_Adder_0_U.ain_s1  <= _111_;
always @(posedge \add_6s_6s_6_2_1_U1.top_add_6s_6s_6_2_1_Adder_0_U.clk )
\add_6s_6s_6_2_1_U1.top_add_6s_6s_6_2_1_Adder_0_U.sum_s1  <= _114_;
always @(posedge \add_6s_6s_6_2_1_U1.top_add_6s_6s_6_2_1_Adder_0_U.clk )
\add_6s_6s_6_2_1_U1.top_add_6s_6s_6_2_1_Adder_0_U.carry_s1  <= _113_;
assign _112_ = \add_6s_6s_6_2_1_U1.top_add_6s_6s_6_2_1_Adder_0_U.ce  ? \add_6s_6s_6_2_1_U1.top_add_6s_6s_6_2_1_Adder_0_U.b [5:3] : \add_6s_6s_6_2_1_U1.top_add_6s_6s_6_2_1_Adder_0_U.bin_s1 ;
assign _111_ = \add_6s_6s_6_2_1_U1.top_add_6s_6s_6_2_1_Adder_0_U.ce  ? \add_6s_6s_6_2_1_U1.top_add_6s_6s_6_2_1_Adder_0_U.a [5:3] : \add_6s_6s_6_2_1_U1.top_add_6s_6s_6_2_1_Adder_0_U.ain_s1 ;
assign _113_ = \add_6s_6s_6_2_1_U1.top_add_6s_6s_6_2_1_Adder_0_U.ce  ? \add_6s_6s_6_2_1_U1.top_add_6s_6s_6_2_1_Adder_0_U.facout_s1  : \add_6s_6s_6_2_1_U1.top_add_6s_6s_6_2_1_Adder_0_U.carry_s1 ;
assign _114_ = \add_6s_6s_6_2_1_U1.top_add_6s_6s_6_2_1_Adder_0_U.ce  ? \add_6s_6s_6_2_1_U1.top_add_6s_6s_6_2_1_Adder_0_U.fas_s1  : \add_6s_6s_6_2_1_U1.top_add_6s_6s_6_2_1_Adder_0_U.sum_s1 ;
assign _115_ = \add_6s_6s_6_2_1_U1.top_add_6s_6s_6_2_1_Adder_0_U.u1.a  + \add_6s_6s_6_2_1_U1.top_add_6s_6s_6_2_1_Adder_0_U.u1.b ;
assign { \add_6s_6s_6_2_1_U1.top_add_6s_6s_6_2_1_Adder_0_U.u1.cout , \add_6s_6s_6_2_1_U1.top_add_6s_6s_6_2_1_Adder_0_U.u1.s  } = _115_ + \add_6s_6s_6_2_1_U1.top_add_6s_6s_6_2_1_Adder_0_U.u1.cin ;
assign _116_ = \add_6s_6s_6_2_1_U1.top_add_6s_6s_6_2_1_Adder_0_U.u2.a  + \add_6s_6s_6_2_1_U1.top_add_6s_6s_6_2_1_Adder_0_U.u2.b ;
assign { \add_6s_6s_6_2_1_U1.top_add_6s_6s_6_2_1_Adder_0_U.u2.cout , \add_6s_6s_6_2_1_U1.top_add_6s_6s_6_2_1_Adder_0_U.u2.s  } = _116_ + \add_6s_6s_6_2_1_U1.top_add_6s_6s_6_2_1_Adder_0_U.u2.cin ;
always @(posedge \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.clk )
\add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.bin_s1  <= _118_;
always @(posedge \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.clk )
\add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.ain_s1  <= _117_;
always @(posedge \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.clk )
\add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.sum_s1  <= _120_;
always @(posedge \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.clk )
\add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.carry_s1  <= _119_;
assign _118_ = \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.ce  ? \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.b [8:4] : \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.bin_s1 ;
assign _117_ = \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.ce  ? \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.a [8:4] : \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.ain_s1 ;
assign _119_ = \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.ce  ? \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.facout_s1  : \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.carry_s1 ;
assign _120_ = \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.ce  ? \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.fas_s1  : \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.sum_s1 ;
assign _121_ = \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.u1.a  + \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.u1.b ;
assign { \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.u1.cout , \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.u1.s  } = _121_ + \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.u1.cin ;
assign _122_ = \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.u2.a  + \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.u2.b ;
assign { \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.u2.cout , \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.u2.s  } = _122_ + \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.u2.cin ;
assign \sub_10s_10ns_10_2_1_U3.top_sub_10s_10ns_10_2_1_Adder_2_U.bin_s0  = ~ \sub_10s_10ns_10_2_1_U3.top_sub_10s_10ns_10_2_1_Adder_2_U.b ;
always @(posedge \sub_10s_10ns_10_2_1_U3.top_sub_10s_10ns_10_2_1_Adder_2_U.clk )
\sub_10s_10ns_10_2_1_U3.top_sub_10s_10ns_10_2_1_Adder_2_U.bin_s1  <= _124_;
always @(posedge \sub_10s_10ns_10_2_1_U3.top_sub_10s_10ns_10_2_1_Adder_2_U.clk )
\sub_10s_10ns_10_2_1_U3.top_sub_10s_10ns_10_2_1_Adder_2_U.ain_s1  <= _123_;
always @(posedge \sub_10s_10ns_10_2_1_U3.top_sub_10s_10ns_10_2_1_Adder_2_U.clk )
\sub_10s_10ns_10_2_1_U3.top_sub_10s_10ns_10_2_1_Adder_2_U.sum_s1  <= _126_;
always @(posedge \sub_10s_10ns_10_2_1_U3.top_sub_10s_10ns_10_2_1_Adder_2_U.clk )
\sub_10s_10ns_10_2_1_U3.top_sub_10s_10ns_10_2_1_Adder_2_U.carry_s1  <= _125_;
assign _124_ = \sub_10s_10ns_10_2_1_U3.top_sub_10s_10ns_10_2_1_Adder_2_U.ce  ? \sub_10s_10ns_10_2_1_U3.top_sub_10s_10ns_10_2_1_Adder_2_U.bin_s0 [9:5] : \sub_10s_10ns_10_2_1_U3.top_sub_10s_10ns_10_2_1_Adder_2_U.bin_s1 ;
assign _123_ = \sub_10s_10ns_10_2_1_U3.top_sub_10s_10ns_10_2_1_Adder_2_U.ce  ? \sub_10s_10ns_10_2_1_U3.top_sub_10s_10ns_10_2_1_Adder_2_U.a [9:5] : \sub_10s_10ns_10_2_1_U3.top_sub_10s_10ns_10_2_1_Adder_2_U.ain_s1 ;
assign _125_ = \sub_10s_10ns_10_2_1_U3.top_sub_10s_10ns_10_2_1_Adder_2_U.ce  ? \sub_10s_10ns_10_2_1_U3.top_sub_10s_10ns_10_2_1_Adder_2_U.facout_s1  : \sub_10s_10ns_10_2_1_U3.top_sub_10s_10ns_10_2_1_Adder_2_U.carry_s1 ;
assign _126_ = \sub_10s_10ns_10_2_1_U3.top_sub_10s_10ns_10_2_1_Adder_2_U.ce  ? \sub_10s_10ns_10_2_1_U3.top_sub_10s_10ns_10_2_1_Adder_2_U.fas_s1  : \sub_10s_10ns_10_2_1_U3.top_sub_10s_10ns_10_2_1_Adder_2_U.sum_s1 ;
assign _127_ = \sub_10s_10ns_10_2_1_U3.top_sub_10s_10ns_10_2_1_Adder_2_U.u1.a  + \sub_10s_10ns_10_2_1_U3.top_sub_10s_10ns_10_2_1_Adder_2_U.u1.b ;
assign { \sub_10s_10ns_10_2_1_U3.top_sub_10s_10ns_10_2_1_Adder_2_U.u1.cout , \sub_10s_10ns_10_2_1_U3.top_sub_10s_10ns_10_2_1_Adder_2_U.u1.s  } = _127_ + \sub_10s_10ns_10_2_1_U3.top_sub_10s_10ns_10_2_1_Adder_2_U.u1.cin ;
assign _128_ = \sub_10s_10ns_10_2_1_U3.top_sub_10s_10ns_10_2_1_Adder_2_U.u2.a  + \sub_10s_10ns_10_2_1_U3.top_sub_10s_10ns_10_2_1_Adder_2_U.u2.b ;
assign { \sub_10s_10ns_10_2_1_U3.top_sub_10s_10ns_10_2_1_Adder_2_U.u2.cout , \sub_10s_10ns_10_2_1_U3.top_sub_10s_10ns_10_2_1_Adder_2_U.u2.s  } = _128_ + \sub_10s_10ns_10_2_1_U3.top_sub_10s_10ns_10_2_1_Adder_2_U.u2.cin ;
assign _129_ = $signed(op_4) > $signed(1'h0);
assign _130_ = $signed(ret_V_5_fu_483_p3) > $signed({ 1'h0, op_7 });
assign _131_ = | op_14[3:0];
always @(posedge ap_clk)
ret_reg_619 <= _024_;
always @(posedge ap_clk)
select_ln850_5_reg_624 <= _025_;
always @(posedge ap_clk)
ret_V_4_reg_748 <= _021_;
always @(posedge ap_clk)
ret_V_14_reg_753 <= _017_;
always @(posedge ap_clk)
ret_V_19_cast_reg_758 <= _019_;
always @(posedge ap_clk)
ret_V_13_reg_701 <= _016_;
always @(posedge ap_clk)
ret_V_12_reg_684 <= _015_;
always @(posedge ap_clk)
ret_V_8_cast_reg_689 <= _022_;
always @(posedge ap_clk)
ret_V_11_reg_587 <= _014_;
always @(posedge ap_clk)
ret_V_reg_592 <= _023_;
always @(posedge ap_clk)
op_25_V_reg_711 <= _013_;
always @(posedge ap_clk)
op_23_V_reg_664 <= _012_;
always @(posedge ap_clk)
op_17_V_reg_765 <= _010_;
always @(posedge ap_clk)
ret_V_2_reg_609 <= _020_;
always @(posedge ap_clk)
icmp_ln886_reg_614 <= _009_;
always @(posedge ap_clk)
sext_ln835_reg_721 <= _026_;
always @(posedge ap_clk)
icmp_ln851_reg_728 <= _008_;
always @(posedge ap_clk)
icmp_ln851_1_reg_743 <= _007_;
always @(posedge ap_clk)
op_21_V_reg_644 <= _011_;
always @(posedge ap_clk)
add_ln69_reg_649 <= _005_;
always @(posedge ap_clk)
ret_V_15_reg_785 <= _018_;
always @(posedge ap_clk)
add_ln69_4_reg_790 <= _003_;
always @(posedge ap_clk)
add_ln69_3_reg_810 <= _002_;
always @(posedge ap_clk)
add_ln69_5_reg_815 <= _004_;
always @(posedge ap_clk)
add_ln691_reg_696 <= _001_;
always @(posedge ap_clk)
add_ln691_1_reg_775 <= _000_;
always @(posedge ap_clk)
ap_CS_fsm <= _006_;
assign _027_ = _030_ ? 2'h2 : 2'h1;
assign _132_ = ap_CS_fsm == 1'h1;
function [24:0] _387_;
input [24:0] a;
input [624:0] b;
input [24:0] s;
case (s)
25'b0000000000000000000000001:
_387_ = b[24:0];
25'b0000000000000000000000010:
_387_ = b[49:25];
25'b0000000000000000000000100:
_387_ = b[74:50];
25'b0000000000000000000001000:
_387_ = b[99:75];
25'b0000000000000000000010000:
_387_ = b[124:100];
25'b0000000000000000000100000:
_387_ = b[149:125];
25'b0000000000000000001000000:
_387_ = b[174:150];
25'b0000000000000000010000000:
_387_ = b[199:175];
25'b0000000000000000100000000:
_387_ = b[224:200];
25'b0000000000000001000000000:
_387_ = b[249:225];
25'b0000000000000010000000000:
_387_ = b[274:250];
25'b0000000000000100000000000:
_387_ = b[299:275];
25'b0000000000001000000000000:
_387_ = b[324:300];
25'b0000000000010000000000000:
_387_ = b[349:325];
25'b0000000000100000000000000:
_387_ = b[374:350];
25'b0000000001000000000000000:
_387_ = b[399:375];
25'b0000000010000000000000000:
_387_ = b[424:400];
25'b0000000100000000000000000:
_387_ = b[449:425];
25'b0000001000000000000000000:
_387_ = b[474:450];
25'b0000010000000000000000000:
_387_ = b[499:475];
25'b0000100000000000000000000:
_387_ = b[524:500];
25'b0001000000000000000000000:
_387_ = b[549:525];
25'b0010000000000000000000000:
_387_ = b[574:550];
25'b0100000000000000000000000:
_387_ = b[599:575];
25'b1000000000000000000000000:
_387_ = b[624:600];
25'b0000000000000000000000000:
_387_ = a;
default:
_387_ = 25'bx;
endcase
endfunction
assign ap_NS_fsm = _387_(25'hxxxxxxx, { 23'h000000, _027_, 600'h000002000002000002000002000002000002000002000002000002000002000002000002000002000002000002000002000002000002000002000002000002000002000002000000000001 }, { _132_, _156_, _155_, _154_, _153_, _152_, _151_, _150_, _149_, _148_, _147_, _146_, _145_, _144_, _143_, _142_, _141_, _140_, _139_, _138_, _137_, _136_, _135_, _134_, _133_ });
assign _133_ = ap_CS_fsm == 25'h1000000;
assign _134_ = ap_CS_fsm == 24'h800000;
assign _135_ = ap_CS_fsm == 23'h400000;
assign _136_ = ap_CS_fsm == 22'h200000;
assign _137_ = ap_CS_fsm == 21'h100000;
assign _138_ = ap_CS_fsm == 20'h80000;
assign _139_ = ap_CS_fsm == 19'h40000;
assign _140_ = ap_CS_fsm == 18'h20000;
assign _141_ = ap_CS_fsm == 17'h10000;
assign _142_ = ap_CS_fsm == 16'h8000;
assign _143_ = ap_CS_fsm == 15'h4000;
assign _144_ = ap_CS_fsm == 14'h2000;
assign _145_ = ap_CS_fsm == 13'h1000;
assign _146_ = ap_CS_fsm == 12'h800;
assign _147_ = ap_CS_fsm == 11'h400;
assign _148_ = ap_CS_fsm == 10'h200;
assign _149_ = ap_CS_fsm == 9'h100;
assign _150_ = ap_CS_fsm == 8'h80;
assign _151_ = ap_CS_fsm == 7'h40;
assign _152_ = ap_CS_fsm == 6'h20;
assign _153_ = ap_CS_fsm == 5'h10;
assign _154_ = ap_CS_fsm == 4'h8;
assign _155_ = ap_CS_fsm == 3'h4;
assign _156_ = ap_CS_fsm == 2'h2;
assign op_31_ap_vld = ap_CS_fsm[24] ? 1'h1 : 1'h0;
assign ap_idle = _029_ ? 1'h1 : 1'h0;
assign _025_ = ap_CS_fsm[4] ? select_ln850_5_fu_266_p3 : select_ln850_5_reg_624;
assign _024_ = ap_CS_fsm[4] ? grp_fu_238_p2 : ret_reg_619;
assign _019_ = ap_CS_fsm[17] ? grp_fu_445_p2[35:4] : ret_V_19_cast_reg_758;
assign _017_ = ap_CS_fsm[17] ? grp_fu_445_p2 : ret_V_14_reg_753;
assign _021_ = ap_CS_fsm[17] ? grp_fu_424_p2 : ret_V_4_reg_748;
assign _016_ = ap_CS_fsm[13] ? ret_V_13_fu_385_p3 : ret_V_13_reg_701;
assign _022_ = ap_CS_fsm[10] ? grp_fu_348_p2[32:1] : ret_V_8_cast_reg_689;
assign _015_ = ap_CS_fsm[10] ? grp_fu_348_p2 : ret_V_12_reg_684;
assign _023_ = ap_CS_fsm[1] ? grp_fu_209_p2[5:1] : ret_V_reg_592;
assign _014_ = ap_CS_fsm[1] ? grp_fu_209_p2 : ret_V_11_reg_587;
assign _013_ = ap_CS_fsm[15] ? grp_fu_395_p2 : op_25_V_reg_711;
assign _012_ = ap_CS_fsm[8] ? grp_fu_327_p2 : op_23_V_reg_664;
assign _010_ = ap_CS_fsm[18] ? op_17_V_fu_498_p2 : op_17_V_reg_765;
assign _009_ = ap_CS_fsm[3] ? icmp_ln886_fu_244_p2 : icmp_ln886_reg_614;
assign _020_ = ap_CS_fsm[3] ? grp_fu_225_p2 : ret_V_2_reg_609;
assign _007_ = ap_CS_fsm[16] ? icmp_ln851_1_fu_455_p2 : icmp_ln851_1_reg_743;
assign _008_ = ap_CS_fsm[16] ? icmp_ln851_fu_418_p2 : icmp_ln851_reg_728;
assign _026_ = ap_CS_fsm[16] ? { op_0[7], op_0[7:5] } : sext_ln835_reg_721;
assign _005_ = ap_CS_fsm[6] ? grp_fu_305_p2 : add_ln69_reg_649;
assign _011_ = ap_CS_fsm[6] ? grp_fu_295_p2[16:6] : op_21_V_reg_644;
assign _003_ = ap_CS_fsm[20] ? grp_fu_516_p2 : add_ln69_4_reg_790;
assign _018_ = ap_CS_fsm[20] ? ret_V_15_fu_534_p3 : ret_V_15_reg_785;
assign _004_ = ap_CS_fsm[22] ? grp_fu_557_p2 : add_ln69_5_reg_815;
assign _002_ = ap_CS_fsm[22] ? grp_fu_549_p2 : add_ln69_3_reg_810;
assign _001_ = ap_CS_fsm[12] ? grp_fu_364_p2 : add_ln691_reg_696;
assign _000_ = _028_ ? grp_fu_504_p2 : add_ln691_1_reg_775;
assign _006_ = ap_rst ? 25'h0000001 : ap_NS_fsm;
assign icmp_ln851_1_fu_455_p2 = _131_ ? 1'h1 : 1'h0;
assign icmp_ln851_fu_418_p2 = _032_ ? 1'h1 : 1'h0;
assign icmp_ln886_fu_244_p2 = _129_ ? 1'h1 : 1'h0;
assign op_17_V_fu_498_p2 = _130_ ? 1'h1 : 1'h0;
assign ret_V_13_fu_385_p3 = ret_V_12_reg_684[33] ? select_ln850_2_fu_379_p3 : ret_V_8_cast_reg_689;
assign ret_V_15_fu_534_p3 = ret_V_14_reg_753[36] ? select_ln850_3_fu_529_p3 : ret_V_19_cast_reg_758;
assign ret_V_5_fu_483_p3 = op_0[7] ? select_ln850_fu_478_p3 : sext_ln835_reg_721;
assign select_ln850_2_fu_379_p3 = op_12[0] ? add_ln691_reg_696 : ret_V_8_cast_reg_689;
assign select_ln850_3_fu_529_p3 = icmp_ln851_1_reg_743 ? add_ln691_1_reg_775 : ret_V_19_cast_reg_758;
assign select_ln850_4_fu_260_p3 = op_2[0] ? ret_V_2_reg_609 : ret_V_reg_592;
assign select_ln850_5_fu_266_p3 = ret_V_11_reg_587[5] ? select_ln850_4_fu_260_p3 : ret_V_reg_592;
assign select_ln850_fu_478_p3 = icmp_ln851_reg_728 ? sext_ln835_reg_721 : ret_V_4_reg_748;
assign ap_CS_fsm_state1 = ap_CS_fsm[0];
assign ap_CS_fsm_state10 = ap_CS_fsm[9];
assign ap_CS_fsm_state11 = ap_CS_fsm[10];
assign ap_CS_fsm_state12 = ap_CS_fsm[11];
assign ap_CS_fsm_state13 = ap_CS_fsm[12];
assign ap_CS_fsm_state14 = ap_CS_fsm[13];
assign ap_CS_fsm_state15 = ap_CS_fsm[14];
assign ap_CS_fsm_state16 = ap_CS_fsm[15];
assign ap_CS_fsm_state17 = ap_CS_fsm[16];
assign ap_CS_fsm_state18 = ap_CS_fsm[17];
assign ap_CS_fsm_state19 = ap_CS_fsm[18];
assign ap_CS_fsm_state2 = ap_CS_fsm[1];
assign ap_CS_fsm_state20 = ap_CS_fsm[19];
assign ap_CS_fsm_state21 = ap_CS_fsm[20];
assign ap_CS_fsm_state22 = ap_CS_fsm[21];
assign ap_CS_fsm_state23 = ap_CS_fsm[22];
assign ap_CS_fsm_state24 = ap_CS_fsm[23];
assign ap_CS_fsm_state25 = ap_CS_fsm[24];
assign ap_CS_fsm_state3 = ap_CS_fsm[2];
assign ap_CS_fsm_state4 = ap_CS_fsm[3];
assign ap_CS_fsm_state5 = ap_CS_fsm[4];
assign ap_CS_fsm_state6 = ap_CS_fsm[5];
assign ap_CS_fsm_state7 = ap_CS_fsm[6];
assign ap_CS_fsm_state8 = ap_CS_fsm[7];
assign ap_CS_fsm_state9 = ap_CS_fsm[8];
assign ap_done = op_31_ap_vld;
assign ap_ready = op_31_ap_vld;
assign grp_fu_209_p0 = { op_8[3], op_8, 1'h0 };
assign grp_fu_209_p1 = { op_2[3], op_2[3], op_2 };
assign grp_fu_238_p0 = { op_4[7], op_4[7], op_4 };
assign grp_fu_238_p1 = { 2'h0, op_6 };
assign grp_fu_295_p0 = { select_ln850_5_reg_624[4], select_ln850_5_reg_624[4], select_ln850_5_reg_624[4], select_ln850_5_reg_624[4], select_ln850_5_reg_624[4], select_ln850_5_reg_624[4], select_ln850_5_reg_624, 6'h00 };
assign grp_fu_295_p1 = { ret_reg_619[9], ret_reg_619, 6'h00 };
assign grp_fu_305_p0 = { 1'h0, op_10 };
assign grp_fu_327_p0 = { 3'h0, add_ln69_reg_649 };
assign grp_fu_327_p1 = { op_21_V_reg_644[10], op_21_V_reg_644 };
assign grp_fu_348_p0 = { op_23_V_reg_664[11], op_23_V_reg_664[11], op_23_V_reg_664[11], op_23_V_reg_664[11], op_23_V_reg_664[11], op_23_V_reg_664[11], op_23_V_reg_664[11], op_23_V_reg_664[11], op_23_V_reg_664[11], op_23_V_reg_664[11], op_23_V_reg_664[11], op_23_V_reg_664[11], op_23_V_reg_664[11], op_23_V_reg_664[11], op_23_V_reg_664[11], op_23_V_reg_664[11], op_23_V_reg_664[11], op_23_V_reg_664[11], op_23_V_reg_664[11], op_23_V_reg_664[11], op_23_V_reg_664[11], op_23_V_reg_664, 1'h0 };
assign grp_fu_348_p1 = { op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12 };
assign grp_fu_395_p1 = { 31'h00000000, icmp_ln886_reg_614 };
assign grp_fu_424_p0 = { op_0[7], op_0[7:5] };
assign grp_fu_445_p0 = { op_25_V_reg_711[31], op_25_V_reg_711, 4'h0 };
assign grp_fu_445_p1 = { op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14 };
assign grp_fu_516_p0 = { 1'h0, op_16 };
assign grp_fu_516_p1 = { 1'h0, op_17_V_reg_765 };
assign grp_fu_549_p1 = { 24'h000000, op_15 };
assign grp_fu_557_p0 = { 3'h0, add_ln69_4_reg_790 };
assign grp_fu_557_p1 = { 1'h0, op_18 };
assign grp_fu_566_p0 = { 27'h0000000, add_ln69_5_reg_815 };
assign icmp_ln886_fu_244_p0 = op_4;
assign op_31 = grp_fu_566_p2;
assign op_9_V_fu_273_p3 = { ret_reg_619, 6'h00 };
assign p_Result_1_fu_471_p3 = op_0[7];
assign p_Result_2_fu_369_p3 = ret_V_12_reg_684[33];
assign p_Result_3_fu_522_p3 = ret_V_14_reg_753[36];
assign p_Result_s_fu_250_p3 = ret_V_11_reg_587[5];
assign ret_V_3_fu_400_p4 = op_0[7:5];
assign rhs_1_fu_284_p3 = { select_ln850_5_reg_624, 6'h00 };
assign rhs_4_fu_434_p3 = { op_25_V_reg_711, 4'h0 };
assign rhs_fu_197_p3 = { op_8, 1'h0 };
assign sext_ln215_fu_230_p0 = op_4;
assign sext_ln703_1_fu_333_p0 = op_12;
assign sext_ln703_2_fu_430_p0 = op_14;
assign sext_ln703_fu_193_p0 = op_2;
assign sext_ln835_fu_410_p1 = { op_0[7], op_0[7:5] };
assign sext_ln886_fu_490_p1 = { ret_V_5_fu_483_p3[3], ret_V_5_fu_483_p3[3], ret_V_5_fu_483_p3[3], ret_V_5_fu_483_p3[3], ret_V_5_fu_483_p3[3], ret_V_5_fu_483_p3 };
assign tmp_3_fu_337_p3 = { op_23_V_reg_664, 1'h0 };
assign trunc_ln851_1_fu_414_p1 = op_0[4:0];
assign trunc_ln851_2_fu_376_p0 = op_12;
assign trunc_ln851_2_fu_376_p1 = op_12[0];
assign trunc_ln851_3_fu_451_p0 = op_14;
assign trunc_ln851_3_fu_451_p1 = op_14[3:0];
assign trunc_ln851_fu_257_p0 = op_2;
assign trunc_ln851_fu_257_p1 = op_2[0];
assign zext_ln886_fu_494_p1 = { 1'h0, op_7 };
assign \sub_10s_10ns_10_2_1_U3.top_sub_10s_10ns_10_2_1_Adder_2_U.ain_s0  = \sub_10s_10ns_10_2_1_U3.top_sub_10s_10ns_10_2_1_Adder_2_U.a ;
assign \sub_10s_10ns_10_2_1_U3.top_sub_10s_10ns_10_2_1_Adder_2_U.s  = { \sub_10s_10ns_10_2_1_U3.top_sub_10s_10ns_10_2_1_Adder_2_U.fas_s2 , \sub_10s_10ns_10_2_1_U3.top_sub_10s_10ns_10_2_1_Adder_2_U.sum_s1  };
assign \sub_10s_10ns_10_2_1_U3.top_sub_10s_10ns_10_2_1_Adder_2_U.u2.a  = \sub_10s_10ns_10_2_1_U3.top_sub_10s_10ns_10_2_1_Adder_2_U.ain_s1 ;
assign \sub_10s_10ns_10_2_1_U3.top_sub_10s_10ns_10_2_1_Adder_2_U.u2.b  = \sub_10s_10ns_10_2_1_U3.top_sub_10s_10ns_10_2_1_Adder_2_U.bin_s1 ;
assign \sub_10s_10ns_10_2_1_U3.top_sub_10s_10ns_10_2_1_Adder_2_U.u2.cin  = \sub_10s_10ns_10_2_1_U3.top_sub_10s_10ns_10_2_1_Adder_2_U.carry_s1 ;
assign \sub_10s_10ns_10_2_1_U3.top_sub_10s_10ns_10_2_1_Adder_2_U.facout_s2  = \sub_10s_10ns_10_2_1_U3.top_sub_10s_10ns_10_2_1_Adder_2_U.u2.cout ;
assign \sub_10s_10ns_10_2_1_U3.top_sub_10s_10ns_10_2_1_Adder_2_U.fas_s2  = \sub_10s_10ns_10_2_1_U3.top_sub_10s_10ns_10_2_1_Adder_2_U.u2.s ;
assign \sub_10s_10ns_10_2_1_U3.top_sub_10s_10ns_10_2_1_Adder_2_U.u1.a  = \sub_10s_10ns_10_2_1_U3.top_sub_10s_10ns_10_2_1_Adder_2_U.a [4:0];
assign \sub_10s_10ns_10_2_1_U3.top_sub_10s_10ns_10_2_1_Adder_2_U.u1.b  = \sub_10s_10ns_10_2_1_U3.top_sub_10s_10ns_10_2_1_Adder_2_U.bin_s0 [4:0];
assign \sub_10s_10ns_10_2_1_U3.top_sub_10s_10ns_10_2_1_Adder_2_U.u1.cin  = 1'h1;
assign \sub_10s_10ns_10_2_1_U3.top_sub_10s_10ns_10_2_1_Adder_2_U.facout_s1  = \sub_10s_10ns_10_2_1_U3.top_sub_10s_10ns_10_2_1_Adder_2_U.u1.cout ;
assign \sub_10s_10ns_10_2_1_U3.top_sub_10s_10ns_10_2_1_Adder_2_U.fas_s1  = \sub_10s_10ns_10_2_1_U3.top_sub_10s_10ns_10_2_1_Adder_2_U.u1.s ;
assign \sub_10s_10ns_10_2_1_U3.top_sub_10s_10ns_10_2_1_Adder_2_U.a  = \sub_10s_10ns_10_2_1_U3.din0 ;
assign \sub_10s_10ns_10_2_1_U3.top_sub_10s_10ns_10_2_1_Adder_2_U.b  = \sub_10s_10ns_10_2_1_U3.din1 ;
assign \sub_10s_10ns_10_2_1_U3.top_sub_10s_10ns_10_2_1_Adder_2_U.ce  = \sub_10s_10ns_10_2_1_U3.ce ;
assign \sub_10s_10ns_10_2_1_U3.top_sub_10s_10ns_10_2_1_Adder_2_U.clk  = \sub_10s_10ns_10_2_1_U3.clk ;
assign \sub_10s_10ns_10_2_1_U3.top_sub_10s_10ns_10_2_1_Adder_2_U.reset  = \sub_10s_10ns_10_2_1_U3.reset ;
assign \sub_10s_10ns_10_2_1_U3.dout  = \sub_10s_10ns_10_2_1_U3.top_sub_10s_10ns_10_2_1_Adder_2_U.s ;
assign \sub_10s_10ns_10_2_1_U3.ce  = 1'h1;
assign \sub_10s_10ns_10_2_1_U3.clk  = ap_clk;
assign \sub_10s_10ns_10_2_1_U3.din0  = { op_4[7], op_4[7], op_4 };
assign \sub_10s_10ns_10_2_1_U3.din1  = { 2'h0, op_6 };
assign grp_fu_238_p2 = \sub_10s_10ns_10_2_1_U3.dout ;
assign \sub_10s_10ns_10_2_1_U3.reset  = ap_rst;
assign \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.ain_s0  = \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.a ;
assign \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.bin_s0  = \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.b ;
assign \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.s  = { \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.fas_s2 , \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.sum_s1  };
assign \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.u2.a  = \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.ain_s1 ;
assign \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.u2.b  = \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.bin_s1 ;
assign \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.u2.cin  = \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.carry_s1 ;
assign \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.facout_s2  = \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.u2.cout ;
assign \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.fas_s2  = \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.u2.s ;
assign \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.u1.a  = \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.a [3:0];
assign \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.u1.b  = \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.b [3:0];
assign \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.u1.cin  = 1'h0;
assign \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.facout_s1  = \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.u1.cout ;
assign \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.fas_s1  = \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.u1.s ;
assign \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.a  = \add_9ns_9ns_9_2_1_U5.din0 ;
assign \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.b  = \add_9ns_9ns_9_2_1_U5.din1 ;
assign \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.ce  = \add_9ns_9ns_9_2_1_U5.ce ;
assign \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.clk  = \add_9ns_9ns_9_2_1_U5.clk ;
assign \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.reset  = \add_9ns_9ns_9_2_1_U5.reset ;
assign \add_9ns_9ns_9_2_1_U5.dout  = \add_9ns_9ns_9_2_1_U5.top_add_9ns_9ns_9_2_1_Adder_4_U.s ;
assign \add_9ns_9ns_9_2_1_U5.ce  = 1'h1;
assign \add_9ns_9ns_9_2_1_U5.clk  = ap_clk;
assign \add_9ns_9ns_9_2_1_U5.din0  = { 1'h0, op_10 };
assign \add_9ns_9ns_9_2_1_U5.din1  = 9'h001;
assign grp_fu_305_p2 = \add_9ns_9ns_9_2_1_U5.dout ;
assign \add_9ns_9ns_9_2_1_U5.reset  = ap_rst;
assign \add_6s_6s_6_2_1_U1.top_add_6s_6s_6_2_1_Adder_0_U.ain_s0  = \add_6s_6s_6_2_1_U1.top_add_6s_6s_6_2_1_Adder_0_U.a ;
assign \add_6s_6s_6_2_1_U1.top_add_6s_6s_6_2_1_Adder_0_U.bin_s0  = \add_6s_6s_6_2_1_U1.top_add_6s_6s_6_2_1_Adder_0_U.b ;
assign \add_6s_6s_6_2_1_U1.top_add_6s_6s_6_2_1_Adder_0_U.s  = { \add_6s_6s_6_2_1_U1.top_add_6s_6s_6_2_1_Adder_0_U.fas_s2 , \add_6s_6s_6_2_1_U1.top_add_6s_6s_6_2_1_Adder_0_U.sum_s1  };
assign \add_6s_6s_6_2_1_U1.top_add_6s_6s_6_2_1_Adder_0_U.u2.a  = \add_6s_6s_6_2_1_U1.top_add_6s_6s_6_2_1_Adder_0_U.ain_s1 ;
assign \add_6s_6s_6_2_1_U1.top_add_6s_6s_6_2_1_Adder_0_U.u2.b  = \add_6s_6s_6_2_1_U1.top_add_6s_6s_6_2_1_Adder_0_U.bin_s1 ;
assign \add_6s_6s_6_2_1_U1.top_add_6s_6s_6_2_1_Adder_0_U.u2.cin  = \add_6s_6s_6_2_1_U1.top_add_6s_6s_6_2_1_Adder_0_U.carry_s1 ;
assign \add_6s_6s_6_2_1_U1.top_add_6s_6s_6_2_1_Adder_0_U.facout_s2  = \add_6s_6s_6_2_1_U1.top_add_6s_6s_6_2_1_Adder_0_U.u2.cout ;
assign \add_6s_6s_6_2_1_U1.top_add_6s_6s_6_2_1_Adder_0_U.fas_s2  = \add_6s_6s_6_2_1_U1.top_add_6s_6s_6_2_1_Adder_0_U.u2.s ;
assign \add_6s_6s_6_2_1_U1.top_add_6s_6s_6_2_1_Adder_0_U.u1.a  = \add_6s_6s_6_2_1_U1.top_add_6s_6s_6_2_1_Adder_0_U.a [2:0];
assign \add_6s_6s_6_2_1_U1.top_add_6s_6s_6_2_1_Adder_0_U.u1.b  = \add_6s_6s_6_2_1_U1.top_add_6s_6s_6_2_1_Adder_0_U.b [2:0];
assign \add_6s_6s_6_2_1_U1.top_add_6s_6s_6_2_1_Adder_0_U.u1.cin  = 1'h0;
assign \add_6s_6s_6_2_1_U1.top_add_6s_6s_6_2_1_Adder_0_U.facout_s1  = \add_6s_6s_6_2_1_U1.top_add_6s_6s_6_2_1_Adder_0_U.u1.cout ;
assign \add_6s_6s_6_2_1_U1.top_add_6s_6s_6_2_1_Adder_0_U.fas_s1  = \add_6s_6s_6_2_1_U1.top_add_6s_6s_6_2_1_Adder_0_U.u1.s ;
assign \add_6s_6s_6_2_1_U1.top_add_6s_6s_6_2_1_Adder_0_U.a  = \add_6s_6s_6_2_1_U1.din0 ;
assign \add_6s_6s_6_2_1_U1.top_add_6s_6s_6_2_1_Adder_0_U.b  = \add_6s_6s_6_2_1_U1.din1 ;
assign \add_6s_6s_6_2_1_U1.top_add_6s_6s_6_2_1_Adder_0_U.ce  = \add_6s_6s_6_2_1_U1.ce ;
assign \add_6s_6s_6_2_1_U1.top_add_6s_6s_6_2_1_Adder_0_U.clk  = \add_6s_6s_6_2_1_U1.clk ;
assign \add_6s_6s_6_2_1_U1.top_add_6s_6s_6_2_1_Adder_0_U.reset  = \add_6s_6s_6_2_1_U1.reset ;
assign \add_6s_6s_6_2_1_U1.dout  = \add_6s_6s_6_2_1_U1.top_add_6s_6s_6_2_1_Adder_0_U.s ;
assign \add_6s_6s_6_2_1_U1.ce  = 1'h1;
assign \add_6s_6s_6_2_1_U1.clk  = ap_clk;
assign \add_6s_6s_6_2_1_U1.din0  = { op_8[3], op_8, 1'h0 };
assign \add_6s_6s_6_2_1_U1.din1  = { op_2[3], op_2[3], op_2 };
assign grp_fu_209_p2 = \add_6s_6s_6_2_1_U1.dout ;
assign \add_6s_6s_6_2_1_U1.reset  = ap_rst;
assign \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.ain_s0  = \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.a ;
assign \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.bin_s0  = \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.b ;
assign \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.s  = { \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.fas_s2 , \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.sum_s1  };
assign \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.u2.a  = \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.ain_s1 ;
assign \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.u2.b  = \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.bin_s1 ;
assign \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.u2.cin  = \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.carry_s1 ;
assign \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.facout_s2  = \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.u2.cout ;
assign \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.fas_s2  = \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.u2.s ;
assign \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.u1.a  = \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.a [1:0];
assign \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.u1.b  = \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.b [1:0];
assign \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.u1.cin  = 1'h0;
assign \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.facout_s1  = \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.u1.cout ;
assign \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.fas_s1  = \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.u1.s ;
assign \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.a  = \add_5ns_5ns_5_2_1_U2.din0 ;
assign \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.b  = \add_5ns_5ns_5_2_1_U2.din1 ;
assign \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.ce  = \add_5ns_5ns_5_2_1_U2.ce ;
assign \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.clk  = \add_5ns_5ns_5_2_1_U2.clk ;
assign \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.reset  = \add_5ns_5ns_5_2_1_U2.reset ;
assign \add_5ns_5ns_5_2_1_U2.dout  = \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.s ;
assign \add_5ns_5ns_5_2_1_U2.ce  = 1'h1;
assign \add_5ns_5ns_5_2_1_U2.clk  = ap_clk;
assign \add_5ns_5ns_5_2_1_U2.din0  = ret_V_reg_592;
assign \add_5ns_5ns_5_2_1_U2.din1  = 5'h01;
assign grp_fu_225_p2 = \add_5ns_5ns_5_2_1_U2.dout ;
assign \add_5ns_5ns_5_2_1_U2.reset  = ap_rst;
assign \add_5ns_5ns_5_2_1_U15.top_add_5ns_5ns_5_2_1_Adder_1_U.ain_s0  = \add_5ns_5ns_5_2_1_U15.top_add_5ns_5ns_5_2_1_Adder_1_U.a ;
assign \add_5ns_5ns_5_2_1_U15.top_add_5ns_5ns_5_2_1_Adder_1_U.bin_s0  = \add_5ns_5ns_5_2_1_U15.top_add_5ns_5ns_5_2_1_Adder_1_U.b ;
assign \add_5ns_5ns_5_2_1_U15.top_add_5ns_5ns_5_2_1_Adder_1_U.s  = { \add_5ns_5ns_5_2_1_U15.top_add_5ns_5ns_5_2_1_Adder_1_U.fas_s2 , \add_5ns_5ns_5_2_1_U15.top_add_5ns_5ns_5_2_1_Adder_1_U.sum_s1  };
assign \add_5ns_5ns_5_2_1_U15.top_add_5ns_5ns_5_2_1_Adder_1_U.u2.a  = \add_5ns_5ns_5_2_1_U15.top_add_5ns_5ns_5_2_1_Adder_1_U.ain_s1 ;
assign \add_5ns_5ns_5_2_1_U15.top_add_5ns_5ns_5_2_1_Adder_1_U.u2.b  = \add_5ns_5ns_5_2_1_U15.top_add_5ns_5ns_5_2_1_Adder_1_U.bin_s1 ;
assign \add_5ns_5ns_5_2_1_U15.top_add_5ns_5ns_5_2_1_Adder_1_U.u2.cin  = \add_5ns_5ns_5_2_1_U15.top_add_5ns_5ns_5_2_1_Adder_1_U.carry_s1 ;
assign \add_5ns_5ns_5_2_1_U15.top_add_5ns_5ns_5_2_1_Adder_1_U.facout_s2  = \add_5ns_5ns_5_2_1_U15.top_add_5ns_5ns_5_2_1_Adder_1_U.u2.cout ;
assign \add_5ns_5ns_5_2_1_U15.top_add_5ns_5ns_5_2_1_Adder_1_U.fas_s2  = \add_5ns_5ns_5_2_1_U15.top_add_5ns_5ns_5_2_1_Adder_1_U.u2.s ;
assign \add_5ns_5ns_5_2_1_U15.top_add_5ns_5ns_5_2_1_Adder_1_U.u1.a  = \add_5ns_5ns_5_2_1_U15.top_add_5ns_5ns_5_2_1_Adder_1_U.a [1:0];
assign \add_5ns_5ns_5_2_1_U15.top_add_5ns_5ns_5_2_1_Adder_1_U.u1.b  = \add_5ns_5ns_5_2_1_U15.top_add_5ns_5ns_5_2_1_Adder_1_U.b [1:0];
assign \add_5ns_5ns_5_2_1_U15.top_add_5ns_5ns_5_2_1_Adder_1_U.u1.cin  = 1'h0;
assign \add_5ns_5ns_5_2_1_U15.top_add_5ns_5ns_5_2_1_Adder_1_U.facout_s1  = \add_5ns_5ns_5_2_1_U15.top_add_5ns_5ns_5_2_1_Adder_1_U.u1.cout ;
assign \add_5ns_5ns_5_2_1_U15.top_add_5ns_5ns_5_2_1_Adder_1_U.fas_s1  = \add_5ns_5ns_5_2_1_U15.top_add_5ns_5ns_5_2_1_Adder_1_U.u1.s ;
assign \add_5ns_5ns_5_2_1_U15.top_add_5ns_5ns_5_2_1_Adder_1_U.a  = \add_5ns_5ns_5_2_1_U15.din0 ;
assign \add_5ns_5ns_5_2_1_U15.top_add_5ns_5ns_5_2_1_Adder_1_U.b  = \add_5ns_5ns_5_2_1_U15.din1 ;
assign \add_5ns_5ns_5_2_1_U15.top_add_5ns_5ns_5_2_1_Adder_1_U.ce  = \add_5ns_5ns_5_2_1_U15.ce ;
assign \add_5ns_5ns_5_2_1_U15.top_add_5ns_5ns_5_2_1_Adder_1_U.clk  = \add_5ns_5ns_5_2_1_U15.clk ;
assign \add_5ns_5ns_5_2_1_U15.top_add_5ns_5ns_5_2_1_Adder_1_U.reset  = \add_5ns_5ns_5_2_1_U15.reset ;
assign \add_5ns_5ns_5_2_1_U15.dout  = \add_5ns_5ns_5_2_1_U15.top_add_5ns_5ns_5_2_1_Adder_1_U.s ;
assign \add_5ns_5ns_5_2_1_U15.ce  = 1'h1;
assign \add_5ns_5ns_5_2_1_U15.clk  = ap_clk;
assign \add_5ns_5ns_5_2_1_U15.din0  = { 3'h0, add_ln69_4_reg_790 };
assign \add_5ns_5ns_5_2_1_U15.din1  = { 1'h0, op_18 };
assign grp_fu_557_p2 = \add_5ns_5ns_5_2_1_U15.dout ;
assign \add_5ns_5ns_5_2_1_U15.reset  = ap_rst;
assign \add_4s_4ns_4_2_1_U10.top_add_4s_4ns_4_2_1_Adder_8_U.ain_s0  = \add_4s_4ns_4_2_1_U10.top_add_4s_4ns_4_2_1_Adder_8_U.a ;
assign \add_4s_4ns_4_2_1_U10.top_add_4s_4ns_4_2_1_Adder_8_U.bin_s0  = \add_4s_4ns_4_2_1_U10.top_add_4s_4ns_4_2_1_Adder_8_U.b ;
assign \add_4s_4ns_4_2_1_U10.top_add_4s_4ns_4_2_1_Adder_8_U.s  = { \add_4s_4ns_4_2_1_U10.top_add_4s_4ns_4_2_1_Adder_8_U.fas_s2 , \add_4s_4ns_4_2_1_U10.top_add_4s_4ns_4_2_1_Adder_8_U.sum_s1  };
assign \add_4s_4ns_4_2_1_U10.top_add_4s_4ns_4_2_1_Adder_8_U.u2.a  = \add_4s_4ns_4_2_1_U10.top_add_4s_4ns_4_2_1_Adder_8_U.ain_s1 ;
assign \add_4s_4ns_4_2_1_U10.top_add_4s_4ns_4_2_1_Adder_8_U.u2.b  = \add_4s_4ns_4_2_1_U10.top_add_4s_4ns_4_2_1_Adder_8_U.bin_s1 ;
assign \add_4s_4ns_4_2_1_U10.top_add_4s_4ns_4_2_1_Adder_8_U.u2.cin  = \add_4s_4ns_4_2_1_U10.top_add_4s_4ns_4_2_1_Adder_8_U.carry_s1 ;
assign \add_4s_4ns_4_2_1_U10.top_add_4s_4ns_4_2_1_Adder_8_U.facout_s2  = \add_4s_4ns_4_2_1_U10.top_add_4s_4ns_4_2_1_Adder_8_U.u2.cout ;
assign \add_4s_4ns_4_2_1_U10.top_add_4s_4ns_4_2_1_Adder_8_U.fas_s2  = \add_4s_4ns_4_2_1_U10.top_add_4s_4ns_4_2_1_Adder_8_U.u2.s ;
assign \add_4s_4ns_4_2_1_U10.top_add_4s_4ns_4_2_1_Adder_8_U.u1.a  = \add_4s_4ns_4_2_1_U10.top_add_4s_4ns_4_2_1_Adder_8_U.a [1:0];
assign \add_4s_4ns_4_2_1_U10.top_add_4s_4ns_4_2_1_Adder_8_U.u1.b  = \add_4s_4ns_4_2_1_U10.top_add_4s_4ns_4_2_1_Adder_8_U.b [1:0];
assign \add_4s_4ns_4_2_1_U10.top_add_4s_4ns_4_2_1_Adder_8_U.u1.cin  = 1'h0;
assign \add_4s_4ns_4_2_1_U10.top_add_4s_4ns_4_2_1_Adder_8_U.facout_s1  = \add_4s_4ns_4_2_1_U10.top_add_4s_4ns_4_2_1_Adder_8_U.u1.cout ;
assign \add_4s_4ns_4_2_1_U10.top_add_4s_4ns_4_2_1_Adder_8_U.fas_s1  = \add_4s_4ns_4_2_1_U10.top_add_4s_4ns_4_2_1_Adder_8_U.u1.s ;
assign \add_4s_4ns_4_2_1_U10.top_add_4s_4ns_4_2_1_Adder_8_U.a  = \add_4s_4ns_4_2_1_U10.din0 ;
assign \add_4s_4ns_4_2_1_U10.top_add_4s_4ns_4_2_1_Adder_8_U.b  = \add_4s_4ns_4_2_1_U10.din1 ;
assign \add_4s_4ns_4_2_1_U10.top_add_4s_4ns_4_2_1_Adder_8_U.ce  = \add_4s_4ns_4_2_1_U10.ce ;
assign \add_4s_4ns_4_2_1_U10.top_add_4s_4ns_4_2_1_Adder_8_U.clk  = \add_4s_4ns_4_2_1_U10.clk ;
assign \add_4s_4ns_4_2_1_U10.top_add_4s_4ns_4_2_1_Adder_8_U.reset  = \add_4s_4ns_4_2_1_U10.reset ;
assign \add_4s_4ns_4_2_1_U10.dout  = \add_4s_4ns_4_2_1_U10.top_add_4s_4ns_4_2_1_Adder_8_U.s ;
assign \add_4s_4ns_4_2_1_U10.ce  = 1'h1;
assign \add_4s_4ns_4_2_1_U10.clk  = ap_clk;
assign \add_4s_4ns_4_2_1_U10.din0  = { op_0[7], op_0[7:5] };
assign \add_4s_4ns_4_2_1_U10.din1  = 4'h1;
assign grp_fu_424_p2 = \add_4s_4ns_4_2_1_U10.dout ;
assign \add_4s_4ns_4_2_1_U10.reset  = ap_rst;
assign \add_37s_37s_37_2_1_U11.top_add_37s_37s_37_2_1_Adder_9_U.ain_s0  = \add_37s_37s_37_2_1_U11.top_add_37s_37s_37_2_1_Adder_9_U.a ;
assign \add_37s_37s_37_2_1_U11.top_add_37s_37s_37_2_1_Adder_9_U.bin_s0  = \add_37s_37s_37_2_1_U11.top_add_37s_37s_37_2_1_Adder_9_U.b ;
assign \add_37s_37s_37_2_1_U11.top_add_37s_37s_37_2_1_Adder_9_U.s  = { \add_37s_37s_37_2_1_U11.top_add_37s_37s_37_2_1_Adder_9_U.fas_s2 , \add_37s_37s_37_2_1_U11.top_add_37s_37s_37_2_1_Adder_9_U.sum_s1  };
assign \add_37s_37s_37_2_1_U11.top_add_37s_37s_37_2_1_Adder_9_U.u2.a  = \add_37s_37s_37_2_1_U11.top_add_37s_37s_37_2_1_Adder_9_U.ain_s1 ;
assign \add_37s_37s_37_2_1_U11.top_add_37s_37s_37_2_1_Adder_9_U.u2.b  = \add_37s_37s_37_2_1_U11.top_add_37s_37s_37_2_1_Adder_9_U.bin_s1 ;
assign \add_37s_37s_37_2_1_U11.top_add_37s_37s_37_2_1_Adder_9_U.u2.cin  = \add_37s_37s_37_2_1_U11.top_add_37s_37s_37_2_1_Adder_9_U.carry_s1 ;
assign \add_37s_37s_37_2_1_U11.top_add_37s_37s_37_2_1_Adder_9_U.facout_s2  = \add_37s_37s_37_2_1_U11.top_add_37s_37s_37_2_1_Adder_9_U.u2.cout ;
assign \add_37s_37s_37_2_1_U11.top_add_37s_37s_37_2_1_Adder_9_U.fas_s2  = \add_37s_37s_37_2_1_U11.top_add_37s_37s_37_2_1_Adder_9_U.u2.s ;
assign \add_37s_37s_37_2_1_U11.top_add_37s_37s_37_2_1_Adder_9_U.u1.a  = \add_37s_37s_37_2_1_U11.top_add_37s_37s_37_2_1_Adder_9_U.a [17:0];
assign \add_37s_37s_37_2_1_U11.top_add_37s_37s_37_2_1_Adder_9_U.u1.b  = \add_37s_37s_37_2_1_U11.top_add_37s_37s_37_2_1_Adder_9_U.b [17:0];
assign \add_37s_37s_37_2_1_U11.top_add_37s_37s_37_2_1_Adder_9_U.u1.cin  = 1'h0;
assign \add_37s_37s_37_2_1_U11.top_add_37s_37s_37_2_1_Adder_9_U.facout_s1  = \add_37s_37s_37_2_1_U11.top_add_37s_37s_37_2_1_Adder_9_U.u1.cout ;
assign \add_37s_37s_37_2_1_U11.top_add_37s_37s_37_2_1_Adder_9_U.fas_s1  = \add_37s_37s_37_2_1_U11.top_add_37s_37s_37_2_1_Adder_9_U.u1.s ;
assign \add_37s_37s_37_2_1_U11.top_add_37s_37s_37_2_1_Adder_9_U.a  = \add_37s_37s_37_2_1_U11.din0 ;
assign \add_37s_37s_37_2_1_U11.top_add_37s_37s_37_2_1_Adder_9_U.b  = \add_37s_37s_37_2_1_U11.din1 ;
assign \add_37s_37s_37_2_1_U11.top_add_37s_37s_37_2_1_Adder_9_U.ce  = \add_37s_37s_37_2_1_U11.ce ;
assign \add_37s_37s_37_2_1_U11.top_add_37s_37s_37_2_1_Adder_9_U.clk  = \add_37s_37s_37_2_1_U11.clk ;
assign \add_37s_37s_37_2_1_U11.top_add_37s_37s_37_2_1_Adder_9_U.reset  = \add_37s_37s_37_2_1_U11.reset ;
assign \add_37s_37s_37_2_1_U11.dout  = \add_37s_37s_37_2_1_U11.top_add_37s_37s_37_2_1_Adder_9_U.s ;
assign \add_37s_37s_37_2_1_U11.ce  = 1'h1;
assign \add_37s_37s_37_2_1_U11.clk  = ap_clk;
assign \add_37s_37s_37_2_1_U11.din0  = { op_25_V_reg_711[31], op_25_V_reg_711, 4'h0 };
assign \add_37s_37s_37_2_1_U11.din1  = { op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14[7], op_14 };
assign grp_fu_445_p2 = \add_37s_37s_37_2_1_U11.dout ;
assign \add_37s_37s_37_2_1_U11.reset  = ap_rst;
assign \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_6_U.ain_s0  = \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_6_U.a ;
assign \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_6_U.bin_s0  = \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_6_U.b ;
assign \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_6_U.s  = { \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_6_U.fas_s2 , \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_6_U.sum_s1  };
assign \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_6_U.u2.a  = \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_6_U.ain_s1 ;
assign \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_6_U.u2.b  = \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_6_U.bin_s1 ;
assign \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_6_U.u2.cin  = \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_6_U.carry_s1 ;
assign \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_6_U.facout_s2  = \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_6_U.u2.cout ;
assign \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_6_U.fas_s2  = \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_6_U.u2.s ;
assign \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_6_U.u1.a  = \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_6_U.a [16:0];
assign \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_6_U.u1.b  = \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_6_U.b [16:0];
assign \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_6_U.u1.cin  = 1'h0;
assign \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_6_U.facout_s1  = \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_6_U.u1.cout ;
assign \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_6_U.fas_s1  = \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_6_U.u1.s ;
assign \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_6_U.a  = \add_34s_34s_34_2_1_U7.din0 ;
assign \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_6_U.b  = \add_34s_34s_34_2_1_U7.din1 ;
assign \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_6_U.ce  = \add_34s_34s_34_2_1_U7.ce ;
assign \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_6_U.clk  = \add_34s_34s_34_2_1_U7.clk ;
assign \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_6_U.reset  = \add_34s_34s_34_2_1_U7.reset ;
assign \add_34s_34s_34_2_1_U7.dout  = \add_34s_34s_34_2_1_U7.top_add_34s_34s_34_2_1_Adder_6_U.s ;
assign \add_34s_34s_34_2_1_U7.ce  = 1'h1;
assign \add_34s_34s_34_2_1_U7.clk  = ap_clk;
assign \add_34s_34s_34_2_1_U7.din0  = { op_23_V_reg_664[11], op_23_V_reg_664[11], op_23_V_reg_664[11], op_23_V_reg_664[11], op_23_V_reg_664[11], op_23_V_reg_664[11], op_23_V_reg_664[11], op_23_V_reg_664[11], op_23_V_reg_664[11], op_23_V_reg_664[11], op_23_V_reg_664[11], op_23_V_reg_664[11], op_23_V_reg_664[11], op_23_V_reg_664[11], op_23_V_reg_664[11], op_23_V_reg_664[11], op_23_V_reg_664[11], op_23_V_reg_664[11], op_23_V_reg_664[11], op_23_V_reg_664[11], op_23_V_reg_664[11], op_23_V_reg_664, 1'h0 };
assign \add_34s_34s_34_2_1_U7.din1  = { op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12 };
assign grp_fu_348_p2 = \add_34s_34s_34_2_1_U7.dout ;
assign \add_34s_34s_34_2_1_U7.reset  = ap_rst;
assign \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s0  = \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.a ;
assign \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s0  = \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.b ;
assign \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.s  = { \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s2 , \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.sum_s1  };
assign \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.a  = \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s1 ;
assign \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.b  = \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s1 ;
assign \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cin  = \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.carry_s1 ;
assign \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.facout_s2  = \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cout ;
assign \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s2  = \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.s ;
assign \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.a  = \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.a [15:0];
assign \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.b  = \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.b [15:0];
assign \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cin  = 1'h0;
assign \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.facout_s1  = \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cout ;
assign \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s1  = \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.s ;
assign \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.a  = \add_32ns_32ns_32_2_1_U9.din0 ;
assign \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.b  = \add_32ns_32ns_32_2_1_U9.din1 ;
assign \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.ce  = \add_32ns_32ns_32_2_1_U9.ce ;
assign \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.clk  = \add_32ns_32ns_32_2_1_U9.clk ;
assign \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.reset  = \add_32ns_32ns_32_2_1_U9.reset ;
assign \add_32ns_32ns_32_2_1_U9.dout  = \add_32ns_32ns_32_2_1_U9.top_add_32ns_32ns_32_2_1_Adder_7_U.s ;
assign \add_32ns_32ns_32_2_1_U9.ce  = 1'h1;
assign \add_32ns_32ns_32_2_1_U9.clk  = ap_clk;
assign \add_32ns_32ns_32_2_1_U9.din0  = ret_V_13_reg_701;
assign \add_32ns_32ns_32_2_1_U9.din1  = { 31'h00000000, icmp_ln886_reg_614 };
assign grp_fu_395_p2 = \add_32ns_32ns_32_2_1_U9.dout ;
assign \add_32ns_32ns_32_2_1_U9.reset  = ap_rst;
assign \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s0  = \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_7_U.a ;
assign \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s0  = \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_7_U.b ;
assign \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_7_U.s  = { \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s2 , \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_7_U.sum_s1  };
assign \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.a  = \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s1 ;
assign \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.b  = \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s1 ;
assign \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cin  = \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_7_U.carry_s1 ;
assign \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_7_U.facout_s2  = \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cout ;
assign \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s2  = \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.s ;
assign \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.a  = \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_7_U.a [15:0];
assign \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.b  = \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_7_U.b [15:0];
assign \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cin  = 1'h0;
assign \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_7_U.facout_s1  = \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cout ;
assign \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s1  = \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.s ;
assign \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_7_U.a  = \add_32ns_32ns_32_2_1_U8.din0 ;
assign \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_7_U.b  = \add_32ns_32ns_32_2_1_U8.din1 ;
assign \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_7_U.ce  = \add_32ns_32ns_32_2_1_U8.ce ;
assign \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_7_U.clk  = \add_32ns_32ns_32_2_1_U8.clk ;
assign \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_7_U.reset  = \add_32ns_32ns_32_2_1_U8.reset ;
assign \add_32ns_32ns_32_2_1_U8.dout  = \add_32ns_32ns_32_2_1_U8.top_add_32ns_32ns_32_2_1_Adder_7_U.s ;
assign \add_32ns_32ns_32_2_1_U8.ce  = 1'h1;
assign \add_32ns_32ns_32_2_1_U8.clk  = ap_clk;
assign \add_32ns_32ns_32_2_1_U8.din0  = ret_V_8_cast_reg_689;
assign \add_32ns_32ns_32_2_1_U8.din1  = 32'd1;
assign grp_fu_364_p2 = \add_32ns_32ns_32_2_1_U8.dout ;
assign \add_32ns_32ns_32_2_1_U8.reset  = ap_rst;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s0  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.a ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s0  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.b ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.s  = { \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s2 , \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.sum_s1  };
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.a  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s1 ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.b  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s1 ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cin  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.carry_s1 ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.facout_s2  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cout ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s2  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.s ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.a  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.a [15:0];
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.b  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.b [15:0];
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cin  = 1'h0;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.facout_s1  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cout ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s1  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.s ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.a  = \add_32ns_32ns_32_2_1_U16.din0 ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.b  = \add_32ns_32ns_32_2_1_U16.din1 ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.ce  = \add_32ns_32ns_32_2_1_U16.ce ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.clk  = \add_32ns_32ns_32_2_1_U16.clk ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.reset  = \add_32ns_32ns_32_2_1_U16.reset ;
assign \add_32ns_32ns_32_2_1_U16.dout  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_7_U.s ;
assign \add_32ns_32ns_32_2_1_U16.ce  = 1'h1;
assign \add_32ns_32ns_32_2_1_U16.clk  = ap_clk;
assign \add_32ns_32ns_32_2_1_U16.din0  = { 27'h0000000, add_ln69_5_reg_815 };
assign \add_32ns_32ns_32_2_1_U16.din1  = add_ln69_3_reg_810;
assign grp_fu_566_p2 = \add_32ns_32ns_32_2_1_U16.dout ;
assign \add_32ns_32ns_32_2_1_U16.reset  = ap_rst;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s0  = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.a ;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s0  = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.b ;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.s  = { \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s2 , \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.sum_s1  };
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.a  = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s1 ;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.b  = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s1 ;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cin  = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.carry_s1 ;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.facout_s2  = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cout ;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s2  = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.s ;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.a  = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.a [15:0];
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.b  = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.b [15:0];
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cin  = 1'h0;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.facout_s1  = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cout ;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s1  = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.s ;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.a  = \add_32ns_32ns_32_2_1_U14.din0 ;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.b  = \add_32ns_32ns_32_2_1_U14.din1 ;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.ce  = \add_32ns_32ns_32_2_1_U14.ce ;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.clk  = \add_32ns_32ns_32_2_1_U14.clk ;
assign \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.reset  = \add_32ns_32ns_32_2_1_U14.reset ;
assign \add_32ns_32ns_32_2_1_U14.dout  = \add_32ns_32ns_32_2_1_U14.top_add_32ns_32ns_32_2_1_Adder_7_U.s ;
assign \add_32ns_32ns_32_2_1_U14.ce  = 1'h1;
assign \add_32ns_32ns_32_2_1_U14.clk  = ap_clk;
assign \add_32ns_32ns_32_2_1_U14.din0  = ret_V_15_reg_785;
assign \add_32ns_32ns_32_2_1_U14.din1  = { 24'h000000, op_15 };
assign grp_fu_549_p2 = \add_32ns_32ns_32_2_1_U14.dout ;
assign \add_32ns_32ns_32_2_1_U14.reset  = ap_rst;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s0  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.a ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s0  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.b ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.s  = { \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s2 , \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.sum_s1  };
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.a  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.ain_s1 ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.b  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.bin_s1 ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cin  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.carry_s1 ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.facout_s2  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.cout ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s2  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.u2.s ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.a  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.a [15:0];
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.b  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.b [15:0];
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cin  = 1'h0;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.facout_s1  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.cout ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.fas_s1  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.u1.s ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.a  = \add_32ns_32ns_32_2_1_U12.din0 ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.b  = \add_32ns_32ns_32_2_1_U12.din1 ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.ce  = \add_32ns_32ns_32_2_1_U12.ce ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.clk  = \add_32ns_32ns_32_2_1_U12.clk ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.reset  = \add_32ns_32ns_32_2_1_U12.reset ;
assign \add_32ns_32ns_32_2_1_U12.dout  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_7_U.s ;
assign \add_32ns_32ns_32_2_1_U12.ce  = 1'h1;
assign \add_32ns_32ns_32_2_1_U12.clk  = ap_clk;
assign \add_32ns_32ns_32_2_1_U12.din0  = ret_V_19_cast_reg_758;
assign \add_32ns_32ns_32_2_1_U12.din1  = 32'd1;
assign grp_fu_504_p2 = \add_32ns_32ns_32_2_1_U12.dout ;
assign \add_32ns_32ns_32_2_1_U12.reset  = ap_rst;
assign \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_10_U.ain_s0  = \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_10_U.a ;
assign \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_10_U.bin_s0  = \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_10_U.b ;
assign \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_10_U.s  = { \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_10_U.fas_s2 , \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_10_U.sum_s1  };
assign \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_10_U.u2.a  = \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_10_U.ain_s1 ;
assign \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_10_U.u2.b  = \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_10_U.bin_s1 ;
assign \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_10_U.u2.cin  = \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_10_U.carry_s1 ;
assign \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_10_U.facout_s2  = \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_10_U.u2.cout ;
assign \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_10_U.fas_s2  = \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_10_U.u2.s ;
assign \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_10_U.u1.a  = \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_10_U.a [0];
assign \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_10_U.u1.b  = \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_10_U.b [0];
assign \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_10_U.u1.cin  = 1'h0;
assign \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_10_U.facout_s1  = \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_10_U.u1.cout ;
assign \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_10_U.fas_s1  = \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_10_U.u1.s ;
assign \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_10_U.a  = \add_2ns_2ns_2_2_1_U13.din0 ;
assign \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_10_U.b  = \add_2ns_2ns_2_2_1_U13.din1 ;
assign \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_10_U.ce  = \add_2ns_2ns_2_2_1_U13.ce ;
assign \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_10_U.clk  = \add_2ns_2ns_2_2_1_U13.clk ;
assign \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_10_U.reset  = \add_2ns_2ns_2_2_1_U13.reset ;
assign \add_2ns_2ns_2_2_1_U13.dout  = \add_2ns_2ns_2_2_1_U13.top_add_2ns_2ns_2_2_1_Adder_10_U.s ;
assign \add_2ns_2ns_2_2_1_U13.ce  = 1'h1;
assign \add_2ns_2ns_2_2_1_U13.clk  = ap_clk;
assign \add_2ns_2ns_2_2_1_U13.din0  = { 1'h0, op_16 };
assign \add_2ns_2ns_2_2_1_U13.din1  = { 1'h0, op_17_V_reg_765 };
assign grp_fu_516_p2 = \add_2ns_2ns_2_2_1_U13.dout ;
assign \add_2ns_2ns_2_2_1_U13.reset  = ap_rst;
assign \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.ain_s0  = \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.a ;
assign \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.bin_s0  = \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.b ;
assign \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.s  = { \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.fas_s2 , \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.sum_s1  };
assign \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.u2.a  = \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.ain_s1 ;
assign \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.u2.b  = \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.bin_s1 ;
assign \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.u2.cin  = \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.carry_s1 ;
assign \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.facout_s2  = \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.u2.cout ;
assign \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.fas_s2  = \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.u2.s ;
assign \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.u1.a  = \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.a [7:0];
assign \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.u1.b  = \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.b [7:0];
assign \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.u1.cin  = 1'h0;
assign \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.facout_s1  = \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.u1.cout ;
assign \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.fas_s1  = \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.u1.s ;
assign \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.a  = \add_17s_17s_17_2_1_U4.din0 ;
assign \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.b  = \add_17s_17s_17_2_1_U4.din1 ;
assign \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.ce  = \add_17s_17s_17_2_1_U4.ce ;
assign \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.clk  = \add_17s_17s_17_2_1_U4.clk ;
assign \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.reset  = \add_17s_17s_17_2_1_U4.reset ;
assign \add_17s_17s_17_2_1_U4.dout  = \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.s ;
assign \add_17s_17s_17_2_1_U4.ce  = 1'h1;
assign \add_17s_17s_17_2_1_U4.clk  = ap_clk;
assign \add_17s_17s_17_2_1_U4.din0  = { select_ln850_5_reg_624[4], select_ln850_5_reg_624[4], select_ln850_5_reg_624[4], select_ln850_5_reg_624[4], select_ln850_5_reg_624[4], select_ln850_5_reg_624[4], select_ln850_5_reg_624, 6'h00 };
assign \add_17s_17s_17_2_1_U4.din1  = { ret_reg_619[9], ret_reg_619, 6'h00 };
assign grp_fu_295_p2 = \add_17s_17s_17_2_1_U4.dout ;
assign \add_17s_17s_17_2_1_U4.reset  = ap_rst;
assign \add_12ns_12s_12_2_1_U6.top_add_12ns_12s_12_2_1_Adder_5_U.ain_s0  = \add_12ns_12s_12_2_1_U6.top_add_12ns_12s_12_2_1_Adder_5_U.a ;
assign \add_12ns_12s_12_2_1_U6.top_add_12ns_12s_12_2_1_Adder_5_U.bin_s0  = \add_12ns_12s_12_2_1_U6.top_add_12ns_12s_12_2_1_Adder_5_U.b ;
assign \add_12ns_12s_12_2_1_U6.top_add_12ns_12s_12_2_1_Adder_5_U.s  = { \add_12ns_12s_12_2_1_U6.top_add_12ns_12s_12_2_1_Adder_5_U.fas_s2 , \add_12ns_12s_12_2_1_U6.top_add_12ns_12s_12_2_1_Adder_5_U.sum_s1  };
assign \add_12ns_12s_12_2_1_U6.top_add_12ns_12s_12_2_1_Adder_5_U.u2.a  = \add_12ns_12s_12_2_1_U6.top_add_12ns_12s_12_2_1_Adder_5_U.ain_s1 ;
assign \add_12ns_12s_12_2_1_U6.top_add_12ns_12s_12_2_1_Adder_5_U.u2.b  = \add_12ns_12s_12_2_1_U6.top_add_12ns_12s_12_2_1_Adder_5_U.bin_s1 ;
assign \add_12ns_12s_12_2_1_U6.top_add_12ns_12s_12_2_1_Adder_5_U.u2.cin  = \add_12ns_12s_12_2_1_U6.top_add_12ns_12s_12_2_1_Adder_5_U.carry_s1 ;
assign \add_12ns_12s_12_2_1_U6.top_add_12ns_12s_12_2_1_Adder_5_U.facout_s2  = \add_12ns_12s_12_2_1_U6.top_add_12ns_12s_12_2_1_Adder_5_U.u2.cout ;
assign \add_12ns_12s_12_2_1_U6.top_add_12ns_12s_12_2_1_Adder_5_U.fas_s2  = \add_12ns_12s_12_2_1_U6.top_add_12ns_12s_12_2_1_Adder_5_U.u2.s ;
assign \add_12ns_12s_12_2_1_U6.top_add_12ns_12s_12_2_1_Adder_5_U.u1.a  = \add_12ns_12s_12_2_1_U6.top_add_12ns_12s_12_2_1_Adder_5_U.a [5:0];
assign \add_12ns_12s_12_2_1_U6.top_add_12ns_12s_12_2_1_Adder_5_U.u1.b  = \add_12ns_12s_12_2_1_U6.top_add_12ns_12s_12_2_1_Adder_5_U.b [5:0];
assign \add_12ns_12s_12_2_1_U6.top_add_12ns_12s_12_2_1_Adder_5_U.u1.cin  = 1'h0;
assign \add_12ns_12s_12_2_1_U6.top_add_12ns_12s_12_2_1_Adder_5_U.facout_s1  = \add_12ns_12s_12_2_1_U6.top_add_12ns_12s_12_2_1_Adder_5_U.u1.cout ;
assign \add_12ns_12s_12_2_1_U6.top_add_12ns_12s_12_2_1_Adder_5_U.fas_s1  = \add_12ns_12s_12_2_1_U6.top_add_12ns_12s_12_2_1_Adder_5_U.u1.s ;
assign \add_12ns_12s_12_2_1_U6.top_add_12ns_12s_12_2_1_Adder_5_U.a  = \add_12ns_12s_12_2_1_U6.din0 ;
assign \add_12ns_12s_12_2_1_U6.top_add_12ns_12s_12_2_1_Adder_5_U.b  = \add_12ns_12s_12_2_1_U6.din1 ;
assign \add_12ns_12s_12_2_1_U6.top_add_12ns_12s_12_2_1_Adder_5_U.ce  = \add_12ns_12s_12_2_1_U6.ce ;
assign \add_12ns_12s_12_2_1_U6.top_add_12ns_12s_12_2_1_Adder_5_U.clk  = \add_12ns_12s_12_2_1_U6.clk ;
assign \add_12ns_12s_12_2_1_U6.top_add_12ns_12s_12_2_1_Adder_5_U.reset  = \add_12ns_12s_12_2_1_U6.reset ;
assign \add_12ns_12s_12_2_1_U6.dout  = \add_12ns_12s_12_2_1_U6.top_add_12ns_12s_12_2_1_Adder_5_U.s ;
assign \add_12ns_12s_12_2_1_U6.ce  = 1'h1;
assign \add_12ns_12s_12_2_1_U6.clk  = ap_clk;
assign \add_12ns_12s_12_2_1_U6.din0  = { 3'h0, add_ln69_reg_649 };
assign \add_12ns_12s_12_2_1_U6.din1  = { op_21_V_reg_644[10], op_21_V_reg_644 };
assign grp_fu_327_p2 = \add_12ns_12s_12_2_1_U6.dout ;
assign \add_12ns_12s_12_2_1_U6.reset  = ap_rst;
endmodule


// Product machine:
module top_A_times_top_B (ap_start, op_0, op_10, op_12, op_14, op_15, op_16, op_18, op_2, op_4, op_6, op_7, op_8, ap_clk, unsafe_signal);
input ap_start;
input [7:0] op_0;
input [7:0] op_10;
input [1:0] op_12;
input [7:0] op_14;
input [7:0] op_15;
input op_16;
input [3:0] op_18;
input [3:0] op_2;
input [7:0] op_4;
input [7:0] op_6;
input [7:0] op_7;
input [3:0] op_8;
input ap_clk;
output unsafe_signal;
reg _setup;
initial _setup = 1'b0;
always @ (posedge ap_clk) _setup <= 1'b1;
reg ap_start_internal;
always @ (posedge ap_clk) if (!_setup) ap_start_internal <= ap_start;
reg [7:0] op_0_internal;
always @ (posedge ap_clk) if (!_setup) op_0_internal <= op_0;
reg [7:0] op_10_internal;
always @ (posedge ap_clk) if (!_setup) op_10_internal <= op_10;
reg [1:0] op_12_internal;
always @ (posedge ap_clk) if (!_setup) op_12_internal <= op_12;
reg [7:0] op_14_internal;
always @ (posedge ap_clk) if (!_setup) op_14_internal <= op_14;
reg [7:0] op_15_internal;
always @ (posedge ap_clk) if (!_setup) op_15_internal <= op_15;
reg op_16_internal;
always @ (posedge ap_clk) if (!_setup) op_16_internal <= op_16;
reg [3:0] op_18_internal;
always @ (posedge ap_clk) if (!_setup) op_18_internal <= op_18;
reg [3:0] op_2_internal;
always @ (posedge ap_clk) if (!_setup) op_2_internal <= op_2;
reg [7:0] op_4_internal;
always @ (posedge ap_clk) if (!_setup) op_4_internal <= op_4;
reg [7:0] op_6_internal;
always @ (posedge ap_clk) if (!_setup) op_6_internal <= op_6;
reg [7:0] op_7_internal;
always @ (posedge ap_clk) if (!_setup) op_7_internal <= op_7;
reg [3:0] op_8_internal;
always @ (posedge ap_clk) if (!_setup) op_8_internal <= op_8;
wire ap_done_A;
wire ap_done_B;
wire ap_done_eq;
assign ap_done_eq = ap_done_A == ap_done_B;
wire ap_idle_A;
wire ap_idle_B;
wire ap_idle_eq;
assign ap_idle_eq = ap_idle_A == ap_idle_B;
wire ap_ready_A;
wire ap_ready_B;
wire ap_ready_eq;
assign ap_ready_eq = ap_ready_A == ap_ready_B;
wire [31:0] op_31_A;
wire [31:0] op_31_B;
wire op_31_eq;
assign op_31_eq = op_31_A == op_31_B;
wire op_31_ap_vld_A;
wire op_31_ap_vld_B;
wire clk_enable_A;
wire clk_enable_B;
assign clk_enable_A = _setup & (~op_31_ap_vld_A | op_31_ap_vld_B);
assign clk_enable_B = _setup;
wire divergent;
assign divergent = ~(ap_done_eq & ap_idle_eq & ap_ready_eq & op_31_eq);
assign unsafe_signal = op_31_ap_vld_A & op_31_ap_vld_B & divergent;
top_A instance_A (
    .ap_clk(ap_clk),
    .clk_enable(clk_enable_A),
    .ap_start(ap_start_internal),
    .op_0(op_0_internal),
    .op_10(op_10_internal),
    .op_12(op_12_internal),
    .op_14(op_14_internal),
    .op_15(op_15_internal),
    .op_16(op_16_internal),
    .op_18(op_18_internal),
    .op_2(op_2_internal),
    .op_4(op_4_internal),
    .op_6(op_6_internal),
    .op_7(op_7_internal),
    .op_8(op_8_internal),
    .ap_done(ap_done_A),
    .ap_idle(ap_idle_A),
    .ap_ready(ap_ready_A),
    .op_31(op_31_A),
    .op_31_ap_vld(op_31_ap_vld_A)
);
top_B instance_B (
    .ap_clk(ap_clk),
    .clk_enable(clk_enable_B),
    .ap_start(ap_start_internal),
    .op_0(op_0_internal),
    .op_10(op_10_internal),
    .op_12(op_12_internal),
    .op_14(op_14_internal),
    .op_15(op_15_internal),
    .op_16(op_16_internal),
    .op_18(op_18_internal),
    .op_2(op_2_internal),
    .op_4(op_4_internal),
    .op_6(op_6_internal),
    .op_7(op_7_internal),
    .op_8(op_8_internal),
    .ap_done(ap_done_B),
    .ap_idle(ap_idle_B),
    .ap_ready(ap_ready_B),
    .op_31(op_31_B),
    .op_31_ap_vld(op_31_ap_vld_B)
);
endmodule
