// Processed by function `construct_kairos` in `verilog_tricks.py`.
// Machine A:
// Processed by function `add_clk_enable_signal` in `verilog_tricks.py`.
// Processed by function `remove_reset_signal` in `verilog_tricks.py`.
module top_A (
  ap_clk,
  ap_start,
  ap_done,
  ap_idle,
  ap_ready,
  op_0,
  op_1,
  op_5,
  op_6,
  op_10,
  op_11,
  op_12,
  op_13,
  op_14,
  op_15,
  op_16,
  op_17,
  op_18,
  op_30,
  op_30_ap_vld,
clk_enable
);
input clk_enable;


input ap_clk;
wire ap_rst;
assign ap_rst = op_30_ap_vld;
input ap_start;
input [1:0] op_0;
input [3:0] op_1;
input [3:0] op_10;
input op_11;
input [3:0] op_12;
input [7:0] op_13;
input [3:0] op_14;
input op_15;
input [15:0] op_16;
input [3:0] op_17;
input op_18;
input [3:0] op_5;
input [7:0] op_6;
output ap_done;
output ap_idle;
output ap_ready;
output [31:0] op_30;
output op_30_ap_vld;


reg [4:0] \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.ain_s1 ;
reg [4:0] \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.bin_s1 ;
reg \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.carry_s1 ;
reg [4:0] \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.sum_s1 ;
reg [4:0] \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.ain_s1 ;
reg [4:0] \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.bin_s1 ;
reg \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.carry_s1 ;
reg [4:0] \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.sum_s1 ;
reg [5:0] \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.ain_s1 ;
reg [5:0] \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.bin_s1 ;
reg \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.carry_s1 ;
reg [5:0] \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.sum_s1 ;
reg [8:0] \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.ain_s1 ;
reg [8:0] \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.bin_s1 ;
reg \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.carry_s1 ;
reg [7:0] \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.sum_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.ain_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.bin_s1 ;
reg \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.carry_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.sum_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.ain_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.bin_s1 ;
reg \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.carry_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.sum_s1 ;
reg [15:0] \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.ain_s1 ;
reg [15:0] \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.bin_s1 ;
reg \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.carry_s1 ;
reg [15:0] \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.sum_s1 ;
reg [15:0] \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.ain_s1 ;
reg [15:0] \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.bin_s1 ;
reg \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.carry_s1 ;
reg [15:0] \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.sum_s1 ;
reg [17:0] \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.ain_s1 ;
reg [17:0] \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.bin_s1 ;
reg \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.carry_s1 ;
reg [16:0] \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.sum_s1 ;
reg [2:0] \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.ain_s1 ;
reg [2:0] \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.bin_s1 ;
reg \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.carry_s1 ;
reg [1:0] \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.sum_s1 ;
reg [2:0] \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.ain_s1 ;
reg [2:0] \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.bin_s1 ;
reg \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.carry_s1 ;
reg [2:0] \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.sum_s1 ;
reg [4:0] \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.ain_s1 ;
reg [4:0] \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.bin_s1 ;
reg \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.carry_s1 ;
reg [3:0] \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.sum_s1 ;
reg [31:0] add_ln691_1_reg_504;
reg [9:0] add_ln691_reg_452;
reg [31:0] add_ln69_1_reg_554;
reg [4:0] add_ln69_2_reg_534;
reg [5:0] add_ln69_3_reg_559;
reg [16:0] add_ln69_reg_529;
reg [20:0] ap_CS_fsm = 21'h000001;
reg icmp_ln851_1_reg_482;
reg icmp_ln851_reg_430;
reg [9:0] op_22_V_reg_467;
reg [31:0] op_28_V_reg_569;
reg [9:0] ret_V_1_reg_457;
reg [34:0] ret_V_2_reg_487;
reg [31:0] ret_V_3_cast_reg_492;
reg [31:0] ret_V_3_reg_524;
reg [11:0] ret_V_reg_435;
reg [8:0] ret_reg_415;
reg [31:0] select_ln1192_reg_574;
reg [8:0] select_ln215_reg_405;
reg [4:0] select_ln69_1_reg_499;
reg [9:0] select_ln69_reg_462;
reg [9:0] sext_ln850_reg_445;
reg [8:0] tmp_1_reg_440;
wire [31:0] _000_;
wire [9:0] _001_;
wire [31:0] _002_;
wire [4:0] _003_;
wire [5:0] _004_;
wire [16:0] _005_;
wire [20:0] _006_;
wire _007_;
wire _008_;
wire [9:0] _009_;
wire [31:0] _010_;
wire [9:0] _011_;
wire [34:0] _012_;
wire [31:0] _013_;
wire [31:0] _014_;
wire [11:0] _015_;
wire [8:0] _016_;
wire [31:0] _017_;
wire [8:0] _018_;
wire [4:0] _019_;
wire [9:0] _020_;
wire [9:0] _021_;
wire [8:0] _022_;
wire [1:0] _023_;
wire _024_;
wire _025_;
wire _026_;
wire _027_;
wire _028_;
wire [4:0] _029_;
wire [4:0] _030_;
wire _031_;
wire [4:0] _032_;
wire [5:0] _033_;
wire [5:0] _034_;
wire [4:0] _035_;
wire [4:0] _036_;
wire _037_;
wire [4:0] _038_;
wire [5:0] _039_;
wire [5:0] _040_;
wire [5:0] _041_;
wire [5:0] _042_;
wire _043_;
wire [5:0] _044_;
wire [6:0] _045_;
wire [6:0] _046_;
wire [8:0] _047_;
wire [8:0] _048_;
wire _049_;
wire [7:0] _050_;
wire [8:0] _051_;
wire [9:0] _052_;
wire [15:0] _053_;
wire [15:0] _054_;
wire _055_;
wire [15:0] _056_;
wire [16:0] _057_;
wire [16:0] _058_;
wire [15:0] _059_;
wire [15:0] _060_;
wire _061_;
wire [15:0] _062_;
wire [16:0] _063_;
wire [16:0] _064_;
wire [15:0] _065_;
wire [15:0] _066_;
wire _067_;
wire [15:0] _068_;
wire [16:0] _069_;
wire [16:0] _070_;
wire [15:0] _071_;
wire [15:0] _072_;
wire _073_;
wire [15:0] _074_;
wire [16:0] _075_;
wire [16:0] _076_;
wire [17:0] _077_;
wire [17:0] _078_;
wire _079_;
wire [16:0] _080_;
wire [17:0] _081_;
wire [18:0] _082_;
wire [2:0] _083_;
wire [2:0] _084_;
wire _085_;
wire [1:0] _086_;
wire [2:0] _087_;
wire [3:0] _088_;
wire [2:0] _089_;
wire [2:0] _090_;
wire _091_;
wire [2:0] _092_;
wire [3:0] _093_;
wire [3:0] _094_;
wire [4:0] _095_;
wire [4:0] _096_;
wire _097_;
wire [3:0] _098_;
wire [4:0] _099_;
wire [5:0] _100_;
wire _101_;
wire _102_;
wire _103_;
wire _104_;
wire _105_;
wire _106_;
wire _107_;
wire _108_;
wire _109_;
wire _110_;
wire _111_;
wire _112_;
wire _113_;
wire _114_;
wire _115_;
wire _116_;
wire _117_;
wire _118_;
wire _119_;
wire _120_;
wire _121_;
wire _122_;
wire _123_;
wire \add_10ns_10ns_10_2_1_U4.ce ;
wire \add_10ns_10ns_10_2_1_U4.clk ;
wire [9:0] \add_10ns_10ns_10_2_1_U4.din0 ;
wire [9:0] \add_10ns_10ns_10_2_1_U4.din1 ;
wire [9:0] \add_10ns_10ns_10_2_1_U4.dout ;
wire \add_10ns_10ns_10_2_1_U4.reset ;
wire [9:0] \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.a ;
wire [9:0] \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.ain_s0 ;
wire [9:0] \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.b ;
wire [9:0] \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.bin_s0 ;
wire \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.ce ;
wire \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.clk ;
wire \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.facout_s1 ;
wire \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.facout_s2 ;
wire [4:0] \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.fas_s1 ;
wire [4:0] \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.fas_s2 ;
wire \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.reset ;
wire [9:0] \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.s ;
wire [4:0] \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.u1.a ;
wire [4:0] \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.u1.b ;
wire \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.u1.cin ;
wire \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.u1.cout ;
wire [4:0] \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.u1.s ;
wire [4:0] \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.u2.a ;
wire [4:0] \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.u2.b ;
wire \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.u2.cin ;
wire \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.u2.cout ;
wire [4:0] \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.u2.s ;
wire \add_10s_10ns_10_2_1_U3.ce ;
wire \add_10s_10ns_10_2_1_U3.clk ;
wire [9:0] \add_10s_10ns_10_2_1_U3.din0 ;
wire [9:0] \add_10s_10ns_10_2_1_U3.din1 ;
wire [9:0] \add_10s_10ns_10_2_1_U3.dout ;
wire \add_10s_10ns_10_2_1_U3.reset ;
wire [9:0] \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.a ;
wire [9:0] \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.ain_s0 ;
wire [9:0] \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.b ;
wire [9:0] \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.bin_s0 ;
wire \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.ce ;
wire \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.clk ;
wire \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.facout_s1 ;
wire \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.facout_s2 ;
wire [4:0] \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.fas_s1 ;
wire [4:0] \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.fas_s2 ;
wire \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.reset ;
wire [9:0] \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.s ;
wire [4:0] \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.u1.a ;
wire [4:0] \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.u1.b ;
wire \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.u1.cin ;
wire \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.u1.cout ;
wire [4:0] \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.u1.s ;
wire [4:0] \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.u2.a ;
wire [4:0] \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.u2.b ;
wire \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.u2.cin ;
wire \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.u2.cout ;
wire [4:0] \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.u2.s ;
wire \add_12ns_12s_12_2_1_U2.ce ;
wire \add_12ns_12s_12_2_1_U2.clk ;
wire [11:0] \add_12ns_12s_12_2_1_U2.din0 ;
wire [11:0] \add_12ns_12s_12_2_1_U2.din1 ;
wire [11:0] \add_12ns_12s_12_2_1_U2.dout ;
wire \add_12ns_12s_12_2_1_U2.reset ;
wire [11:0] \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.a ;
wire [11:0] \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.ain_s0 ;
wire [11:0] \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.b ;
wire [11:0] \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.bin_s0 ;
wire \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.ce ;
wire \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.clk ;
wire \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.facout_s1 ;
wire \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.facout_s2 ;
wire [5:0] \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.fas_s1 ;
wire [5:0] \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.fas_s2 ;
wire \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.reset ;
wire [11:0] \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.s ;
wire [5:0] \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.u1.a ;
wire [5:0] \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.u1.b ;
wire \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.u1.cin ;
wire \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.u1.cout ;
wire [5:0] \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.u1.s ;
wire [5:0] \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.u2.a ;
wire [5:0] \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.u2.b ;
wire \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.u2.cin ;
wire \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.u2.cout ;
wire [5:0] \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.u2.s ;
wire \add_17s_17s_17_2_1_U7.ce ;
wire \add_17s_17s_17_2_1_U7.clk ;
wire [16:0] \add_17s_17s_17_2_1_U7.din0 ;
wire [16:0] \add_17s_17s_17_2_1_U7.din1 ;
wire [16:0] \add_17s_17s_17_2_1_U7.dout ;
wire \add_17s_17s_17_2_1_U7.reset ;
wire [16:0] \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.a ;
wire [16:0] \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.ain_s0 ;
wire [16:0] \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.b ;
wire [16:0] \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.bin_s0 ;
wire \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.ce ;
wire \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.clk ;
wire \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.facout_s1 ;
wire \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.facout_s2 ;
wire [7:0] \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.fas_s1 ;
wire [8:0] \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.fas_s2 ;
wire \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.reset ;
wire [16:0] \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.s ;
wire [7:0] \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.u1.a ;
wire [7:0] \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.u1.b ;
wire \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.u1.cin ;
wire \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.u1.cout ;
wire [7:0] \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.u1.s ;
wire [8:0] \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.u2.a ;
wire [8:0] \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.u2.b ;
wire \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.u2.cin ;
wire \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.u2.cout ;
wire [8:0] \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.u2.s ;
wire \add_32ns_32ns_32_2_1_U12.ce ;
wire \add_32ns_32ns_32_2_1_U12.clk ;
wire [31:0] \add_32ns_32ns_32_2_1_U12.din0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U12.din1 ;
wire [31:0] \add_32ns_32ns_32_2_1_U12.dout ;
wire \add_32ns_32ns_32_2_1_U12.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.a ;
wire [31:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.ain_s0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.b ;
wire [31:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.bin_s0 ;
wire \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.ce ;
wire \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.clk ;
wire \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.facout_s1 ;
wire \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.facout_s2 ;
wire [15:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.fas_s1 ;
wire [15:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.fas_s2 ;
wire \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.b ;
wire \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.cin ;
wire \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.b ;
wire \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.cin ;
wire \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.s ;
wire \add_32ns_32ns_32_2_1_U6.ce ;
wire \add_32ns_32ns_32_2_1_U6.clk ;
wire [31:0] \add_32ns_32ns_32_2_1_U6.din0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U6.din1 ;
wire [31:0] \add_32ns_32ns_32_2_1_U6.dout ;
wire \add_32ns_32ns_32_2_1_U6.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.a ;
wire [31:0] \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.ain_s0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.b ;
wire [31:0] \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.bin_s0 ;
wire \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.ce ;
wire \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.clk ;
wire \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.facout_s1 ;
wire \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.facout_s2 ;
wire [15:0] \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.fas_s1 ;
wire [15:0] \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.fas_s2 ;
wire \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.b ;
wire \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.cin ;
wire \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.b ;
wire \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.cin ;
wire \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.s ;
wire \add_32s_32ns_32_2_1_U11.ce ;
wire \add_32s_32ns_32_2_1_U11.clk ;
wire [31:0] \add_32s_32ns_32_2_1_U11.din0 ;
wire [31:0] \add_32s_32ns_32_2_1_U11.din1 ;
wire [31:0] \add_32s_32ns_32_2_1_U11.dout ;
wire \add_32s_32ns_32_2_1_U11.reset ;
wire [31:0] \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.a ;
wire [31:0] \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.ain_s0 ;
wire [31:0] \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.b ;
wire [31:0] \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.bin_s0 ;
wire \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.ce ;
wire \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.clk ;
wire \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.facout_s1 ;
wire \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.facout_s2 ;
wire [15:0] \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.fas_s1 ;
wire [15:0] \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.fas_s2 ;
wire \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.reset ;
wire [31:0] \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.s ;
wire [15:0] \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.u1.a ;
wire [15:0] \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.u1.b ;
wire \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.u1.cin ;
wire \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.u1.cout ;
wire [15:0] \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.u1.s ;
wire [15:0] \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.u2.a ;
wire [15:0] \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.u2.b ;
wire \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.u2.cin ;
wire \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.u2.cout ;
wire [15:0] \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.u2.s ;
wire \add_32s_32ns_32_2_1_U9.ce ;
wire \add_32s_32ns_32_2_1_U9.clk ;
wire [31:0] \add_32s_32ns_32_2_1_U9.din0 ;
wire [31:0] \add_32s_32ns_32_2_1_U9.din1 ;
wire [31:0] \add_32s_32ns_32_2_1_U9.dout ;
wire \add_32s_32ns_32_2_1_U9.reset ;
wire [31:0] \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.a ;
wire [31:0] \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.ain_s0 ;
wire [31:0] \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.b ;
wire [31:0] \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.bin_s0 ;
wire \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.ce ;
wire \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.clk ;
wire \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.facout_s1 ;
wire \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.facout_s2 ;
wire [15:0] \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.fas_s1 ;
wire [15:0] \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.fas_s2 ;
wire \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.reset ;
wire [31:0] \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.s ;
wire [15:0] \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.u1.a ;
wire [15:0] \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.u1.b ;
wire \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.u1.cin ;
wire \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.u1.cout ;
wire [15:0] \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.u1.s ;
wire [15:0] \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.u2.a ;
wire [15:0] \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.u2.b ;
wire \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.u2.cin ;
wire \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.u2.cout ;
wire [15:0] \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.u2.s ;
wire \add_35s_35s_35_2_1_U5.ce ;
wire \add_35s_35s_35_2_1_U5.clk ;
wire [34:0] \add_35s_35s_35_2_1_U5.din0 ;
wire [34:0] \add_35s_35s_35_2_1_U5.din1 ;
wire [34:0] \add_35s_35s_35_2_1_U5.dout ;
wire \add_35s_35s_35_2_1_U5.reset ;
wire [34:0] \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.a ;
wire [34:0] \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.ain_s0 ;
wire [34:0] \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.b ;
wire [34:0] \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.bin_s0 ;
wire \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.ce ;
wire \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.clk ;
wire \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.facout_s1 ;
wire \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.facout_s2 ;
wire [16:0] \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.fas_s1 ;
wire [17:0] \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.fas_s2 ;
wire \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.reset ;
wire [34:0] \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.s ;
wire [16:0] \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.u1.a ;
wire [16:0] \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.u1.b ;
wire \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.u1.cin ;
wire \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.u1.cout ;
wire [16:0] \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.u1.s ;
wire [17:0] \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.u2.a ;
wire [17:0] \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.u2.b ;
wire \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.u2.cin ;
wire \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.u2.cout ;
wire [17:0] \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.u2.s ;
wire \add_5ns_5ns_5_2_1_U8.ce ;
wire \add_5ns_5ns_5_2_1_U8.clk ;
wire [4:0] \add_5ns_5ns_5_2_1_U8.din0 ;
wire [4:0] \add_5ns_5ns_5_2_1_U8.din1 ;
wire [4:0] \add_5ns_5ns_5_2_1_U8.dout ;
wire \add_5ns_5ns_5_2_1_U8.reset ;
wire [4:0] \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.a ;
wire [4:0] \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.ain_s0 ;
wire [4:0] \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.b ;
wire [4:0] \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.bin_s0 ;
wire \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.ce ;
wire \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.clk ;
wire \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.facout_s1 ;
wire \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.facout_s2 ;
wire [1:0] \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.fas_s1 ;
wire [2:0] \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.fas_s2 ;
wire \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.reset ;
wire [4:0] \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.s ;
wire [1:0] \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.u1.a ;
wire [1:0] \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.u1.b ;
wire \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.u1.cin ;
wire \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.u1.cout ;
wire [1:0] \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.u1.s ;
wire [2:0] \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.u2.a ;
wire [2:0] \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.u2.b ;
wire \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.u2.cin ;
wire \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.u2.cout ;
wire [2:0] \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.u2.s ;
wire \add_6s_6s_6_2_1_U10.ce ;
wire \add_6s_6s_6_2_1_U10.clk ;
wire [5:0] \add_6s_6s_6_2_1_U10.din0 ;
wire [5:0] \add_6s_6s_6_2_1_U10.din1 ;
wire [5:0] \add_6s_6s_6_2_1_U10.dout ;
wire \add_6s_6s_6_2_1_U10.reset ;
wire [5:0] \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.a ;
wire [5:0] \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.ain_s0 ;
wire [5:0] \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.b ;
wire [5:0] \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.bin_s0 ;
wire \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.ce ;
wire \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.clk ;
wire \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.facout_s1 ;
wire \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.facout_s2 ;
wire [2:0] \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.fas_s1 ;
wire [2:0] \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.fas_s2 ;
wire \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.reset ;
wire [5:0] \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.s ;
wire [2:0] \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.u1.a ;
wire [2:0] \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.u1.b ;
wire \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.u1.cin ;
wire \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.u1.cout ;
wire [2:0] \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.u1.s ;
wire [2:0] \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.u2.a ;
wire [2:0] \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.u2.b ;
wire \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.u2.cin ;
wire \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.u2.cout ;
wire [2:0] \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.u2.s ;
wire \add_9s_9ns_9_2_1_U1.ce ;
wire \add_9s_9ns_9_2_1_U1.clk ;
wire [8:0] \add_9s_9ns_9_2_1_U1.din0 ;
wire [8:0] \add_9s_9ns_9_2_1_U1.din1 ;
wire [8:0] \add_9s_9ns_9_2_1_U1.dout ;
wire \add_9s_9ns_9_2_1_U1.reset ;
wire [8:0] \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.a ;
wire [8:0] \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.ain_s0 ;
wire [8:0] \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.b ;
wire [8:0] \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.bin_s0 ;
wire \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.ce ;
wire \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.clk ;
wire \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.facout_s1 ;
wire \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.facout_s2 ;
wire [3:0] \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.fas_s1 ;
wire [4:0] \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.fas_s2 ;
wire \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.reset ;
wire [8:0] \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.s ;
wire [3:0] \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.u1.a ;
wire [3:0] \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.u1.b ;
wire \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.u1.cin ;
wire \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.u1.cout ;
wire [3:0] \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.u1.s ;
wire [4:0] \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.u2.a ;
wire [4:0] \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.u2.b ;
wire \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.u2.cin ;
wire \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.u2.cout ;
wire [4:0] \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.u2.s ;
wire ap_CS_fsm_state1;
wire ap_CS_fsm_state10;
wire ap_CS_fsm_state11;
wire ap_CS_fsm_state12;
wire ap_CS_fsm_state13;
wire ap_CS_fsm_state14;
wire ap_CS_fsm_state15;
wire ap_CS_fsm_state16;
wire ap_CS_fsm_state17;
wire ap_CS_fsm_state18;
wire ap_CS_fsm_state19;
wire ap_CS_fsm_state2;
wire ap_CS_fsm_state20;
wire ap_CS_fsm_state21;
wire ap_CS_fsm_state3;
wire ap_CS_fsm_state4;
wire ap_CS_fsm_state5;
wire ap_CS_fsm_state6;
wire ap_CS_fsm_state7;
wire ap_CS_fsm_state8;
wire ap_CS_fsm_state9;
wire [20:0] ap_NS_fsm;
wire ap_clk;
wire ap_done;
wire ap_idle;
wire ap_ready;
wire ap_rst;
wire ap_start;
wire [8:0] grp_fu_185_p0;
wire [8:0] grp_fu_185_p2;
wire [11:0] grp_fu_201_p0;
wire [11:0] grp_fu_201_p1;
wire [11:0] grp_fu_201_p2;
wire [9:0] grp_fu_230_p0;
wire [9:0] grp_fu_230_p2;
wire [9:0] grp_fu_263_p2;
wire [34:0] grp_fu_282_p0;
wire [34:0] grp_fu_282_p1;
wire [34:0] grp_fu_282_p2;
wire [31:0] grp_fu_308_p2;
wire [16:0] grp_fu_333_p0;
wire [16:0] grp_fu_333_p1;
wire [16:0] grp_fu_333_p2;
wire [4:0] grp_fu_339_p0;
wire [4:0] grp_fu_339_p2;
wire [31:0] grp_fu_370_p0;
wire [31:0] grp_fu_370_p2;
wire [5:0] grp_fu_378_p0;
wire [5:0] grp_fu_378_p1;
wire [5:0] grp_fu_378_p2;
wire [31:0] grp_fu_387_p0;
wire [31:0] grp_fu_387_p2;
wire [31:0] grp_fu_400_p2;
wire icmp_ln851_1_fu_292_p2;
wire icmp_ln851_fu_211_p2;
wire [1:0] op_0;
wire [3:0] op_1;
wire [3:0] op_10;
wire op_11;
wire [3:0] op_12;
wire [7:0] op_13;
wire [3:0] op_14;
wire op_15;
wire [15:0] op_16;
wire [3:0] op_17;
wire op_18;
wire [31:0] op_30;
wire op_30_ap_vld;
wire [3:0] op_5;
wire [7:0] op_6;
wire op_8_V_fu_169_p1;
wire p_Result_1_fu_344_p3;
wire p_Result_s_fu_236_p3;
wire [9:0] ret_V_1_fu_248_p3;
wire [31:0] ret_V_3_fu_356_p3;
wire [31:0] select_ln1192_fu_392_p3;
wire [8:0] select_ln215_fu_173_p3;
wire [4:0] select_ln69_1_fu_313_p3;
wire [9:0] select_ln69_fu_255_p3;
wire [31:0] select_ln850_1_fu_351_p3;
wire [9:0] select_ln850_fu_243_p3;
wire [3:0] sext_ln1192_fu_190_p0;
wire [3:0] sext_ln703_fu_267_p0;
wire [9:0] sext_ln850_fu_227_p1;
wire [11:0] tmp_fu_271_p3;
wire [3:0] trunc_ln851_1_fu_288_p0;
wire [1:0] trunc_ln851_1_fu_288_p1;
wire [3:0] trunc_ln851_fu_207_p0;
wire [2:0] trunc_ln851_fu_207_p1;


assign _024_ = ap_CS_fsm[13] & icmp_ln851_1_reg_482;
assign _025_ = icmp_ln851_reg_430 & ap_CS_fsm[6];
assign _026_ = _028_ & ap_CS_fsm[0];
assign _027_ = ap_start & ap_CS_fsm[0];
assign _028_ = ~ ap_start;
always @(posedge \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.clk )
\add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.bin_s1  <= _030_;
always @(posedge \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.clk )
\add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.ain_s1  <= _029_;
always @(posedge \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.clk )
\add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.sum_s1  <= _032_;
always @(posedge \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.clk )
\add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.carry_s1  <= _031_;
assign _030_ = \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.ce  ? \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.b [9:5] : \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.bin_s1 ;
assign _029_ = \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.ce  ? \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.a [9:5] : \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.ain_s1 ;
assign _031_ = \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.ce  ? \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.facout_s1  : \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.carry_s1 ;
assign _032_ = \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.ce  ? \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.fas_s1  : \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.sum_s1 ;
assign _033_ = \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.u1.a  + \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.u1.b ;
assign { \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.u1.cout , \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.u1.s  } = _033_ + \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.u1.cin ;
assign _034_ = \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.u2.a  + \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.u2.b ;
assign { \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.u2.cout , \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.u2.s  } = _034_ + \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.u2.cin ;
always @(posedge \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.clk )
\add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.bin_s1  <= _036_;
always @(posedge \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.clk )
\add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.ain_s1  <= _035_;
always @(posedge \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.clk )
\add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.sum_s1  <= _038_;
always @(posedge \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.clk )
\add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.carry_s1  <= _037_;
assign _036_ = \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.ce  ? \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.b [9:5] : \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.bin_s1 ;
assign _035_ = \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.ce  ? \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.a [9:5] : \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.ain_s1 ;
assign _037_ = \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.ce  ? \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.facout_s1  : \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.carry_s1 ;
assign _038_ = \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.ce  ? \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.fas_s1  : \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.sum_s1 ;
assign _039_ = \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.u1.a  + \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.u1.b ;
assign { \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.u1.cout , \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.u1.s  } = _039_ + \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.u1.cin ;
assign _040_ = \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.u2.a  + \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.u2.b ;
assign { \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.u2.cout , \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.u2.s  } = _040_ + \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.u2.cin ;
always @(posedge \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.clk )
\add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.bin_s1  <= _042_;
always @(posedge \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.clk )
\add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.ain_s1  <= _041_;
always @(posedge \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.clk )
\add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.sum_s1  <= _044_;
always @(posedge \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.clk )
\add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.carry_s1  <= _043_;
assign _042_ = \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.ce  ? \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.b [11:6] : \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.bin_s1 ;
assign _041_ = \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.ce  ? \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.a [11:6] : \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.ain_s1 ;
assign _043_ = \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.ce  ? \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.facout_s1  : \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.carry_s1 ;
assign _044_ = \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.ce  ? \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.fas_s1  : \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.sum_s1 ;
assign _045_ = \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.u1.a  + \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.u1.b ;
assign { \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.u1.cout , \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.u1.s  } = _045_ + \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.u1.cin ;
assign _046_ = \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.u2.a  + \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.u2.b ;
assign { \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.u2.cout , \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.u2.s  } = _046_ + \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.u2.cin ;
always @(posedge \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.clk )
\add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.bin_s1  <= _048_;
always @(posedge \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.clk )
\add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.ain_s1  <= _047_;
always @(posedge \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.clk )
\add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.sum_s1  <= _050_;
always @(posedge \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.clk )
\add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.carry_s1  <= _049_;
assign _048_ = \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.ce  ? \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.b [16:8] : \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.bin_s1 ;
assign _047_ = \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.ce  ? \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.a [16:8] : \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.ain_s1 ;
assign _049_ = \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.ce  ? \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.facout_s1  : \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.carry_s1 ;
assign _050_ = \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.ce  ? \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.fas_s1  : \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.sum_s1 ;
assign _051_ = \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.u1.a  + \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.u1.b ;
assign { \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.u1.cout , \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.u1.s  } = _051_ + \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.u1.cin ;
assign _052_ = \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.u2.a  + \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.u2.b ;
assign { \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.u2.cout , \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.u2.s  } = _052_ + \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.u2.cin ;
always @(posedge \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.clk )
\add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.bin_s1  <= _054_;
always @(posedge \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.clk )
\add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.ain_s1  <= _053_;
always @(posedge \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.clk )
\add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.sum_s1  <= _056_;
always @(posedge \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.clk )
\add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.carry_s1  <= _055_;
assign _054_ = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.ce  ? \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.b [31:16] : \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.bin_s1 ;
assign _053_ = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.ce  ? \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.a [31:16] : \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.ain_s1 ;
assign _055_ = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.ce  ? \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.facout_s1  : \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.carry_s1 ;
assign _056_ = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.ce  ? \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.fas_s1  : \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.sum_s1 ;
assign _057_ = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.a  + \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.b ;
assign { \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.cout , \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.s  } = _057_ + \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.cin ;
assign _058_ = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.a  + \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.b ;
assign { \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.cout , \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.s  } = _058_ + \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.cin ;
always @(posedge \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.clk )
\add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.bin_s1  <= _060_;
always @(posedge \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.clk )
\add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.ain_s1  <= _059_;
always @(posedge \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.clk )
\add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.sum_s1  <= _062_;
always @(posedge \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.clk )
\add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.carry_s1  <= _061_;
assign _060_ = \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.ce  ? \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.b [31:16] : \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.bin_s1 ;
assign _059_ = \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.ce  ? \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.a [31:16] : \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.ain_s1 ;
assign _061_ = \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.ce  ? \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.facout_s1  : \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.carry_s1 ;
assign _062_ = \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.ce  ? \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.fas_s1  : \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.sum_s1 ;
assign _063_ = \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.a  + \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.b ;
assign { \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.cout , \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.s  } = _063_ + \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.cin ;
assign _064_ = \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.a  + \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.b ;
assign { \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.cout , \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.s  } = _064_ + \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.cin ;
always @(posedge \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.clk )
\add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.bin_s1  <= _066_;
always @(posedge \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.clk )
\add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.ain_s1  <= _065_;
always @(posedge \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.clk )
\add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.sum_s1  <= _068_;
always @(posedge \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.clk )
\add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.carry_s1  <= _067_;
assign _066_ = \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.ce  ? \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.b [31:16] : \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.bin_s1 ;
assign _065_ = \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.ce  ? \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.a [31:16] : \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.ain_s1 ;
assign _067_ = \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.ce  ? \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.facout_s1  : \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.carry_s1 ;
assign _068_ = \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.ce  ? \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.fas_s1  : \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.sum_s1 ;
assign _069_ = \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.u1.a  + \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.u1.b ;
assign { \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.u1.cout , \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.u1.s  } = _069_ + \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.u1.cin ;
assign _070_ = \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.u2.a  + \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.u2.b ;
assign { \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.u2.cout , \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.u2.s  } = _070_ + \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.u2.cin ;
always @(posedge \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.clk )
\add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.bin_s1  <= _072_;
always @(posedge \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.clk )
\add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.ain_s1  <= _071_;
always @(posedge \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.clk )
\add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.sum_s1  <= _074_;
always @(posedge \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.clk )
\add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.carry_s1  <= _073_;
assign _072_ = \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.ce  ? \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.b [31:16] : \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.bin_s1 ;
assign _071_ = \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.ce  ? \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.a [31:16] : \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.ain_s1 ;
assign _073_ = \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.ce  ? \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.facout_s1  : \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.carry_s1 ;
assign _074_ = \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.ce  ? \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.fas_s1  : \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.sum_s1 ;
assign _075_ = \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.u1.a  + \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.u1.b ;
assign { \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.u1.cout , \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.u1.s  } = _075_ + \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.u1.cin ;
assign _076_ = \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.u2.a  + \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.u2.b ;
assign { \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.u2.cout , \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.u2.s  } = _076_ + \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.u2.cin ;
always @(posedge \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.clk )
\add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.bin_s1  <= _078_;
always @(posedge \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.clk )
\add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.ain_s1  <= _077_;
always @(posedge \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.clk )
\add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.sum_s1  <= _080_;
always @(posedge \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.clk )
\add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.carry_s1  <= _079_;
assign _078_ = \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.ce  ? \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.b [34:17] : \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.bin_s1 ;
assign _077_ = \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.ce  ? \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.a [34:17] : \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.ain_s1 ;
assign _079_ = \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.ce  ? \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.facout_s1  : \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.carry_s1 ;
assign _080_ = \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.ce  ? \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.fas_s1  : \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.sum_s1 ;
assign _081_ = \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.u1.a  + \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.u1.b ;
assign { \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.u1.cout , \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.u1.s  } = _081_ + \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.u1.cin ;
assign _082_ = \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.u2.a  + \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.u2.b ;
assign { \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.u2.cout , \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.u2.s  } = _082_ + \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.u2.cin ;
always @(posedge \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.clk )
\add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.bin_s1  <= _084_;
always @(posedge \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.clk )
\add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.ain_s1  <= _083_;
always @(posedge \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.clk )
\add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.sum_s1  <= _086_;
always @(posedge \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.clk )
\add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.carry_s1  <= _085_;
assign _084_ = \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.ce  ? \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.b [4:2] : \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.bin_s1 ;
assign _083_ = \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.ce  ? \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.a [4:2] : \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.ain_s1 ;
assign _085_ = \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.ce  ? \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.facout_s1  : \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.carry_s1 ;
assign _086_ = \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.ce  ? \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.fas_s1  : \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.sum_s1 ;
assign _087_ = \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.u1.a  + \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.u1.b ;
assign { \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.u1.cout , \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.u1.s  } = _087_ + \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.u1.cin ;
assign _088_ = \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.u2.a  + \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.u2.b ;
assign { \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.u2.cout , \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.u2.s  } = _088_ + \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.u2.cin ;
always @(posedge \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.clk )
\add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.bin_s1  <= _090_;
always @(posedge \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.clk )
\add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.ain_s1  <= _089_;
always @(posedge \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.clk )
\add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.sum_s1  <= _092_;
always @(posedge \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.clk )
\add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.carry_s1  <= _091_;
assign _090_ = \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.ce  ? \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.b [5:3] : \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.bin_s1 ;
assign _089_ = \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.ce  ? \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.a [5:3] : \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.ain_s1 ;
assign _091_ = \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.ce  ? \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.facout_s1  : \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.carry_s1 ;
assign _092_ = \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.ce  ? \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.fas_s1  : \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.sum_s1 ;
assign _093_ = \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.u1.a  + \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.u1.b ;
assign { \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.u1.cout , \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.u1.s  } = _093_ + \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.u1.cin ;
assign _094_ = \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.u2.a  + \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.u2.b ;
assign { \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.u2.cout , \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.u2.s  } = _094_ + \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.u2.cin ;
always @(posedge \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.clk )
\add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.bin_s1  <= _096_;
always @(posedge \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.clk )
\add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.ain_s1  <= _095_;
always @(posedge \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.clk )
\add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.sum_s1  <= _098_;
always @(posedge \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.clk )
\add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.carry_s1  <= _097_;
assign _096_ = \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.ce  ? \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.b [8:4] : \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.bin_s1 ;
assign _095_ = \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.ce  ? \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.a [8:4] : \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.ain_s1 ;
assign _097_ = \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.ce  ? \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.facout_s1  : \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.carry_s1 ;
assign _098_ = \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.ce  ? \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.fas_s1  : \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.sum_s1 ;
assign _099_ = \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.u1.a  + \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.u1.b ;
assign { \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.u1.cout , \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.u1.s  } = _099_ + \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.u1.cin ;
assign _100_ = \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.u2.a  + \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.u2.b ;
assign { \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.u2.cout , \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.u2.s  } = _100_ + \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.u2.cin ;
assign _101_ = | op_12[1:0];
assign _102_ = | op_10[2:0];
always @(posedge ap_clk)
sext_ln850_reg_445 <= _021_;
always @(posedge ap_clk)
select_ln69_1_reg_499 <= _019_;
always @(posedge ap_clk)
select_ln215_reg_405 <= _018_;
always @(posedge ap_clk)
ret_reg_415 <= _016_;
always @(posedge ap_clk)
ret_V_reg_435 <= _015_;
always @(posedge ap_clk)
tmp_1_reg_440 <= _022_;
always @(posedge ap_clk)
ret_V_2_reg_487 <= _012_;
always @(posedge ap_clk)
ret_V_3_cast_reg_492 <= _013_;
always @(posedge ap_clk)
ret_V_1_reg_457 <= _011_;
always @(posedge ap_clk)
select_ln69_reg_462 <= _020_;
always @(posedge ap_clk)
op_28_V_reg_569 <= _010_;
always @(posedge ap_clk)
select_ln1192_reg_574 <= _017_;
always @(posedge ap_clk)
op_22_V_reg_467 <= _009_;
always @(posedge ap_clk)
icmp_ln851_reg_430 <= _008_;
always @(posedge ap_clk)
icmp_ln851_1_reg_482 <= _007_;
always @(posedge ap_clk)
ret_V_3_reg_524 <= _014_;
always @(posedge ap_clk)
add_ln69_reg_529 <= _005_;
always @(posedge ap_clk)
add_ln69_2_reg_534 <= _003_;
always @(posedge ap_clk)
add_ln69_1_reg_554 <= _002_;
always @(posedge ap_clk)
add_ln69_3_reg_559 <= _004_;
always @(posedge ap_clk)
add_ln691_reg_452 <= _001_;
always @(posedge ap_clk)
add_ln691_1_reg_504 <= _000_;
always @(posedge ap_clk)
ap_CS_fsm <= _006_;
assign _023_ = _027_ ? 2'h2 : 2'h1;
assign _103_ = ap_CS_fsm == 1'h1;
function [20:0] _300_;
input [20:0] a;
input [440:0] b;
input [20:0] s;
case (s)
21'b000000000000000000001:
_300_ = b[20:0];
21'b000000000000000000010:
_300_ = b[41:21];
21'b000000000000000000100:
_300_ = b[62:42];
21'b000000000000000001000:
_300_ = b[83:63];
21'b000000000000000010000:
_300_ = b[104:84];
21'b000000000000000100000:
_300_ = b[125:105];
21'b000000000000001000000:
_300_ = b[146:126];
21'b000000000000010000000:
_300_ = b[167:147];
21'b000000000000100000000:
_300_ = b[188:168];
21'b000000000001000000000:
_300_ = b[209:189];
21'b000000000010000000000:
_300_ = b[230:210];
21'b000000000100000000000:
_300_ = b[251:231];
21'b000000001000000000000:
_300_ = b[272:252];
21'b000000010000000000000:
_300_ = b[293:273];
21'b000000100000000000000:
_300_ = b[314:294];
21'b000001000000000000000:
_300_ = b[335:315];
21'b000010000000000000000:
_300_ = b[356:336];
21'b000100000000000000000:
_300_ = b[377:357];
21'b001000000000000000000:
_300_ = b[398:378];
21'b010000000000000000000:
_300_ = b[419:399];
21'b100000000000000000000:
_300_ = b[440:420];
21'b000000000000000000000:
_300_ = a;
default:
_300_ = 21'bx;
endcase
endfunction
assign ap_NS_fsm = _300_(21'hxxxxxx, { 19'h00000, _023_, 420'h000020000200002000020000200002000020000200002000020000200002000020000200002000020000200002000020000000001 }, { _103_, _123_, _122_, _121_, _120_, _119_, _118_, _117_, _116_, _115_, _114_, _113_, _112_, _111_, _110_, _109_, _108_, _107_, _106_, _105_, _104_ });
assign _104_ = ap_CS_fsm == 21'h100000;
assign _105_ = ap_CS_fsm == 20'h80000;
assign _106_ = ap_CS_fsm == 19'h40000;
assign _107_ = ap_CS_fsm == 18'h20000;
assign _108_ = ap_CS_fsm == 17'h10000;
assign _109_ = ap_CS_fsm == 16'h8000;
assign _110_ = ap_CS_fsm == 15'h4000;
assign _111_ = ap_CS_fsm == 14'h2000;
assign _112_ = ap_CS_fsm == 13'h1000;
assign _113_ = ap_CS_fsm == 12'h800;
assign _114_ = ap_CS_fsm == 11'h400;
assign _115_ = ap_CS_fsm == 10'h200;
assign _116_ = ap_CS_fsm == 9'h100;
assign _117_ = ap_CS_fsm == 8'h80;
assign _118_ = ap_CS_fsm == 7'h40;
assign _119_ = ap_CS_fsm == 6'h20;
assign _120_ = ap_CS_fsm == 5'h10;
assign _121_ = ap_CS_fsm == 4'h8;
assign _122_ = ap_CS_fsm == 3'h4;
assign _123_ = ap_CS_fsm == 2'h2;
assign op_30_ap_vld = ap_CS_fsm[20] ? 1'h1 : 1'h0;
assign ap_idle = _026_ ? 1'h1 : 1'h0;
assign _021_ = ap_CS_fsm[5] ? { tmp_1_reg_440[8], tmp_1_reg_440 } : sext_ln850_reg_445;
assign _019_ = ap_CS_fsm[12] ? select_ln69_1_fu_313_p3 : select_ln69_1_reg_499;
assign _018_ = ap_CS_fsm[0] ? select_ln215_fu_173_p3 : select_ln215_reg_405;
assign _016_ = ap_CS_fsm[2] ? grp_fu_185_p2 : ret_reg_415;
assign _022_ = ap_CS_fsm[4] ? grp_fu_201_p2[11:3] : tmp_1_reg_440;
assign _015_ = ap_CS_fsm[4] ? grp_fu_201_p2 : ret_V_reg_435;
assign _013_ = ap_CS_fsm[11] ? grp_fu_282_p2[33:2] : ret_V_3_cast_reg_492;
assign _012_ = ap_CS_fsm[11] ? grp_fu_282_p2 : ret_V_2_reg_487;
assign _020_ = ap_CS_fsm[7] ? select_ln69_fu_255_p3 : select_ln69_reg_462;
assign _011_ = ap_CS_fsm[7] ? ret_V_1_fu_248_p3 : ret_V_1_reg_457;
assign _017_ = ap_CS_fsm[18] ? select_ln1192_fu_392_p3 : select_ln1192_reg_574;
assign _010_ = ap_CS_fsm[18] ? grp_fu_387_p2 : op_28_V_reg_569;
assign _009_ = ap_CS_fsm[9] ? grp_fu_263_p2 : op_22_V_reg_467;
assign _008_ = ap_CS_fsm[3] ? icmp_ln851_fu_211_p2 : icmp_ln851_reg_430;
assign _007_ = ap_CS_fsm[10] ? icmp_ln851_1_fu_292_p2 : icmp_ln851_1_reg_482;
assign _003_ = ap_CS_fsm[14] ? grp_fu_339_p2 : add_ln69_2_reg_534;
assign _005_ = ap_CS_fsm[14] ? grp_fu_333_p2 : add_ln69_reg_529;
assign _014_ = ap_CS_fsm[14] ? ret_V_3_fu_356_p3 : ret_V_3_reg_524;
assign _004_ = ap_CS_fsm[16] ? grp_fu_378_p2 : add_ln69_3_reg_559;
assign _002_ = ap_CS_fsm[16] ? grp_fu_370_p2 : add_ln69_1_reg_554;
assign _001_ = _025_ ? grp_fu_230_p2 : add_ln691_reg_452;
assign _000_ = _024_ ? grp_fu_308_p2 : add_ln691_1_reg_504;
assign _006_ = ap_rst ? 21'h000001 : ap_NS_fsm;
assign icmp_ln851_1_fu_292_p2 = _101_ ? 1'h1 : 1'h0;
assign icmp_ln851_fu_211_p2 = _102_ ? 1'h1 : 1'h0;
assign ret_V_1_fu_248_p3 = ret_V_reg_435[11] ? select_ln850_fu_243_p3 : sext_ln850_reg_445;
assign ret_V_3_fu_356_p3 = ret_V_2_reg_487[34] ? select_ln850_1_fu_351_p3 : ret_V_3_cast_reg_492;
assign select_ln1192_fu_392_p3 = op_18 ? 32'd4294967295 : 32'd0;
assign select_ln215_fu_173_p3 = op_5[0] ? 9'h1ff : 9'h000;
assign select_ln69_1_fu_313_p3 = op_15 ? 5'h1f : 5'h00;
assign select_ln69_fu_255_p3 = op_11 ? 10'h3ff : 10'h000;
assign select_ln850_1_fu_351_p3 = icmp_ln851_1_reg_482 ? add_ln691_1_reg_504 : ret_V_3_cast_reg_492;
assign select_ln850_fu_243_p3 = icmp_ln851_reg_430 ? add_ln691_reg_452 : sext_ln850_reg_445;
assign ap_CS_fsm_state1 = ap_CS_fsm[0];
assign ap_CS_fsm_state10 = ap_CS_fsm[9];
assign ap_CS_fsm_state11 = ap_CS_fsm[10];
assign ap_CS_fsm_state12 = ap_CS_fsm[11];
assign ap_CS_fsm_state13 = ap_CS_fsm[12];
assign ap_CS_fsm_state14 = ap_CS_fsm[13];
assign ap_CS_fsm_state15 = ap_CS_fsm[14];
assign ap_CS_fsm_state16 = ap_CS_fsm[15];
assign ap_CS_fsm_state17 = ap_CS_fsm[16];
assign ap_CS_fsm_state18 = ap_CS_fsm[17];
assign ap_CS_fsm_state19 = ap_CS_fsm[18];
assign ap_CS_fsm_state2 = ap_CS_fsm[1];
assign ap_CS_fsm_state20 = ap_CS_fsm[19];
assign ap_CS_fsm_state21 = ap_CS_fsm[20];
assign ap_CS_fsm_state3 = ap_CS_fsm[2];
assign ap_CS_fsm_state4 = ap_CS_fsm[3];
assign ap_CS_fsm_state5 = ap_CS_fsm[4];
assign ap_CS_fsm_state6 = ap_CS_fsm[5];
assign ap_CS_fsm_state7 = ap_CS_fsm[6];
assign ap_CS_fsm_state8 = ap_CS_fsm[7];
assign ap_CS_fsm_state9 = ap_CS_fsm[8];
assign ap_done = op_30_ap_vld;
assign ap_ready = op_30_ap_vld;
assign grp_fu_185_p0 = { op_6[7], op_6 };
assign grp_fu_201_p0 = { ret_reg_415, 3'h0 };
assign grp_fu_201_p1 = { op_10[3], op_10[3], op_10[3], op_10[3], op_10[3], op_10[3], op_10[3], op_10[3], op_10 };
assign grp_fu_230_p0 = { tmp_1_reg_440[8], tmp_1_reg_440 };
assign grp_fu_282_p0 = { op_22_V_reg_467[9], op_22_V_reg_467[9], op_22_V_reg_467[9], op_22_V_reg_467[9], op_22_V_reg_467[9], op_22_V_reg_467[9], op_22_V_reg_467[9], op_22_V_reg_467[9], op_22_V_reg_467[9], op_22_V_reg_467[9], op_22_V_reg_467[9], op_22_V_reg_467[9], op_22_V_reg_467[9], op_22_V_reg_467[9], op_22_V_reg_467[9], op_22_V_reg_467[9], op_22_V_reg_467[9], op_22_V_reg_467[9], op_22_V_reg_467[9], op_22_V_reg_467[9], op_22_V_reg_467[9], op_22_V_reg_467[9], op_22_V_reg_467[9], op_22_V_reg_467, 2'h0 };
assign grp_fu_282_p1 = { op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12 };
assign grp_fu_333_p0 = { op_16[15], op_16 };
assign grp_fu_333_p1 = { op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13 };
assign grp_fu_339_p0 = { 1'h0, op_14 };
assign grp_fu_370_p0 = { add_ln69_reg_529[16], add_ln69_reg_529[16], add_ln69_reg_529[16], add_ln69_reg_529[16], add_ln69_reg_529[16], add_ln69_reg_529[16], add_ln69_reg_529[16], add_ln69_reg_529[16], add_ln69_reg_529[16], add_ln69_reg_529[16], add_ln69_reg_529[16], add_ln69_reg_529[16], add_ln69_reg_529[16], add_ln69_reg_529[16], add_ln69_reg_529[16], add_ln69_reg_529 };
assign grp_fu_378_p0 = { add_ln69_2_reg_534[4], add_ln69_2_reg_534 };
assign grp_fu_378_p1 = { op_17[3], op_17[3], op_17 };
assign grp_fu_387_p0 = { add_ln69_3_reg_559[5], add_ln69_3_reg_559[5], add_ln69_3_reg_559[5], add_ln69_3_reg_559[5], add_ln69_3_reg_559[5], add_ln69_3_reg_559[5], add_ln69_3_reg_559[5], add_ln69_3_reg_559[5], add_ln69_3_reg_559[5], add_ln69_3_reg_559[5], add_ln69_3_reg_559[5], add_ln69_3_reg_559[5], add_ln69_3_reg_559[5], add_ln69_3_reg_559[5], add_ln69_3_reg_559[5], add_ln69_3_reg_559[5], add_ln69_3_reg_559[5], add_ln69_3_reg_559[5], add_ln69_3_reg_559[5], add_ln69_3_reg_559[5], add_ln69_3_reg_559[5], add_ln69_3_reg_559[5], add_ln69_3_reg_559[5], add_ln69_3_reg_559[5], add_ln69_3_reg_559[5], add_ln69_3_reg_559[5], add_ln69_3_reg_559 };
assign op_30 = grp_fu_400_p2;
assign op_8_V_fu_169_p1 = op_5[0];
assign p_Result_1_fu_344_p3 = ret_V_2_reg_487[34];
assign p_Result_s_fu_236_p3 = ret_V_reg_435[11];
assign sext_ln1192_fu_190_p0 = op_10;
assign sext_ln703_fu_267_p0 = op_12;
assign sext_ln850_fu_227_p1 = { tmp_1_reg_440[8], tmp_1_reg_440 };
assign tmp_fu_271_p3 = { op_22_V_reg_467, 2'h0 };
assign trunc_ln851_1_fu_288_p0 = op_12;
assign trunc_ln851_1_fu_288_p1 = op_12[1:0];
assign trunc_ln851_fu_207_p0 = op_10;
assign trunc_ln851_fu_207_p1 = op_10[2:0];
assign \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.ain_s0  = \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.a ;
assign \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.bin_s0  = \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.b ;
assign \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.s  = { \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.fas_s2 , \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.sum_s1  };
assign \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.u2.a  = \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.ain_s1 ;
assign \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.u2.b  = \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.bin_s1 ;
assign \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.u2.cin  = \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.carry_s1 ;
assign \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.facout_s2  = \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.u2.cout ;
assign \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.fas_s2  = \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.u2.s ;
assign \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.u1.a  = \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.a [3:0];
assign \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.u1.b  = \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.b [3:0];
assign \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.u1.cin  = 1'h0;
assign \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.facout_s1  = \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.u1.cout ;
assign \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.fas_s1  = \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.u1.s ;
assign \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.a  = \add_9s_9ns_9_2_1_U1.din0 ;
assign \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.b  = \add_9s_9ns_9_2_1_U1.din1 ;
assign \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.ce  = \add_9s_9ns_9_2_1_U1.ce ;
assign \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.clk  = \add_9s_9ns_9_2_1_U1.clk ;
assign \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.reset  = \add_9s_9ns_9_2_1_U1.reset ;
assign \add_9s_9ns_9_2_1_U1.dout  = \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.s ;
assign \add_9s_9ns_9_2_1_U1.ce  = 1'h1;
assign \add_9s_9ns_9_2_1_U1.clk  = ap_clk;
assign \add_9s_9ns_9_2_1_U1.din0  = { op_6[7], op_6 };
assign \add_9s_9ns_9_2_1_U1.din1  = select_ln215_reg_405;
assign grp_fu_185_p2 = \add_9s_9ns_9_2_1_U1.dout ;
assign \add_9s_9ns_9_2_1_U1.reset  = ap_rst;
assign \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.ain_s0  = \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.a ;
assign \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.bin_s0  = \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.b ;
assign \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.s  = { \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.fas_s2 , \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.sum_s1  };
assign \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.u2.a  = \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.ain_s1 ;
assign \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.u2.b  = \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.bin_s1 ;
assign \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.u2.cin  = \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.carry_s1 ;
assign \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.facout_s2  = \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.u2.cout ;
assign \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.fas_s2  = \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.u2.s ;
assign \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.u1.a  = \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.a [2:0];
assign \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.u1.b  = \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.b [2:0];
assign \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.u1.cin  = 1'h0;
assign \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.facout_s1  = \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.u1.cout ;
assign \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.fas_s1  = \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.u1.s ;
assign \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.a  = \add_6s_6s_6_2_1_U10.din0 ;
assign \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.b  = \add_6s_6s_6_2_1_U10.din1 ;
assign \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.ce  = \add_6s_6s_6_2_1_U10.ce ;
assign \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.clk  = \add_6s_6s_6_2_1_U10.clk ;
assign \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.reset  = \add_6s_6s_6_2_1_U10.reset ;
assign \add_6s_6s_6_2_1_U10.dout  = \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.s ;
assign \add_6s_6s_6_2_1_U10.ce  = 1'h1;
assign \add_6s_6s_6_2_1_U10.clk  = ap_clk;
assign \add_6s_6s_6_2_1_U10.din0  = { add_ln69_2_reg_534[4], add_ln69_2_reg_534 };
assign \add_6s_6s_6_2_1_U10.din1  = { op_17[3], op_17[3], op_17 };
assign grp_fu_378_p2 = \add_6s_6s_6_2_1_U10.dout ;
assign \add_6s_6s_6_2_1_U10.reset  = ap_rst;
assign \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.ain_s0  = \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.a ;
assign \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.bin_s0  = \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.b ;
assign \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.s  = { \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.fas_s2 , \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.sum_s1  };
assign \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.u2.a  = \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.ain_s1 ;
assign \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.u2.b  = \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.bin_s1 ;
assign \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.u2.cin  = \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.carry_s1 ;
assign \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.facout_s2  = \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.u2.cout ;
assign \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.fas_s2  = \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.u2.s ;
assign \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.u1.a  = \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.a [1:0];
assign \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.u1.b  = \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.b [1:0];
assign \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.u1.cin  = 1'h0;
assign \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.facout_s1  = \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.u1.cout ;
assign \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.fas_s1  = \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.u1.s ;
assign \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.a  = \add_5ns_5ns_5_2_1_U8.din0 ;
assign \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.b  = \add_5ns_5ns_5_2_1_U8.din1 ;
assign \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.ce  = \add_5ns_5ns_5_2_1_U8.ce ;
assign \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.clk  = \add_5ns_5ns_5_2_1_U8.clk ;
assign \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.reset  = \add_5ns_5ns_5_2_1_U8.reset ;
assign \add_5ns_5ns_5_2_1_U8.dout  = \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.s ;
assign \add_5ns_5ns_5_2_1_U8.ce  = 1'h1;
assign \add_5ns_5ns_5_2_1_U8.clk  = ap_clk;
assign \add_5ns_5ns_5_2_1_U8.din0  = { 1'h0, op_14 };
assign \add_5ns_5ns_5_2_1_U8.din1  = select_ln69_1_reg_499;
assign grp_fu_339_p2 = \add_5ns_5ns_5_2_1_U8.dout ;
assign \add_5ns_5ns_5_2_1_U8.reset  = ap_rst;
assign \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.ain_s0  = \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.a ;
assign \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.bin_s0  = \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.b ;
assign \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.s  = { \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.fas_s2 , \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.sum_s1  };
assign \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.u2.a  = \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.ain_s1 ;
assign \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.u2.b  = \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.bin_s1 ;
assign \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.u2.cin  = \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.carry_s1 ;
assign \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.facout_s2  = \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.u2.cout ;
assign \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.fas_s2  = \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.u2.s ;
assign \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.u1.a  = \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.a [16:0];
assign \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.u1.b  = \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.b [16:0];
assign \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.u1.cin  = 1'h0;
assign \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.facout_s1  = \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.u1.cout ;
assign \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.fas_s1  = \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.u1.s ;
assign \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.a  = \add_35s_35s_35_2_1_U5.din0 ;
assign \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.b  = \add_35s_35s_35_2_1_U5.din1 ;
assign \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.ce  = \add_35s_35s_35_2_1_U5.ce ;
assign \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.clk  = \add_35s_35s_35_2_1_U5.clk ;
assign \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.reset  = \add_35s_35s_35_2_1_U5.reset ;
assign \add_35s_35s_35_2_1_U5.dout  = \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.s ;
assign \add_35s_35s_35_2_1_U5.ce  = 1'h1;
assign \add_35s_35s_35_2_1_U5.clk  = ap_clk;
assign \add_35s_35s_35_2_1_U5.din0  = { op_22_V_reg_467[9], op_22_V_reg_467[9], op_22_V_reg_467[9], op_22_V_reg_467[9], op_22_V_reg_467[9], op_22_V_reg_467[9], op_22_V_reg_467[9], op_22_V_reg_467[9], op_22_V_reg_467[9], op_22_V_reg_467[9], op_22_V_reg_467[9], op_22_V_reg_467[9], op_22_V_reg_467[9], op_22_V_reg_467[9], op_22_V_reg_467[9], op_22_V_reg_467[9], op_22_V_reg_467[9], op_22_V_reg_467[9], op_22_V_reg_467[9], op_22_V_reg_467[9], op_22_V_reg_467[9], op_22_V_reg_467[9], op_22_V_reg_467[9], op_22_V_reg_467, 2'h0 };
assign \add_35s_35s_35_2_1_U5.din1  = { op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12 };
assign grp_fu_282_p2 = \add_35s_35s_35_2_1_U5.dout ;
assign \add_35s_35s_35_2_1_U5.reset  = ap_rst;
assign \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.ain_s0  = \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.a ;
assign \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.bin_s0  = \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.b ;
assign \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.s  = { \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.fas_s2 , \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.sum_s1  };
assign \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.u2.a  = \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.ain_s1 ;
assign \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.u2.b  = \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.bin_s1 ;
assign \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.u2.cin  = \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.carry_s1 ;
assign \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.facout_s2  = \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.u2.cout ;
assign \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.fas_s2  = \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.u2.s ;
assign \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.u1.a  = \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.a [15:0];
assign \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.u1.b  = \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.b [15:0];
assign \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.u1.cin  = 1'h0;
assign \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.facout_s1  = \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.u1.cout ;
assign \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.fas_s1  = \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.u1.s ;
assign \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.a  = \add_32s_32ns_32_2_1_U9.din0 ;
assign \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.b  = \add_32s_32ns_32_2_1_U9.din1 ;
assign \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.ce  = \add_32s_32ns_32_2_1_U9.ce ;
assign \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.clk  = \add_32s_32ns_32_2_1_U9.clk ;
assign \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.reset  = \add_32s_32ns_32_2_1_U9.reset ;
assign \add_32s_32ns_32_2_1_U9.dout  = \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.s ;
assign \add_32s_32ns_32_2_1_U9.ce  = 1'h1;
assign \add_32s_32ns_32_2_1_U9.clk  = ap_clk;
assign \add_32s_32ns_32_2_1_U9.din0  = { add_ln69_reg_529[16], add_ln69_reg_529[16], add_ln69_reg_529[16], add_ln69_reg_529[16], add_ln69_reg_529[16], add_ln69_reg_529[16], add_ln69_reg_529[16], add_ln69_reg_529[16], add_ln69_reg_529[16], add_ln69_reg_529[16], add_ln69_reg_529[16], add_ln69_reg_529[16], add_ln69_reg_529[16], add_ln69_reg_529[16], add_ln69_reg_529[16], add_ln69_reg_529 };
assign \add_32s_32ns_32_2_1_U9.din1  = ret_V_3_reg_524;
assign grp_fu_370_p2 = \add_32s_32ns_32_2_1_U9.dout ;
assign \add_32s_32ns_32_2_1_U9.reset  = ap_rst;
assign \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.ain_s0  = \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.a ;
assign \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.bin_s0  = \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.b ;
assign \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.s  = { \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.fas_s2 , \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.sum_s1  };
assign \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.u2.a  = \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.ain_s1 ;
assign \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.u2.b  = \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.bin_s1 ;
assign \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.u2.cin  = \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.carry_s1 ;
assign \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.facout_s2  = \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.u2.cout ;
assign \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.fas_s2  = \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.u2.s ;
assign \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.u1.a  = \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.a [15:0];
assign \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.u1.b  = \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.b [15:0];
assign \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.u1.cin  = 1'h0;
assign \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.facout_s1  = \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.u1.cout ;
assign \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.fas_s1  = \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.u1.s ;
assign \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.a  = \add_32s_32ns_32_2_1_U11.din0 ;
assign \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.b  = \add_32s_32ns_32_2_1_U11.din1 ;
assign \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.ce  = \add_32s_32ns_32_2_1_U11.ce ;
assign \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.clk  = \add_32s_32ns_32_2_1_U11.clk ;
assign \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.reset  = \add_32s_32ns_32_2_1_U11.reset ;
assign \add_32s_32ns_32_2_1_U11.dout  = \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.s ;
assign \add_32s_32ns_32_2_1_U11.ce  = 1'h1;
assign \add_32s_32ns_32_2_1_U11.clk  = ap_clk;
assign \add_32s_32ns_32_2_1_U11.din0  = { add_ln69_3_reg_559[5], add_ln69_3_reg_559[5], add_ln69_3_reg_559[5], add_ln69_3_reg_559[5], add_ln69_3_reg_559[5], add_ln69_3_reg_559[5], add_ln69_3_reg_559[5], add_ln69_3_reg_559[5], add_ln69_3_reg_559[5], add_ln69_3_reg_559[5], add_ln69_3_reg_559[5], add_ln69_3_reg_559[5], add_ln69_3_reg_559[5], add_ln69_3_reg_559[5], add_ln69_3_reg_559[5], add_ln69_3_reg_559[5], add_ln69_3_reg_559[5], add_ln69_3_reg_559[5], add_ln69_3_reg_559[5], add_ln69_3_reg_559[5], add_ln69_3_reg_559[5], add_ln69_3_reg_559[5], add_ln69_3_reg_559[5], add_ln69_3_reg_559[5], add_ln69_3_reg_559[5], add_ln69_3_reg_559[5], add_ln69_3_reg_559 };
assign \add_32s_32ns_32_2_1_U11.din1  = add_ln69_1_reg_554;
assign grp_fu_387_p2 = \add_32s_32ns_32_2_1_U11.dout ;
assign \add_32s_32ns_32_2_1_U11.reset  = ap_rst;
assign \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.ain_s0  = \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.a ;
assign \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.bin_s0  = \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.b ;
assign \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.s  = { \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.fas_s2 , \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.sum_s1  };
assign \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.a  = \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.ain_s1 ;
assign \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.b  = \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.bin_s1 ;
assign \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.cin  = \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.carry_s1 ;
assign \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.facout_s2  = \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.cout ;
assign \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.fas_s2  = \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.s ;
assign \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.a  = \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.a [15:0];
assign \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.b  = \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.b [15:0];
assign \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.cin  = 1'h0;
assign \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.facout_s1  = \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.cout ;
assign \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.fas_s1  = \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.s ;
assign \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.a  = \add_32ns_32ns_32_2_1_U6.din0 ;
assign \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.b  = \add_32ns_32ns_32_2_1_U6.din1 ;
assign \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.ce  = \add_32ns_32ns_32_2_1_U6.ce ;
assign \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.clk  = \add_32ns_32ns_32_2_1_U6.clk ;
assign \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.reset  = \add_32ns_32ns_32_2_1_U6.reset ;
assign \add_32ns_32ns_32_2_1_U6.dout  = \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.s ;
assign \add_32ns_32ns_32_2_1_U6.ce  = 1'h1;
assign \add_32ns_32ns_32_2_1_U6.clk  = ap_clk;
assign \add_32ns_32ns_32_2_1_U6.din0  = ret_V_3_cast_reg_492;
assign \add_32ns_32ns_32_2_1_U6.din1  = 32'd1;
assign grp_fu_308_p2 = \add_32ns_32ns_32_2_1_U6.dout ;
assign \add_32ns_32ns_32_2_1_U6.reset  = ap_rst;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.ain_s0  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.a ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.bin_s0  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.b ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.s  = { \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.fas_s2 , \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.sum_s1  };
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.a  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.ain_s1 ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.b  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.bin_s1 ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.cin  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.carry_s1 ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.facout_s2  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.cout ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.fas_s2  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.s ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.a  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.a [15:0];
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.b  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.b [15:0];
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.cin  = 1'h0;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.facout_s1  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.cout ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.fas_s1  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.s ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.a  = \add_32ns_32ns_32_2_1_U12.din0 ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.b  = \add_32ns_32ns_32_2_1_U12.din1 ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.ce  = \add_32ns_32ns_32_2_1_U12.ce ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.clk  = \add_32ns_32ns_32_2_1_U12.clk ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.reset  = \add_32ns_32ns_32_2_1_U12.reset ;
assign \add_32ns_32ns_32_2_1_U12.dout  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.s ;
assign \add_32ns_32ns_32_2_1_U12.ce  = 1'h1;
assign \add_32ns_32ns_32_2_1_U12.clk  = ap_clk;
assign \add_32ns_32ns_32_2_1_U12.din0  = op_28_V_reg_569;
assign \add_32ns_32ns_32_2_1_U12.din1  = select_ln1192_reg_574;
assign grp_fu_400_p2 = \add_32ns_32ns_32_2_1_U12.dout ;
assign \add_32ns_32ns_32_2_1_U12.reset  = ap_rst;
assign \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.ain_s0  = \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.a ;
assign \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.bin_s0  = \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.b ;
assign \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.s  = { \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.fas_s2 , \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.sum_s1  };
assign \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.u2.a  = \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.ain_s1 ;
assign \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.u2.b  = \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.bin_s1 ;
assign \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.u2.cin  = \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.carry_s1 ;
assign \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.facout_s2  = \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.u2.cout ;
assign \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.fas_s2  = \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.u2.s ;
assign \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.u1.a  = \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.a [7:0];
assign \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.u1.b  = \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.b [7:0];
assign \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.u1.cin  = 1'h0;
assign \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.facout_s1  = \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.u1.cout ;
assign \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.fas_s1  = \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.u1.s ;
assign \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.a  = \add_17s_17s_17_2_1_U7.din0 ;
assign \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.b  = \add_17s_17s_17_2_1_U7.din1 ;
assign \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.ce  = \add_17s_17s_17_2_1_U7.ce ;
assign \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.clk  = \add_17s_17s_17_2_1_U7.clk ;
assign \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.reset  = \add_17s_17s_17_2_1_U7.reset ;
assign \add_17s_17s_17_2_1_U7.dout  = \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.s ;
assign \add_17s_17s_17_2_1_U7.ce  = 1'h1;
assign \add_17s_17s_17_2_1_U7.clk  = ap_clk;
assign \add_17s_17s_17_2_1_U7.din0  = { op_16[15], op_16 };
assign \add_17s_17s_17_2_1_U7.din1  = { op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13 };
assign grp_fu_333_p2 = \add_17s_17s_17_2_1_U7.dout ;
assign \add_17s_17s_17_2_1_U7.reset  = ap_rst;
assign \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.ain_s0  = \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.a ;
assign \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.bin_s0  = \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.b ;
assign \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.s  = { \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.fas_s2 , \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.sum_s1  };
assign \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.u2.a  = \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.ain_s1 ;
assign \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.u2.b  = \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.bin_s1 ;
assign \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.u2.cin  = \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.carry_s1 ;
assign \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.facout_s2  = \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.u2.cout ;
assign \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.fas_s2  = \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.u2.s ;
assign \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.u1.a  = \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.a [5:0];
assign \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.u1.b  = \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.b [5:0];
assign \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.u1.cin  = 1'h0;
assign \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.facout_s1  = \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.u1.cout ;
assign \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.fas_s1  = \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.u1.s ;
assign \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.a  = \add_12ns_12s_12_2_1_U2.din0 ;
assign \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.b  = \add_12ns_12s_12_2_1_U2.din1 ;
assign \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.ce  = \add_12ns_12s_12_2_1_U2.ce ;
assign \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.clk  = \add_12ns_12s_12_2_1_U2.clk ;
assign \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.reset  = \add_12ns_12s_12_2_1_U2.reset ;
assign \add_12ns_12s_12_2_1_U2.dout  = \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.s ;
assign \add_12ns_12s_12_2_1_U2.ce  = 1'h1;
assign \add_12ns_12s_12_2_1_U2.clk  = ap_clk;
assign \add_12ns_12s_12_2_1_U2.din0  = { ret_reg_415, 3'h0 };
assign \add_12ns_12s_12_2_1_U2.din1  = { op_10[3], op_10[3], op_10[3], op_10[3], op_10[3], op_10[3], op_10[3], op_10[3], op_10 };
assign grp_fu_201_p2 = \add_12ns_12s_12_2_1_U2.dout ;
assign \add_12ns_12s_12_2_1_U2.reset  = ap_rst;
assign \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.ain_s0  = \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.a ;
assign \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.bin_s0  = \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.b ;
assign \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.s  = { \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.fas_s2 , \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.sum_s1  };
assign \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.u2.a  = \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.ain_s1 ;
assign \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.u2.b  = \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.bin_s1 ;
assign \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.u2.cin  = \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.carry_s1 ;
assign \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.facout_s2  = \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.u2.cout ;
assign \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.fas_s2  = \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.u2.s ;
assign \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.u1.a  = \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.a [4:0];
assign \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.u1.b  = \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.b [4:0];
assign \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.u1.cin  = 1'h0;
assign \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.facout_s1  = \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.u1.cout ;
assign \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.fas_s1  = \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.u1.s ;
assign \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.a  = \add_10s_10ns_10_2_1_U3.din0 ;
assign \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.b  = \add_10s_10ns_10_2_1_U3.din1 ;
assign \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.ce  = \add_10s_10ns_10_2_1_U3.ce ;
assign \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.clk  = \add_10s_10ns_10_2_1_U3.clk ;
assign \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.reset  = \add_10s_10ns_10_2_1_U3.reset ;
assign \add_10s_10ns_10_2_1_U3.dout  = \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.s ;
assign \add_10s_10ns_10_2_1_U3.ce  = 1'h1;
assign \add_10s_10ns_10_2_1_U3.clk  = ap_clk;
assign \add_10s_10ns_10_2_1_U3.din0  = { tmp_1_reg_440[8], tmp_1_reg_440 };
assign \add_10s_10ns_10_2_1_U3.din1  = 10'h001;
assign grp_fu_230_p2 = \add_10s_10ns_10_2_1_U3.dout ;
assign \add_10s_10ns_10_2_1_U3.reset  = ap_rst;
assign \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.ain_s0  = \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.a ;
assign \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.bin_s0  = \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.b ;
assign \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.s  = { \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.fas_s2 , \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.sum_s1  };
assign \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.u2.a  = \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.ain_s1 ;
assign \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.u2.b  = \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.bin_s1 ;
assign \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.u2.cin  = \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.carry_s1 ;
assign \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.facout_s2  = \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.u2.cout ;
assign \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.fas_s2  = \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.u2.s ;
assign \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.u1.a  = \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.a [4:0];
assign \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.u1.b  = \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.b [4:0];
assign \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.u1.cin  = 1'h0;
assign \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.facout_s1  = \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.u1.cout ;
assign \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.fas_s1  = \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.u1.s ;
assign \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.a  = \add_10ns_10ns_10_2_1_U4.din0 ;
assign \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.b  = \add_10ns_10ns_10_2_1_U4.din1 ;
assign \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.ce  = \add_10ns_10ns_10_2_1_U4.ce ;
assign \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.clk  = \add_10ns_10ns_10_2_1_U4.clk ;
assign \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.reset  = \add_10ns_10ns_10_2_1_U4.reset ;
assign \add_10ns_10ns_10_2_1_U4.dout  = \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.s ;
assign \add_10ns_10ns_10_2_1_U4.ce  = 1'h1;
assign \add_10ns_10ns_10_2_1_U4.clk  = ap_clk;
assign \add_10ns_10ns_10_2_1_U4.din0  = ret_V_1_reg_457;
assign \add_10ns_10ns_10_2_1_U4.din1  = select_ln69_reg_462;
assign grp_fu_263_p2 = \add_10ns_10ns_10_2_1_U4.dout ;
assign \add_10ns_10ns_10_2_1_U4.reset  = ap_rst;
endmodule


// Machine B:
// Processed by function `add_clk_enable_signal` in `verilog_tricks.py`.
// Processed by function `remove_reset_signal` in `verilog_tricks.py`.
module top_B (
  ap_clk,
  ap_start,
  ap_done,
  ap_idle,
  ap_ready,
  op_0,
  op_1,
  op_5,
  op_6,
  op_10,
  op_11,
  op_12,
  op_13,
  op_14,
  op_15,
  op_16,
  op_17,
  op_18,
  op_30,
  op_30_ap_vld,
clk_enable
);
input clk_enable;


input ap_clk;
wire ap_rst;
assign ap_rst = op_30_ap_vld;
input ap_start;
input [1:0] op_0;
input [3:0] op_1;
input [3:0] op_10;
input op_11;
input [3:0] op_12;
input [7:0] op_13;
input [3:0] op_14;
input op_15;
input [15:0] op_16;
input [3:0] op_17;
input op_18;
input [3:0] op_5;
input [7:0] op_6;
output ap_done;
output ap_idle;
output ap_ready;
output [31:0] op_30;
output op_30_ap_vld;


reg [4:0] \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.ain_s1 ;
reg [4:0] \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.bin_s1 ;
reg \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.carry_s1 ;
reg [4:0] \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.sum_s1 ;
reg [4:0] \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.ain_s1 ;
reg [4:0] \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.bin_s1 ;
reg \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.carry_s1 ;
reg [4:0] \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.sum_s1 ;
reg [5:0] \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.ain_s1 ;
reg [5:0] \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.bin_s1 ;
reg \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.carry_s1 ;
reg [5:0] \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.sum_s1 ;
reg [8:0] \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.ain_s1 ;
reg [8:0] \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.bin_s1 ;
reg \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.carry_s1 ;
reg [7:0] \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.sum_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.ain_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.bin_s1 ;
reg \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.carry_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.sum_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.ain_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.bin_s1 ;
reg \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.carry_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.sum_s1 ;
reg [15:0] \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.ain_s1 ;
reg [15:0] \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.bin_s1 ;
reg \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.carry_s1 ;
reg [15:0] \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.sum_s1 ;
reg [15:0] \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.ain_s1 ;
reg [15:0] \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.bin_s1 ;
reg \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.carry_s1 ;
reg [15:0] \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.sum_s1 ;
reg [17:0] \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.ain_s1 ;
reg [17:0] \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.bin_s1 ;
reg \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.carry_s1 ;
reg [16:0] \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.sum_s1 ;
reg [2:0] \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.ain_s1 ;
reg [2:0] \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.bin_s1 ;
reg \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.carry_s1 ;
reg [1:0] \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.sum_s1 ;
reg [2:0] \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.ain_s1 ;
reg [2:0] \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.bin_s1 ;
reg \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.carry_s1 ;
reg [2:0] \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.sum_s1 ;
reg [4:0] \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.ain_s1 ;
reg [4:0] \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.bin_s1 ;
reg \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.carry_s1 ;
reg [3:0] \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.sum_s1 ;
reg [31:0] add_ln691_1_reg_504;
reg [9:0] add_ln691_reg_452;
reg [31:0] add_ln69_1_reg_554;
reg [4:0] add_ln69_2_reg_534;
reg [5:0] add_ln69_3_reg_559;
reg [16:0] add_ln69_reg_529;
reg [20:0] ap_CS_fsm = 21'h000001;
reg icmp_ln851_1_reg_482;
reg icmp_ln851_reg_430;
reg [9:0] op_22_V_reg_467;
reg [31:0] op_28_V_reg_569;
reg [9:0] ret_V_1_reg_457;
reg [34:0] ret_V_2_reg_487;
reg [31:0] ret_V_3_cast_reg_492;
reg [31:0] ret_V_3_reg_524;
reg [11:0] ret_V_reg_435;
reg [8:0] ret_reg_415;
reg [31:0] select_ln1192_reg_574;
reg [8:0] select_ln215_reg_405;
reg [4:0] select_ln69_1_reg_499;
reg [9:0] select_ln69_reg_462;
reg [9:0] sext_ln850_reg_445;
reg [8:0] tmp_1_reg_440;
wire [31:0] _000_;
wire [9:0] _001_;
wire [31:0] _002_;
wire [4:0] _003_;
wire [5:0] _004_;
wire [16:0] _005_;
wire [20:0] _006_;
wire _007_;
wire _008_;
wire [9:0] _009_;
wire [31:0] _010_;
wire [9:0] _011_;
wire [34:0] _012_;
wire [31:0] _013_;
wire [31:0] _014_;
wire [11:0] _015_;
wire [8:0] _016_;
wire [31:0] _017_;
wire [8:0] _018_;
wire [4:0] _019_;
wire [9:0] _020_;
wire [9:0] _021_;
wire [8:0] _022_;
wire [1:0] _023_;
wire _024_;
wire _025_;
wire _026_;
wire _027_;
wire _028_;
wire [4:0] _029_;
wire [4:0] _030_;
wire _031_;
wire [4:0] _032_;
wire [5:0] _033_;
wire [5:0] _034_;
wire [4:0] _035_;
wire [4:0] _036_;
wire _037_;
wire [4:0] _038_;
wire [5:0] _039_;
wire [5:0] _040_;
wire [5:0] _041_;
wire [5:0] _042_;
wire _043_;
wire [5:0] _044_;
wire [6:0] _045_;
wire [6:0] _046_;
wire [8:0] _047_;
wire [8:0] _048_;
wire _049_;
wire [7:0] _050_;
wire [8:0] _051_;
wire [9:0] _052_;
wire [15:0] _053_;
wire [15:0] _054_;
wire _055_;
wire [15:0] _056_;
wire [16:0] _057_;
wire [16:0] _058_;
wire [15:0] _059_;
wire [15:0] _060_;
wire _061_;
wire [15:0] _062_;
wire [16:0] _063_;
wire [16:0] _064_;
wire [15:0] _065_;
wire [15:0] _066_;
wire _067_;
wire [15:0] _068_;
wire [16:0] _069_;
wire [16:0] _070_;
wire [15:0] _071_;
wire [15:0] _072_;
wire _073_;
wire [15:0] _074_;
wire [16:0] _075_;
wire [16:0] _076_;
wire [17:0] _077_;
wire [17:0] _078_;
wire _079_;
wire [16:0] _080_;
wire [17:0] _081_;
wire [18:0] _082_;
wire [2:0] _083_;
wire [2:0] _084_;
wire _085_;
wire [1:0] _086_;
wire [2:0] _087_;
wire [3:0] _088_;
wire [2:0] _089_;
wire [2:0] _090_;
wire _091_;
wire [2:0] _092_;
wire [3:0] _093_;
wire [3:0] _094_;
wire [4:0] _095_;
wire [4:0] _096_;
wire _097_;
wire [3:0] _098_;
wire [4:0] _099_;
wire [5:0] _100_;
wire _101_;
wire _102_;
wire _103_;
wire _104_;
wire _105_;
wire _106_;
wire _107_;
wire _108_;
wire _109_;
wire _110_;
wire _111_;
wire _112_;
wire _113_;
wire _114_;
wire _115_;
wire _116_;
wire _117_;
wire _118_;
wire _119_;
wire _120_;
wire _121_;
wire _122_;
wire _123_;
wire \add_10ns_10ns_10_2_1_U4.ce ;
wire \add_10ns_10ns_10_2_1_U4.clk ;
wire [9:0] \add_10ns_10ns_10_2_1_U4.din0 ;
wire [9:0] \add_10ns_10ns_10_2_1_U4.din1 ;
wire [9:0] \add_10ns_10ns_10_2_1_U4.dout ;
wire \add_10ns_10ns_10_2_1_U4.reset ;
wire [9:0] \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.a ;
wire [9:0] \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.ain_s0 ;
wire [9:0] \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.b ;
wire [9:0] \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.bin_s0 ;
wire \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.ce ;
wire \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.clk ;
wire \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.facout_s1 ;
wire \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.facout_s2 ;
wire [4:0] \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.fas_s1 ;
wire [4:0] \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.fas_s2 ;
wire \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.reset ;
wire [9:0] \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.s ;
wire [4:0] \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.u1.a ;
wire [4:0] \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.u1.b ;
wire \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.u1.cin ;
wire \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.u1.cout ;
wire [4:0] \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.u1.s ;
wire [4:0] \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.u2.a ;
wire [4:0] \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.u2.b ;
wire \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.u2.cin ;
wire \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.u2.cout ;
wire [4:0] \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.u2.s ;
wire \add_10s_10ns_10_2_1_U3.ce ;
wire \add_10s_10ns_10_2_1_U3.clk ;
wire [9:0] \add_10s_10ns_10_2_1_U3.din0 ;
wire [9:0] \add_10s_10ns_10_2_1_U3.din1 ;
wire [9:0] \add_10s_10ns_10_2_1_U3.dout ;
wire \add_10s_10ns_10_2_1_U3.reset ;
wire [9:0] \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.a ;
wire [9:0] \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.ain_s0 ;
wire [9:0] \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.b ;
wire [9:0] \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.bin_s0 ;
wire \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.ce ;
wire \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.clk ;
wire \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.facout_s1 ;
wire \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.facout_s2 ;
wire [4:0] \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.fas_s1 ;
wire [4:0] \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.fas_s2 ;
wire \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.reset ;
wire [9:0] \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.s ;
wire [4:0] \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.u1.a ;
wire [4:0] \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.u1.b ;
wire \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.u1.cin ;
wire \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.u1.cout ;
wire [4:0] \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.u1.s ;
wire [4:0] \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.u2.a ;
wire [4:0] \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.u2.b ;
wire \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.u2.cin ;
wire \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.u2.cout ;
wire [4:0] \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.u2.s ;
wire \add_12ns_12s_12_2_1_U2.ce ;
wire \add_12ns_12s_12_2_1_U2.clk ;
wire [11:0] \add_12ns_12s_12_2_1_U2.din0 ;
wire [11:0] \add_12ns_12s_12_2_1_U2.din1 ;
wire [11:0] \add_12ns_12s_12_2_1_U2.dout ;
wire \add_12ns_12s_12_2_1_U2.reset ;
wire [11:0] \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.a ;
wire [11:0] \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.ain_s0 ;
wire [11:0] \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.b ;
wire [11:0] \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.bin_s0 ;
wire \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.ce ;
wire \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.clk ;
wire \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.facout_s1 ;
wire \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.facout_s2 ;
wire [5:0] \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.fas_s1 ;
wire [5:0] \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.fas_s2 ;
wire \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.reset ;
wire [11:0] \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.s ;
wire [5:0] \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.u1.a ;
wire [5:0] \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.u1.b ;
wire \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.u1.cin ;
wire \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.u1.cout ;
wire [5:0] \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.u1.s ;
wire [5:0] \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.u2.a ;
wire [5:0] \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.u2.b ;
wire \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.u2.cin ;
wire \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.u2.cout ;
wire [5:0] \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.u2.s ;
wire \add_17s_17s_17_2_1_U7.ce ;
wire \add_17s_17s_17_2_1_U7.clk ;
wire [16:0] \add_17s_17s_17_2_1_U7.din0 ;
wire [16:0] \add_17s_17s_17_2_1_U7.din1 ;
wire [16:0] \add_17s_17s_17_2_1_U7.dout ;
wire \add_17s_17s_17_2_1_U7.reset ;
wire [16:0] \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.a ;
wire [16:0] \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.ain_s0 ;
wire [16:0] \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.b ;
wire [16:0] \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.bin_s0 ;
wire \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.ce ;
wire \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.clk ;
wire \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.facout_s1 ;
wire \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.facout_s2 ;
wire [7:0] \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.fas_s1 ;
wire [8:0] \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.fas_s2 ;
wire \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.reset ;
wire [16:0] \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.s ;
wire [7:0] \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.u1.a ;
wire [7:0] \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.u1.b ;
wire \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.u1.cin ;
wire \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.u1.cout ;
wire [7:0] \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.u1.s ;
wire [8:0] \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.u2.a ;
wire [8:0] \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.u2.b ;
wire \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.u2.cin ;
wire \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.u2.cout ;
wire [8:0] \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.u2.s ;
wire \add_32ns_32ns_32_2_1_U12.ce ;
wire \add_32ns_32ns_32_2_1_U12.clk ;
wire [31:0] \add_32ns_32ns_32_2_1_U12.din0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U12.din1 ;
wire [31:0] \add_32ns_32ns_32_2_1_U12.dout ;
wire \add_32ns_32ns_32_2_1_U12.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.a ;
wire [31:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.ain_s0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.b ;
wire [31:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.bin_s0 ;
wire \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.ce ;
wire \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.clk ;
wire \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.facout_s1 ;
wire \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.facout_s2 ;
wire [15:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.fas_s1 ;
wire [15:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.fas_s2 ;
wire \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.b ;
wire \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.cin ;
wire \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.b ;
wire \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.cin ;
wire \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.s ;
wire \add_32ns_32ns_32_2_1_U6.ce ;
wire \add_32ns_32ns_32_2_1_U6.clk ;
wire [31:0] \add_32ns_32ns_32_2_1_U6.din0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U6.din1 ;
wire [31:0] \add_32ns_32ns_32_2_1_U6.dout ;
wire \add_32ns_32ns_32_2_1_U6.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.a ;
wire [31:0] \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.ain_s0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.b ;
wire [31:0] \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.bin_s0 ;
wire \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.ce ;
wire \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.clk ;
wire \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.facout_s1 ;
wire \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.facout_s2 ;
wire [15:0] \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.fas_s1 ;
wire [15:0] \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.fas_s2 ;
wire \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.b ;
wire \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.cin ;
wire \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.b ;
wire \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.cin ;
wire \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.s ;
wire \add_32s_32ns_32_2_1_U11.ce ;
wire \add_32s_32ns_32_2_1_U11.clk ;
wire [31:0] \add_32s_32ns_32_2_1_U11.din0 ;
wire [31:0] \add_32s_32ns_32_2_1_U11.din1 ;
wire [31:0] \add_32s_32ns_32_2_1_U11.dout ;
wire \add_32s_32ns_32_2_1_U11.reset ;
wire [31:0] \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.a ;
wire [31:0] \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.ain_s0 ;
wire [31:0] \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.b ;
wire [31:0] \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.bin_s0 ;
wire \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.ce ;
wire \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.clk ;
wire \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.facout_s1 ;
wire \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.facout_s2 ;
wire [15:0] \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.fas_s1 ;
wire [15:0] \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.fas_s2 ;
wire \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.reset ;
wire [31:0] \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.s ;
wire [15:0] \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.u1.a ;
wire [15:0] \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.u1.b ;
wire \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.u1.cin ;
wire \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.u1.cout ;
wire [15:0] \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.u1.s ;
wire [15:0] \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.u2.a ;
wire [15:0] \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.u2.b ;
wire \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.u2.cin ;
wire \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.u2.cout ;
wire [15:0] \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.u2.s ;
wire \add_32s_32ns_32_2_1_U9.ce ;
wire \add_32s_32ns_32_2_1_U9.clk ;
wire [31:0] \add_32s_32ns_32_2_1_U9.din0 ;
wire [31:0] \add_32s_32ns_32_2_1_U9.din1 ;
wire [31:0] \add_32s_32ns_32_2_1_U9.dout ;
wire \add_32s_32ns_32_2_1_U9.reset ;
wire [31:0] \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.a ;
wire [31:0] \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.ain_s0 ;
wire [31:0] \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.b ;
wire [31:0] \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.bin_s0 ;
wire \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.ce ;
wire \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.clk ;
wire \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.facout_s1 ;
wire \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.facout_s2 ;
wire [15:0] \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.fas_s1 ;
wire [15:0] \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.fas_s2 ;
wire \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.reset ;
wire [31:0] \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.s ;
wire [15:0] \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.u1.a ;
wire [15:0] \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.u1.b ;
wire \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.u1.cin ;
wire \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.u1.cout ;
wire [15:0] \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.u1.s ;
wire [15:0] \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.u2.a ;
wire [15:0] \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.u2.b ;
wire \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.u2.cin ;
wire \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.u2.cout ;
wire [15:0] \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.u2.s ;
wire \add_35s_35s_35_2_1_U5.ce ;
wire \add_35s_35s_35_2_1_U5.clk ;
wire [34:0] \add_35s_35s_35_2_1_U5.din0 ;
wire [34:0] \add_35s_35s_35_2_1_U5.din1 ;
wire [34:0] \add_35s_35s_35_2_1_U5.dout ;
wire \add_35s_35s_35_2_1_U5.reset ;
wire [34:0] \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.a ;
wire [34:0] \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.ain_s0 ;
wire [34:0] \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.b ;
wire [34:0] \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.bin_s0 ;
wire \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.ce ;
wire \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.clk ;
wire \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.facout_s1 ;
wire \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.facout_s2 ;
wire [16:0] \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.fas_s1 ;
wire [17:0] \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.fas_s2 ;
wire \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.reset ;
wire [34:0] \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.s ;
wire [16:0] \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.u1.a ;
wire [16:0] \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.u1.b ;
wire \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.u1.cin ;
wire \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.u1.cout ;
wire [16:0] \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.u1.s ;
wire [17:0] \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.u2.a ;
wire [17:0] \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.u2.b ;
wire \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.u2.cin ;
wire \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.u2.cout ;
wire [17:0] \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.u2.s ;
wire \add_5ns_5ns_5_2_1_U8.ce ;
wire \add_5ns_5ns_5_2_1_U8.clk ;
wire [4:0] \add_5ns_5ns_5_2_1_U8.din0 ;
wire [4:0] \add_5ns_5ns_5_2_1_U8.din1 ;
wire [4:0] \add_5ns_5ns_5_2_1_U8.dout ;
wire \add_5ns_5ns_5_2_1_U8.reset ;
wire [4:0] \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.a ;
wire [4:0] \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.ain_s0 ;
wire [4:0] \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.b ;
wire [4:0] \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.bin_s0 ;
wire \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.ce ;
wire \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.clk ;
wire \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.facout_s1 ;
wire \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.facout_s2 ;
wire [1:0] \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.fas_s1 ;
wire [2:0] \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.fas_s2 ;
wire \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.reset ;
wire [4:0] \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.s ;
wire [1:0] \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.u1.a ;
wire [1:0] \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.u1.b ;
wire \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.u1.cin ;
wire \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.u1.cout ;
wire [1:0] \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.u1.s ;
wire [2:0] \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.u2.a ;
wire [2:0] \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.u2.b ;
wire \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.u2.cin ;
wire \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.u2.cout ;
wire [2:0] \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.u2.s ;
wire \add_6s_6s_6_2_1_U10.ce ;
wire \add_6s_6s_6_2_1_U10.clk ;
wire [5:0] \add_6s_6s_6_2_1_U10.din0 ;
wire [5:0] \add_6s_6s_6_2_1_U10.din1 ;
wire [5:0] \add_6s_6s_6_2_1_U10.dout ;
wire \add_6s_6s_6_2_1_U10.reset ;
wire [5:0] \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.a ;
wire [5:0] \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.ain_s0 ;
wire [5:0] \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.b ;
wire [5:0] \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.bin_s0 ;
wire \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.ce ;
wire \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.clk ;
wire \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.facout_s1 ;
wire \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.facout_s2 ;
wire [2:0] \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.fas_s1 ;
wire [2:0] \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.fas_s2 ;
wire \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.reset ;
wire [5:0] \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.s ;
wire [2:0] \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.u1.a ;
wire [2:0] \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.u1.b ;
wire \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.u1.cin ;
wire \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.u1.cout ;
wire [2:0] \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.u1.s ;
wire [2:0] \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.u2.a ;
wire [2:0] \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.u2.b ;
wire \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.u2.cin ;
wire \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.u2.cout ;
wire [2:0] \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.u2.s ;
wire \add_9s_9ns_9_2_1_U1.ce ;
wire \add_9s_9ns_9_2_1_U1.clk ;
wire [8:0] \add_9s_9ns_9_2_1_U1.din0 ;
wire [8:0] \add_9s_9ns_9_2_1_U1.din1 ;
wire [8:0] \add_9s_9ns_9_2_1_U1.dout ;
wire \add_9s_9ns_9_2_1_U1.reset ;
wire [8:0] \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.a ;
wire [8:0] \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.ain_s0 ;
wire [8:0] \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.b ;
wire [8:0] \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.bin_s0 ;
wire \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.ce ;
wire \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.clk ;
wire \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.facout_s1 ;
wire \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.facout_s2 ;
wire [3:0] \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.fas_s1 ;
wire [4:0] \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.fas_s2 ;
wire \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.reset ;
wire [8:0] \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.s ;
wire [3:0] \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.u1.a ;
wire [3:0] \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.u1.b ;
wire \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.u1.cin ;
wire \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.u1.cout ;
wire [3:0] \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.u1.s ;
wire [4:0] \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.u2.a ;
wire [4:0] \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.u2.b ;
wire \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.u2.cin ;
wire \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.u2.cout ;
wire [4:0] \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.u2.s ;
wire ap_CS_fsm_state1;
wire ap_CS_fsm_state10;
wire ap_CS_fsm_state11;
wire ap_CS_fsm_state12;
wire ap_CS_fsm_state13;
wire ap_CS_fsm_state14;
wire ap_CS_fsm_state15;
wire ap_CS_fsm_state16;
wire ap_CS_fsm_state17;
wire ap_CS_fsm_state18;
wire ap_CS_fsm_state19;
wire ap_CS_fsm_state2;
wire ap_CS_fsm_state20;
wire ap_CS_fsm_state21;
wire ap_CS_fsm_state3;
wire ap_CS_fsm_state4;
wire ap_CS_fsm_state5;
wire ap_CS_fsm_state6;
wire ap_CS_fsm_state7;
wire ap_CS_fsm_state8;
wire ap_CS_fsm_state9;
wire [20:0] ap_NS_fsm;
wire ap_clk;
wire ap_done;
wire ap_idle;
wire ap_ready;
wire ap_rst;
wire ap_start;
wire [8:0] grp_fu_185_p0;
wire [8:0] grp_fu_185_p2;
wire [11:0] grp_fu_201_p0;
wire [11:0] grp_fu_201_p1;
wire [11:0] grp_fu_201_p2;
wire [9:0] grp_fu_230_p0;
wire [9:0] grp_fu_230_p2;
wire [9:0] grp_fu_263_p2;
wire [34:0] grp_fu_282_p0;
wire [34:0] grp_fu_282_p1;
wire [34:0] grp_fu_282_p2;
wire [31:0] grp_fu_308_p2;
wire [16:0] grp_fu_333_p0;
wire [16:0] grp_fu_333_p1;
wire [16:0] grp_fu_333_p2;
wire [4:0] grp_fu_339_p0;
wire [4:0] grp_fu_339_p2;
wire [31:0] grp_fu_370_p0;
wire [31:0] grp_fu_370_p2;
wire [5:0] grp_fu_378_p0;
wire [5:0] grp_fu_378_p1;
wire [5:0] grp_fu_378_p2;
wire [31:0] grp_fu_387_p0;
wire [31:0] grp_fu_387_p2;
wire [31:0] grp_fu_400_p2;
wire icmp_ln851_1_fu_292_p2;
wire icmp_ln851_fu_211_p2;
wire [1:0] op_0;
wire [3:0] op_1;
wire [3:0] op_10;
wire op_11;
wire [3:0] op_12;
wire [7:0] op_13;
wire [3:0] op_14;
wire op_15;
wire [15:0] op_16;
wire [3:0] op_17;
wire op_18;
wire [31:0] op_30;
wire op_30_ap_vld;
wire [3:0] op_5;
wire [7:0] op_6;
wire op_8_V_fu_169_p1;
wire p_Result_1_fu_344_p3;
wire p_Result_s_fu_236_p3;
wire [9:0] ret_V_1_fu_248_p3;
wire [31:0] ret_V_3_fu_356_p3;
wire [31:0] select_ln1192_fu_392_p3;
wire [8:0] select_ln215_fu_173_p3;
wire [4:0] select_ln69_1_fu_313_p3;
wire [9:0] select_ln69_fu_255_p3;
wire [31:0] select_ln850_1_fu_351_p3;
wire [9:0] select_ln850_fu_243_p3;
wire [3:0] sext_ln1192_fu_190_p0;
wire [3:0] sext_ln703_fu_267_p0;
wire [9:0] sext_ln850_fu_227_p1;
wire [11:0] tmp_fu_271_p3;
wire [3:0] trunc_ln851_1_fu_288_p0;
wire [1:0] trunc_ln851_1_fu_288_p1;
wire [3:0] trunc_ln851_fu_207_p0;
wire [2:0] trunc_ln851_fu_207_p1;


assign _024_ = ap_CS_fsm[13] & icmp_ln851_1_reg_482;
assign _025_ = icmp_ln851_reg_430 & ap_CS_fsm[6];
assign _026_ = _028_ & ap_CS_fsm[0];
assign _027_ = ap_start & ap_CS_fsm[0];
assign _028_ = ~ ap_start;
always @(posedge \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.clk )
\add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.bin_s1  <= _030_;
always @(posedge \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.clk )
\add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.ain_s1  <= _029_;
always @(posedge \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.clk )
\add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.sum_s1  <= _032_;
always @(posedge \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.clk )
\add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.carry_s1  <= _031_;
assign _030_ = \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.ce  ? \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.b [9:5] : \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.bin_s1 ;
assign _029_ = \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.ce  ? \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.a [9:5] : \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.ain_s1 ;
assign _031_ = \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.ce  ? \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.facout_s1  : \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.carry_s1 ;
assign _032_ = \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.ce  ? \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.fas_s1  : \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.sum_s1 ;
assign _033_ = \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.u1.a  + \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.u1.b ;
assign { \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.u1.cout , \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.u1.s  } = _033_ + \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.u1.cin ;
assign _034_ = \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.u2.a  + \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.u2.b ;
assign { \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.u2.cout , \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.u2.s  } = _034_ + \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.u2.cin ;
always @(posedge \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.clk )
\add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.bin_s1  <= _036_;
always @(posedge \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.clk )
\add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.ain_s1  <= _035_;
always @(posedge \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.clk )
\add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.sum_s1  <= _038_;
always @(posedge \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.clk )
\add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.carry_s1  <= _037_;
assign _036_ = \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.ce  ? \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.b [9:5] : \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.bin_s1 ;
assign _035_ = \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.ce  ? \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.a [9:5] : \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.ain_s1 ;
assign _037_ = \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.ce  ? \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.facout_s1  : \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.carry_s1 ;
assign _038_ = \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.ce  ? \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.fas_s1  : \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.sum_s1 ;
assign _039_ = \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.u1.a  + \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.u1.b ;
assign { \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.u1.cout , \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.u1.s  } = _039_ + \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.u1.cin ;
assign _040_ = \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.u2.a  + \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.u2.b ;
assign { \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.u2.cout , \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.u2.s  } = _040_ + \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.u2.cin ;
always @(posedge \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.clk )
\add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.bin_s1  <= _042_;
always @(posedge \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.clk )
\add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.ain_s1  <= _041_;
always @(posedge \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.clk )
\add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.sum_s1  <= _044_;
always @(posedge \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.clk )
\add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.carry_s1  <= _043_;
assign _042_ = \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.ce  ? \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.b [11:6] : \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.bin_s1 ;
assign _041_ = \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.ce  ? \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.a [11:6] : \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.ain_s1 ;
assign _043_ = \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.ce  ? \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.facout_s1  : \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.carry_s1 ;
assign _044_ = \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.ce  ? \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.fas_s1  : \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.sum_s1 ;
assign _045_ = \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.u1.a  + \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.u1.b ;
assign { \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.u1.cout , \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.u1.s  } = _045_ + \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.u1.cin ;
assign _046_ = \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.u2.a  + \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.u2.b ;
assign { \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.u2.cout , \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.u2.s  } = _046_ + \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.u2.cin ;
always @(posedge \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.clk )
\add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.bin_s1  <= _048_;
always @(posedge \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.clk )
\add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.ain_s1  <= _047_;
always @(posedge \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.clk )
\add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.sum_s1  <= _050_;
always @(posedge \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.clk )
\add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.carry_s1  <= _049_;
assign _048_ = \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.ce  ? \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.b [16:8] : \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.bin_s1 ;
assign _047_ = \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.ce  ? \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.a [16:8] : \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.ain_s1 ;
assign _049_ = \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.ce  ? \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.facout_s1  : \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.carry_s1 ;
assign _050_ = \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.ce  ? \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.fas_s1  : \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.sum_s1 ;
assign _051_ = \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.u1.a  + \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.u1.b ;
assign { \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.u1.cout , \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.u1.s  } = _051_ + \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.u1.cin ;
assign _052_ = \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.u2.a  + \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.u2.b ;
assign { \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.u2.cout , \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.u2.s  } = _052_ + \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.u2.cin ;
always @(posedge \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.clk )
\add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.bin_s1  <= _054_;
always @(posedge \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.clk )
\add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.ain_s1  <= _053_;
always @(posedge \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.clk )
\add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.sum_s1  <= _056_;
always @(posedge \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.clk )
\add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.carry_s1  <= _055_;
assign _054_ = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.ce  ? \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.b [31:16] : \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.bin_s1 ;
assign _053_ = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.ce  ? \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.a [31:16] : \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.ain_s1 ;
assign _055_ = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.ce  ? \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.facout_s1  : \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.carry_s1 ;
assign _056_ = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.ce  ? \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.fas_s1  : \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.sum_s1 ;
assign _057_ = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.a  + \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.b ;
assign { \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.cout , \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.s  } = _057_ + \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.cin ;
assign _058_ = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.a  + \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.b ;
assign { \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.cout , \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.s  } = _058_ + \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.cin ;
always @(posedge \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.clk )
\add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.bin_s1  <= _060_;
always @(posedge \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.clk )
\add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.ain_s1  <= _059_;
always @(posedge \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.clk )
\add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.sum_s1  <= _062_;
always @(posedge \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.clk )
\add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.carry_s1  <= _061_;
assign _060_ = \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.ce  ? \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.b [31:16] : \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.bin_s1 ;
assign _059_ = \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.ce  ? \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.a [31:16] : \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.ain_s1 ;
assign _061_ = \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.ce  ? \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.facout_s1  : \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.carry_s1 ;
assign _062_ = \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.ce  ? \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.fas_s1  : \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.sum_s1 ;
assign _063_ = \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.a  + \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.b ;
assign { \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.cout , \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.s  } = _063_ + \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.cin ;
assign _064_ = \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.a  + \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.b ;
assign { \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.cout , \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.s  } = _064_ + \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.cin ;
always @(posedge \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.clk )
\add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.bin_s1  <= _066_;
always @(posedge \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.clk )
\add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.ain_s1  <= _065_;
always @(posedge \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.clk )
\add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.sum_s1  <= _068_;
always @(posedge \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.clk )
\add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.carry_s1  <= _067_;
assign _066_ = \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.ce  ? \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.b [31:16] : \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.bin_s1 ;
assign _065_ = \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.ce  ? \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.a [31:16] : \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.ain_s1 ;
assign _067_ = \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.ce  ? \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.facout_s1  : \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.carry_s1 ;
assign _068_ = \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.ce  ? \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.fas_s1  : \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.sum_s1 ;
assign _069_ = \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.u1.a  + \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.u1.b ;
assign { \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.u1.cout , \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.u1.s  } = _069_ + \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.u1.cin ;
assign _070_ = \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.u2.a  + \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.u2.b ;
assign { \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.u2.cout , \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.u2.s  } = _070_ + \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.u2.cin ;
always @(posedge \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.clk )
\add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.bin_s1  <= _072_;
always @(posedge \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.clk )
\add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.ain_s1  <= _071_;
always @(posedge \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.clk )
\add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.sum_s1  <= _074_;
always @(posedge \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.clk )
\add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.carry_s1  <= _073_;
assign _072_ = \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.ce  ? \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.b [31:16] : \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.bin_s1 ;
assign _071_ = \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.ce  ? \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.a [31:16] : \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.ain_s1 ;
assign _073_ = \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.ce  ? \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.facout_s1  : \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.carry_s1 ;
assign _074_ = \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.ce  ? \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.fas_s1  : \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.sum_s1 ;
assign _075_ = \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.u1.a  + \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.u1.b ;
assign { \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.u1.cout , \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.u1.s  } = _075_ + \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.u1.cin ;
assign _076_ = \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.u2.a  + \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.u2.b ;
assign { \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.u2.cout , \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.u2.s  } = _076_ + \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.u2.cin ;
always @(posedge \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.clk )
\add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.bin_s1  <= _078_;
always @(posedge \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.clk )
\add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.ain_s1  <= _077_;
always @(posedge \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.clk )
\add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.sum_s1  <= _080_;
always @(posedge \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.clk )
\add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.carry_s1  <= _079_;
assign _078_ = \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.ce  ? \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.b [34:17] : \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.bin_s1 ;
assign _077_ = \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.ce  ? \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.a [34:17] : \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.ain_s1 ;
assign _079_ = \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.ce  ? \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.facout_s1  : \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.carry_s1 ;
assign _080_ = \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.ce  ? \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.fas_s1  : \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.sum_s1 ;
assign _081_ = \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.u1.a  + \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.u1.b ;
assign { \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.u1.cout , \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.u1.s  } = _081_ + \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.u1.cin ;
assign _082_ = \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.u2.a  + \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.u2.b ;
assign { \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.u2.cout , \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.u2.s  } = _082_ + \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.u2.cin ;
always @(posedge \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.clk )
\add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.bin_s1  <= _084_;
always @(posedge \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.clk )
\add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.ain_s1  <= _083_;
always @(posedge \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.clk )
\add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.sum_s1  <= _086_;
always @(posedge \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.clk )
\add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.carry_s1  <= _085_;
assign _084_ = \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.ce  ? \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.b [4:2] : \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.bin_s1 ;
assign _083_ = \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.ce  ? \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.a [4:2] : \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.ain_s1 ;
assign _085_ = \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.ce  ? \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.facout_s1  : \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.carry_s1 ;
assign _086_ = \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.ce  ? \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.fas_s1  : \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.sum_s1 ;
assign _087_ = \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.u1.a  + \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.u1.b ;
assign { \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.u1.cout , \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.u1.s  } = _087_ + \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.u1.cin ;
assign _088_ = \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.u2.a  + \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.u2.b ;
assign { \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.u2.cout , \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.u2.s  } = _088_ + \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.u2.cin ;
always @(posedge \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.clk )
\add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.bin_s1  <= _090_;
always @(posedge \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.clk )
\add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.ain_s1  <= _089_;
always @(posedge \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.clk )
\add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.sum_s1  <= _092_;
always @(posedge \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.clk )
\add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.carry_s1  <= _091_;
assign _090_ = \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.ce  ? \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.b [5:3] : \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.bin_s1 ;
assign _089_ = \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.ce  ? \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.a [5:3] : \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.ain_s1 ;
assign _091_ = \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.ce  ? \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.facout_s1  : \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.carry_s1 ;
assign _092_ = \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.ce  ? \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.fas_s1  : \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.sum_s1 ;
assign _093_ = \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.u1.a  + \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.u1.b ;
assign { \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.u1.cout , \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.u1.s  } = _093_ + \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.u1.cin ;
assign _094_ = \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.u2.a  + \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.u2.b ;
assign { \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.u2.cout , \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.u2.s  } = _094_ + \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.u2.cin ;
always @(posedge \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.clk )
\add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.bin_s1  <= _096_;
always @(posedge \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.clk )
\add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.ain_s1  <= _095_;
always @(posedge \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.clk )
\add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.sum_s1  <= _098_;
always @(posedge \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.clk )
\add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.carry_s1  <= _097_;
assign _096_ = \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.ce  ? \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.b [8:4] : \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.bin_s1 ;
assign _095_ = \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.ce  ? \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.a [8:4] : \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.ain_s1 ;
assign _097_ = \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.ce  ? \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.facout_s1  : \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.carry_s1 ;
assign _098_ = \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.ce  ? \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.fas_s1  : \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.sum_s1 ;
assign _099_ = \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.u1.a  + \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.u1.b ;
assign { \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.u1.cout , \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.u1.s  } = _099_ + \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.u1.cin ;
assign _100_ = \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.u2.a  + \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.u2.b ;
assign { \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.u2.cout , \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.u2.s  } = _100_ + \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.u2.cin ;
assign _101_ = | op_12[1:0];
assign _102_ = | op_10[2:0];
always @(posedge ap_clk)
sext_ln850_reg_445 <= _021_;
always @(posedge ap_clk)
select_ln69_1_reg_499 <= _019_;
always @(posedge ap_clk)
select_ln215_reg_405 <= _018_;
always @(posedge ap_clk)
ret_reg_415 <= _016_;
always @(posedge ap_clk)
ret_V_reg_435 <= _015_;
always @(posedge ap_clk)
tmp_1_reg_440 <= _022_;
always @(posedge ap_clk)
ret_V_2_reg_487 <= _012_;
always @(posedge ap_clk)
ret_V_3_cast_reg_492 <= _013_;
always @(posedge ap_clk)
ret_V_1_reg_457 <= _011_;
always @(posedge ap_clk)
select_ln69_reg_462 <= _020_;
always @(posedge ap_clk)
op_28_V_reg_569 <= _010_;
always @(posedge ap_clk)
select_ln1192_reg_574 <= _017_;
always @(posedge ap_clk)
op_22_V_reg_467 <= _009_;
always @(posedge ap_clk)
icmp_ln851_reg_430 <= _008_;
always @(posedge ap_clk)
icmp_ln851_1_reg_482 <= _007_;
always @(posedge ap_clk)
ret_V_3_reg_524 <= _014_;
always @(posedge ap_clk)
add_ln69_reg_529 <= _005_;
always @(posedge ap_clk)
add_ln69_2_reg_534 <= _003_;
always @(posedge ap_clk)
add_ln69_1_reg_554 <= _002_;
always @(posedge ap_clk)
add_ln69_3_reg_559 <= _004_;
always @(posedge ap_clk)
add_ln691_reg_452 <= _001_;
always @(posedge ap_clk)
add_ln691_1_reg_504 <= _000_;
always @(posedge ap_clk)
ap_CS_fsm <= _006_;
assign _023_ = _027_ ? 2'h2 : 2'h1;
assign _103_ = ap_CS_fsm == 1'h1;
function [20:0] _300_;
input [20:0] a;
input [440:0] b;
input [20:0] s;
case (s)
21'b000000000000000000001:
_300_ = b[20:0];
21'b000000000000000000010:
_300_ = b[41:21];
21'b000000000000000000100:
_300_ = b[62:42];
21'b000000000000000001000:
_300_ = b[83:63];
21'b000000000000000010000:
_300_ = b[104:84];
21'b000000000000000100000:
_300_ = b[125:105];
21'b000000000000001000000:
_300_ = b[146:126];
21'b000000000000010000000:
_300_ = b[167:147];
21'b000000000000100000000:
_300_ = b[188:168];
21'b000000000001000000000:
_300_ = b[209:189];
21'b000000000010000000000:
_300_ = b[230:210];
21'b000000000100000000000:
_300_ = b[251:231];
21'b000000001000000000000:
_300_ = b[272:252];
21'b000000010000000000000:
_300_ = b[293:273];
21'b000000100000000000000:
_300_ = b[314:294];
21'b000001000000000000000:
_300_ = b[335:315];
21'b000010000000000000000:
_300_ = b[356:336];
21'b000100000000000000000:
_300_ = b[377:357];
21'b001000000000000000000:
_300_ = b[398:378];
21'b010000000000000000000:
_300_ = b[419:399];
21'b100000000000000000000:
_300_ = b[440:420];
21'b000000000000000000000:
_300_ = a;
default:
_300_ = 21'bx;
endcase
endfunction
assign ap_NS_fsm = _300_(21'hxxxxxx, { 19'h00000, _023_, 420'h000020000200002000020000200002000020000200002000020000200002000020000200002000020000200002000020000000001 }, { _103_, _123_, _122_, _121_, _120_, _119_, _118_, _117_, _116_, _115_, _114_, _113_, _112_, _111_, _110_, _109_, _108_, _107_, _106_, _105_, _104_ });
assign _104_ = ap_CS_fsm == 21'h100000;
assign _105_ = ap_CS_fsm == 20'h80000;
assign _106_ = ap_CS_fsm == 19'h40000;
assign _107_ = ap_CS_fsm == 18'h20000;
assign _108_ = ap_CS_fsm == 17'h10000;
assign _109_ = ap_CS_fsm == 16'h8000;
assign _110_ = ap_CS_fsm == 15'h4000;
assign _111_ = ap_CS_fsm == 14'h2000;
assign _112_ = ap_CS_fsm == 13'h1000;
assign _113_ = ap_CS_fsm == 12'h800;
assign _114_ = ap_CS_fsm == 11'h400;
assign _115_ = ap_CS_fsm == 10'h200;
assign _116_ = ap_CS_fsm == 9'h100;
assign _117_ = ap_CS_fsm == 8'h80;
assign _118_ = ap_CS_fsm == 7'h40;
assign _119_ = ap_CS_fsm == 6'h20;
assign _120_ = ap_CS_fsm == 5'h10;
assign _121_ = ap_CS_fsm == 4'h8;
assign _122_ = ap_CS_fsm == 3'h4;
assign _123_ = ap_CS_fsm == 2'h2;
assign op_30_ap_vld = ap_CS_fsm[20] ? 1'h1 : 1'h0;
assign ap_idle = _026_ ? 1'h1 : 1'h0;
assign _021_ = ap_CS_fsm[5] ? { tmp_1_reg_440[8], tmp_1_reg_440 } : sext_ln850_reg_445;
assign _019_ = ap_CS_fsm[12] ? select_ln69_1_fu_313_p3 : select_ln69_1_reg_499;
assign _018_ = ap_CS_fsm[0] ? select_ln215_fu_173_p3 : select_ln215_reg_405;
assign _016_ = ap_CS_fsm[2] ? grp_fu_185_p2 : ret_reg_415;
assign _022_ = ap_CS_fsm[4] ? grp_fu_201_p2[11:3] : tmp_1_reg_440;
assign _015_ = ap_CS_fsm[4] ? grp_fu_201_p2 : ret_V_reg_435;
assign _013_ = ap_CS_fsm[11] ? grp_fu_282_p2[33:2] : ret_V_3_cast_reg_492;
assign _012_ = ap_CS_fsm[11] ? grp_fu_282_p2 : ret_V_2_reg_487;
assign _020_ = ap_CS_fsm[7] ? select_ln69_fu_255_p3 : select_ln69_reg_462;
assign _011_ = ap_CS_fsm[7] ? ret_V_1_fu_248_p3 : ret_V_1_reg_457;
assign _017_ = ap_CS_fsm[18] ? select_ln1192_fu_392_p3 : select_ln1192_reg_574;
assign _010_ = ap_CS_fsm[18] ? grp_fu_387_p2 : op_28_V_reg_569;
assign _009_ = ap_CS_fsm[9] ? grp_fu_263_p2 : op_22_V_reg_467;
assign _008_ = ap_CS_fsm[3] ? icmp_ln851_fu_211_p2 : icmp_ln851_reg_430;
assign _007_ = ap_CS_fsm[10] ? icmp_ln851_1_fu_292_p2 : icmp_ln851_1_reg_482;
assign _003_ = ap_CS_fsm[14] ? grp_fu_339_p2 : add_ln69_2_reg_534;
assign _005_ = ap_CS_fsm[14] ? grp_fu_333_p2 : add_ln69_reg_529;
assign _014_ = ap_CS_fsm[14] ? ret_V_3_fu_356_p3 : ret_V_3_reg_524;
assign _004_ = ap_CS_fsm[16] ? grp_fu_378_p2 : add_ln69_3_reg_559;
assign _002_ = ap_CS_fsm[16] ? grp_fu_370_p2 : add_ln69_1_reg_554;
assign _001_ = _025_ ? grp_fu_230_p2 : add_ln691_reg_452;
assign _000_ = _024_ ? grp_fu_308_p2 : add_ln691_1_reg_504;
assign _006_ = ap_rst ? 21'h000001 : ap_NS_fsm;
assign icmp_ln851_1_fu_292_p2 = _101_ ? 1'h1 : 1'h0;
assign icmp_ln851_fu_211_p2 = _102_ ? 1'h1 : 1'h0;
assign ret_V_1_fu_248_p3 = ret_V_reg_435[11] ? select_ln850_fu_243_p3 : sext_ln850_reg_445;
assign ret_V_3_fu_356_p3 = ret_V_2_reg_487[34] ? select_ln850_1_fu_351_p3 : ret_V_3_cast_reg_492;
assign select_ln1192_fu_392_p3 = op_18 ? 32'd4294967295 : 32'd0;
assign select_ln215_fu_173_p3 = op_5[0] ? 9'h1ff : 9'h000;
assign select_ln69_1_fu_313_p3 = op_15 ? 5'h1f : 5'h00;
assign select_ln69_fu_255_p3 = op_11 ? 10'h3ff : 10'h000;
assign select_ln850_1_fu_351_p3 = icmp_ln851_1_reg_482 ? add_ln691_1_reg_504 : ret_V_3_cast_reg_492;
assign select_ln850_fu_243_p3 = icmp_ln851_reg_430 ? add_ln691_reg_452 : sext_ln850_reg_445;
assign ap_CS_fsm_state1 = ap_CS_fsm[0];
assign ap_CS_fsm_state10 = ap_CS_fsm[9];
assign ap_CS_fsm_state11 = ap_CS_fsm[10];
assign ap_CS_fsm_state12 = ap_CS_fsm[11];
assign ap_CS_fsm_state13 = ap_CS_fsm[12];
assign ap_CS_fsm_state14 = ap_CS_fsm[13];
assign ap_CS_fsm_state15 = ap_CS_fsm[14];
assign ap_CS_fsm_state16 = ap_CS_fsm[15];
assign ap_CS_fsm_state17 = ap_CS_fsm[16];
assign ap_CS_fsm_state18 = ap_CS_fsm[17];
assign ap_CS_fsm_state19 = ap_CS_fsm[18];
assign ap_CS_fsm_state2 = ap_CS_fsm[1];
assign ap_CS_fsm_state20 = ap_CS_fsm[19];
assign ap_CS_fsm_state21 = ap_CS_fsm[20];
assign ap_CS_fsm_state3 = ap_CS_fsm[2];
assign ap_CS_fsm_state4 = ap_CS_fsm[3];
assign ap_CS_fsm_state5 = ap_CS_fsm[4];
assign ap_CS_fsm_state6 = ap_CS_fsm[5];
assign ap_CS_fsm_state7 = ap_CS_fsm[6];
assign ap_CS_fsm_state8 = ap_CS_fsm[7];
assign ap_CS_fsm_state9 = ap_CS_fsm[8];
assign ap_done = op_30_ap_vld;
assign ap_ready = op_30_ap_vld;
assign grp_fu_185_p0 = { op_6[7], op_6 };
assign grp_fu_201_p0 = { ret_reg_415, 3'h0 };
assign grp_fu_201_p1 = { op_10[3], op_10[3], op_10[3], op_10[3], op_10[3], op_10[3], op_10[3], op_10[3], op_10 };
assign grp_fu_230_p0 = { tmp_1_reg_440[8], tmp_1_reg_440 };
assign grp_fu_282_p0 = { op_22_V_reg_467[9], op_22_V_reg_467[9], op_22_V_reg_467[9], op_22_V_reg_467[9], op_22_V_reg_467[9], op_22_V_reg_467[9], op_22_V_reg_467[9], op_22_V_reg_467[9], op_22_V_reg_467[9], op_22_V_reg_467[9], op_22_V_reg_467[9], op_22_V_reg_467[9], op_22_V_reg_467[9], op_22_V_reg_467[9], op_22_V_reg_467[9], op_22_V_reg_467[9], op_22_V_reg_467[9], op_22_V_reg_467[9], op_22_V_reg_467[9], op_22_V_reg_467[9], op_22_V_reg_467[9], op_22_V_reg_467[9], op_22_V_reg_467[9], op_22_V_reg_467, 2'h0 };
assign grp_fu_282_p1 = { op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12 };
assign grp_fu_333_p0 = { op_16[15], op_16 };
assign grp_fu_333_p1 = { op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13 };
assign grp_fu_339_p0 = { 1'h0, op_14 };
assign grp_fu_370_p0 = { add_ln69_reg_529[16], add_ln69_reg_529[16], add_ln69_reg_529[16], add_ln69_reg_529[16], add_ln69_reg_529[16], add_ln69_reg_529[16], add_ln69_reg_529[16], add_ln69_reg_529[16], add_ln69_reg_529[16], add_ln69_reg_529[16], add_ln69_reg_529[16], add_ln69_reg_529[16], add_ln69_reg_529[16], add_ln69_reg_529[16], add_ln69_reg_529[16], add_ln69_reg_529 };
assign grp_fu_378_p0 = { add_ln69_2_reg_534[4], add_ln69_2_reg_534 };
assign grp_fu_378_p1 = { op_17[3], op_17[3], op_17 };
assign grp_fu_387_p0 = { add_ln69_3_reg_559[5], add_ln69_3_reg_559[5], add_ln69_3_reg_559[5], add_ln69_3_reg_559[5], add_ln69_3_reg_559[5], add_ln69_3_reg_559[5], add_ln69_3_reg_559[5], add_ln69_3_reg_559[5], add_ln69_3_reg_559[5], add_ln69_3_reg_559[5], add_ln69_3_reg_559[5], add_ln69_3_reg_559[5], add_ln69_3_reg_559[5], add_ln69_3_reg_559[5], add_ln69_3_reg_559[5], add_ln69_3_reg_559[5], add_ln69_3_reg_559[5], add_ln69_3_reg_559[5], add_ln69_3_reg_559[5], add_ln69_3_reg_559[5], add_ln69_3_reg_559[5], add_ln69_3_reg_559[5], add_ln69_3_reg_559[5], add_ln69_3_reg_559[5], add_ln69_3_reg_559[5], add_ln69_3_reg_559[5], add_ln69_3_reg_559 };
assign op_30 = grp_fu_400_p2;
assign op_8_V_fu_169_p1 = op_5[0];
assign p_Result_1_fu_344_p3 = ret_V_2_reg_487[34];
assign p_Result_s_fu_236_p3 = ret_V_reg_435[11];
assign sext_ln1192_fu_190_p0 = op_10;
assign sext_ln703_fu_267_p0 = op_12;
assign sext_ln850_fu_227_p1 = { tmp_1_reg_440[8], tmp_1_reg_440 };
assign tmp_fu_271_p3 = { op_22_V_reg_467, 2'h0 };
assign trunc_ln851_1_fu_288_p0 = op_12;
assign trunc_ln851_1_fu_288_p1 = op_12[1:0];
assign trunc_ln851_fu_207_p0 = op_10;
assign trunc_ln851_fu_207_p1 = op_10[2:0];
assign \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.ain_s0  = \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.a ;
assign \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.bin_s0  = \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.b ;
assign \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.s  = { \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.fas_s2 , \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.sum_s1  };
assign \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.u2.a  = \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.ain_s1 ;
assign \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.u2.b  = \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.bin_s1 ;
assign \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.u2.cin  = \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.carry_s1 ;
assign \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.facout_s2  = \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.u2.cout ;
assign \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.fas_s2  = \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.u2.s ;
assign \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.u1.a  = \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.a [3:0];
assign \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.u1.b  = \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.b [3:0];
assign \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.u1.cin  = 1'h0;
assign \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.facout_s1  = \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.u1.cout ;
assign \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.fas_s1  = \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.u1.s ;
assign \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.a  = \add_9s_9ns_9_2_1_U1.din0 ;
assign \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.b  = \add_9s_9ns_9_2_1_U1.din1 ;
assign \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.ce  = \add_9s_9ns_9_2_1_U1.ce ;
assign \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.clk  = \add_9s_9ns_9_2_1_U1.clk ;
assign \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.reset  = \add_9s_9ns_9_2_1_U1.reset ;
assign \add_9s_9ns_9_2_1_U1.dout  = \add_9s_9ns_9_2_1_U1.top_add_9s_9ns_9_2_1_Adder_0_U.s ;
assign \add_9s_9ns_9_2_1_U1.ce  = 1'h1;
assign \add_9s_9ns_9_2_1_U1.clk  = ap_clk;
assign \add_9s_9ns_9_2_1_U1.din0  = { op_6[7], op_6 };
assign \add_9s_9ns_9_2_1_U1.din1  = select_ln215_reg_405;
assign grp_fu_185_p2 = \add_9s_9ns_9_2_1_U1.dout ;
assign \add_9s_9ns_9_2_1_U1.reset  = ap_rst;
assign \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.ain_s0  = \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.a ;
assign \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.bin_s0  = \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.b ;
assign \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.s  = { \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.fas_s2 , \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.sum_s1  };
assign \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.u2.a  = \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.ain_s1 ;
assign \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.u2.b  = \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.bin_s1 ;
assign \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.u2.cin  = \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.carry_s1 ;
assign \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.facout_s2  = \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.u2.cout ;
assign \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.fas_s2  = \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.u2.s ;
assign \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.u1.a  = \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.a [2:0];
assign \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.u1.b  = \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.b [2:0];
assign \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.u1.cin  = 1'h0;
assign \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.facout_s1  = \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.u1.cout ;
assign \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.fas_s1  = \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.u1.s ;
assign \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.a  = \add_6s_6s_6_2_1_U10.din0 ;
assign \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.b  = \add_6s_6s_6_2_1_U10.din1 ;
assign \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.ce  = \add_6s_6s_6_2_1_U10.ce ;
assign \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.clk  = \add_6s_6s_6_2_1_U10.clk ;
assign \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.reset  = \add_6s_6s_6_2_1_U10.reset ;
assign \add_6s_6s_6_2_1_U10.dout  = \add_6s_6s_6_2_1_U10.top_add_6s_6s_6_2_1_Adder_9_U.s ;
assign \add_6s_6s_6_2_1_U10.ce  = 1'h1;
assign \add_6s_6s_6_2_1_U10.clk  = ap_clk;
assign \add_6s_6s_6_2_1_U10.din0  = { add_ln69_2_reg_534[4], add_ln69_2_reg_534 };
assign \add_6s_6s_6_2_1_U10.din1  = { op_17[3], op_17[3], op_17 };
assign grp_fu_378_p2 = \add_6s_6s_6_2_1_U10.dout ;
assign \add_6s_6s_6_2_1_U10.reset  = ap_rst;
assign \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.ain_s0  = \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.a ;
assign \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.bin_s0  = \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.b ;
assign \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.s  = { \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.fas_s2 , \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.sum_s1  };
assign \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.u2.a  = \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.ain_s1 ;
assign \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.u2.b  = \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.bin_s1 ;
assign \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.u2.cin  = \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.carry_s1 ;
assign \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.facout_s2  = \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.u2.cout ;
assign \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.fas_s2  = \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.u2.s ;
assign \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.u1.a  = \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.a [1:0];
assign \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.u1.b  = \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.b [1:0];
assign \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.u1.cin  = 1'h0;
assign \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.facout_s1  = \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.u1.cout ;
assign \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.fas_s1  = \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.u1.s ;
assign \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.a  = \add_5ns_5ns_5_2_1_U8.din0 ;
assign \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.b  = \add_5ns_5ns_5_2_1_U8.din1 ;
assign \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.ce  = \add_5ns_5ns_5_2_1_U8.ce ;
assign \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.clk  = \add_5ns_5ns_5_2_1_U8.clk ;
assign \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.reset  = \add_5ns_5ns_5_2_1_U8.reset ;
assign \add_5ns_5ns_5_2_1_U8.dout  = \add_5ns_5ns_5_2_1_U8.top_add_5ns_5ns_5_2_1_Adder_7_U.s ;
assign \add_5ns_5ns_5_2_1_U8.ce  = 1'h1;
assign \add_5ns_5ns_5_2_1_U8.clk  = ap_clk;
assign \add_5ns_5ns_5_2_1_U8.din0  = { 1'h0, op_14 };
assign \add_5ns_5ns_5_2_1_U8.din1  = select_ln69_1_reg_499;
assign grp_fu_339_p2 = \add_5ns_5ns_5_2_1_U8.dout ;
assign \add_5ns_5ns_5_2_1_U8.reset  = ap_rst;
assign \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.ain_s0  = \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.a ;
assign \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.bin_s0  = \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.b ;
assign \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.s  = { \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.fas_s2 , \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.sum_s1  };
assign \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.u2.a  = \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.ain_s1 ;
assign \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.u2.b  = \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.bin_s1 ;
assign \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.u2.cin  = \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.carry_s1 ;
assign \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.facout_s2  = \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.u2.cout ;
assign \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.fas_s2  = \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.u2.s ;
assign \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.u1.a  = \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.a [16:0];
assign \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.u1.b  = \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.b [16:0];
assign \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.u1.cin  = 1'h0;
assign \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.facout_s1  = \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.u1.cout ;
assign \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.fas_s1  = \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.u1.s ;
assign \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.a  = \add_35s_35s_35_2_1_U5.din0 ;
assign \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.b  = \add_35s_35s_35_2_1_U5.din1 ;
assign \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.ce  = \add_35s_35s_35_2_1_U5.ce ;
assign \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.clk  = \add_35s_35s_35_2_1_U5.clk ;
assign \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.reset  = \add_35s_35s_35_2_1_U5.reset ;
assign \add_35s_35s_35_2_1_U5.dout  = \add_35s_35s_35_2_1_U5.top_add_35s_35s_35_2_1_Adder_4_U.s ;
assign \add_35s_35s_35_2_1_U5.ce  = 1'h1;
assign \add_35s_35s_35_2_1_U5.clk  = ap_clk;
assign \add_35s_35s_35_2_1_U5.din0  = { op_22_V_reg_467[9], op_22_V_reg_467[9], op_22_V_reg_467[9], op_22_V_reg_467[9], op_22_V_reg_467[9], op_22_V_reg_467[9], op_22_V_reg_467[9], op_22_V_reg_467[9], op_22_V_reg_467[9], op_22_V_reg_467[9], op_22_V_reg_467[9], op_22_V_reg_467[9], op_22_V_reg_467[9], op_22_V_reg_467[9], op_22_V_reg_467[9], op_22_V_reg_467[9], op_22_V_reg_467[9], op_22_V_reg_467[9], op_22_V_reg_467[9], op_22_V_reg_467[9], op_22_V_reg_467[9], op_22_V_reg_467[9], op_22_V_reg_467[9], op_22_V_reg_467, 2'h0 };
assign \add_35s_35s_35_2_1_U5.din1  = { op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12[3], op_12 };
assign grp_fu_282_p2 = \add_35s_35s_35_2_1_U5.dout ;
assign \add_35s_35s_35_2_1_U5.reset  = ap_rst;
assign \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.ain_s0  = \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.a ;
assign \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.bin_s0  = \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.b ;
assign \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.s  = { \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.fas_s2 , \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.sum_s1  };
assign \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.u2.a  = \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.ain_s1 ;
assign \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.u2.b  = \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.bin_s1 ;
assign \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.u2.cin  = \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.carry_s1 ;
assign \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.facout_s2  = \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.u2.cout ;
assign \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.fas_s2  = \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.u2.s ;
assign \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.u1.a  = \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.a [15:0];
assign \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.u1.b  = \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.b [15:0];
assign \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.u1.cin  = 1'h0;
assign \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.facout_s1  = \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.u1.cout ;
assign \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.fas_s1  = \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.u1.s ;
assign \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.a  = \add_32s_32ns_32_2_1_U9.din0 ;
assign \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.b  = \add_32s_32ns_32_2_1_U9.din1 ;
assign \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.ce  = \add_32s_32ns_32_2_1_U9.ce ;
assign \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.clk  = \add_32s_32ns_32_2_1_U9.clk ;
assign \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.reset  = \add_32s_32ns_32_2_1_U9.reset ;
assign \add_32s_32ns_32_2_1_U9.dout  = \add_32s_32ns_32_2_1_U9.top_add_32s_32ns_32_2_1_Adder_8_U.s ;
assign \add_32s_32ns_32_2_1_U9.ce  = 1'h1;
assign \add_32s_32ns_32_2_1_U9.clk  = ap_clk;
assign \add_32s_32ns_32_2_1_U9.din0  = { add_ln69_reg_529[16], add_ln69_reg_529[16], add_ln69_reg_529[16], add_ln69_reg_529[16], add_ln69_reg_529[16], add_ln69_reg_529[16], add_ln69_reg_529[16], add_ln69_reg_529[16], add_ln69_reg_529[16], add_ln69_reg_529[16], add_ln69_reg_529[16], add_ln69_reg_529[16], add_ln69_reg_529[16], add_ln69_reg_529[16], add_ln69_reg_529[16], add_ln69_reg_529 };
assign \add_32s_32ns_32_2_1_U9.din1  = ret_V_3_reg_524;
assign grp_fu_370_p2 = \add_32s_32ns_32_2_1_U9.dout ;
assign \add_32s_32ns_32_2_1_U9.reset  = ap_rst;
assign \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.ain_s0  = \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.a ;
assign \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.bin_s0  = \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.b ;
assign \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.s  = { \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.fas_s2 , \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.sum_s1  };
assign \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.u2.a  = \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.ain_s1 ;
assign \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.u2.b  = \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.bin_s1 ;
assign \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.u2.cin  = \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.carry_s1 ;
assign \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.facout_s2  = \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.u2.cout ;
assign \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.fas_s2  = \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.u2.s ;
assign \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.u1.a  = \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.a [15:0];
assign \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.u1.b  = \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.b [15:0];
assign \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.u1.cin  = 1'h0;
assign \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.facout_s1  = \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.u1.cout ;
assign \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.fas_s1  = \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.u1.s ;
assign \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.a  = \add_32s_32ns_32_2_1_U11.din0 ;
assign \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.b  = \add_32s_32ns_32_2_1_U11.din1 ;
assign \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.ce  = \add_32s_32ns_32_2_1_U11.ce ;
assign \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.clk  = \add_32s_32ns_32_2_1_U11.clk ;
assign \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.reset  = \add_32s_32ns_32_2_1_U11.reset ;
assign \add_32s_32ns_32_2_1_U11.dout  = \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_8_U.s ;
assign \add_32s_32ns_32_2_1_U11.ce  = 1'h1;
assign \add_32s_32ns_32_2_1_U11.clk  = ap_clk;
assign \add_32s_32ns_32_2_1_U11.din0  = { add_ln69_3_reg_559[5], add_ln69_3_reg_559[5], add_ln69_3_reg_559[5], add_ln69_3_reg_559[5], add_ln69_3_reg_559[5], add_ln69_3_reg_559[5], add_ln69_3_reg_559[5], add_ln69_3_reg_559[5], add_ln69_3_reg_559[5], add_ln69_3_reg_559[5], add_ln69_3_reg_559[5], add_ln69_3_reg_559[5], add_ln69_3_reg_559[5], add_ln69_3_reg_559[5], add_ln69_3_reg_559[5], add_ln69_3_reg_559[5], add_ln69_3_reg_559[5], add_ln69_3_reg_559[5], add_ln69_3_reg_559[5], add_ln69_3_reg_559[5], add_ln69_3_reg_559[5], add_ln69_3_reg_559[5], add_ln69_3_reg_559[5], add_ln69_3_reg_559[5], add_ln69_3_reg_559[5], add_ln69_3_reg_559[5], add_ln69_3_reg_559 };
assign \add_32s_32ns_32_2_1_U11.din1  = add_ln69_1_reg_554;
assign grp_fu_387_p2 = \add_32s_32ns_32_2_1_U11.dout ;
assign \add_32s_32ns_32_2_1_U11.reset  = ap_rst;
assign \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.ain_s0  = \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.a ;
assign \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.bin_s0  = \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.b ;
assign \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.s  = { \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.fas_s2 , \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.sum_s1  };
assign \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.a  = \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.ain_s1 ;
assign \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.b  = \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.bin_s1 ;
assign \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.cin  = \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.carry_s1 ;
assign \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.facout_s2  = \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.cout ;
assign \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.fas_s2  = \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.s ;
assign \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.a  = \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.a [15:0];
assign \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.b  = \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.b [15:0];
assign \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.cin  = 1'h0;
assign \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.facout_s1  = \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.cout ;
assign \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.fas_s1  = \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.s ;
assign \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.a  = \add_32ns_32ns_32_2_1_U6.din0 ;
assign \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.b  = \add_32ns_32ns_32_2_1_U6.din1 ;
assign \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.ce  = \add_32ns_32ns_32_2_1_U6.ce ;
assign \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.clk  = \add_32ns_32ns_32_2_1_U6.clk ;
assign \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.reset  = \add_32ns_32ns_32_2_1_U6.reset ;
assign \add_32ns_32ns_32_2_1_U6.dout  = \add_32ns_32ns_32_2_1_U6.top_add_32ns_32ns_32_2_1_Adder_5_U.s ;
assign \add_32ns_32ns_32_2_1_U6.ce  = 1'h1;
assign \add_32ns_32ns_32_2_1_U6.clk  = ap_clk;
assign \add_32ns_32ns_32_2_1_U6.din0  = ret_V_3_cast_reg_492;
assign \add_32ns_32ns_32_2_1_U6.din1  = 32'd1;
assign grp_fu_308_p2 = \add_32ns_32ns_32_2_1_U6.dout ;
assign \add_32ns_32ns_32_2_1_U6.reset  = ap_rst;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.ain_s0  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.a ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.bin_s0  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.b ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.s  = { \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.fas_s2 , \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.sum_s1  };
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.a  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.ain_s1 ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.b  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.bin_s1 ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.cin  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.carry_s1 ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.facout_s2  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.cout ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.fas_s2  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.u2.s ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.a  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.a [15:0];
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.b  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.b [15:0];
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.cin  = 1'h0;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.facout_s1  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.cout ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.fas_s1  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.u1.s ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.a  = \add_32ns_32ns_32_2_1_U12.din0 ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.b  = \add_32ns_32ns_32_2_1_U12.din1 ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.ce  = \add_32ns_32ns_32_2_1_U12.ce ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.clk  = \add_32ns_32ns_32_2_1_U12.clk ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.reset  = \add_32ns_32ns_32_2_1_U12.reset ;
assign \add_32ns_32ns_32_2_1_U12.dout  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_5_U.s ;
assign \add_32ns_32ns_32_2_1_U12.ce  = 1'h1;
assign \add_32ns_32ns_32_2_1_U12.clk  = ap_clk;
assign \add_32ns_32ns_32_2_1_U12.din0  = op_28_V_reg_569;
assign \add_32ns_32ns_32_2_1_U12.din1  = select_ln1192_reg_574;
assign grp_fu_400_p2 = \add_32ns_32ns_32_2_1_U12.dout ;
assign \add_32ns_32ns_32_2_1_U12.reset  = ap_rst;
assign \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.ain_s0  = \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.a ;
assign \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.bin_s0  = \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.b ;
assign \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.s  = { \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.fas_s2 , \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.sum_s1  };
assign \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.u2.a  = \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.ain_s1 ;
assign \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.u2.b  = \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.bin_s1 ;
assign \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.u2.cin  = \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.carry_s1 ;
assign \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.facout_s2  = \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.u2.cout ;
assign \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.fas_s2  = \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.u2.s ;
assign \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.u1.a  = \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.a [7:0];
assign \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.u1.b  = \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.b [7:0];
assign \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.u1.cin  = 1'h0;
assign \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.facout_s1  = \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.u1.cout ;
assign \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.fas_s1  = \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.u1.s ;
assign \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.a  = \add_17s_17s_17_2_1_U7.din0 ;
assign \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.b  = \add_17s_17s_17_2_1_U7.din1 ;
assign \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.ce  = \add_17s_17s_17_2_1_U7.ce ;
assign \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.clk  = \add_17s_17s_17_2_1_U7.clk ;
assign \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.reset  = \add_17s_17s_17_2_1_U7.reset ;
assign \add_17s_17s_17_2_1_U7.dout  = \add_17s_17s_17_2_1_U7.top_add_17s_17s_17_2_1_Adder_6_U.s ;
assign \add_17s_17s_17_2_1_U7.ce  = 1'h1;
assign \add_17s_17s_17_2_1_U7.clk  = ap_clk;
assign \add_17s_17s_17_2_1_U7.din0  = { op_16[15], op_16 };
assign \add_17s_17s_17_2_1_U7.din1  = { op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13[7], op_13 };
assign grp_fu_333_p2 = \add_17s_17s_17_2_1_U7.dout ;
assign \add_17s_17s_17_2_1_U7.reset  = ap_rst;
assign \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.ain_s0  = \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.a ;
assign \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.bin_s0  = \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.b ;
assign \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.s  = { \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.fas_s2 , \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.sum_s1  };
assign \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.u2.a  = \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.ain_s1 ;
assign \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.u2.b  = \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.bin_s1 ;
assign \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.u2.cin  = \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.carry_s1 ;
assign \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.facout_s2  = \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.u2.cout ;
assign \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.fas_s2  = \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.u2.s ;
assign \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.u1.a  = \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.a [5:0];
assign \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.u1.b  = \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.b [5:0];
assign \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.u1.cin  = 1'h0;
assign \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.facout_s1  = \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.u1.cout ;
assign \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.fas_s1  = \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.u1.s ;
assign \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.a  = \add_12ns_12s_12_2_1_U2.din0 ;
assign \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.b  = \add_12ns_12s_12_2_1_U2.din1 ;
assign \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.ce  = \add_12ns_12s_12_2_1_U2.ce ;
assign \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.clk  = \add_12ns_12s_12_2_1_U2.clk ;
assign \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.reset  = \add_12ns_12s_12_2_1_U2.reset ;
assign \add_12ns_12s_12_2_1_U2.dout  = \add_12ns_12s_12_2_1_U2.top_add_12ns_12s_12_2_1_Adder_1_U.s ;
assign \add_12ns_12s_12_2_1_U2.ce  = 1'h1;
assign \add_12ns_12s_12_2_1_U2.clk  = ap_clk;
assign \add_12ns_12s_12_2_1_U2.din0  = { ret_reg_415, 3'h0 };
assign \add_12ns_12s_12_2_1_U2.din1  = { op_10[3], op_10[3], op_10[3], op_10[3], op_10[3], op_10[3], op_10[3], op_10[3], op_10 };
assign grp_fu_201_p2 = \add_12ns_12s_12_2_1_U2.dout ;
assign \add_12ns_12s_12_2_1_U2.reset  = ap_rst;
assign \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.ain_s0  = \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.a ;
assign \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.bin_s0  = \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.b ;
assign \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.s  = { \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.fas_s2 , \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.sum_s1  };
assign \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.u2.a  = \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.ain_s1 ;
assign \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.u2.b  = \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.bin_s1 ;
assign \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.u2.cin  = \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.carry_s1 ;
assign \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.facout_s2  = \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.u2.cout ;
assign \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.fas_s2  = \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.u2.s ;
assign \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.u1.a  = \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.a [4:0];
assign \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.u1.b  = \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.b [4:0];
assign \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.u1.cin  = 1'h0;
assign \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.facout_s1  = \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.u1.cout ;
assign \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.fas_s1  = \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.u1.s ;
assign \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.a  = \add_10s_10ns_10_2_1_U3.din0 ;
assign \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.b  = \add_10s_10ns_10_2_1_U3.din1 ;
assign \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.ce  = \add_10s_10ns_10_2_1_U3.ce ;
assign \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.clk  = \add_10s_10ns_10_2_1_U3.clk ;
assign \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.reset  = \add_10s_10ns_10_2_1_U3.reset ;
assign \add_10s_10ns_10_2_1_U3.dout  = \add_10s_10ns_10_2_1_U3.top_add_10s_10ns_10_2_1_Adder_2_U.s ;
assign \add_10s_10ns_10_2_1_U3.ce  = 1'h1;
assign \add_10s_10ns_10_2_1_U3.clk  = ap_clk;
assign \add_10s_10ns_10_2_1_U3.din0  = { tmp_1_reg_440[8], tmp_1_reg_440 };
assign \add_10s_10ns_10_2_1_U3.din1  = 10'h001;
assign grp_fu_230_p2 = \add_10s_10ns_10_2_1_U3.dout ;
assign \add_10s_10ns_10_2_1_U3.reset  = ap_rst;
assign \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.ain_s0  = \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.a ;
assign \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.bin_s0  = \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.b ;
assign \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.s  = { \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.fas_s2 , \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.sum_s1  };
assign \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.u2.a  = \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.ain_s1 ;
assign \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.u2.b  = \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.bin_s1 ;
assign \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.u2.cin  = \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.carry_s1 ;
assign \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.facout_s2  = \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.u2.cout ;
assign \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.fas_s2  = \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.u2.s ;
assign \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.u1.a  = \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.a [4:0];
assign \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.u1.b  = \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.b [4:0];
assign \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.u1.cin  = 1'h0;
assign \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.facout_s1  = \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.u1.cout ;
assign \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.fas_s1  = \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.u1.s ;
assign \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.a  = \add_10ns_10ns_10_2_1_U4.din0 ;
assign \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.b  = \add_10ns_10ns_10_2_1_U4.din1 ;
assign \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.ce  = \add_10ns_10ns_10_2_1_U4.ce ;
assign \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.clk  = \add_10ns_10ns_10_2_1_U4.clk ;
assign \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.reset  = \add_10ns_10ns_10_2_1_U4.reset ;
assign \add_10ns_10ns_10_2_1_U4.dout  = \add_10ns_10ns_10_2_1_U4.top_add_10ns_10ns_10_2_1_Adder_3_U.s ;
assign \add_10ns_10ns_10_2_1_U4.ce  = 1'h1;
assign \add_10ns_10ns_10_2_1_U4.clk  = ap_clk;
assign \add_10ns_10ns_10_2_1_U4.din0  = ret_V_1_reg_457;
assign \add_10ns_10ns_10_2_1_U4.din1  = select_ln69_reg_462;
assign grp_fu_263_p2 = \add_10ns_10ns_10_2_1_U4.dout ;
assign \add_10ns_10ns_10_2_1_U4.reset  = ap_rst;
endmodule


// Product machine:
module top_A_times_top_B (ap_start, op_0, op_1, op_10, op_11, op_12, op_13, op_14, op_15, op_16, op_17, op_18, op_5, op_6, ap_clk, unsafe_signal);
input ap_start;
input [1:0] op_0;
input [3:0] op_1;
input [3:0] op_10;
input op_11;
input [3:0] op_12;
input [7:0] op_13;
input [3:0] op_14;
input op_15;
input [15:0] op_16;
input [3:0] op_17;
input op_18;
input [3:0] op_5;
input [7:0] op_6;
input ap_clk;
output unsafe_signal;
reg _setup;
initial _setup = 1'b0;
always @ (posedge ap_clk) _setup <= 1'b1;
reg ap_start_internal;
always @ (posedge ap_clk) if (!_setup) ap_start_internal <= ap_start;
reg [1:0] op_0_internal;
always @ (posedge ap_clk) if (!_setup) op_0_internal <= op_0;
reg [3:0] op_1_internal;
always @ (posedge ap_clk) if (!_setup) op_1_internal <= op_1;
reg [3:0] op_10_internal;
always @ (posedge ap_clk) if (!_setup) op_10_internal <= op_10;
reg op_11_internal;
always @ (posedge ap_clk) if (!_setup) op_11_internal <= op_11;
reg [3:0] op_12_internal;
always @ (posedge ap_clk) if (!_setup) op_12_internal <= op_12;
reg [7:0] op_13_internal;
always @ (posedge ap_clk) if (!_setup) op_13_internal <= op_13;
reg [3:0] op_14_internal;
always @ (posedge ap_clk) if (!_setup) op_14_internal <= op_14;
reg op_15_internal;
always @ (posedge ap_clk) if (!_setup) op_15_internal <= op_15;
reg [15:0] op_16_internal;
always @ (posedge ap_clk) if (!_setup) op_16_internal <= op_16;
reg [3:0] op_17_internal;
always @ (posedge ap_clk) if (!_setup) op_17_internal <= op_17;
reg op_18_internal;
always @ (posedge ap_clk) if (!_setup) op_18_internal <= op_18;
reg [3:0] op_5_internal;
always @ (posedge ap_clk) if (!_setup) op_5_internal <= op_5;
reg [7:0] op_6_internal;
always @ (posedge ap_clk) if (!_setup) op_6_internal <= op_6;
wire ap_done_A;
wire ap_done_B;
wire ap_done_eq;
assign ap_done_eq = ap_done_A == ap_done_B;
wire ap_idle_A;
wire ap_idle_B;
wire ap_idle_eq;
assign ap_idle_eq = ap_idle_A == ap_idle_B;
wire ap_ready_A;
wire ap_ready_B;
wire ap_ready_eq;
assign ap_ready_eq = ap_ready_A == ap_ready_B;
wire [31:0] op_30_A;
wire [31:0] op_30_B;
wire op_30_eq;
assign op_30_eq = op_30_A == op_30_B;
wire op_30_ap_vld_A;
wire op_30_ap_vld_B;
wire clk_enable_A;
wire clk_enable_B;
assign clk_enable_A = _setup & (~op_30_ap_vld_A | op_30_ap_vld_B);
assign clk_enable_B = _setup;
wire divergent;
assign divergent = ~(ap_done_eq & ap_idle_eq & ap_ready_eq & op_30_eq);
assign unsafe_signal = op_30_ap_vld_A & op_30_ap_vld_B & divergent;
top_A instance_A (
    .ap_clk(ap_clk),
    .clk_enable(clk_enable_A),
    .ap_start(ap_start_internal),
    .op_0(op_0_internal),
    .op_1(op_1_internal),
    .op_10(op_10_internal),
    .op_11(op_11_internal),
    .op_12(op_12_internal),
    .op_13(op_13_internal),
    .op_14(op_14_internal),
    .op_15(op_15_internal),
    .op_16(op_16_internal),
    .op_17(op_17_internal),
    .op_18(op_18_internal),
    .op_5(op_5_internal),
    .op_6(op_6_internal),
    .ap_done(ap_done_A),
    .ap_idle(ap_idle_A),
    .ap_ready(ap_ready_A),
    .op_30(op_30_A),
    .op_30_ap_vld(op_30_ap_vld_A)
);
top_B instance_B (
    .ap_clk(ap_clk),
    .clk_enable(clk_enable_B),
    .ap_start(ap_start_internal),
    .op_0(op_0_internal),
    .op_1(op_1_internal),
    .op_10(op_10_internal),
    .op_11(op_11_internal),
    .op_12(op_12_internal),
    .op_13(op_13_internal),
    .op_14(op_14_internal),
    .op_15(op_15_internal),
    .op_16(op_16_internal),
    .op_17(op_17_internal),
    .op_18(op_18_internal),
    .op_5(op_5_internal),
    .op_6(op_6_internal),
    .ap_done(ap_done_B),
    .ap_idle(ap_idle_B),
    .ap_ready(ap_ready_B),
    .op_30(op_30_B),
    .op_30_ap_vld(op_30_ap_vld_B)
);
endmodule
