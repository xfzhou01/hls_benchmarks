// Processed by function `construct_kairos` in `verilog_tricks.py`.
// Machine A:
// Processed by function `add_clk_enable_signal` in `verilog_tricks.py`.
// Processed by function `remove_reset_signal` in `verilog_tricks.py`.
module top_A (
  ap_clk,
  ap_start,
  ap_done,
  ap_idle,
  ap_ready,
  op_0,
  op_1,
  op_2,
  op_3,
  op_7,
  op_8,
  op_10,
  op_12,
  op_13,
  op_14,
  op_28,
  op_28_ap_vld,
clk_enable
);
input clk_enable;


input ap_clk;
wire ap_rst;
assign ap_rst = op_28_ap_vld;
input ap_start;
input [1:0] op_0;
input [3:0] op_1;
input [3:0] op_10;
input [1:0] op_12;
input [3:0] op_13;
input [7:0] op_14;
input [7:0] op_2;
input [15:0] op_3;
input [1:0] op_7;
input [1:0] op_8;
output ap_done;
output ap_idle;
output ap_ready;
output [31:0] op_28;
output op_28_ap_vld;


reg Range1_all_ones_reg_1030;
reg Range1_all_zeros_reg_1037;
reg Range2_all_ones_reg_1025;
reg [4:0] \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.ain_s1 ;
reg [4:0] \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.bin_s1 ;
reg \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.carry_s1 ;
reg [4:0] \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.sum_s1 ;
reg [7:0] \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.ain_s1 ;
reg [7:0] \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.bin_s1 ;
reg \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.carry_s1 ;
reg [6:0] \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.sum_s1 ;
reg [8:0] \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.ain_s1 ;
reg [8:0] \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.bin_s1 ;
reg \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.carry_s1 ;
reg [7:0] \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.sum_s1 ;
reg \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.ain_s1 ;
reg \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.bin_s1 ;
reg \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.carry_s1 ;
reg \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.sum_s1 ;
reg \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.ain_s1 ;
reg \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.bin_s1 ;
reg \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.carry_s1 ;
reg \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.sum_s1 ;
reg \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.ain_s1 ;
reg \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.bin_s1 ;
reg \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.carry_s1 ;
reg \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.sum_s1 ;
reg [1:0] \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.ain_s1 ;
reg [1:0] \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.bin_s1 ;
reg \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.carry_s1 ;
reg \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.sum_s1 ;
reg [1:0] \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.ain_s1 ;
reg [1:0] \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.bin_s1 ;
reg \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.carry_s1 ;
reg \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.sum_s1 ;
reg [1:0] \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.ain_s1 ;
reg [1:0] \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.bin_s1 ;
reg \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.carry_s1 ;
reg [1:0] \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.sum_s1 ;
reg [2:0] \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.ain_s1 ;
reg [2:0] \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.bin_s1 ;
reg \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.carry_s1 ;
reg [1:0] \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.sum_s1 ;
reg [2:0] \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.ain_s1 ;
reg [2:0] \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.bin_s1 ;
reg \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.carry_s1 ;
reg [2:0] \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.sum_s1 ;
reg [2:0] \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.ain_s1 ;
reg [2:0] \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.bin_s1 ;
reg \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.carry_s1 ;
reg [2:0] \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.sum_s1 ;
reg [2:0] \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.ain_s1 ;
reg [2:0] \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.bin_s1 ;
reg \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.carry_s1 ;
reg [2:0] \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.sum_s1 ;
reg [2:0] \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.ain_s1 ;
reg [2:0] \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.bin_s1 ;
reg \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.carry_s1 ;
reg [2:0] \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.sum_s1 ;
reg [2:0] \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.ain_s1 ;
reg [2:0] \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.bin_s1 ;
reg \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.carry_s1 ;
reg [2:0] \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.sum_s1 ;
reg [5:0] add_ln691_1_reg_1284;
reg [5:0] add_ln691_2_reg_1375;
reg [1:0] add_ln691_reg_1237;
reg [5:0] add_ln69_2_reg_1314;
reg [3:0] add_ln69_reg_1207;
reg and_ln384_reg_1370;
reg and_ln414_reg_1047;
reg and_ln786_reg_1104;
reg [29:0] ap_CS_fsm = 30'h00000001;
reg carry_1_reg_1081;
reg deleted_zeros_reg_1098;
reg [14:0] empty_reg_1093;
reg icmp_ln414_reg_1020;
reg icmp_ln768_reg_1340;
reg icmp_ln786_reg_1345;
reg icmp_ln851_1_reg_1015;
reg icmp_ln851_2_reg_1127;
reg icmp_ln851_3_reg_1262;
reg icmp_ln851_reg_1137;
reg lhs_V_1_reg_1247;
reg newsignbit_reg_1326;
reg [4:0] op_22_V_reg_1242;
reg [5:0] op_25_V_reg_1350;
reg [1:0] op_5_V_reg_1152;
reg or_ln340_reg_1132;
reg or_ln785_1_reg_1358;
reg p_Result_10_reg_981;
reg p_Result_11_reg_994;
reg p_Result_12_reg_1068;
reg p_Result_13_reg_1319;
reg [4:0] p_Result_1_reg_1009;
reg [3:0] p_Result_s_reg_1004;
reg [1:0] p_Val2_1_reg_989;
reg [1:0] p_Val2_2_reg_1062;
reg [8:0] ret_V_17_reg_976;
reg [15:0] ret_V_18_reg_1110;
reg [2:0] ret_V_19_reg_1157;
reg [7:0] ret_V_20_reg_959;
reg [1:0] ret_V_21_cast_reg_1200;
reg [1:0] ret_V_21_reg_1052;
reg [2:0] ret_V_23_reg_1195;
reg [16:0] ret_V_24_reg_1232;
reg [9:0] ret_V_26_reg_1267;
reg [5:0] ret_V_27_reg_1289;
reg [5:0] ret_V_28_reg_1380;
reg [2:0] ret_V_3_reg_1147;
reg [1:0] ret_V_4_cast_reg_964;
reg [1:0] ret_V_6_reg_1042;
reg [2:0] ret_V_reg_1115;
reg [5:0] select_ln1192_reg_1385;
reg [1:0] select_ln340_reg_1142;
reg [5:0] select_ln69_reg_1309;
reg [5:0] sext_ln850_reg_1277;
reg [2:0] \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.ain_s1 ;
reg [2:0] \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.bin_s1 ;
reg \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.carry_s1 ;
reg [1:0] \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.sum_s1 ;
reg [4:0] \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.ain_s1 ;
reg [4:0] \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.bin_s1 ;
reg \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.carry_s1 ;
reg [3:0] \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.sum_s1 ;
reg [3:0] tmp_2_reg_1334;
reg [4:0] tmp_3_reg_1272;
reg [1:0] trunc_ln414_reg_999;
reg [1:0] trunc_ln728_reg_1165;
reg [1:0] trunc_ln851_1_reg_971;
reg [12:0] trunc_ln851_reg_1122;
reg underflow_1_reg_1364;
reg xor_ln416_reg_1075;
wire _000_;
wire _001_;
wire _002_;
wire [5:0] _003_;
wire [5:0] _004_;
wire [1:0] _005_;
wire [5:0] _006_;
wire [3:0] _007_;
wire _008_;
wire _009_;
wire _010_;
wire [29:0] _011_;
wire _012_;
wire _013_;
wire [14:0] _014_;
wire _015_;
wire _016_;
wire _017_;
wire _018_;
wire _019_;
wire _020_;
wire _021_;
wire _022_;
wire _023_;
wire [4:0] _024_;
wire [5:0] _025_;
wire [1:0] _026_;
wire _027_;
wire _028_;
wire _029_;
wire _030_;
wire _031_;
wire _032_;
wire [4:0] _033_;
wire [3:0] _034_;
wire [1:0] _035_;
wire [1:0] _036_;
wire [8:0] _037_;
wire [15:0] _038_;
wire [2:0] _039_;
wire [7:0] _040_;
wire [1:0] _041_;
wire [1:0] _042_;
wire [2:0] _043_;
wire [16:0] _044_;
wire [9:0] _045_;
wire [5:0] _046_;
wire [5:0] _047_;
wire [2:0] _048_;
wire [1:0] _049_;
wire [1:0] _050_;
wire [2:0] _051_;
wire [5:0] _052_;
wire [1:0] _053_;
wire [1:0] _054_;
wire [5:0] _055_;
wire [3:0] _056_;
wire [4:0] _057_;
wire [1:0] _058_;
wire [1:0] _059_;
wire [1:0] _060_;
wire [12:0] _061_;
wire _062_;
wire _063_;
wire [1:0] _064_;
wire _065_;
wire _066_;
wire _067_;
wire _068_;
wire _069_;
wire _070_;
wire _071_;
wire _072_;
wire _073_;
wire _074_;
wire _075_;
wire [4:0] _076_;
wire [4:0] _077_;
wire _078_;
wire [4:0] _079_;
wire [5:0] _080_;
wire [5:0] _081_;
wire [7:0] _082_;
wire [7:0] _083_;
wire _084_;
wire [6:0] _085_;
wire [7:0] _086_;
wire [8:0] _087_;
wire [8:0] _088_;
wire [8:0] _089_;
wire _090_;
wire [7:0] _091_;
wire [8:0] _092_;
wire [9:0] _093_;
wire _094_;
wire _095_;
wire _096_;
wire _097_;
wire [1:0] _098_;
wire [1:0] _099_;
wire _100_;
wire _101_;
wire _102_;
wire _103_;
wire [1:0] _104_;
wire [1:0] _105_;
wire _106_;
wire _107_;
wire _108_;
wire _109_;
wire [1:0] _110_;
wire [1:0] _111_;
wire [1:0] _112_;
wire [1:0] _113_;
wire _114_;
wire _115_;
wire [1:0] _116_;
wire [2:0] _117_;
wire [1:0] _118_;
wire [1:0] _119_;
wire _120_;
wire _121_;
wire [1:0] _122_;
wire [2:0] _123_;
wire [1:0] _124_;
wire [1:0] _125_;
wire _126_;
wire [1:0] _127_;
wire [2:0] _128_;
wire [2:0] _129_;
wire [2:0] _130_;
wire [2:0] _131_;
wire _132_;
wire [1:0] _133_;
wire [2:0] _134_;
wire [3:0] _135_;
wire [2:0] _136_;
wire [2:0] _137_;
wire _138_;
wire [2:0] _139_;
wire [3:0] _140_;
wire [3:0] _141_;
wire [2:0] _142_;
wire [2:0] _143_;
wire _144_;
wire [2:0] _145_;
wire [3:0] _146_;
wire [3:0] _147_;
wire [2:0] _148_;
wire [2:0] _149_;
wire _150_;
wire [2:0] _151_;
wire [3:0] _152_;
wire [3:0] _153_;
wire [2:0] _154_;
wire [2:0] _155_;
wire _156_;
wire [2:0] _157_;
wire [3:0] _158_;
wire [3:0] _159_;
wire [2:0] _160_;
wire [2:0] _161_;
wire _162_;
wire [2:0] _163_;
wire [3:0] _164_;
wire [3:0] _165_;
wire [2:0] _166_;
wire [2:0] _167_;
wire _168_;
wire [1:0] _169_;
wire [2:0] _170_;
wire [3:0] _171_;
wire [4:0] _172_;
wire [4:0] _173_;
wire _174_;
wire [3:0] _175_;
wire [4:0] _176_;
wire [5:0] _177_;
wire _178_;
wire _179_;
wire _180_;
wire _181_;
wire _182_;
wire _183_;
wire _184_;
wire _185_;
wire _186_;
wire _187_;
wire _188_;
wire _189_;
wire _190_;
wire _191_;
wire _192_;
wire _193_;
wire _194_;
wire _195_;
wire _196_;
wire _197_;
wire _198_;
wire _199_;
wire _200_;
wire _201_;
wire _202_;
wire _203_;
wire _204_;
wire _205_;
wire _206_;
wire _207_;
wire _208_;
wire _209_;
wire _210_;
wire _211_;
wire _212_;
wire _213_;
wire Range1_all_ones_fu_329_p2;
wire Range1_all_zeros_fu_334_p2;
wire Range2_all_ones_fu_324_p2;
wire \add_10ns_10s_10_2_1_U11.ce ;
wire \add_10ns_10s_10_2_1_U11.clk ;
wire [9:0] \add_10ns_10s_10_2_1_U11.din0 ;
wire [9:0] \add_10ns_10s_10_2_1_U11.din1 ;
wire [9:0] \add_10ns_10s_10_2_1_U11.dout ;
wire \add_10ns_10s_10_2_1_U11.reset ;
wire [9:0] \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.a ;
wire [9:0] \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.ain_s0 ;
wire [9:0] \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.b ;
wire [9:0] \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.bin_s0 ;
wire \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.ce ;
wire \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.clk ;
wire \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.facout_s1 ;
wire \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.facout_s2 ;
wire [4:0] \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.fas_s1 ;
wire [4:0] \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.fas_s2 ;
wire \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.reset ;
wire [9:0] \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.s ;
wire [4:0] \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.u1.a ;
wire [4:0] \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.u1.b ;
wire \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.u1.cin ;
wire \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.u1.cout ;
wire [4:0] \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.u1.s ;
wire [4:0] \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.u2.a ;
wire [4:0] \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.u2.b ;
wire \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.u2.cin ;
wire \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.u2.cout ;
wire [4:0] \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.u2.s ;
wire \add_15ns_15ns_15_2_1_U6.ce ;
wire \add_15ns_15ns_15_2_1_U6.clk ;
wire [14:0] \add_15ns_15ns_15_2_1_U6.din0 ;
wire [14:0] \add_15ns_15ns_15_2_1_U6.din1 ;
wire [14:0] \add_15ns_15ns_15_2_1_U6.dout ;
wire \add_15ns_15ns_15_2_1_U6.reset ;
wire [14:0] \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.a ;
wire [14:0] \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.ain_s0 ;
wire [14:0] \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.b ;
wire [14:0] \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.bin_s0 ;
wire \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.ce ;
wire \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.clk ;
wire \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.facout_s1 ;
wire \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.facout_s2 ;
wire [6:0] \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.fas_s1 ;
wire [7:0] \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.fas_s2 ;
wire \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.reset ;
wire [14:0] \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.s ;
wire [6:0] \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.u1.a ;
wire [6:0] \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.u1.b ;
wire \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.u1.cin ;
wire \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.u1.cout ;
wire [6:0] \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.u1.s ;
wire [7:0] \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.u2.a ;
wire [7:0] \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.u2.b ;
wire \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.u2.cin ;
wire \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.u2.cout ;
wire [7:0] \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.u2.s ;
wire \add_17s_17s_17_2_1_U8.ce ;
wire \add_17s_17s_17_2_1_U8.clk ;
wire [16:0] \add_17s_17s_17_2_1_U8.din0 ;
wire [16:0] \add_17s_17s_17_2_1_U8.din1 ;
wire [16:0] \add_17s_17s_17_2_1_U8.dout ;
wire \add_17s_17s_17_2_1_U8.reset ;
wire [16:0] \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.a ;
wire [16:0] \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.ain_s0 ;
wire [16:0] \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.b ;
wire [16:0] \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.bin_s0 ;
wire \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.ce ;
wire \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.clk ;
wire \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.facout_s1 ;
wire \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.facout_s2 ;
wire [7:0] \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.fas_s1 ;
wire [8:0] \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.fas_s2 ;
wire \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.reset ;
wire [16:0] \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.s ;
wire [7:0] \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.u1.a ;
wire [7:0] \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.u1.b ;
wire \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.u1.cin ;
wire \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.u1.cout ;
wire [7:0] \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.u1.s ;
wire [8:0] \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.u2.a ;
wire [8:0] \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.u2.b ;
wire \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.u2.cin ;
wire \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.u2.cout ;
wire [8:0] \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.u2.s ;
wire \add_2ns_2ns_2_2_1_U2.ce ;
wire \add_2ns_2ns_2_2_1_U2.clk ;
wire [1:0] \add_2ns_2ns_2_2_1_U2.din0 ;
wire [1:0] \add_2ns_2ns_2_2_1_U2.din1 ;
wire [1:0] \add_2ns_2ns_2_2_1_U2.dout ;
wire \add_2ns_2ns_2_2_1_U2.reset ;
wire [1:0] \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.a ;
wire [1:0] \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.ain_s0 ;
wire [1:0] \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.b ;
wire [1:0] \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.bin_s0 ;
wire \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.ce ;
wire \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.clk ;
wire \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.facout_s1 ;
wire \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.facout_s2 ;
wire \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.fas_s1 ;
wire \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.fas_s2 ;
wire \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.reset ;
wire [1:0] \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.s ;
wire \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.a ;
wire \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.b ;
wire \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.cin ;
wire \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.cout ;
wire \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.s ;
wire \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.a ;
wire \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.b ;
wire \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.cin ;
wire \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.cout ;
wire \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.s ;
wire \add_2ns_2ns_2_2_1_U3.ce ;
wire \add_2ns_2ns_2_2_1_U3.clk ;
wire [1:0] \add_2ns_2ns_2_2_1_U3.din0 ;
wire [1:0] \add_2ns_2ns_2_2_1_U3.din1 ;
wire [1:0] \add_2ns_2ns_2_2_1_U3.dout ;
wire \add_2ns_2ns_2_2_1_U3.reset ;
wire [1:0] \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.a ;
wire [1:0] \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.ain_s0 ;
wire [1:0] \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.b ;
wire [1:0] \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.bin_s0 ;
wire \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.ce ;
wire \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.clk ;
wire \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.facout_s1 ;
wire \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.facout_s2 ;
wire \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.fas_s1 ;
wire \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.fas_s2 ;
wire \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.reset ;
wire [1:0] \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.s ;
wire \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.a ;
wire \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.b ;
wire \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.cin ;
wire \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.cout ;
wire \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.s ;
wire \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.a ;
wire \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.b ;
wire \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.cin ;
wire \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.cout ;
wire \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.s ;
wire \add_2ns_2ns_2_2_1_U9.ce ;
wire \add_2ns_2ns_2_2_1_U9.clk ;
wire [1:0] \add_2ns_2ns_2_2_1_U9.din0 ;
wire [1:0] \add_2ns_2ns_2_2_1_U9.din1 ;
wire [1:0] \add_2ns_2ns_2_2_1_U9.dout ;
wire \add_2ns_2ns_2_2_1_U9.reset ;
wire [1:0] \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.a ;
wire [1:0] \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.ain_s0 ;
wire [1:0] \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.b ;
wire [1:0] \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.bin_s0 ;
wire \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.ce ;
wire \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.clk ;
wire \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.facout_s1 ;
wire \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.facout_s2 ;
wire \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.fas_s1 ;
wire \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.fas_s2 ;
wire \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.reset ;
wire [1:0] \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.s ;
wire \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.a ;
wire \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.b ;
wire \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.cin ;
wire \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.cout ;
wire \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.s ;
wire \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.a ;
wire \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.b ;
wire \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.cin ;
wire \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.cout ;
wire \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.s ;
wire \add_3ns_3ns_3_2_1_U4.ce ;
wire \add_3ns_3ns_3_2_1_U4.clk ;
wire [2:0] \add_3ns_3ns_3_2_1_U4.din0 ;
wire [2:0] \add_3ns_3ns_3_2_1_U4.din1 ;
wire [2:0] \add_3ns_3ns_3_2_1_U4.dout ;
wire \add_3ns_3ns_3_2_1_U4.reset ;
wire [2:0] \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.a ;
wire [2:0] \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.ain_s0 ;
wire [2:0] \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.b ;
wire [2:0] \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.bin_s0 ;
wire \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.ce ;
wire \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.clk ;
wire \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.facout_s1 ;
wire \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.facout_s2 ;
wire \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.fas_s1 ;
wire [1:0] \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.fas_s2 ;
wire \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.reset ;
wire [2:0] \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.s ;
wire \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.u1.a ;
wire \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.u1.b ;
wire \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.u1.cin ;
wire \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.u1.cout ;
wire \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.u1.s ;
wire [1:0] \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.u2.a ;
wire [1:0] \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.u2.b ;
wire \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.u2.cin ;
wire \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.u2.cout ;
wire [1:0] \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.u2.s ;
wire \add_3s_3s_3_2_1_U5.ce ;
wire \add_3s_3s_3_2_1_U5.clk ;
wire [2:0] \add_3s_3s_3_2_1_U5.din0 ;
wire [2:0] \add_3s_3s_3_2_1_U5.din1 ;
wire [2:0] \add_3s_3s_3_2_1_U5.dout ;
wire \add_3s_3s_3_2_1_U5.reset ;
wire [2:0] \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.a ;
wire [2:0] \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.ain_s0 ;
wire [2:0] \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.b ;
wire [2:0] \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.bin_s0 ;
wire \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.ce ;
wire \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.clk ;
wire \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.facout_s1 ;
wire \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.facout_s2 ;
wire \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.fas_s1 ;
wire [1:0] \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.fas_s2 ;
wire \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.reset ;
wire [2:0] \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.s ;
wire \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.u1.a ;
wire \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.u1.b ;
wire \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.u1.cin ;
wire \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.u1.cout ;
wire \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.u1.s ;
wire [1:0] \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.u2.a ;
wire [1:0] \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.u2.b ;
wire \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.u2.cin ;
wire \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.u2.cout ;
wire [1:0] \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.u2.s ;
wire \add_4s_4ns_4_2_1_U7.ce ;
wire \add_4s_4ns_4_2_1_U7.clk ;
wire [3:0] \add_4s_4ns_4_2_1_U7.din0 ;
wire [3:0] \add_4s_4ns_4_2_1_U7.din1 ;
wire [3:0] \add_4s_4ns_4_2_1_U7.dout ;
wire \add_4s_4ns_4_2_1_U7.reset ;
wire [3:0] \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.a ;
wire [3:0] \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.ain_s0 ;
wire [3:0] \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.b ;
wire [3:0] \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.bin_s0 ;
wire \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.ce ;
wire \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.clk ;
wire \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.facout_s1 ;
wire \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.facout_s2 ;
wire [1:0] \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.fas_s1 ;
wire [1:0] \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.fas_s2 ;
wire \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.reset ;
wire [3:0] \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.s ;
wire [1:0] \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.u1.a ;
wire [1:0] \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.u1.b ;
wire \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.u1.cin ;
wire \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.u1.cout ;
wire [1:0] \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.u1.s ;
wire [1:0] \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.u2.a ;
wire [1:0] \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.u2.b ;
wire \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.u2.cin ;
wire \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.u2.cout ;
wire [1:0] \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.u2.s ;
wire \add_5s_5s_5_2_1_U10.ce ;
wire \add_5s_5s_5_2_1_U10.clk ;
wire [4:0] \add_5s_5s_5_2_1_U10.din0 ;
wire [4:0] \add_5s_5s_5_2_1_U10.din1 ;
wire [4:0] \add_5s_5s_5_2_1_U10.dout ;
wire \add_5s_5s_5_2_1_U10.reset ;
wire [4:0] \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.a ;
wire [4:0] \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.ain_s0 ;
wire [4:0] \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.b ;
wire [4:0] \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.bin_s0 ;
wire \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.ce ;
wire \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.clk ;
wire \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.facout_s1 ;
wire \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.facout_s2 ;
wire [1:0] \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.fas_s1 ;
wire [2:0] \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.fas_s2 ;
wire \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.reset ;
wire [4:0] \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.s ;
wire [1:0] \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.u1.a ;
wire [1:0] \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.u1.b ;
wire \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.u1.cin ;
wire \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.u1.cout ;
wire [1:0] \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.u1.s ;
wire [2:0] \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.u2.a ;
wire [2:0] \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.u2.b ;
wire \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.u2.cin ;
wire \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.u2.cout ;
wire [2:0] \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.u2.s ;
wire \add_6ns_6ns_6_2_1_U15.ce ;
wire \add_6ns_6ns_6_2_1_U15.clk ;
wire [5:0] \add_6ns_6ns_6_2_1_U15.din0 ;
wire [5:0] \add_6ns_6ns_6_2_1_U15.din1 ;
wire [5:0] \add_6ns_6ns_6_2_1_U15.dout ;
wire \add_6ns_6ns_6_2_1_U15.reset ;
wire [5:0] \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.a ;
wire [5:0] \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.ain_s0 ;
wire [5:0] \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.b ;
wire [5:0] \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.bin_s0 ;
wire \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.ce ;
wire \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.clk ;
wire \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.facout_s1 ;
wire \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.facout_s2 ;
wire [2:0] \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.fas_s1 ;
wire [2:0] \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.fas_s2 ;
wire \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.reset ;
wire [5:0] \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.s ;
wire [2:0] \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.u1.a ;
wire [2:0] \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.u1.b ;
wire \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.u1.cin ;
wire \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.u1.cout ;
wire [2:0] \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.u1.s ;
wire [2:0] \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.u2.a ;
wire [2:0] \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.u2.b ;
wire \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.u2.cin ;
wire \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.u2.cout ;
wire [2:0] \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.u2.s ;
wire \add_6ns_6ns_6_2_1_U16.ce ;
wire \add_6ns_6ns_6_2_1_U16.clk ;
wire [5:0] \add_6ns_6ns_6_2_1_U16.din0 ;
wire [5:0] \add_6ns_6ns_6_2_1_U16.din1 ;
wire [5:0] \add_6ns_6ns_6_2_1_U16.dout ;
wire \add_6ns_6ns_6_2_1_U16.reset ;
wire [5:0] \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.a ;
wire [5:0] \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.ain_s0 ;
wire [5:0] \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.b ;
wire [5:0] \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.bin_s0 ;
wire \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.ce ;
wire \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.clk ;
wire \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.facout_s1 ;
wire \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.facout_s2 ;
wire [2:0] \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.fas_s1 ;
wire [2:0] \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.fas_s2 ;
wire \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.reset ;
wire [5:0] \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.s ;
wire [2:0] \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.u1.a ;
wire [2:0] \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.u1.b ;
wire \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.u1.cin ;
wire \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.u1.cout ;
wire [2:0] \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.u1.s ;
wire [2:0] \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.u2.a ;
wire [2:0] \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.u2.b ;
wire \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.u2.cin ;
wire \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.u2.cout ;
wire [2:0] \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.u2.s ;
wire \add_6ns_6ns_6_2_1_U17.ce ;
wire \add_6ns_6ns_6_2_1_U17.clk ;
wire [5:0] \add_6ns_6ns_6_2_1_U17.din0 ;
wire [5:0] \add_6ns_6ns_6_2_1_U17.din1 ;
wire [5:0] \add_6ns_6ns_6_2_1_U17.dout ;
wire \add_6ns_6ns_6_2_1_U17.reset ;
wire [5:0] \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.a ;
wire [5:0] \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.ain_s0 ;
wire [5:0] \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.b ;
wire [5:0] \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.bin_s0 ;
wire \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.ce ;
wire \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.clk ;
wire \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.facout_s1 ;
wire \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.facout_s2 ;
wire [2:0] \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.fas_s1 ;
wire [2:0] \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.fas_s2 ;
wire \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.reset ;
wire [5:0] \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.s ;
wire [2:0] \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.u1.a ;
wire [2:0] \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.u1.b ;
wire \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.u1.cin ;
wire \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.u1.cout ;
wire [2:0] \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.u1.s ;
wire [2:0] \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.u2.a ;
wire [2:0] \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.u2.b ;
wire \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.u2.cin ;
wire \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.u2.cout ;
wire [2:0] \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.u2.s ;
wire \add_6ns_6s_6_2_1_U13.ce ;
wire \add_6ns_6s_6_2_1_U13.clk ;
wire [5:0] \add_6ns_6s_6_2_1_U13.din0 ;
wire [5:0] \add_6ns_6s_6_2_1_U13.din1 ;
wire [5:0] \add_6ns_6s_6_2_1_U13.dout ;
wire \add_6ns_6s_6_2_1_U13.reset ;
wire [5:0] \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.a ;
wire [5:0] \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.ain_s0 ;
wire [5:0] \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.b ;
wire [5:0] \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.bin_s0 ;
wire \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.ce ;
wire \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.clk ;
wire \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.facout_s1 ;
wire \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.facout_s2 ;
wire [2:0] \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.fas_s1 ;
wire [2:0] \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.fas_s2 ;
wire \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.reset ;
wire [5:0] \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.s ;
wire [2:0] \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.u1.a ;
wire [2:0] \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.u1.b ;
wire \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.u1.cin ;
wire \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.u1.cout ;
wire [2:0] \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.u1.s ;
wire [2:0] \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.u2.a ;
wire [2:0] \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.u2.b ;
wire \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.u2.cin ;
wire \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.u2.cout ;
wire [2:0] \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.u2.s ;
wire \add_6s_6ns_6_2_1_U12.ce ;
wire \add_6s_6ns_6_2_1_U12.clk ;
wire [5:0] \add_6s_6ns_6_2_1_U12.din0 ;
wire [5:0] \add_6s_6ns_6_2_1_U12.din1 ;
wire [5:0] \add_6s_6ns_6_2_1_U12.dout ;
wire \add_6s_6ns_6_2_1_U12.reset ;
wire [5:0] \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.a ;
wire [5:0] \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.ain_s0 ;
wire [5:0] \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.b ;
wire [5:0] \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.bin_s0 ;
wire \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.ce ;
wire \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.clk ;
wire \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.facout_s1 ;
wire \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.facout_s2 ;
wire [2:0] \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.fas_s1 ;
wire [2:0] \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.fas_s2 ;
wire \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.reset ;
wire [5:0] \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.s ;
wire [2:0] \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.u1.a ;
wire [2:0] \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.u1.b ;
wire \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.u1.cin ;
wire \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.u1.cout ;
wire [2:0] \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.u1.s ;
wire [2:0] \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.u2.a ;
wire [2:0] \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.u2.b ;
wire \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.u2.cin ;
wire \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.u2.cout ;
wire [2:0] \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.u2.s ;
wire and_ln384_fu_881_p2;
wire and_ln414_fu_339_p2;
wire and_ln780_fu_409_p2;
wire and_ln781_fu_498_p2;
wire and_ln785_1_fu_534_p2;
wire and_ln785_fu_525_p2;
wire and_ln786_fu_420_p2;
wire and_ln850_fu_774_p2;
wire ap_CS_fsm_state1;
wire ap_CS_fsm_state10;
wire ap_CS_fsm_state11;
wire ap_CS_fsm_state12;
wire ap_CS_fsm_state13;
wire ap_CS_fsm_state14;
wire ap_CS_fsm_state15;
wire ap_CS_fsm_state16;
wire ap_CS_fsm_state17;
wire ap_CS_fsm_state18;
wire ap_CS_fsm_state19;
wire ap_CS_fsm_state2;
wire ap_CS_fsm_state20;
wire ap_CS_fsm_state21;
wire ap_CS_fsm_state22;
wire ap_CS_fsm_state23;
wire ap_CS_fsm_state24;
wire ap_CS_fsm_state25;
wire ap_CS_fsm_state26;
wire ap_CS_fsm_state27;
wire ap_CS_fsm_state28;
wire ap_CS_fsm_state29;
wire ap_CS_fsm_state3;
wire ap_CS_fsm_state30;
wire ap_CS_fsm_state4;
wire ap_CS_fsm_state5;
wire ap_CS_fsm_state6;
wire ap_CS_fsm_state7;
wire ap_CS_fsm_state8;
wire ap_CS_fsm_state9;
wire [29:0] ap_NS_fsm;
wire ap_clk;
wire ap_done;
wire ap_idle;
wire ap_ready;
wire ap_rst;
wire ap_start;
wire carry_1_fu_383_p2;
wire deleted_ones_fu_414_p3;
wire deleted_zeros_fu_391_p3;
wire [15:0] empty_fu_387_p0;
wire [14:0] empty_fu_387_p1;
wire [8:0] grp_fu_221_p0;
wire [8:0] grp_fu_221_p1;
wire [8:0] grp_fu_221_p2;
wire [1:0] grp_fu_314_p2;
wire [1:0] grp_fu_365_p1;
wire [1:0] grp_fu_365_p2;
wire [2:0] grp_fu_493_p2;
wire [2:0] grp_fu_578_p0;
wire [2:0] grp_fu_578_p1;
wire [2:0] grp_fu_578_p2;
wire [14:0] grp_fu_591_p0;
wire [14:0] grp_fu_591_p2;
wire [3:0] grp_fu_600_p0;
wire [3:0] grp_fu_600_p1;
wire [3:0] grp_fu_600_p2;
wire [16:0] grp_fu_633_p0;
wire [16:0] grp_fu_633_p1;
wire [16:0] grp_fu_633_p2;
wire [1:0] grp_fu_639_p2;
wire [4:0] grp_fu_647_p0;
wire [4:0] grp_fu_647_p1;
wire [4:0] grp_fu_647_p2;
wire [9:0] grp_fu_692_p0;
wire [9:0] grp_fu_692_p1;
wire [9:0] grp_fu_692_p2;
wire [5:0] grp_fu_721_p0;
wire [5:0] grp_fu_721_p2;
wire [5:0] grp_fu_749_p1;
wire [5:0] grp_fu_749_p2;
wire [4:0] grp_fu_793_p0;
wire [4:0] grp_fu_793_p1;
wire [4:0] grp_fu_793_p2;
wire [5:0] grp_fu_829_p2;
wire [5:0] grp_fu_862_p2;
wire [5:0] grp_fu_935_p2;
wire icmp_ln414_fu_319_p2;
wire icmp_ln768_fu_833_p2;
wire icmp_ln786_fu_838_p2;
wire icmp_ln851_1_fu_309_p2;
wire icmp_ln851_2_fu_456_p2;
wire icmp_ln851_3_fu_702_p2;
wire icmp_ln851_fu_488_p2;
wire [15:0] lhs_1_fu_425_p3;
wire lhs_V_1_fu_676_p2;
wire [4:0] lhs_fu_205_p3;
wire neg_src_fu_508_p2;
wire newsignbit_fu_815_p1;
wire [1:0] op_0;
wire [3:0] op_1;
wire [3:0] op_10;
wire [1:0] op_12;
wire [3:0] op_13;
wire [7:0] op_14;
wire op_19_V_fu_902_p3;
wire [7:0] op_2;
wire [31:0] op_28;
wire op_28_ap_vld;
wire [15:0] op_3;
wire [1:0] op_5_V_fu_539_p3;
wire [1:0] op_7;
wire [1:0] op_8;
wire or_ln340_1_fu_897_p2;
wire or_ln340_2_fu_513_p2;
wire or_ln340_fu_483_p2;
wire or_ln384_fu_876_p2;
wire or_ln388_fu_867_p2;
wire or_ln785_1_fu_843_p2;
wire or_ln785_2_fu_529_p2;
wire or_ln785_fu_467_p2;
wire or_ln786_fu_852_p2;
wire overflow_1_fu_892_p2;
wire overflow_fu_477_p2;
wire p_Result_2_fu_343_p3;
wire p_Result_3_fu_762_p3;
wire p_Result_5_fu_653_p3;
wire p_Result_8_fu_727_p3;
wire p_Result_9_fu_908_p3;
wire p_Result_s_16_fu_545_p3;
wire [15:0] ret_V_18_fu_432_p1;
wire [15:0] ret_V_18_fu_432_p2;
wire [2:0] ret_V_19_fu_557_p3;
wire [7:0] ret_V_20_fu_239_p1;
wire [7:0] ret_V_20_fu_239_p2;
wire [1:0] ret_V_21_fu_355_p3;
wire ret_V_22_fu_780_p2;
wire [1:0] ret_V_25_fu_665_p3;
wire [5:0] ret_V_27_fu_739_p3;
wire [5:0] ret_V_28_fu_920_p3;
wire ret_V_8_fu_754_p3;
wire [15:0] rhs_3_fu_622_p3;
wire [3:0] rhs_fu_227_p3;
wire [5:0] select_ln1192_fu_927_p3;
wire [1:0] select_ln340_fu_518_p3;
wire [1:0] select_ln69_fu_799_p3;
wire [1:0] select_ln850_1_fu_350_p3;
wire [1:0] select_ln850_2_fu_660_p3;
wire [5:0] select_ln850_3_fu_734_p3;
wire [5:0] select_ln850_4_fu_915_p3;
wire [2:0] select_ln850_fu_552_p3;
wire [7:0] sext_ln1192_2_fu_681_p0;
wire [15:0] sext_ln1192_fu_619_p0;
wire [7:0] sext_ln1195_fu_235_p1;
wire [7:0] sext_ln703_fu_217_p0;
wire [5:0] sext_ln850_fu_718_p1;
wire \sub_5s_5s_5_2_1_U14.ce ;
wire \sub_5s_5s_5_2_1_U14.clk ;
wire [4:0] \sub_5s_5s_5_2_1_U14.din0 ;
wire [4:0] \sub_5s_5s_5_2_1_U14.din1 ;
wire [4:0] \sub_5s_5s_5_2_1_U14.dout ;
wire \sub_5s_5s_5_2_1_U14.reset ;
wire [4:0] \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.a ;
wire [4:0] \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.ain_s0 ;
wire [4:0] \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.b ;
wire [4:0] \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.bin_s0 ;
wire \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.ce ;
wire \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.clk ;
wire \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.facout_s1 ;
wire \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.facout_s2 ;
wire [1:0] \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.fas_s1 ;
wire [2:0] \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.fas_s2 ;
wire \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.reset ;
wire [4:0] \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.s ;
wire [1:0] \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.u1.a ;
wire [1:0] \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.u1.b ;
wire \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.u1.cin ;
wire \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.u1.cout ;
wire [1:0] \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.u1.s ;
wire [2:0] \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.u2.a ;
wire [2:0] \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.u2.b ;
wire \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.u2.cin ;
wire \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.u2.cout ;
wire [2:0] \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.u2.s ;
wire \sub_9s_9s_9_2_1_U1.ce ;
wire \sub_9s_9s_9_2_1_U1.clk ;
wire [8:0] \sub_9s_9s_9_2_1_U1.din0 ;
wire [8:0] \sub_9s_9s_9_2_1_U1.din1 ;
wire [8:0] \sub_9s_9s_9_2_1_U1.dout ;
wire \sub_9s_9s_9_2_1_U1.reset ;
wire [8:0] \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.a ;
wire [8:0] \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.ain_s0 ;
wire [8:0] \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.b ;
wire [8:0] \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.bin_s0 ;
wire \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.ce ;
wire \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.clk ;
wire \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.facout_s1 ;
wire \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.facout_s2 ;
wire [3:0] \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.fas_s1 ;
wire [4:0] \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.fas_s2 ;
wire \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.reset ;
wire [8:0] \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.s ;
wire [3:0] \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.u1.a ;
wire [3:0] \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.u1.b ;
wire \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.u1.cin ;
wire \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.u1.cout ;
wire [3:0] \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.u1.s ;
wire [4:0] \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.u2.a ;
wire [4:0] \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.u2.b ;
wire \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.u2.cin ;
wire \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.u2.cout ;
wire [4:0] \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.u2.s ;
wire tmp_fu_396_p3;
wire [1:0] trunc_ln414_fu_285_p1;
wire [1:0] trunc_ln728_fu_564_p1;
wire [1:0] trunc_ln851_1_fu_255_p1;
wire trunc_ln851_2_fu_770_p1;
wire [15:0] trunc_ln851_3_fu_452_p0;
wire [12:0] trunc_ln851_3_fu_452_p1;
wire [7:0] trunc_ln851_4_fu_698_p0;
wire [4:0] trunc_ln851_4_fu_698_p1;
wire [12:0] trunc_ln851_fu_448_p1;
wire underflow_1_fu_857_p2;
wire xor_ln384_fu_871_p2;
wire xor_ln416_fu_378_p2;
wire xor_ln780_fu_403_p2;
wire xor_ln781_fu_502_p2;
wire xor_ln785_1_fu_472_p2;
wire xor_ln785_2_fu_887_p2;
wire xor_ln785_fu_462_p2;
wire xor_ln786_fu_847_p2;
wire [2:0] zext_ln886_fu_672_p1;


assign _065_ = icmp_ln851_3_reg_1262 & ap_CS_fsm[19];
assign _066_ = lhs_V_1_reg_1247 & ap_CS_fsm[26];
assign _067_ = ap_CS_fsm[15] & icmp_ln851_2_reg_1127;
assign _068_ = _070_ & ap_CS_fsm[0];
assign _069_ = ap_start & ap_CS_fsm[0];
assign and_ln384_fu_881_p2 = or_ln388_fu_867_p2 & or_ln384_fu_876_p2;
assign and_ln414_fu_339_p2 = p_Result_10_reg_981 & icmp_ln414_reg_1020;
assign and_ln780_fu_409_p2 = xor_ln780_fu_403_p2 & Range2_all_ones_reg_1025;
assign and_ln781_fu_498_p2 = carry_1_reg_1081 & Range1_all_ones_reg_1030;
assign and_ln785_1_fu_534_p2 = or_ln785_2_fu_529_p2 & and_ln786_reg_1104;
assign and_ln785_fu_525_p2 = xor_ln416_reg_1075 & deleted_zeros_reg_1098;
assign and_ln786_fu_420_p2 = p_Result_12_reg_1068 & deleted_ones_fu_414_p3;
assign and_ln850_fu_774_p2 = op_8[0] & op_8[1];
assign carry_1_fu_383_p2 = xor_ln416_reg_1075 & p_Result_11_reg_994;
assign neg_src_fu_508_p2 = xor_ln781_fu_502_p2 & p_Result_10_reg_981;
assign overflow_1_fu_892_p2 = xor_ln785_2_fu_887_p2 & or_ln785_1_reg_1358;
assign overflow_fu_477_p2 = xor_ln785_1_fu_472_p2 & or_ln785_fu_467_p2;
assign underflow_1_fu_857_p2 = p_Result_13_reg_1319 & or_ln786_fu_852_p2;
assign xor_ln384_fu_871_p2 = ~ or_ln785_1_reg_1358;
assign xor_ln780_fu_403_p2 = ~ ret_V_17_reg_976[4];
assign xor_ln781_fu_502_p2 = ~ and_ln781_fu_498_p2;
assign xor_ln785_2_fu_887_p2 = ~ p_Result_13_reg_1319;
assign xor_ln785_fu_462_p2 = ~ deleted_zeros_reg_1098;
assign xor_ln785_1_fu_472_p2 = ~ p_Result_10_reg_981;
assign xor_ln786_fu_847_p2 = ~ newsignbit_reg_1326;
assign xor_ln416_fu_378_p2 = ~ p_Result_12_reg_1068;
assign _070_ = ~ ap_start;
assign _071_ = p_Result_1_reg_1009 == 5'h1f;
assign _072_ = ! p_Result_1_reg_1009;
assign _073_ = p_Result_s_reg_1004 == 4'hf;
assign _074_ = ! trunc_ln851_1_reg_971;
assign _075_ = ! trunc_ln851_reg_1122;
always @(posedge \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.clk )
\add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.bin_s1  <= _077_;
always @(posedge \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.clk )
\add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.ain_s1  <= _076_;
always @(posedge \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.clk )
\add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.sum_s1  <= _079_;
always @(posedge \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.clk )
\add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.carry_s1  <= _078_;
assign _077_ = \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.ce  ? \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.b [9:5] : \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.bin_s1 ;
assign _076_ = \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.ce  ? \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.a [9:5] : \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.ain_s1 ;
assign _078_ = \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.ce  ? \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.facout_s1  : \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.carry_s1 ;
assign _079_ = \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.ce  ? \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.fas_s1  : \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.sum_s1 ;
assign _080_ = \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.u1.a  + \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.u1.b ;
assign { \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.u1.cout , \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.u1.s  } = _080_ + \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.u1.cin ;
assign _081_ = \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.u2.a  + \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.u2.b ;
assign { \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.u2.cout , \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.u2.s  } = _081_ + \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.u2.cin ;
always @(posedge \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.clk )
\add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.bin_s1  <= _083_;
always @(posedge \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.clk )
\add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.ain_s1  <= _082_;
always @(posedge \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.clk )
\add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.sum_s1  <= _085_;
always @(posedge \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.clk )
\add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.carry_s1  <= _084_;
assign _083_ = \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.ce  ? \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.b [14:7] : \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.bin_s1 ;
assign _082_ = \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.ce  ? \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.a [14:7] : \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.ain_s1 ;
assign _084_ = \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.ce  ? \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.facout_s1  : \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.carry_s1 ;
assign _085_ = \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.ce  ? \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.fas_s1  : \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.sum_s1 ;
assign _086_ = \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.u1.a  + \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.u1.b ;
assign { \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.u1.cout , \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.u1.s  } = _086_ + \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.u1.cin ;
assign _087_ = \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.u2.a  + \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.u2.b ;
assign { \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.u2.cout , \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.u2.s  } = _087_ + \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.u2.cin ;
always @(posedge \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.clk )
\add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.bin_s1  <= _089_;
always @(posedge \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.clk )
\add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.ain_s1  <= _088_;
always @(posedge \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.clk )
\add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.sum_s1  <= _091_;
always @(posedge \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.clk )
\add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.carry_s1  <= _090_;
assign _089_ = \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.ce  ? \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.b [16:8] : \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.bin_s1 ;
assign _088_ = \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.ce  ? \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.a [16:8] : \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.ain_s1 ;
assign _090_ = \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.ce  ? \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.facout_s1  : \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.carry_s1 ;
assign _091_ = \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.ce  ? \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.fas_s1  : \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.sum_s1 ;
assign _092_ = \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.u1.a  + \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.u1.b ;
assign { \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.u1.cout , \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.u1.s  } = _092_ + \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.u1.cin ;
assign _093_ = \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.u2.a  + \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.u2.b ;
assign { \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.u2.cout , \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.u2.s  } = _093_ + \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.u2.cin ;
always @(posedge \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.clk )
\add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.bin_s1  <= _095_;
always @(posedge \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.clk )
\add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.ain_s1  <= _094_;
always @(posedge \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.clk )
\add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.sum_s1  <= _097_;
always @(posedge \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.clk )
\add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.carry_s1  <= _096_;
assign _095_ = \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.ce  ? \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.b [1] : \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.bin_s1 ;
assign _094_ = \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.ce  ? \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.a [1] : \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.ain_s1 ;
assign _096_ = \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.ce  ? \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.facout_s1  : \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.carry_s1 ;
assign _097_ = \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.ce  ? \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.fas_s1  : \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.sum_s1 ;
assign _098_ = \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.a  + \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.b ;
assign { \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.cout , \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.s  } = _098_ + \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.cin ;
assign _099_ = \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.a  + \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.b ;
assign { \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.cout , \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.s  } = _099_ + \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.cin ;
always @(posedge \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.clk )
\add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.bin_s1  <= _101_;
always @(posedge \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.clk )
\add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.ain_s1  <= _100_;
always @(posedge \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.clk )
\add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.sum_s1  <= _103_;
always @(posedge \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.clk )
\add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.carry_s1  <= _102_;
assign _101_ = \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.ce  ? \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.b [1] : \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.bin_s1 ;
assign _100_ = \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.ce  ? \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.a [1] : \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.ain_s1 ;
assign _102_ = \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.ce  ? \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.facout_s1  : \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.carry_s1 ;
assign _103_ = \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.ce  ? \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.fas_s1  : \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.sum_s1 ;
assign _104_ = \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.a  + \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.b ;
assign { \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.cout , \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.s  } = _104_ + \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.cin ;
assign _105_ = \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.a  + \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.b ;
assign { \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.cout , \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.s  } = _105_ + \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.cin ;
always @(posedge \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.clk )
\add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.bin_s1  <= _107_;
always @(posedge \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.clk )
\add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.ain_s1  <= _106_;
always @(posedge \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.clk )
\add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.sum_s1  <= _109_;
always @(posedge \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.clk )
\add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.carry_s1  <= _108_;
assign _107_ = \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.ce  ? \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.b [1] : \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.bin_s1 ;
assign _106_ = \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.ce  ? \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.a [1] : \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.ain_s1 ;
assign _108_ = \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.ce  ? \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.facout_s1  : \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.carry_s1 ;
assign _109_ = \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.ce  ? \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.fas_s1  : \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.sum_s1 ;
assign _110_ = \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.a  + \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.b ;
assign { \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.cout , \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.s  } = _110_ + \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.cin ;
assign _111_ = \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.a  + \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.b ;
assign { \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.cout , \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.s  } = _111_ + \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.cin ;
always @(posedge \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.clk )
\add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.bin_s1  <= _113_;
always @(posedge \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.clk )
\add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.ain_s1  <= _112_;
always @(posedge \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.clk )
\add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.sum_s1  <= _115_;
always @(posedge \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.clk )
\add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.carry_s1  <= _114_;
assign _113_ = \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.ce  ? \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.b [2:1] : \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.bin_s1 ;
assign _112_ = \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.ce  ? \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.a [2:1] : \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.ain_s1 ;
assign _114_ = \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.ce  ? \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.facout_s1  : \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.carry_s1 ;
assign _115_ = \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.ce  ? \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.fas_s1  : \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.sum_s1 ;
assign _116_ = \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.u1.a  + \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.u1.b ;
assign { \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.u1.cout , \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.u1.s  } = _116_ + \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.u1.cin ;
assign _117_ = \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.u2.a  + \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.u2.b ;
assign { \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.u2.cout , \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.u2.s  } = _117_ + \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.u2.cin ;
always @(posedge \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.clk )
\add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.bin_s1  <= _119_;
always @(posedge \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.clk )
\add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.ain_s1  <= _118_;
always @(posedge \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.clk )
\add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.sum_s1  <= _121_;
always @(posedge \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.clk )
\add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.carry_s1  <= _120_;
assign _119_ = \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.ce  ? \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.b [2:1] : \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.bin_s1 ;
assign _118_ = \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.ce  ? \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.a [2:1] : \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.ain_s1 ;
assign _120_ = \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.ce  ? \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.facout_s1  : \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.carry_s1 ;
assign _121_ = \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.ce  ? \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.fas_s1  : \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.sum_s1 ;
assign _122_ = \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.u1.a  + \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.u1.b ;
assign { \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.u1.cout , \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.u1.s  } = _122_ + \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.u1.cin ;
assign _123_ = \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.u2.a  + \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.u2.b ;
assign { \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.u2.cout , \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.u2.s  } = _123_ + \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.u2.cin ;
always @(posedge \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.clk )
\add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.bin_s1  <= _125_;
always @(posedge \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.clk )
\add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.ain_s1  <= _124_;
always @(posedge \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.clk )
\add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.sum_s1  <= _127_;
always @(posedge \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.clk )
\add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.carry_s1  <= _126_;
assign _125_ = \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.ce  ? \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.b [3:2] : \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.bin_s1 ;
assign _124_ = \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.ce  ? \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.a [3:2] : \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.ain_s1 ;
assign _126_ = \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.ce  ? \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.facout_s1  : \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.carry_s1 ;
assign _127_ = \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.ce  ? \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.fas_s1  : \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.sum_s1 ;
assign _128_ = \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.u1.a  + \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.u1.b ;
assign { \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.u1.cout , \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.u1.s  } = _128_ + \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.u1.cin ;
assign _129_ = \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.u2.a  + \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.u2.b ;
assign { \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.u2.cout , \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.u2.s  } = _129_ + \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.u2.cin ;
always @(posedge \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.clk )
\add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.bin_s1  <= _131_;
always @(posedge \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.clk )
\add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.ain_s1  <= _130_;
always @(posedge \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.clk )
\add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.sum_s1  <= _133_;
always @(posedge \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.clk )
\add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.carry_s1  <= _132_;
assign _131_ = \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.ce  ? \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.b [4:2] : \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.bin_s1 ;
assign _130_ = \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.ce  ? \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.a [4:2] : \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.ain_s1 ;
assign _132_ = \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.ce  ? \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.facout_s1  : \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.carry_s1 ;
assign _133_ = \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.ce  ? \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.fas_s1  : \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.sum_s1 ;
assign _134_ = \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.u1.a  + \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.u1.b ;
assign { \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.u1.cout , \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.u1.s  } = _134_ + \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.u1.cin ;
assign _135_ = \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.u2.a  + \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.u2.b ;
assign { \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.u2.cout , \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.u2.s  } = _135_ + \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.u2.cin ;
always @(posedge \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.clk )
\add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.bin_s1  <= _137_;
always @(posedge \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.clk )
\add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.ain_s1  <= _136_;
always @(posedge \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.clk )
\add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.sum_s1  <= _139_;
always @(posedge \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.clk )
\add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.carry_s1  <= _138_;
assign _137_ = \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.ce  ? \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.b [5:3] : \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.bin_s1 ;
assign _136_ = \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.ce  ? \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.a [5:3] : \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.ain_s1 ;
assign _138_ = \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.ce  ? \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.facout_s1  : \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.carry_s1 ;
assign _139_ = \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.ce  ? \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.fas_s1  : \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.sum_s1 ;
assign _140_ = \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.u1.a  + \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.u1.b ;
assign { \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.u1.cout , \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.u1.s  } = _140_ + \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.u1.cin ;
assign _141_ = \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.u2.a  + \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.u2.b ;
assign { \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.u2.cout , \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.u2.s  } = _141_ + \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.u2.cin ;
always @(posedge \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.clk )
\add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.bin_s1  <= _143_;
always @(posedge \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.clk )
\add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.ain_s1  <= _142_;
always @(posedge \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.clk )
\add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.sum_s1  <= _145_;
always @(posedge \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.clk )
\add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.carry_s1  <= _144_;
assign _143_ = \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.ce  ? \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.b [5:3] : \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.bin_s1 ;
assign _142_ = \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.ce  ? \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.a [5:3] : \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.ain_s1 ;
assign _144_ = \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.ce  ? \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.facout_s1  : \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.carry_s1 ;
assign _145_ = \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.ce  ? \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.fas_s1  : \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.sum_s1 ;
assign _146_ = \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.u1.a  + \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.u1.b ;
assign { \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.u1.cout , \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.u1.s  } = _146_ + \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.u1.cin ;
assign _147_ = \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.u2.a  + \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.u2.b ;
assign { \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.u2.cout , \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.u2.s  } = _147_ + \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.u2.cin ;
always @(posedge \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.clk )
\add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.bin_s1  <= _149_;
always @(posedge \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.clk )
\add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.ain_s1  <= _148_;
always @(posedge \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.clk )
\add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.sum_s1  <= _151_;
always @(posedge \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.clk )
\add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.carry_s1  <= _150_;
assign _149_ = \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.ce  ? \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.b [5:3] : \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.bin_s1 ;
assign _148_ = \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.ce  ? \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.a [5:3] : \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.ain_s1 ;
assign _150_ = \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.ce  ? \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.facout_s1  : \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.carry_s1 ;
assign _151_ = \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.ce  ? \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.fas_s1  : \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.sum_s1 ;
assign _152_ = \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.u1.a  + \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.u1.b ;
assign { \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.u1.cout , \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.u1.s  } = _152_ + \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.u1.cin ;
assign _153_ = \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.u2.a  + \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.u2.b ;
assign { \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.u2.cout , \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.u2.s  } = _153_ + \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.u2.cin ;
always @(posedge \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.clk )
\add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.bin_s1  <= _155_;
always @(posedge \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.clk )
\add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.ain_s1  <= _154_;
always @(posedge \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.clk )
\add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.sum_s1  <= _157_;
always @(posedge \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.clk )
\add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.carry_s1  <= _156_;
assign _155_ = \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.ce  ? \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.b [5:3] : \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.bin_s1 ;
assign _154_ = \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.ce  ? \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.a [5:3] : \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.ain_s1 ;
assign _156_ = \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.ce  ? \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.facout_s1  : \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.carry_s1 ;
assign _157_ = \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.ce  ? \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.fas_s1  : \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.sum_s1 ;
assign _158_ = \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.u1.a  + \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.u1.b ;
assign { \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.u1.cout , \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.u1.s  } = _158_ + \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.u1.cin ;
assign _159_ = \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.u2.a  + \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.u2.b ;
assign { \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.u2.cout , \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.u2.s  } = _159_ + \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.u2.cin ;
always @(posedge \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.clk )
\add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.bin_s1  <= _161_;
always @(posedge \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.clk )
\add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.ain_s1  <= _160_;
always @(posedge \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.clk )
\add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.sum_s1  <= _163_;
always @(posedge \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.clk )
\add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.carry_s1  <= _162_;
assign _161_ = \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.ce  ? \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.b [5:3] : \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.bin_s1 ;
assign _160_ = \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.ce  ? \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.a [5:3] : \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.ain_s1 ;
assign _162_ = \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.ce  ? \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.facout_s1  : \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.carry_s1 ;
assign _163_ = \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.ce  ? \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.fas_s1  : \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.sum_s1 ;
assign _164_ = \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.u1.a  + \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.u1.b ;
assign { \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.u1.cout , \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.u1.s  } = _164_ + \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.u1.cin ;
assign _165_ = \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.u2.a  + \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.u2.b ;
assign { \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.u2.cout , \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.u2.s  } = _165_ + \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.u2.cin ;
assign \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.bin_s0  = ~ \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.b ;
always @(posedge \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.clk )
\sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.bin_s1  <= _167_;
always @(posedge \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.clk )
\sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.ain_s1  <= _166_;
always @(posedge \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.clk )
\sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.sum_s1  <= _169_;
always @(posedge \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.clk )
\sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.carry_s1  <= _168_;
assign _167_ = \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.ce  ? \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.bin_s0 [4:2] : \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.bin_s1 ;
assign _166_ = \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.ce  ? \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.a [4:2] : \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.ain_s1 ;
assign _168_ = \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.ce  ? \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.facout_s1  : \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.carry_s1 ;
assign _169_ = \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.ce  ? \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.fas_s1  : \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.sum_s1 ;
assign _170_ = \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.u1.a  + \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.u1.b ;
assign { \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.u1.cout , \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.u1.s  } = _170_ + \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.u1.cin ;
assign _171_ = \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.u2.a  + \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.u2.b ;
assign { \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.u2.cout , \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.u2.s  } = _171_ + \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.u2.cin ;
assign \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.bin_s0  = ~ \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.b ;
always @(posedge \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.clk )
\sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.bin_s1  <= _173_;
always @(posedge \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.clk )
\sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.ain_s1  <= _172_;
always @(posedge \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.clk )
\sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.sum_s1  <= _175_;
always @(posedge \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.clk )
\sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.carry_s1  <= _174_;
assign _173_ = \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.ce  ? \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.bin_s0 [8:4] : \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.bin_s1 ;
assign _172_ = \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.ce  ? \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.a [8:4] : \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.ain_s1 ;
assign _174_ = \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.ce  ? \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.facout_s1  : \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.carry_s1 ;
assign _175_ = \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.ce  ? \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.fas_s1  : \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.sum_s1 ;
assign _176_ = \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.u1.a  + \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.u1.b ;
assign { \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.u1.cout , \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.u1.s  } = _176_ + \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.u1.cin ;
assign _177_ = \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.u2.a  + \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.u2.b ;
assign { \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.u2.cout , \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.u2.s  } = _177_ + \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.u2.cin ;
assign _178_ = $signed(ret_V_19_reg_1157) > $signed({ 1'h0, ret_V_25_fu_665_p3 });
assign _179_ = | trunc_ln414_reg_999;
assign _180_ = | tmp_2_reg_1334;
assign _181_ = tmp_2_reg_1334 != 4'hf;
assign _182_ = | op_3[12:0];
assign _183_ = | op_14[4:0];
assign or_ln340_1_fu_897_p2 = underflow_1_reg_1364 | overflow_1_fu_892_p2;
assign or_ln340_2_fu_513_p2 = or_ln340_reg_1132 | neg_src_fu_508_p2;
assign or_ln340_fu_483_p2 = overflow_fu_477_p2 | and_ln786_reg_1104;
assign or_ln384_fu_876_p2 = xor_ln384_fu_871_p2 | p_Result_13_reg_1319;
assign or_ln388_fu_867_p2 = underflow_1_reg_1364 | newsignbit_reg_1326;
assign or_ln785_1_fu_843_p2 = newsignbit_reg_1326 | icmp_ln768_reg_1340;
assign or_ln785_2_fu_529_p2 = p_Result_10_reg_981 | and_ln785_fu_525_p2;
assign or_ln785_fu_467_p2 = xor_ln785_fu_462_p2 | p_Result_12_reg_1068;
assign or_ln786_fu_852_p2 = xor_ln786_fu_847_p2 | icmp_ln786_reg_1345;
assign ret_V_18_fu_432_p2 = op_3 | { op_1, 12'h000 };
assign ret_V_20_fu_239_p2 = $signed({ op_7, 2'h0 }) | $signed(op_2);
always @(posedge ap_clk)
select_ln69_reg_1309[5:2] <= 4'h0;
always @(posedge ap_clk)
xor_ln416_reg_1075 <= _063_;
always @(posedge ap_clk)
sext_ln850_reg_1277 <= _055_;
always @(posedge ap_clk)
select_ln340_reg_1142 <= _053_;
always @(posedge ap_clk)
ret_V_3_reg_1147 <= _048_;
always @(posedge ap_clk)
ret_V_28_reg_1380 <= _047_;
always @(posedge ap_clk)
select_ln1192_reg_1385 <= _052_;
always @(posedge ap_clk)
ret_V_27_reg_1289 <= _046_;
always @(posedge ap_clk)
ret_V_26_reg_1267 <= _045_;
always @(posedge ap_clk)
tmp_3_reg_1272 <= _057_;
always @(posedge ap_clk)
ret_V_20_reg_959 <= _040_;
always @(posedge ap_clk)
ret_V_4_cast_reg_964 <= _049_;
always @(posedge ap_clk)
trunc_ln851_1_reg_971 <= _060_;
always @(posedge ap_clk)
p_Val2_2_reg_1062 <= _036_;
always @(posedge ap_clk)
p_Result_12_reg_1068 <= _031_;
always @(posedge ap_clk)
or_ln785_1_reg_1358 <= _028_;
always @(posedge ap_clk)
underflow_1_reg_1364 <= _062_;
always @(posedge ap_clk)
op_5_V_reg_1152 <= _026_;
always @(posedge ap_clk)
ret_V_19_reg_1157 <= _039_;
always @(posedge ap_clk)
trunc_ln728_reg_1165 <= _059_;
always @(posedge ap_clk)
ret_V_24_reg_1232 <= _044_;
always @(posedge ap_clk)
op_22_V_reg_1242 <= _024_;
always @(posedge ap_clk)
p_Result_13_reg_1319 <= _032_;
always @(posedge ap_clk)
newsignbit_reg_1326 <= _023_;
always @(posedge ap_clk)
tmp_2_reg_1334 <= _056_;
always @(posedge ap_clk)
or_ln340_reg_1132 <= _027_;
always @(posedge ap_clk)
icmp_ln851_reg_1137 <= _021_;
always @(posedge ap_clk)
lhs_V_1_reg_1247 <= _022_;
always @(posedge ap_clk)
icmp_ln851_3_reg_1262 <= _020_;
always @(posedge ap_clk)
ret_V_17_reg_976 <= _037_;
always @(posedge ap_clk)
p_Result_10_reg_981 <= _029_;
always @(posedge ap_clk)
p_Val2_1_reg_989 <= _035_;
always @(posedge ap_clk)
p_Result_11_reg_994 <= _030_;
always @(posedge ap_clk)
trunc_ln414_reg_999 <= _058_;
always @(posedge ap_clk)
p_Result_s_reg_1004 <= _034_;
always @(posedge ap_clk)
p_Result_1_reg_1009 <= _033_;
always @(posedge ap_clk)
icmp_ln851_1_reg_1015 <= _018_;
always @(posedge ap_clk)
icmp_ln768_reg_1340 <= _016_;
always @(posedge ap_clk)
icmp_ln786_reg_1345 <= _017_;
always @(posedge ap_clk)
op_25_V_reg_1350 <= _025_;
always @(posedge ap_clk)
carry_1_reg_1081 <= _012_;
always @(posedge ap_clk)
empty_reg_1093 <= _014_;
always @(posedge ap_clk)
deleted_zeros_reg_1098 <= _013_;
always @(posedge ap_clk)
and_ln786_reg_1104 <= _010_;
always @(posedge ap_clk)
ret_V_18_reg_1110 <= _038_;
always @(posedge ap_clk)
ret_V_reg_1115 <= _051_;
always @(posedge ap_clk)
trunc_ln851_reg_1122 <= _061_;
always @(posedge ap_clk)
icmp_ln851_2_reg_1127 <= _019_;
always @(posedge ap_clk)
and_ln414_reg_1047 <= _009_;
always @(posedge ap_clk)
ret_V_21_reg_1052 <= _042_;
always @(posedge ap_clk)
and_ln384_reg_1370 <= _008_;
always @(posedge ap_clk)
ret_V_23_reg_1195 <= _043_;
always @(posedge ap_clk)
ret_V_21_cast_reg_1200 <= _041_;
always @(posedge ap_clk)
add_ln69_reg_1207 <= _007_;
always @(posedge ap_clk)
select_ln69_reg_1309[1:0] <= _054_;
always @(posedge ap_clk)
add_ln69_2_reg_1314 <= _006_;
always @(posedge ap_clk)
add_ln691_reg_1237 <= _005_;
always @(posedge ap_clk)
add_ln691_2_reg_1375 <= _004_;
always @(posedge ap_clk)
add_ln691_1_reg_1284 <= _003_;
always @(posedge ap_clk)
icmp_ln414_reg_1020 <= _015_;
always @(posedge ap_clk)
Range2_all_ones_reg_1025 <= _002_;
always @(posedge ap_clk)
Range1_all_ones_reg_1030 <= _000_;
always @(posedge ap_clk)
Range1_all_zeros_reg_1037 <= _001_;
always @(posedge ap_clk)
ret_V_6_reg_1042 <= _050_;
always @(posedge ap_clk)
ap_CS_fsm <= _011_;
assign _064_ = _069_ ? 2'h2 : 2'h1;
assign _184_ = ap_CS_fsm == 1'h1;
function [29:0] _536_;
input [29:0] a;
input [899:0] b;
input [29:0] s;
case (s)
30'b000000000000000000000000000001:
_536_ = b[29:0];
30'b000000000000000000000000000010:
_536_ = b[59:30];
30'b000000000000000000000000000100:
_536_ = b[89:60];
30'b000000000000000000000000001000:
_536_ = b[119:90];
30'b000000000000000000000000010000:
_536_ = b[149:120];
30'b000000000000000000000000100000:
_536_ = b[179:150];
30'b000000000000000000000001000000:
_536_ = b[209:180];
30'b000000000000000000000010000000:
_536_ = b[239:210];
30'b000000000000000000000100000000:
_536_ = b[269:240];
30'b000000000000000000001000000000:
_536_ = b[299:270];
30'b000000000000000000010000000000:
_536_ = b[329:300];
30'b000000000000000000100000000000:
_536_ = b[359:330];
30'b000000000000000001000000000000:
_536_ = b[389:360];
30'b000000000000000010000000000000:
_536_ = b[419:390];
30'b000000000000000100000000000000:
_536_ = b[449:420];
30'b000000000000001000000000000000:
_536_ = b[479:450];
30'b000000000000010000000000000000:
_536_ = b[509:480];
30'b000000000000100000000000000000:
_536_ = b[539:510];
30'b000000000001000000000000000000:
_536_ = b[569:540];
30'b000000000010000000000000000000:
_536_ = b[599:570];
30'b000000000100000000000000000000:
_536_ = b[629:600];
30'b000000001000000000000000000000:
_536_ = b[659:630];
30'b000000010000000000000000000000:
_536_ = b[689:660];
30'b000000100000000000000000000000:
_536_ = b[719:690];
30'b000001000000000000000000000000:
_536_ = b[749:720];
30'b000010000000000000000000000000:
_536_ = b[779:750];
30'b000100000000000000000000000000:
_536_ = b[809:780];
30'b001000000000000000000000000000:
_536_ = b[839:810];
30'b010000000000000000000000000000:
_536_ = b[869:840];
30'b100000000000000000000000000000:
_536_ = b[899:870];
30'b000000000000000000000000000000:
_536_ = a;
default:
_536_ = 30'bx;
endcase
endfunction
assign ap_NS_fsm = _536_(30'hxxxxxxxx, { 28'h0000000, _064_, 870'h00000004000000200000010000000800000040000002000000100000008000000400000020000001000000080000004000000200000010000000800000040000002000000100000008000000400000020000001000000080000004000000200000010000000800000000000001 }, { _184_, _213_, _212_, _211_, _210_, _209_, _208_, _207_, _206_, _205_, _204_, _203_, _202_, _201_, _200_, _199_, _198_, _197_, _196_, _195_, _194_, _193_, _192_, _191_, _190_, _189_, _188_, _187_, _186_, _185_ });
assign _185_ = ap_CS_fsm == 30'h20000000;
assign _186_ = ap_CS_fsm == 29'h10000000;
assign _187_ = ap_CS_fsm == 28'h8000000;
assign _188_ = ap_CS_fsm == 27'h4000000;
assign _189_ = ap_CS_fsm == 26'h2000000;
assign _190_ = ap_CS_fsm == 25'h1000000;
assign _191_ = ap_CS_fsm == 24'h800000;
assign _192_ = ap_CS_fsm == 23'h400000;
assign _193_ = ap_CS_fsm == 22'h200000;
assign _194_ = ap_CS_fsm == 21'h100000;
assign _195_ = ap_CS_fsm == 20'h80000;
assign _196_ = ap_CS_fsm == 19'h40000;
assign _197_ = ap_CS_fsm == 18'h20000;
assign _198_ = ap_CS_fsm == 17'h10000;
assign _199_ = ap_CS_fsm == 16'h8000;
assign _200_ = ap_CS_fsm == 15'h4000;
assign _201_ = ap_CS_fsm == 14'h2000;
assign _202_ = ap_CS_fsm == 13'h1000;
assign _203_ = ap_CS_fsm == 12'h800;
assign _204_ = ap_CS_fsm == 11'h400;
assign _205_ = ap_CS_fsm == 10'h200;
assign _206_ = ap_CS_fsm == 9'h100;
assign _207_ = ap_CS_fsm == 8'h80;
assign _208_ = ap_CS_fsm == 7'h40;
assign _209_ = ap_CS_fsm == 6'h20;
assign _210_ = ap_CS_fsm == 5'h10;
assign _211_ = ap_CS_fsm == 4'h8;
assign _212_ = ap_CS_fsm == 3'h4;
assign _213_ = ap_CS_fsm == 2'h2;
assign op_28_ap_vld = ap_CS_fsm[29] ? 1'h1 : 1'h0;
assign ap_idle = _068_ ? 1'h1 : 1'h0;
assign _063_ = ap_CS_fsm[6] ? xor_ln416_fu_378_p2 : xor_ln416_reg_1075;
assign _055_ = ap_CS_fsm[18] ? { tmp_3_reg_1272[4], tmp_3_reg_1272 } : sext_ln850_reg_1277;
assign _048_ = ap_CS_fsm[10] ? grp_fu_493_p2 : ret_V_3_reg_1147;
assign _053_ = ap_CS_fsm[10] ? select_ln340_fu_518_p3 : select_ln340_reg_1142;
assign _052_ = ap_CS_fsm[27] ? select_ln1192_fu_927_p3 : select_ln1192_reg_1385;
assign _047_ = ap_CS_fsm[27] ? ret_V_28_fu_920_p3 : ret_V_28_reg_1380;
assign _046_ = ap_CS_fsm[20] ? ret_V_27_fu_739_p3 : ret_V_27_reg_1289;
assign _057_ = ap_CS_fsm[17] ? grp_fu_692_p2[9:5] : tmp_3_reg_1272;
assign _045_ = ap_CS_fsm[17] ? grp_fu_692_p2 : ret_V_26_reg_1267;
assign _060_ = ap_CS_fsm[0] ? ret_V_20_fu_239_p2[1:0] : trunc_ln851_1_reg_971;
assign _049_ = ap_CS_fsm[0] ? ret_V_20_fu_239_p2[3:2] : ret_V_4_cast_reg_964;
assign _040_ = ap_CS_fsm[0] ? ret_V_20_fu_239_p2 : ret_V_20_reg_959;
assign _031_ = ap_CS_fsm[5] ? grp_fu_365_p2[1] : p_Result_12_reg_1068;
assign _036_ = ap_CS_fsm[5] ? grp_fu_365_p2 : p_Val2_2_reg_1062;
assign _062_ = ap_CS_fsm[25] ? underflow_1_fu_857_p2 : underflow_1_reg_1364;
assign _028_ = ap_CS_fsm[25] ? or_ln785_1_fu_843_p2 : or_ln785_1_reg_1358;
assign _059_ = ap_CS_fsm[11] ? ret_V_19_fu_557_p3[1:0] : trunc_ln728_reg_1165;
assign _039_ = ap_CS_fsm[11] ? ret_V_19_fu_557_p3 : ret_V_19_reg_1157;
assign _026_ = ap_CS_fsm[11] ? op_5_V_fu_539_p3 : op_5_V_reg_1152;
assign _024_ = ap_CS_fsm[15] ? grp_fu_647_p2 : op_22_V_reg_1242;
assign _044_ = ap_CS_fsm[15] ? grp_fu_633_p2 : ret_V_24_reg_1232;
assign _056_ = ap_CS_fsm[23] ? grp_fu_793_p2[4:1] : tmp_2_reg_1334;
assign _023_ = ap_CS_fsm[23] ? grp_fu_793_p2[0] : newsignbit_reg_1326;
assign _032_ = ap_CS_fsm[23] ? grp_fu_793_p2[4] : p_Result_13_reg_1319;
assign _021_ = ap_CS_fsm[9] ? icmp_ln851_fu_488_p2 : icmp_ln851_reg_1137;
assign _027_ = ap_CS_fsm[9] ? or_ln340_fu_483_p2 : or_ln340_reg_1132;
assign _020_ = ap_CS_fsm[16] ? icmp_ln851_3_fu_702_p2 : icmp_ln851_3_reg_1262;
assign _022_ = ap_CS_fsm[16] ? lhs_V_1_fu_676_p2 : lhs_V_1_reg_1247;
assign _018_ = ap_CS_fsm[1] ? icmp_ln851_1_fu_309_p2 : icmp_ln851_1_reg_1015;
assign _033_ = ap_CS_fsm[1] ? grp_fu_221_p2[8:4] : p_Result_1_reg_1009;
assign _034_ = ap_CS_fsm[1] ? grp_fu_221_p2[8:5] : p_Result_s_reg_1004;
assign _058_ = ap_CS_fsm[1] ? grp_fu_221_p2[1:0] : trunc_ln414_reg_999;
assign _030_ = ap_CS_fsm[1] ? grp_fu_221_p2[3] : p_Result_11_reg_994;
assign _035_ = ap_CS_fsm[1] ? grp_fu_221_p2[3:2] : p_Val2_1_reg_989;
assign _029_ = ap_CS_fsm[1] ? grp_fu_221_p2[8] : p_Result_10_reg_981;
assign _037_ = ap_CS_fsm[1] ? grp_fu_221_p2 : ret_V_17_reg_976;
assign _025_ = ap_CS_fsm[24] ? grp_fu_829_p2 : op_25_V_reg_1350;
assign _017_ = ap_CS_fsm[24] ? icmp_ln786_fu_838_p2 : icmp_ln786_reg_1345;
assign _016_ = ap_CS_fsm[24] ? icmp_ln768_fu_833_p2 : icmp_ln768_reg_1340;
assign _012_ = ap_CS_fsm[7] ? carry_1_fu_383_p2 : carry_1_reg_1081;
assign _019_ = ap_CS_fsm[8] ? icmp_ln851_2_fu_456_p2 : icmp_ln851_2_reg_1127;
assign _061_ = ap_CS_fsm[8] ? ret_V_18_fu_432_p2[12:0] : trunc_ln851_reg_1122;
assign _051_ = ap_CS_fsm[8] ? ret_V_18_fu_432_p2[15:13] : ret_V_reg_1115;
assign _038_ = ap_CS_fsm[8] ? ret_V_18_fu_432_p2 : ret_V_18_reg_1110;
assign _010_ = ap_CS_fsm[8] ? and_ln786_fu_420_p2 : and_ln786_reg_1104;
assign _013_ = ap_CS_fsm[8] ? deleted_zeros_fu_391_p3 : deleted_zeros_reg_1098;
assign _014_ = ap_CS_fsm[8] ? op_3[14:0] : empty_reg_1093;
assign _042_ = ap_CS_fsm[3] ? ret_V_21_fu_355_p3 : ret_V_21_reg_1052;
assign _009_ = ap_CS_fsm[3] ? and_ln414_fu_339_p2 : and_ln414_reg_1047;
assign _008_ = ap_CS_fsm[26] ? and_ln384_fu_881_p2 : and_ln384_reg_1370;
assign _007_ = ap_CS_fsm[13] ? grp_fu_600_p2 : add_ln69_reg_1207;
assign _041_ = ap_CS_fsm[13] ? grp_fu_591_p2[14:13] : ret_V_21_cast_reg_1200;
assign _043_ = ap_CS_fsm[13] ? grp_fu_578_p2 : ret_V_23_reg_1195;
assign _006_ = ap_CS_fsm[22] ? grp_fu_749_p2 : add_ln69_2_reg_1314;
assign _054_ = ap_CS_fsm[22] ? select_ln69_fu_799_p3 : select_ln69_reg_1309[1:0];
assign _005_ = _067_ ? grp_fu_639_p2 : add_ln691_reg_1237;
assign _004_ = _066_ ? grp_fu_862_p2 : add_ln691_2_reg_1375;
assign _003_ = _065_ ? grp_fu_721_p2 : add_ln691_1_reg_1284;
assign _050_ = ap_CS_fsm[2] ? grp_fu_314_p2 : ret_V_6_reg_1042;
assign _001_ = ap_CS_fsm[2] ? Range1_all_zeros_fu_334_p2 : Range1_all_zeros_reg_1037;
assign _000_ = ap_CS_fsm[2] ? Range1_all_ones_fu_329_p2 : Range1_all_ones_reg_1030;
assign _002_ = ap_CS_fsm[2] ? Range2_all_ones_fu_324_p2 : Range2_all_ones_reg_1025;
assign _015_ = ap_CS_fsm[2] ? icmp_ln414_fu_319_p2 : icmp_ln414_reg_1020;
assign _011_ = ap_rst ? 30'h00000001 : ap_NS_fsm;
assign Range1_all_ones_fu_329_p2 = _071_ ? 1'h1 : 1'h0;
assign Range1_all_zeros_fu_334_p2 = _072_ ? 1'h1 : 1'h0;
assign Range2_all_ones_fu_324_p2 = _073_ ? 1'h1 : 1'h0;
assign deleted_ones_fu_414_p3 = carry_1_reg_1081 ? and_ln780_fu_409_p2 : Range1_all_ones_reg_1030;
assign deleted_zeros_fu_391_p3 = carry_1_reg_1081 ? Range1_all_ones_reg_1030 : Range1_all_zeros_reg_1037;
assign icmp_ln414_fu_319_p2 = _179_ ? 1'h1 : 1'h0;
assign icmp_ln768_fu_833_p2 = _180_ ? 1'h1 : 1'h0;
assign icmp_ln786_fu_838_p2 = _181_ ? 1'h1 : 1'h0;
assign icmp_ln851_1_fu_309_p2 = _074_ ? 1'h1 : 1'h0;
assign icmp_ln851_2_fu_456_p2 = _182_ ? 1'h1 : 1'h0;
assign icmp_ln851_3_fu_702_p2 = _183_ ? 1'h1 : 1'h0;
assign icmp_ln851_fu_488_p2 = _075_ ? 1'h1 : 1'h0;
assign lhs_V_1_fu_676_p2 = _178_ ? 1'h1 : 1'h0;
assign op_19_V_fu_902_p3 = or_ln340_1_fu_897_p2 ? and_ln384_reg_1370 : newsignbit_reg_1326;
assign op_5_V_fu_539_p3 = and_ln785_1_fu_534_p2 ? p_Val2_2_reg_1062 : select_ln340_reg_1142;
assign ret_V_19_fu_557_p3 = ret_V_18_reg_1110[15] ? select_ln850_fu_552_p3 : ret_V_reg_1115;
assign ret_V_21_fu_355_p3 = ret_V_20_reg_959[7] ? select_ln850_1_fu_350_p3 : ret_V_4_cast_reg_964;
assign ret_V_25_fu_665_p3 = ret_V_24_reg_1232[16] ? select_ln850_2_fu_660_p3 : ret_V_21_cast_reg_1200;
assign ret_V_27_fu_739_p3 = ret_V_26_reg_1267[9] ? select_ln850_3_fu_734_p3 : sext_ln850_reg_1277;
assign ret_V_28_fu_920_p3 = op_25_V_reg_1350[5] ? select_ln850_4_fu_915_p3 : { 1'h0, op_25_V_reg_1350[4:0] };
assign select_ln1192_fu_927_p3 = op_19_V_fu_902_p3 ? 6'h3f : 6'h00;
assign select_ln340_fu_518_p3 = or_ln340_2_fu_513_p2 ? 2'h0 : p_Val2_2_reg_1062;
assign select_ln69_fu_799_p3 = ret_V_22_fu_780_p2 ? 2'h2 : 2'h1;
assign select_ln850_1_fu_350_p3 = icmp_ln851_1_reg_1015 ? ret_V_4_cast_reg_964 : ret_V_6_reg_1042;
assign select_ln850_2_fu_660_p3 = icmp_ln851_2_reg_1127 ? add_ln691_reg_1237 : ret_V_21_cast_reg_1200;
assign select_ln850_3_fu_734_p3 = icmp_ln851_3_reg_1262 ? add_ln691_1_reg_1284 : sext_ln850_reg_1277;
assign select_ln850_4_fu_915_p3 = lhs_V_1_reg_1247 ? add_ln691_2_reg_1375 : { 1'h1, op_25_V_reg_1350[4:0] };
assign select_ln850_fu_552_p3 = icmp_ln851_reg_1137 ? ret_V_reg_1115 : ret_V_3_reg_1147;
assign ret_V_22_fu_780_p2 = op_8[1] ^ and_ln850_fu_774_p2;
assign ap_CS_fsm_state1 = ap_CS_fsm[0];
assign ap_CS_fsm_state10 = ap_CS_fsm[9];
assign ap_CS_fsm_state11 = ap_CS_fsm[10];
assign ap_CS_fsm_state12 = ap_CS_fsm[11];
assign ap_CS_fsm_state13 = ap_CS_fsm[12];
assign ap_CS_fsm_state14 = ap_CS_fsm[13];
assign ap_CS_fsm_state15 = ap_CS_fsm[14];
assign ap_CS_fsm_state16 = ap_CS_fsm[15];
assign ap_CS_fsm_state17 = ap_CS_fsm[16];
assign ap_CS_fsm_state18 = ap_CS_fsm[17];
assign ap_CS_fsm_state19 = ap_CS_fsm[18];
assign ap_CS_fsm_state2 = ap_CS_fsm[1];
assign ap_CS_fsm_state20 = ap_CS_fsm[19];
assign ap_CS_fsm_state21 = ap_CS_fsm[20];
assign ap_CS_fsm_state22 = ap_CS_fsm[21];
assign ap_CS_fsm_state23 = ap_CS_fsm[22];
assign ap_CS_fsm_state24 = ap_CS_fsm[23];
assign ap_CS_fsm_state25 = ap_CS_fsm[24];
assign ap_CS_fsm_state26 = ap_CS_fsm[25];
assign ap_CS_fsm_state27 = ap_CS_fsm[26];
assign ap_CS_fsm_state28 = ap_CS_fsm[27];
assign ap_CS_fsm_state29 = ap_CS_fsm[28];
assign ap_CS_fsm_state3 = ap_CS_fsm[2];
assign ap_CS_fsm_state30 = ap_CS_fsm[29];
assign ap_CS_fsm_state4 = ap_CS_fsm[3];
assign ap_CS_fsm_state5 = ap_CS_fsm[4];
assign ap_CS_fsm_state6 = ap_CS_fsm[5];
assign ap_CS_fsm_state7 = ap_CS_fsm[6];
assign ap_CS_fsm_state8 = ap_CS_fsm[7];
assign ap_CS_fsm_state9 = ap_CS_fsm[8];
assign ap_done = op_28_ap_vld;
assign ap_ready = op_28_ap_vld;
assign empty_fu_387_p0 = op_3;
assign empty_fu_387_p1 = op_3[14:0];
assign grp_fu_221_p0 = { op_1[3], op_1[3], op_1[3], op_1[3], op_1, 1'h0 };
assign grp_fu_221_p1 = { op_2[7], op_2 };
assign grp_fu_365_p1 = { 1'h0, and_ln414_reg_1047 };
assign grp_fu_578_p0 = { op_5_V_reg_1152[1], op_5_V_reg_1152 };
assign grp_fu_578_p1 = { op_0[1], op_0 };
assign grp_fu_591_p0 = { trunc_ln728_reg_1165, 13'h0000 };
assign grp_fu_600_p0 = { ret_V_19_reg_1157[2], ret_V_19_reg_1157 };
assign grp_fu_600_p1 = { 2'h0, op_12 };
assign grp_fu_633_p0 = { ret_V_19_reg_1157[2], ret_V_19_reg_1157, 13'h0000 };
assign grp_fu_633_p1 = { op_3[15], op_3 };
assign grp_fu_647_p0 = { add_ln69_reg_1207[3], add_ln69_reg_1207 };
assign grp_fu_647_p1 = { ret_V_23_reg_1195[2], ret_V_23_reg_1195[2], ret_V_23_reg_1195 };
assign grp_fu_692_p0 = { op_22_V_reg_1242, 5'h00 };
assign grp_fu_692_p1 = { op_14[7], op_14[7], op_14 };
assign grp_fu_721_p0 = { tmp_3_reg_1272[4], tmp_3_reg_1272 };
assign grp_fu_749_p1 = { ret_V_21_reg_1052[1], ret_V_21_reg_1052[1], ret_V_21_reg_1052[1], ret_V_21_reg_1052[1], ret_V_21_reg_1052 };
assign grp_fu_793_p0 = { ret_V_19_reg_1157[2], ret_V_19_reg_1157[2], ret_V_19_reg_1157 };
assign grp_fu_793_p1 = { op_13[3], op_13 };
assign lhs_1_fu_425_p3 = { op_1, 12'h000 };
assign lhs_fu_205_p3 = { op_1, 1'h0 };
assign newsignbit_fu_815_p1 = grp_fu_793_p2[0];
assign op_28 = { grp_fu_935_p2[5], grp_fu_935_p2[5], grp_fu_935_p2[5], grp_fu_935_p2[5], grp_fu_935_p2[5], grp_fu_935_p2[5], grp_fu_935_p2[5], grp_fu_935_p2[5], grp_fu_935_p2[5], grp_fu_935_p2[5], grp_fu_935_p2[5], grp_fu_935_p2[5], grp_fu_935_p2[5], grp_fu_935_p2[5], grp_fu_935_p2[5], grp_fu_935_p2[5], grp_fu_935_p2[5], grp_fu_935_p2[5], grp_fu_935_p2[5], grp_fu_935_p2[5], grp_fu_935_p2[5], grp_fu_935_p2[5], grp_fu_935_p2[5], grp_fu_935_p2[5], grp_fu_935_p2[5], grp_fu_935_p2[5], grp_fu_935_p2 };
assign p_Result_2_fu_343_p3 = ret_V_20_reg_959[7];
assign p_Result_3_fu_762_p3 = op_8[1];
assign p_Result_5_fu_653_p3 = ret_V_24_reg_1232[16];
assign p_Result_8_fu_727_p3 = ret_V_26_reg_1267[9];
assign p_Result_9_fu_908_p3 = op_25_V_reg_1350[5];
assign p_Result_s_16_fu_545_p3 = ret_V_18_reg_1110[15];
assign ret_V_18_fu_432_p1 = op_3;
assign ret_V_20_fu_239_p1 = op_2;
assign ret_V_8_fu_754_p3 = op_8[1];
assign rhs_3_fu_622_p3 = { ret_V_19_reg_1157, 13'h0000 };
assign rhs_fu_227_p3 = { op_7, 2'h0 };
assign sext_ln1192_2_fu_681_p0 = op_14;
assign sext_ln1192_fu_619_p0 = op_3;
assign sext_ln1195_fu_235_p1 = { op_7[1], op_7[1], op_7[1], op_7[1], op_7, 2'h0 };
assign sext_ln703_fu_217_p0 = op_2;
assign sext_ln850_fu_718_p1 = { tmp_3_reg_1272[4], tmp_3_reg_1272 };
assign tmp_fu_396_p3 = ret_V_17_reg_976[4];
assign trunc_ln414_fu_285_p1 = grp_fu_221_p2[1:0];
assign trunc_ln728_fu_564_p1 = ret_V_19_fu_557_p3[1:0];
assign trunc_ln851_1_fu_255_p1 = ret_V_20_fu_239_p2[1:0];
assign trunc_ln851_2_fu_770_p1 = op_8[0];
assign trunc_ln851_3_fu_452_p0 = op_3;
assign trunc_ln851_3_fu_452_p1 = op_3[12:0];
assign trunc_ln851_4_fu_698_p0 = op_14;
assign trunc_ln851_4_fu_698_p1 = op_14[4:0];
assign trunc_ln851_fu_448_p1 = ret_V_18_fu_432_p2[12:0];
assign zext_ln886_fu_672_p1 = { 1'h0, ret_V_25_fu_665_p3 };
assign \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.ain_s0  = \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.a ;
assign \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.s  = { \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.fas_s2 , \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.sum_s1  };
assign \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.u2.a  = \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.ain_s1 ;
assign \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.u2.b  = \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.bin_s1 ;
assign \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.u2.cin  = \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.carry_s1 ;
assign \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.facout_s2  = \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.u2.cout ;
assign \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.fas_s2  = \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.u2.s ;
assign \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.u1.a  = \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.a [3:0];
assign \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.u1.b  = \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.bin_s0 [3:0];
assign \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.u1.cin  = 1'h1;
assign \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.facout_s1  = \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.u1.cout ;
assign \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.fas_s1  = \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.u1.s ;
assign \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.a  = \sub_9s_9s_9_2_1_U1.din0 ;
assign \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.b  = \sub_9s_9s_9_2_1_U1.din1 ;
assign \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.ce  = \sub_9s_9s_9_2_1_U1.ce ;
assign \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.clk  = \sub_9s_9s_9_2_1_U1.clk ;
assign \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.reset  = \sub_9s_9s_9_2_1_U1.reset ;
assign \sub_9s_9s_9_2_1_U1.dout  = \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.s ;
assign \sub_9s_9s_9_2_1_U1.ce  = 1'h1;
assign \sub_9s_9s_9_2_1_U1.clk  = ap_clk;
assign \sub_9s_9s_9_2_1_U1.din0  = { op_1[3], op_1[3], op_1[3], op_1[3], op_1, 1'h0 };
assign \sub_9s_9s_9_2_1_U1.din1  = { op_2[7], op_2 };
assign grp_fu_221_p2 = \sub_9s_9s_9_2_1_U1.dout ;
assign \sub_9s_9s_9_2_1_U1.reset  = ap_rst;
assign \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.ain_s0  = \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.a ;
assign \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.s  = { \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.fas_s2 , \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.sum_s1  };
assign \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.u2.a  = \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.ain_s1 ;
assign \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.u2.b  = \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.bin_s1 ;
assign \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.u2.cin  = \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.carry_s1 ;
assign \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.facout_s2  = \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.u2.cout ;
assign \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.fas_s2  = \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.u2.s ;
assign \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.u1.a  = \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.a [1:0];
assign \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.u1.b  = \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.bin_s0 [1:0];
assign \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.u1.cin  = 1'h1;
assign \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.facout_s1  = \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.u1.cout ;
assign \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.fas_s1  = \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.u1.s ;
assign \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.a  = \sub_5s_5s_5_2_1_U14.din0 ;
assign \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.b  = \sub_5s_5s_5_2_1_U14.din1 ;
assign \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.ce  = \sub_5s_5s_5_2_1_U14.ce ;
assign \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.clk  = \sub_5s_5s_5_2_1_U14.clk ;
assign \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.reset  = \sub_5s_5s_5_2_1_U14.reset ;
assign \sub_5s_5s_5_2_1_U14.dout  = \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.s ;
assign \sub_5s_5s_5_2_1_U14.ce  = 1'h1;
assign \sub_5s_5s_5_2_1_U14.clk  = ap_clk;
assign \sub_5s_5s_5_2_1_U14.din0  = { ret_V_19_reg_1157[2], ret_V_19_reg_1157[2], ret_V_19_reg_1157 };
assign \sub_5s_5s_5_2_1_U14.din1  = { op_13[3], op_13 };
assign grp_fu_793_p2 = \sub_5s_5s_5_2_1_U14.dout ;
assign \sub_5s_5s_5_2_1_U14.reset  = ap_rst;
assign \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.ain_s0  = \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.a ;
assign \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.bin_s0  = \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.b ;
assign \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.s  = { \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.fas_s2 , \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.sum_s1  };
assign \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.u2.a  = \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.ain_s1 ;
assign \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.u2.b  = \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.bin_s1 ;
assign \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.u2.cin  = \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.carry_s1 ;
assign \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.facout_s2  = \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.u2.cout ;
assign \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.fas_s2  = \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.u2.s ;
assign \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.u1.a  = \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.a [2:0];
assign \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.u1.b  = \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.b [2:0];
assign \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.u1.cin  = 1'h0;
assign \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.facout_s1  = \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.u1.cout ;
assign \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.fas_s1  = \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.u1.s ;
assign \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.a  = \add_6s_6ns_6_2_1_U12.din0 ;
assign \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.b  = \add_6s_6ns_6_2_1_U12.din1 ;
assign \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.ce  = \add_6s_6ns_6_2_1_U12.ce ;
assign \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.clk  = \add_6s_6ns_6_2_1_U12.clk ;
assign \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.reset  = \add_6s_6ns_6_2_1_U12.reset ;
assign \add_6s_6ns_6_2_1_U12.dout  = \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.s ;
assign \add_6s_6ns_6_2_1_U12.ce  = 1'h1;
assign \add_6s_6ns_6_2_1_U12.clk  = ap_clk;
assign \add_6s_6ns_6_2_1_U12.din0  = { tmp_3_reg_1272[4], tmp_3_reg_1272 };
assign \add_6s_6ns_6_2_1_U12.din1  = 6'h01;
assign grp_fu_721_p2 = \add_6s_6ns_6_2_1_U12.dout ;
assign \add_6s_6ns_6_2_1_U12.reset  = ap_rst;
assign \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.ain_s0  = \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.a ;
assign \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.bin_s0  = \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.b ;
assign \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.s  = { \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.fas_s2 , \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.sum_s1  };
assign \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.u2.a  = \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.ain_s1 ;
assign \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.u2.b  = \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.bin_s1 ;
assign \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.u2.cin  = \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.carry_s1 ;
assign \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.facout_s2  = \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.u2.cout ;
assign \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.fas_s2  = \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.u2.s ;
assign \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.u1.a  = \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.a [2:0];
assign \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.u1.b  = \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.b [2:0];
assign \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.u1.cin  = 1'h0;
assign \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.facout_s1  = \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.u1.cout ;
assign \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.fas_s1  = \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.u1.s ;
assign \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.a  = \add_6ns_6s_6_2_1_U13.din0 ;
assign \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.b  = \add_6ns_6s_6_2_1_U13.din1 ;
assign \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.ce  = \add_6ns_6s_6_2_1_U13.ce ;
assign \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.clk  = \add_6ns_6s_6_2_1_U13.clk ;
assign \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.reset  = \add_6ns_6s_6_2_1_U13.reset ;
assign \add_6ns_6s_6_2_1_U13.dout  = \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.s ;
assign \add_6ns_6s_6_2_1_U13.ce  = 1'h1;
assign \add_6ns_6s_6_2_1_U13.clk  = ap_clk;
assign \add_6ns_6s_6_2_1_U13.din0  = ret_V_27_reg_1289;
assign \add_6ns_6s_6_2_1_U13.din1  = { ret_V_21_reg_1052[1], ret_V_21_reg_1052[1], ret_V_21_reg_1052[1], ret_V_21_reg_1052[1], ret_V_21_reg_1052 };
assign grp_fu_749_p2 = \add_6ns_6s_6_2_1_U13.dout ;
assign \add_6ns_6s_6_2_1_U13.reset  = ap_rst;
assign \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.ain_s0  = \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.a ;
assign \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.bin_s0  = \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.b ;
assign \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.s  = { \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.fas_s2 , \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.sum_s1  };
assign \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.u2.a  = \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.ain_s1 ;
assign \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.u2.b  = \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.bin_s1 ;
assign \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.u2.cin  = \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.carry_s1 ;
assign \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.facout_s2  = \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.u2.cout ;
assign \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.fas_s2  = \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.u2.s ;
assign \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.u1.a  = \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.a [2:0];
assign \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.u1.b  = \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.b [2:0];
assign \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.u1.cin  = 1'h0;
assign \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.facout_s1  = \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.u1.cout ;
assign \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.fas_s1  = \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.u1.s ;
assign \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.a  = \add_6ns_6ns_6_2_1_U17.din0 ;
assign \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.b  = \add_6ns_6ns_6_2_1_U17.din1 ;
assign \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.ce  = \add_6ns_6ns_6_2_1_U17.ce ;
assign \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.clk  = \add_6ns_6ns_6_2_1_U17.clk ;
assign \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.reset  = \add_6ns_6ns_6_2_1_U17.reset ;
assign \add_6ns_6ns_6_2_1_U17.dout  = \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.s ;
assign \add_6ns_6ns_6_2_1_U17.ce  = 1'h1;
assign \add_6ns_6ns_6_2_1_U17.clk  = ap_clk;
assign \add_6ns_6ns_6_2_1_U17.din0  = ret_V_28_reg_1380;
assign \add_6ns_6ns_6_2_1_U17.din1  = select_ln1192_reg_1385;
assign grp_fu_935_p2 = \add_6ns_6ns_6_2_1_U17.dout ;
assign \add_6ns_6ns_6_2_1_U17.reset  = ap_rst;
assign \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.ain_s0  = \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.a ;
assign \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.bin_s0  = \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.b ;
assign \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.s  = { \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.fas_s2 , \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.sum_s1  };
assign \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.u2.a  = \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.ain_s1 ;
assign \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.u2.b  = \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.bin_s1 ;
assign \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.u2.cin  = \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.carry_s1 ;
assign \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.facout_s2  = \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.u2.cout ;
assign \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.fas_s2  = \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.u2.s ;
assign \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.u1.a  = \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.a [2:0];
assign \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.u1.b  = \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.b [2:0];
assign \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.u1.cin  = 1'h0;
assign \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.facout_s1  = \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.u1.cout ;
assign \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.fas_s1  = \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.u1.s ;
assign \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.a  = \add_6ns_6ns_6_2_1_U16.din0 ;
assign \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.b  = \add_6ns_6ns_6_2_1_U16.din1 ;
assign \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.ce  = \add_6ns_6ns_6_2_1_U16.ce ;
assign \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.clk  = \add_6ns_6ns_6_2_1_U16.clk ;
assign \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.reset  = \add_6ns_6ns_6_2_1_U16.reset ;
assign \add_6ns_6ns_6_2_1_U16.dout  = \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.s ;
assign \add_6ns_6ns_6_2_1_U16.ce  = 1'h1;
assign \add_6ns_6ns_6_2_1_U16.clk  = ap_clk;
assign \add_6ns_6ns_6_2_1_U16.din0  = op_25_V_reg_1350;
assign \add_6ns_6ns_6_2_1_U16.din1  = 6'h01;
assign grp_fu_862_p2 = \add_6ns_6ns_6_2_1_U16.dout ;
assign \add_6ns_6ns_6_2_1_U16.reset  = ap_rst;
assign \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.ain_s0  = \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.a ;
assign \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.bin_s0  = \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.b ;
assign \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.s  = { \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.fas_s2 , \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.sum_s1  };
assign \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.u2.a  = \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.ain_s1 ;
assign \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.u2.b  = \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.bin_s1 ;
assign \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.u2.cin  = \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.carry_s1 ;
assign \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.facout_s2  = \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.u2.cout ;
assign \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.fas_s2  = \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.u2.s ;
assign \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.u1.a  = \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.a [2:0];
assign \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.u1.b  = \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.b [2:0];
assign \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.u1.cin  = 1'h0;
assign \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.facout_s1  = \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.u1.cout ;
assign \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.fas_s1  = \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.u1.s ;
assign \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.a  = \add_6ns_6ns_6_2_1_U15.din0 ;
assign \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.b  = \add_6ns_6ns_6_2_1_U15.din1 ;
assign \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.ce  = \add_6ns_6ns_6_2_1_U15.ce ;
assign \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.clk  = \add_6ns_6ns_6_2_1_U15.clk ;
assign \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.reset  = \add_6ns_6ns_6_2_1_U15.reset ;
assign \add_6ns_6ns_6_2_1_U15.dout  = \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.s ;
assign \add_6ns_6ns_6_2_1_U15.ce  = 1'h1;
assign \add_6ns_6ns_6_2_1_U15.clk  = ap_clk;
assign \add_6ns_6ns_6_2_1_U15.din0  = add_ln69_2_reg_1314;
assign \add_6ns_6ns_6_2_1_U15.din1  = select_ln69_reg_1309;
assign grp_fu_829_p2 = \add_6ns_6ns_6_2_1_U15.dout ;
assign \add_6ns_6ns_6_2_1_U15.reset  = ap_rst;
assign \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.ain_s0  = \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.a ;
assign \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.bin_s0  = \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.b ;
assign \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.s  = { \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.fas_s2 , \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.sum_s1  };
assign \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.u2.a  = \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.ain_s1 ;
assign \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.u2.b  = \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.bin_s1 ;
assign \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.u2.cin  = \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.carry_s1 ;
assign \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.facout_s2  = \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.u2.cout ;
assign \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.fas_s2  = \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.u2.s ;
assign \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.u1.a  = \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.a [1:0];
assign \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.u1.b  = \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.b [1:0];
assign \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.u1.cin  = 1'h0;
assign \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.facout_s1  = \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.u1.cout ;
assign \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.fas_s1  = \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.u1.s ;
assign \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.a  = \add_5s_5s_5_2_1_U10.din0 ;
assign \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.b  = \add_5s_5s_5_2_1_U10.din1 ;
assign \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.ce  = \add_5s_5s_5_2_1_U10.ce ;
assign \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.clk  = \add_5s_5s_5_2_1_U10.clk ;
assign \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.reset  = \add_5s_5s_5_2_1_U10.reset ;
assign \add_5s_5s_5_2_1_U10.dout  = \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.s ;
assign \add_5s_5s_5_2_1_U10.ce  = 1'h1;
assign \add_5s_5s_5_2_1_U10.clk  = ap_clk;
assign \add_5s_5s_5_2_1_U10.din0  = { add_ln69_reg_1207[3], add_ln69_reg_1207 };
assign \add_5s_5s_5_2_1_U10.din1  = { ret_V_23_reg_1195[2], ret_V_23_reg_1195[2], ret_V_23_reg_1195 };
assign grp_fu_647_p2 = \add_5s_5s_5_2_1_U10.dout ;
assign \add_5s_5s_5_2_1_U10.reset  = ap_rst;
assign \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.ain_s0  = \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.a ;
assign \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.bin_s0  = \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.b ;
assign \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.s  = { \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.fas_s2 , \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.sum_s1  };
assign \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.u2.a  = \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.ain_s1 ;
assign \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.u2.b  = \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.bin_s1 ;
assign \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.u2.cin  = \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.carry_s1 ;
assign \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.facout_s2  = \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.u2.cout ;
assign \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.fas_s2  = \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.u2.s ;
assign \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.u1.a  = \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.a [1:0];
assign \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.u1.b  = \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.b [1:0];
assign \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.u1.cin  = 1'h0;
assign \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.facout_s1  = \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.u1.cout ;
assign \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.fas_s1  = \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.u1.s ;
assign \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.a  = \add_4s_4ns_4_2_1_U7.din0 ;
assign \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.b  = \add_4s_4ns_4_2_1_U7.din1 ;
assign \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.ce  = \add_4s_4ns_4_2_1_U7.ce ;
assign \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.clk  = \add_4s_4ns_4_2_1_U7.clk ;
assign \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.reset  = \add_4s_4ns_4_2_1_U7.reset ;
assign \add_4s_4ns_4_2_1_U7.dout  = \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.s ;
assign \add_4s_4ns_4_2_1_U7.ce  = 1'h1;
assign \add_4s_4ns_4_2_1_U7.clk  = ap_clk;
assign \add_4s_4ns_4_2_1_U7.din0  = { ret_V_19_reg_1157[2], ret_V_19_reg_1157 };
assign \add_4s_4ns_4_2_1_U7.din1  = { 2'h0, op_12 };
assign grp_fu_600_p2 = \add_4s_4ns_4_2_1_U7.dout ;
assign \add_4s_4ns_4_2_1_U7.reset  = ap_rst;
assign \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.ain_s0  = \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.a ;
assign \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.bin_s0  = \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.b ;
assign \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.s  = { \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.fas_s2 , \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.sum_s1  };
assign \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.u2.a  = \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.ain_s1 ;
assign \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.u2.b  = \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.bin_s1 ;
assign \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.u2.cin  = \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.carry_s1 ;
assign \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.facout_s2  = \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.u2.cout ;
assign \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.fas_s2  = \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.u2.s ;
assign \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.u1.a  = \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.a [0];
assign \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.u1.b  = \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.b [0];
assign \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.u1.cin  = 1'h0;
assign \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.facout_s1  = \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.u1.cout ;
assign \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.fas_s1  = \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.u1.s ;
assign \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.a  = \add_3s_3s_3_2_1_U5.din0 ;
assign \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.b  = \add_3s_3s_3_2_1_U5.din1 ;
assign \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.ce  = \add_3s_3s_3_2_1_U5.ce ;
assign \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.clk  = \add_3s_3s_3_2_1_U5.clk ;
assign \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.reset  = \add_3s_3s_3_2_1_U5.reset ;
assign \add_3s_3s_3_2_1_U5.dout  = \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.s ;
assign \add_3s_3s_3_2_1_U5.ce  = 1'h1;
assign \add_3s_3s_3_2_1_U5.clk  = ap_clk;
assign \add_3s_3s_3_2_1_U5.din0  = { op_5_V_reg_1152[1], op_5_V_reg_1152 };
assign \add_3s_3s_3_2_1_U5.din1  = { op_0[1], op_0 };
assign grp_fu_578_p2 = \add_3s_3s_3_2_1_U5.dout ;
assign \add_3s_3s_3_2_1_U5.reset  = ap_rst;
assign \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.ain_s0  = \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.a ;
assign \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.bin_s0  = \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.b ;
assign \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.s  = { \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.fas_s2 , \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.sum_s1  };
assign \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.u2.a  = \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.ain_s1 ;
assign \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.u2.b  = \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.bin_s1 ;
assign \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.u2.cin  = \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.carry_s1 ;
assign \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.facout_s2  = \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.u2.cout ;
assign \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.fas_s2  = \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.u2.s ;
assign \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.u1.a  = \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.a [0];
assign \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.u1.b  = \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.b [0];
assign \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.u1.cin  = 1'h0;
assign \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.facout_s1  = \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.u1.cout ;
assign \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.fas_s1  = \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.u1.s ;
assign \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.a  = \add_3ns_3ns_3_2_1_U4.din0 ;
assign \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.b  = \add_3ns_3ns_3_2_1_U4.din1 ;
assign \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.ce  = \add_3ns_3ns_3_2_1_U4.ce ;
assign \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.clk  = \add_3ns_3ns_3_2_1_U4.clk ;
assign \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.reset  = \add_3ns_3ns_3_2_1_U4.reset ;
assign \add_3ns_3ns_3_2_1_U4.dout  = \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.s ;
assign \add_3ns_3ns_3_2_1_U4.ce  = 1'h1;
assign \add_3ns_3ns_3_2_1_U4.clk  = ap_clk;
assign \add_3ns_3ns_3_2_1_U4.din0  = ret_V_reg_1115;
assign \add_3ns_3ns_3_2_1_U4.din1  = 3'h1;
assign grp_fu_493_p2 = \add_3ns_3ns_3_2_1_U4.dout ;
assign \add_3ns_3ns_3_2_1_U4.reset  = ap_rst;
assign \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.ain_s0  = \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.a ;
assign \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.bin_s0  = \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.b ;
assign \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.s  = { \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.fas_s2 , \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.sum_s1  };
assign \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.a  = \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.ain_s1 ;
assign \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.b  = \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.bin_s1 ;
assign \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.cin  = \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.carry_s1 ;
assign \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.facout_s2  = \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.cout ;
assign \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.fas_s2  = \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.s ;
assign \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.a  = \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.a [0];
assign \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.b  = \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.b [0];
assign \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.cin  = 1'h0;
assign \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.facout_s1  = \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.cout ;
assign \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.fas_s1  = \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.s ;
assign \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.a  = \add_2ns_2ns_2_2_1_U9.din0 ;
assign \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.b  = \add_2ns_2ns_2_2_1_U9.din1 ;
assign \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.ce  = \add_2ns_2ns_2_2_1_U9.ce ;
assign \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.clk  = \add_2ns_2ns_2_2_1_U9.clk ;
assign \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.reset  = \add_2ns_2ns_2_2_1_U9.reset ;
assign \add_2ns_2ns_2_2_1_U9.dout  = \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.s ;
assign \add_2ns_2ns_2_2_1_U9.ce  = 1'h1;
assign \add_2ns_2ns_2_2_1_U9.clk  = ap_clk;
assign \add_2ns_2ns_2_2_1_U9.din0  = ret_V_21_cast_reg_1200;
assign \add_2ns_2ns_2_2_1_U9.din1  = 2'h1;
assign grp_fu_639_p2 = \add_2ns_2ns_2_2_1_U9.dout ;
assign \add_2ns_2ns_2_2_1_U9.reset  = ap_rst;
assign \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.ain_s0  = \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.a ;
assign \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.bin_s0  = \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.b ;
assign \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.s  = { \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.fas_s2 , \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.sum_s1  };
assign \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.a  = \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.ain_s1 ;
assign \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.b  = \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.bin_s1 ;
assign \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.cin  = \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.carry_s1 ;
assign \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.facout_s2  = \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.cout ;
assign \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.fas_s2  = \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.s ;
assign \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.a  = \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.a [0];
assign \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.b  = \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.b [0];
assign \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.cin  = 1'h0;
assign \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.facout_s1  = \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.cout ;
assign \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.fas_s1  = \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.s ;
assign \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.a  = \add_2ns_2ns_2_2_1_U3.din0 ;
assign \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.b  = \add_2ns_2ns_2_2_1_U3.din1 ;
assign \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.ce  = \add_2ns_2ns_2_2_1_U3.ce ;
assign \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.clk  = \add_2ns_2ns_2_2_1_U3.clk ;
assign \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.reset  = \add_2ns_2ns_2_2_1_U3.reset ;
assign \add_2ns_2ns_2_2_1_U3.dout  = \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.s ;
assign \add_2ns_2ns_2_2_1_U3.ce  = 1'h1;
assign \add_2ns_2ns_2_2_1_U3.clk  = ap_clk;
assign \add_2ns_2ns_2_2_1_U3.din0  = p_Val2_1_reg_989;
assign \add_2ns_2ns_2_2_1_U3.din1  = { 1'h0, and_ln414_reg_1047 };
assign grp_fu_365_p2 = \add_2ns_2ns_2_2_1_U3.dout ;
assign \add_2ns_2ns_2_2_1_U3.reset  = ap_rst;
assign \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.ain_s0  = \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.a ;
assign \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.bin_s0  = \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.b ;
assign \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.s  = { \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.fas_s2 , \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.sum_s1  };
assign \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.a  = \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.ain_s1 ;
assign \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.b  = \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.bin_s1 ;
assign \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.cin  = \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.carry_s1 ;
assign \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.facout_s2  = \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.cout ;
assign \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.fas_s2  = \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.s ;
assign \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.a  = \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.a [0];
assign \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.b  = \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.b [0];
assign \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.cin  = 1'h0;
assign \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.facout_s1  = \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.cout ;
assign \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.fas_s1  = \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.s ;
assign \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.a  = \add_2ns_2ns_2_2_1_U2.din0 ;
assign \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.b  = \add_2ns_2ns_2_2_1_U2.din1 ;
assign \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.ce  = \add_2ns_2ns_2_2_1_U2.ce ;
assign \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.clk  = \add_2ns_2ns_2_2_1_U2.clk ;
assign \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.reset  = \add_2ns_2ns_2_2_1_U2.reset ;
assign \add_2ns_2ns_2_2_1_U2.dout  = \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.s ;
assign \add_2ns_2ns_2_2_1_U2.ce  = 1'h1;
assign \add_2ns_2ns_2_2_1_U2.clk  = ap_clk;
assign \add_2ns_2ns_2_2_1_U2.din0  = ret_V_4_cast_reg_964;
assign \add_2ns_2ns_2_2_1_U2.din1  = 2'h1;
assign grp_fu_314_p2 = \add_2ns_2ns_2_2_1_U2.dout ;
assign \add_2ns_2ns_2_2_1_U2.reset  = ap_rst;
assign \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.ain_s0  = \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.a ;
assign \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.bin_s0  = \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.b ;
assign \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.s  = { \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.fas_s2 , \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.sum_s1  };
assign \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.u2.a  = \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.ain_s1 ;
assign \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.u2.b  = \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.bin_s1 ;
assign \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.u2.cin  = \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.carry_s1 ;
assign \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.facout_s2  = \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.u2.cout ;
assign \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.fas_s2  = \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.u2.s ;
assign \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.u1.a  = \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.a [7:0];
assign \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.u1.b  = \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.b [7:0];
assign \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.u1.cin  = 1'h0;
assign \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.facout_s1  = \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.u1.cout ;
assign \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.fas_s1  = \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.u1.s ;
assign \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.a  = \add_17s_17s_17_2_1_U8.din0 ;
assign \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.b  = \add_17s_17s_17_2_1_U8.din1 ;
assign \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.ce  = \add_17s_17s_17_2_1_U8.ce ;
assign \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.clk  = \add_17s_17s_17_2_1_U8.clk ;
assign \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.reset  = \add_17s_17s_17_2_1_U8.reset ;
assign \add_17s_17s_17_2_1_U8.dout  = \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.s ;
assign \add_17s_17s_17_2_1_U8.ce  = 1'h1;
assign \add_17s_17s_17_2_1_U8.clk  = ap_clk;
assign \add_17s_17s_17_2_1_U8.din0  = { ret_V_19_reg_1157[2], ret_V_19_reg_1157, 13'h0000 };
assign \add_17s_17s_17_2_1_U8.din1  = { op_3[15], op_3 };
assign grp_fu_633_p2 = \add_17s_17s_17_2_1_U8.dout ;
assign \add_17s_17s_17_2_1_U8.reset  = ap_rst;
assign \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.ain_s0  = \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.a ;
assign \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.bin_s0  = \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.b ;
assign \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.s  = { \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.fas_s2 , \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.sum_s1  };
assign \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.u2.a  = \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.ain_s1 ;
assign \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.u2.b  = \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.bin_s1 ;
assign \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.u2.cin  = \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.carry_s1 ;
assign \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.facout_s2  = \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.u2.cout ;
assign \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.fas_s2  = \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.u2.s ;
assign \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.u1.a  = \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.a [6:0];
assign \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.u1.b  = \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.b [6:0];
assign \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.u1.cin  = 1'h0;
assign \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.facout_s1  = \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.u1.cout ;
assign \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.fas_s1  = \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.u1.s ;
assign \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.a  = \add_15ns_15ns_15_2_1_U6.din0 ;
assign \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.b  = \add_15ns_15ns_15_2_1_U6.din1 ;
assign \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.ce  = \add_15ns_15ns_15_2_1_U6.ce ;
assign \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.clk  = \add_15ns_15ns_15_2_1_U6.clk ;
assign \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.reset  = \add_15ns_15ns_15_2_1_U6.reset ;
assign \add_15ns_15ns_15_2_1_U6.dout  = \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.s ;
assign \add_15ns_15ns_15_2_1_U6.ce  = 1'h1;
assign \add_15ns_15ns_15_2_1_U6.clk  = ap_clk;
assign \add_15ns_15ns_15_2_1_U6.din0  = { trunc_ln728_reg_1165, 13'h0000 };
assign \add_15ns_15ns_15_2_1_U6.din1  = empty_reg_1093;
assign grp_fu_591_p2 = \add_15ns_15ns_15_2_1_U6.dout ;
assign \add_15ns_15ns_15_2_1_U6.reset  = ap_rst;
assign \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.ain_s0  = \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.a ;
assign \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.bin_s0  = \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.b ;
assign \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.s  = { \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.fas_s2 , \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.sum_s1  };
assign \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.u2.a  = \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.ain_s1 ;
assign \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.u2.b  = \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.bin_s1 ;
assign \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.u2.cin  = \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.carry_s1 ;
assign \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.facout_s2  = \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.u2.cout ;
assign \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.fas_s2  = \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.u2.s ;
assign \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.u1.a  = \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.a [4:0];
assign \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.u1.b  = \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.b [4:0];
assign \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.u1.cin  = 1'h0;
assign \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.facout_s1  = \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.u1.cout ;
assign \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.fas_s1  = \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.u1.s ;
assign \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.a  = \add_10ns_10s_10_2_1_U11.din0 ;
assign \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.b  = \add_10ns_10s_10_2_1_U11.din1 ;
assign \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.ce  = \add_10ns_10s_10_2_1_U11.ce ;
assign \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.clk  = \add_10ns_10s_10_2_1_U11.clk ;
assign \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.reset  = \add_10ns_10s_10_2_1_U11.reset ;
assign \add_10ns_10s_10_2_1_U11.dout  = \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.s ;
assign \add_10ns_10s_10_2_1_U11.ce  = 1'h1;
assign \add_10ns_10s_10_2_1_U11.clk  = ap_clk;
assign \add_10ns_10s_10_2_1_U11.din0  = { op_22_V_reg_1242, 5'h00 };
assign \add_10ns_10s_10_2_1_U11.din1  = { op_14[7], op_14[7], op_14 };
assign grp_fu_692_p2 = \add_10ns_10s_10_2_1_U11.dout ;
assign \add_10ns_10s_10_2_1_U11.reset  = ap_rst;
endmodule


// Machine B:
// Processed by function `add_clk_enable_signal` in `verilog_tricks.py`.
// Processed by function `remove_reset_signal` in `verilog_tricks.py`.
module top_B (
  ap_clk,
  ap_start,
  ap_done,
  ap_idle,
  ap_ready,
  op_0,
  op_1,
  op_2,
  op_3,
  op_7,
  op_8,
  op_10,
  op_12,
  op_13,
  op_14,
  op_28,
  op_28_ap_vld,
clk_enable
);
input clk_enable;


input ap_clk;
wire ap_rst;
assign ap_rst = op_28_ap_vld;
input ap_start;
input [1:0] op_0;
input [3:0] op_1;
input [3:0] op_10;
input [1:0] op_12;
input [3:0] op_13;
input [7:0] op_14;
input [7:0] op_2;
input [15:0] op_3;
input [1:0] op_7;
input [1:0] op_8;
output ap_done;
output ap_idle;
output ap_ready;
output [31:0] op_28;
output op_28_ap_vld;


reg Range1_all_ones_reg_1030;
reg Range1_all_zeros_reg_1037;
reg Range2_all_ones_reg_1025;
reg [4:0] \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.ain_s1 ;
reg [4:0] \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.bin_s1 ;
reg \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.carry_s1 ;
reg [4:0] \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.sum_s1 ;
reg [7:0] \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.ain_s1 ;
reg [7:0] \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.bin_s1 ;
reg \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.carry_s1 ;
reg [6:0] \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.sum_s1 ;
reg [8:0] \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.ain_s1 ;
reg [8:0] \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.bin_s1 ;
reg \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.carry_s1 ;
reg [7:0] \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.sum_s1 ;
reg \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.ain_s1 ;
reg \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.bin_s1 ;
reg \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.carry_s1 ;
reg \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.sum_s1 ;
reg \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.ain_s1 ;
reg \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.bin_s1 ;
reg \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.carry_s1 ;
reg \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.sum_s1 ;
reg \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.ain_s1 ;
reg \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.bin_s1 ;
reg \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.carry_s1 ;
reg \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.sum_s1 ;
reg [1:0] \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.ain_s1 ;
reg [1:0] \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.bin_s1 ;
reg \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.carry_s1 ;
reg \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.sum_s1 ;
reg [1:0] \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.ain_s1 ;
reg [1:0] \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.bin_s1 ;
reg \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.carry_s1 ;
reg \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.sum_s1 ;
reg [1:0] \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.ain_s1 ;
reg [1:0] \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.bin_s1 ;
reg \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.carry_s1 ;
reg [1:0] \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.sum_s1 ;
reg [2:0] \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.ain_s1 ;
reg [2:0] \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.bin_s1 ;
reg \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.carry_s1 ;
reg [1:0] \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.sum_s1 ;
reg [2:0] \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.ain_s1 ;
reg [2:0] \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.bin_s1 ;
reg \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.carry_s1 ;
reg [2:0] \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.sum_s1 ;
reg [2:0] \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.ain_s1 ;
reg [2:0] \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.bin_s1 ;
reg \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.carry_s1 ;
reg [2:0] \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.sum_s1 ;
reg [2:0] \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.ain_s1 ;
reg [2:0] \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.bin_s1 ;
reg \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.carry_s1 ;
reg [2:0] \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.sum_s1 ;
reg [2:0] \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.ain_s1 ;
reg [2:0] \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.bin_s1 ;
reg \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.carry_s1 ;
reg [2:0] \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.sum_s1 ;
reg [2:0] \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.ain_s1 ;
reg [2:0] \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.bin_s1 ;
reg \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.carry_s1 ;
reg [2:0] \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.sum_s1 ;
reg [5:0] add_ln691_1_reg_1284;
reg [5:0] add_ln691_2_reg_1375;
reg [1:0] add_ln691_reg_1237;
reg [5:0] add_ln69_2_reg_1314;
reg [3:0] add_ln69_reg_1207;
reg and_ln384_reg_1370;
reg and_ln414_reg_1047;
reg and_ln786_reg_1104;
reg [29:0] ap_CS_fsm = 30'h00000001;
reg carry_1_reg_1081;
reg deleted_zeros_reg_1098;
reg [14:0] empty_reg_1093;
reg icmp_ln414_reg_1020;
reg icmp_ln768_reg_1340;
reg icmp_ln786_reg_1345;
reg icmp_ln851_1_reg_1015;
reg icmp_ln851_2_reg_1127;
reg icmp_ln851_3_reg_1262;
reg icmp_ln851_reg_1137;
reg lhs_V_1_reg_1247;
reg newsignbit_reg_1326;
reg [4:0] op_22_V_reg_1242;
reg [5:0] op_25_V_reg_1350;
reg [1:0] op_5_V_reg_1152;
reg or_ln340_reg_1132;
reg or_ln785_1_reg_1358;
reg p_Result_10_reg_981;
reg p_Result_11_reg_994;
reg p_Result_12_reg_1068;
reg p_Result_13_reg_1319;
reg [4:0] p_Result_1_reg_1009;
reg [3:0] p_Result_s_reg_1004;
reg [1:0] p_Val2_1_reg_989;
reg [1:0] p_Val2_2_reg_1062;
reg [8:0] ret_V_17_reg_976;
reg [15:0] ret_V_18_reg_1110;
reg [2:0] ret_V_19_reg_1157;
reg [7:0] ret_V_20_reg_959;
reg [1:0] ret_V_21_cast_reg_1200;
reg [1:0] ret_V_21_reg_1052;
reg [2:0] ret_V_23_reg_1195;
reg [16:0] ret_V_24_reg_1232;
reg [9:0] ret_V_26_reg_1267;
reg [5:0] ret_V_27_reg_1289;
reg [5:0] ret_V_28_reg_1380;
reg [2:0] ret_V_3_reg_1147;
reg [1:0] ret_V_4_cast_reg_964;
reg [1:0] ret_V_6_reg_1042;
reg [2:0] ret_V_reg_1115;
reg [5:0] select_ln1192_reg_1385;
reg [1:0] select_ln340_reg_1142;
reg [5:0] select_ln69_reg_1309;
reg [5:0] sext_ln850_reg_1277;
reg [2:0] \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.ain_s1 ;
reg [2:0] \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.bin_s1 ;
reg \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.carry_s1 ;
reg [1:0] \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.sum_s1 ;
reg [4:0] \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.ain_s1 ;
reg [4:0] \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.bin_s1 ;
reg \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.carry_s1 ;
reg [3:0] \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.sum_s1 ;
reg [3:0] tmp_2_reg_1334;
reg [4:0] tmp_3_reg_1272;
reg [1:0] trunc_ln414_reg_999;
reg [1:0] trunc_ln728_reg_1165;
reg [1:0] trunc_ln851_1_reg_971;
reg [12:0] trunc_ln851_reg_1122;
reg underflow_1_reg_1364;
reg xor_ln416_reg_1075;
wire _000_;
wire _001_;
wire _002_;
wire [5:0] _003_;
wire [5:0] _004_;
wire [1:0] _005_;
wire [5:0] _006_;
wire [3:0] _007_;
wire _008_;
wire _009_;
wire _010_;
wire [29:0] _011_;
wire _012_;
wire _013_;
wire [14:0] _014_;
wire _015_;
wire _016_;
wire _017_;
wire _018_;
wire _019_;
wire _020_;
wire _021_;
wire _022_;
wire _023_;
wire [4:0] _024_;
wire [5:0] _025_;
wire [1:0] _026_;
wire _027_;
wire _028_;
wire _029_;
wire _030_;
wire _031_;
wire _032_;
wire [4:0] _033_;
wire [3:0] _034_;
wire [1:0] _035_;
wire [1:0] _036_;
wire [8:0] _037_;
wire [15:0] _038_;
wire [2:0] _039_;
wire [7:0] _040_;
wire [1:0] _041_;
wire [1:0] _042_;
wire [2:0] _043_;
wire [16:0] _044_;
wire [9:0] _045_;
wire [5:0] _046_;
wire [5:0] _047_;
wire [2:0] _048_;
wire [1:0] _049_;
wire [1:0] _050_;
wire [2:0] _051_;
wire [5:0] _052_;
wire [1:0] _053_;
wire [1:0] _054_;
wire [5:0] _055_;
wire [3:0] _056_;
wire [4:0] _057_;
wire [1:0] _058_;
wire [1:0] _059_;
wire [1:0] _060_;
wire [12:0] _061_;
wire _062_;
wire _063_;
wire [1:0] _064_;
wire _065_;
wire _066_;
wire _067_;
wire _068_;
wire _069_;
wire _070_;
wire _071_;
wire _072_;
wire _073_;
wire _074_;
wire _075_;
wire [4:0] _076_;
wire [4:0] _077_;
wire _078_;
wire [4:0] _079_;
wire [5:0] _080_;
wire [5:0] _081_;
wire [7:0] _082_;
wire [7:0] _083_;
wire _084_;
wire [6:0] _085_;
wire [7:0] _086_;
wire [8:0] _087_;
wire [8:0] _088_;
wire [8:0] _089_;
wire _090_;
wire [7:0] _091_;
wire [8:0] _092_;
wire [9:0] _093_;
wire _094_;
wire _095_;
wire _096_;
wire _097_;
wire [1:0] _098_;
wire [1:0] _099_;
wire _100_;
wire _101_;
wire _102_;
wire _103_;
wire [1:0] _104_;
wire [1:0] _105_;
wire _106_;
wire _107_;
wire _108_;
wire _109_;
wire [1:0] _110_;
wire [1:0] _111_;
wire [1:0] _112_;
wire [1:0] _113_;
wire _114_;
wire _115_;
wire [1:0] _116_;
wire [2:0] _117_;
wire [1:0] _118_;
wire [1:0] _119_;
wire _120_;
wire _121_;
wire [1:0] _122_;
wire [2:0] _123_;
wire [1:0] _124_;
wire [1:0] _125_;
wire _126_;
wire [1:0] _127_;
wire [2:0] _128_;
wire [2:0] _129_;
wire [2:0] _130_;
wire [2:0] _131_;
wire _132_;
wire [1:0] _133_;
wire [2:0] _134_;
wire [3:0] _135_;
wire [2:0] _136_;
wire [2:0] _137_;
wire _138_;
wire [2:0] _139_;
wire [3:0] _140_;
wire [3:0] _141_;
wire [2:0] _142_;
wire [2:0] _143_;
wire _144_;
wire [2:0] _145_;
wire [3:0] _146_;
wire [3:0] _147_;
wire [2:0] _148_;
wire [2:0] _149_;
wire _150_;
wire [2:0] _151_;
wire [3:0] _152_;
wire [3:0] _153_;
wire [2:0] _154_;
wire [2:0] _155_;
wire _156_;
wire [2:0] _157_;
wire [3:0] _158_;
wire [3:0] _159_;
wire [2:0] _160_;
wire [2:0] _161_;
wire _162_;
wire [2:0] _163_;
wire [3:0] _164_;
wire [3:0] _165_;
wire [2:0] _166_;
wire [2:0] _167_;
wire _168_;
wire [1:0] _169_;
wire [2:0] _170_;
wire [3:0] _171_;
wire [4:0] _172_;
wire [4:0] _173_;
wire _174_;
wire [3:0] _175_;
wire [4:0] _176_;
wire [5:0] _177_;
wire _178_;
wire _179_;
wire _180_;
wire _181_;
wire _182_;
wire _183_;
wire _184_;
wire _185_;
wire _186_;
wire _187_;
wire _188_;
wire _189_;
wire _190_;
wire _191_;
wire _192_;
wire _193_;
wire _194_;
wire _195_;
wire _196_;
wire _197_;
wire _198_;
wire _199_;
wire _200_;
wire _201_;
wire _202_;
wire _203_;
wire _204_;
wire _205_;
wire _206_;
wire _207_;
wire _208_;
wire _209_;
wire _210_;
wire _211_;
wire _212_;
wire _213_;
wire Range1_all_ones_fu_329_p2;
wire Range1_all_zeros_fu_334_p2;
wire Range2_all_ones_fu_324_p2;
wire \add_10ns_10s_10_2_1_U11.ce ;
wire \add_10ns_10s_10_2_1_U11.clk ;
wire [9:0] \add_10ns_10s_10_2_1_U11.din0 ;
wire [9:0] \add_10ns_10s_10_2_1_U11.din1 ;
wire [9:0] \add_10ns_10s_10_2_1_U11.dout ;
wire \add_10ns_10s_10_2_1_U11.reset ;
wire [9:0] \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.a ;
wire [9:0] \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.ain_s0 ;
wire [9:0] \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.b ;
wire [9:0] \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.bin_s0 ;
wire \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.ce ;
wire \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.clk ;
wire \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.facout_s1 ;
wire \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.facout_s2 ;
wire [4:0] \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.fas_s1 ;
wire [4:0] \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.fas_s2 ;
wire \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.reset ;
wire [9:0] \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.s ;
wire [4:0] \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.u1.a ;
wire [4:0] \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.u1.b ;
wire \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.u1.cin ;
wire \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.u1.cout ;
wire [4:0] \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.u1.s ;
wire [4:0] \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.u2.a ;
wire [4:0] \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.u2.b ;
wire \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.u2.cin ;
wire \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.u2.cout ;
wire [4:0] \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.u2.s ;
wire \add_15ns_15ns_15_2_1_U6.ce ;
wire \add_15ns_15ns_15_2_1_U6.clk ;
wire [14:0] \add_15ns_15ns_15_2_1_U6.din0 ;
wire [14:0] \add_15ns_15ns_15_2_1_U6.din1 ;
wire [14:0] \add_15ns_15ns_15_2_1_U6.dout ;
wire \add_15ns_15ns_15_2_1_U6.reset ;
wire [14:0] \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.a ;
wire [14:0] \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.ain_s0 ;
wire [14:0] \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.b ;
wire [14:0] \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.bin_s0 ;
wire \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.ce ;
wire \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.clk ;
wire \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.facout_s1 ;
wire \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.facout_s2 ;
wire [6:0] \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.fas_s1 ;
wire [7:0] \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.fas_s2 ;
wire \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.reset ;
wire [14:0] \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.s ;
wire [6:0] \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.u1.a ;
wire [6:0] \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.u1.b ;
wire \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.u1.cin ;
wire \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.u1.cout ;
wire [6:0] \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.u1.s ;
wire [7:0] \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.u2.a ;
wire [7:0] \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.u2.b ;
wire \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.u2.cin ;
wire \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.u2.cout ;
wire [7:0] \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.u2.s ;
wire \add_17s_17s_17_2_1_U8.ce ;
wire \add_17s_17s_17_2_1_U8.clk ;
wire [16:0] \add_17s_17s_17_2_1_U8.din0 ;
wire [16:0] \add_17s_17s_17_2_1_U8.din1 ;
wire [16:0] \add_17s_17s_17_2_1_U8.dout ;
wire \add_17s_17s_17_2_1_U8.reset ;
wire [16:0] \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.a ;
wire [16:0] \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.ain_s0 ;
wire [16:0] \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.b ;
wire [16:0] \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.bin_s0 ;
wire \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.ce ;
wire \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.clk ;
wire \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.facout_s1 ;
wire \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.facout_s2 ;
wire [7:0] \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.fas_s1 ;
wire [8:0] \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.fas_s2 ;
wire \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.reset ;
wire [16:0] \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.s ;
wire [7:0] \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.u1.a ;
wire [7:0] \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.u1.b ;
wire \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.u1.cin ;
wire \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.u1.cout ;
wire [7:0] \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.u1.s ;
wire [8:0] \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.u2.a ;
wire [8:0] \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.u2.b ;
wire \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.u2.cin ;
wire \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.u2.cout ;
wire [8:0] \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.u2.s ;
wire \add_2ns_2ns_2_2_1_U2.ce ;
wire \add_2ns_2ns_2_2_1_U2.clk ;
wire [1:0] \add_2ns_2ns_2_2_1_U2.din0 ;
wire [1:0] \add_2ns_2ns_2_2_1_U2.din1 ;
wire [1:0] \add_2ns_2ns_2_2_1_U2.dout ;
wire \add_2ns_2ns_2_2_1_U2.reset ;
wire [1:0] \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.a ;
wire [1:0] \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.ain_s0 ;
wire [1:0] \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.b ;
wire [1:0] \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.bin_s0 ;
wire \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.ce ;
wire \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.clk ;
wire \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.facout_s1 ;
wire \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.facout_s2 ;
wire \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.fas_s1 ;
wire \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.fas_s2 ;
wire \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.reset ;
wire [1:0] \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.s ;
wire \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.a ;
wire \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.b ;
wire \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.cin ;
wire \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.cout ;
wire \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.s ;
wire \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.a ;
wire \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.b ;
wire \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.cin ;
wire \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.cout ;
wire \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.s ;
wire \add_2ns_2ns_2_2_1_U3.ce ;
wire \add_2ns_2ns_2_2_1_U3.clk ;
wire [1:0] \add_2ns_2ns_2_2_1_U3.din0 ;
wire [1:0] \add_2ns_2ns_2_2_1_U3.din1 ;
wire [1:0] \add_2ns_2ns_2_2_1_U3.dout ;
wire \add_2ns_2ns_2_2_1_U3.reset ;
wire [1:0] \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.a ;
wire [1:0] \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.ain_s0 ;
wire [1:0] \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.b ;
wire [1:0] \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.bin_s0 ;
wire \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.ce ;
wire \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.clk ;
wire \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.facout_s1 ;
wire \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.facout_s2 ;
wire \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.fas_s1 ;
wire \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.fas_s2 ;
wire \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.reset ;
wire [1:0] \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.s ;
wire \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.a ;
wire \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.b ;
wire \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.cin ;
wire \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.cout ;
wire \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.s ;
wire \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.a ;
wire \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.b ;
wire \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.cin ;
wire \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.cout ;
wire \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.s ;
wire \add_2ns_2ns_2_2_1_U9.ce ;
wire \add_2ns_2ns_2_2_1_U9.clk ;
wire [1:0] \add_2ns_2ns_2_2_1_U9.din0 ;
wire [1:0] \add_2ns_2ns_2_2_1_U9.din1 ;
wire [1:0] \add_2ns_2ns_2_2_1_U9.dout ;
wire \add_2ns_2ns_2_2_1_U9.reset ;
wire [1:0] \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.a ;
wire [1:0] \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.ain_s0 ;
wire [1:0] \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.b ;
wire [1:0] \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.bin_s0 ;
wire \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.ce ;
wire \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.clk ;
wire \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.facout_s1 ;
wire \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.facout_s2 ;
wire \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.fas_s1 ;
wire \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.fas_s2 ;
wire \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.reset ;
wire [1:0] \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.s ;
wire \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.a ;
wire \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.b ;
wire \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.cin ;
wire \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.cout ;
wire \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.s ;
wire \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.a ;
wire \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.b ;
wire \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.cin ;
wire \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.cout ;
wire \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.s ;
wire \add_3ns_3ns_3_2_1_U4.ce ;
wire \add_3ns_3ns_3_2_1_U4.clk ;
wire [2:0] \add_3ns_3ns_3_2_1_U4.din0 ;
wire [2:0] \add_3ns_3ns_3_2_1_U4.din1 ;
wire [2:0] \add_3ns_3ns_3_2_1_U4.dout ;
wire \add_3ns_3ns_3_2_1_U4.reset ;
wire [2:0] \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.a ;
wire [2:0] \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.ain_s0 ;
wire [2:0] \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.b ;
wire [2:0] \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.bin_s0 ;
wire \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.ce ;
wire \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.clk ;
wire \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.facout_s1 ;
wire \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.facout_s2 ;
wire \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.fas_s1 ;
wire [1:0] \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.fas_s2 ;
wire \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.reset ;
wire [2:0] \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.s ;
wire \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.u1.a ;
wire \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.u1.b ;
wire \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.u1.cin ;
wire \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.u1.cout ;
wire \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.u1.s ;
wire [1:0] \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.u2.a ;
wire [1:0] \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.u2.b ;
wire \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.u2.cin ;
wire \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.u2.cout ;
wire [1:0] \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.u2.s ;
wire \add_3s_3s_3_2_1_U5.ce ;
wire \add_3s_3s_3_2_1_U5.clk ;
wire [2:0] \add_3s_3s_3_2_1_U5.din0 ;
wire [2:0] \add_3s_3s_3_2_1_U5.din1 ;
wire [2:0] \add_3s_3s_3_2_1_U5.dout ;
wire \add_3s_3s_3_2_1_U5.reset ;
wire [2:0] \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.a ;
wire [2:0] \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.ain_s0 ;
wire [2:0] \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.b ;
wire [2:0] \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.bin_s0 ;
wire \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.ce ;
wire \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.clk ;
wire \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.facout_s1 ;
wire \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.facout_s2 ;
wire \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.fas_s1 ;
wire [1:0] \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.fas_s2 ;
wire \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.reset ;
wire [2:0] \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.s ;
wire \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.u1.a ;
wire \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.u1.b ;
wire \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.u1.cin ;
wire \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.u1.cout ;
wire \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.u1.s ;
wire [1:0] \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.u2.a ;
wire [1:0] \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.u2.b ;
wire \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.u2.cin ;
wire \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.u2.cout ;
wire [1:0] \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.u2.s ;
wire \add_4s_4ns_4_2_1_U7.ce ;
wire \add_4s_4ns_4_2_1_U7.clk ;
wire [3:0] \add_4s_4ns_4_2_1_U7.din0 ;
wire [3:0] \add_4s_4ns_4_2_1_U7.din1 ;
wire [3:0] \add_4s_4ns_4_2_1_U7.dout ;
wire \add_4s_4ns_4_2_1_U7.reset ;
wire [3:0] \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.a ;
wire [3:0] \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.ain_s0 ;
wire [3:0] \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.b ;
wire [3:0] \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.bin_s0 ;
wire \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.ce ;
wire \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.clk ;
wire \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.facout_s1 ;
wire \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.facout_s2 ;
wire [1:0] \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.fas_s1 ;
wire [1:0] \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.fas_s2 ;
wire \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.reset ;
wire [3:0] \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.s ;
wire [1:0] \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.u1.a ;
wire [1:0] \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.u1.b ;
wire \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.u1.cin ;
wire \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.u1.cout ;
wire [1:0] \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.u1.s ;
wire [1:0] \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.u2.a ;
wire [1:0] \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.u2.b ;
wire \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.u2.cin ;
wire \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.u2.cout ;
wire [1:0] \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.u2.s ;
wire \add_5s_5s_5_2_1_U10.ce ;
wire \add_5s_5s_5_2_1_U10.clk ;
wire [4:0] \add_5s_5s_5_2_1_U10.din0 ;
wire [4:0] \add_5s_5s_5_2_1_U10.din1 ;
wire [4:0] \add_5s_5s_5_2_1_U10.dout ;
wire \add_5s_5s_5_2_1_U10.reset ;
wire [4:0] \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.a ;
wire [4:0] \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.ain_s0 ;
wire [4:0] \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.b ;
wire [4:0] \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.bin_s0 ;
wire \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.ce ;
wire \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.clk ;
wire \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.facout_s1 ;
wire \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.facout_s2 ;
wire [1:0] \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.fas_s1 ;
wire [2:0] \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.fas_s2 ;
wire \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.reset ;
wire [4:0] \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.s ;
wire [1:0] \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.u1.a ;
wire [1:0] \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.u1.b ;
wire \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.u1.cin ;
wire \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.u1.cout ;
wire [1:0] \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.u1.s ;
wire [2:0] \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.u2.a ;
wire [2:0] \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.u2.b ;
wire \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.u2.cin ;
wire \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.u2.cout ;
wire [2:0] \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.u2.s ;
wire \add_6ns_6ns_6_2_1_U15.ce ;
wire \add_6ns_6ns_6_2_1_U15.clk ;
wire [5:0] \add_6ns_6ns_6_2_1_U15.din0 ;
wire [5:0] \add_6ns_6ns_6_2_1_U15.din1 ;
wire [5:0] \add_6ns_6ns_6_2_1_U15.dout ;
wire \add_6ns_6ns_6_2_1_U15.reset ;
wire [5:0] \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.a ;
wire [5:0] \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.ain_s0 ;
wire [5:0] \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.b ;
wire [5:0] \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.bin_s0 ;
wire \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.ce ;
wire \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.clk ;
wire \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.facout_s1 ;
wire \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.facout_s2 ;
wire [2:0] \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.fas_s1 ;
wire [2:0] \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.fas_s2 ;
wire \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.reset ;
wire [5:0] \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.s ;
wire [2:0] \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.u1.a ;
wire [2:0] \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.u1.b ;
wire \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.u1.cin ;
wire \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.u1.cout ;
wire [2:0] \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.u1.s ;
wire [2:0] \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.u2.a ;
wire [2:0] \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.u2.b ;
wire \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.u2.cin ;
wire \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.u2.cout ;
wire [2:0] \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.u2.s ;
wire \add_6ns_6ns_6_2_1_U16.ce ;
wire \add_6ns_6ns_6_2_1_U16.clk ;
wire [5:0] \add_6ns_6ns_6_2_1_U16.din0 ;
wire [5:0] \add_6ns_6ns_6_2_1_U16.din1 ;
wire [5:0] \add_6ns_6ns_6_2_1_U16.dout ;
wire \add_6ns_6ns_6_2_1_U16.reset ;
wire [5:0] \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.a ;
wire [5:0] \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.ain_s0 ;
wire [5:0] \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.b ;
wire [5:0] \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.bin_s0 ;
wire \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.ce ;
wire \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.clk ;
wire \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.facout_s1 ;
wire \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.facout_s2 ;
wire [2:0] \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.fas_s1 ;
wire [2:0] \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.fas_s2 ;
wire \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.reset ;
wire [5:0] \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.s ;
wire [2:0] \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.u1.a ;
wire [2:0] \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.u1.b ;
wire \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.u1.cin ;
wire \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.u1.cout ;
wire [2:0] \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.u1.s ;
wire [2:0] \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.u2.a ;
wire [2:0] \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.u2.b ;
wire \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.u2.cin ;
wire \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.u2.cout ;
wire [2:0] \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.u2.s ;
wire \add_6ns_6ns_6_2_1_U17.ce ;
wire \add_6ns_6ns_6_2_1_U17.clk ;
wire [5:0] \add_6ns_6ns_6_2_1_U17.din0 ;
wire [5:0] \add_6ns_6ns_6_2_1_U17.din1 ;
wire [5:0] \add_6ns_6ns_6_2_1_U17.dout ;
wire \add_6ns_6ns_6_2_1_U17.reset ;
wire [5:0] \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.a ;
wire [5:0] \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.ain_s0 ;
wire [5:0] \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.b ;
wire [5:0] \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.bin_s0 ;
wire \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.ce ;
wire \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.clk ;
wire \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.facout_s1 ;
wire \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.facout_s2 ;
wire [2:0] \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.fas_s1 ;
wire [2:0] \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.fas_s2 ;
wire \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.reset ;
wire [5:0] \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.s ;
wire [2:0] \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.u1.a ;
wire [2:0] \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.u1.b ;
wire \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.u1.cin ;
wire \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.u1.cout ;
wire [2:0] \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.u1.s ;
wire [2:0] \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.u2.a ;
wire [2:0] \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.u2.b ;
wire \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.u2.cin ;
wire \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.u2.cout ;
wire [2:0] \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.u2.s ;
wire \add_6ns_6s_6_2_1_U13.ce ;
wire \add_6ns_6s_6_2_1_U13.clk ;
wire [5:0] \add_6ns_6s_6_2_1_U13.din0 ;
wire [5:0] \add_6ns_6s_6_2_1_U13.din1 ;
wire [5:0] \add_6ns_6s_6_2_1_U13.dout ;
wire \add_6ns_6s_6_2_1_U13.reset ;
wire [5:0] \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.a ;
wire [5:0] \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.ain_s0 ;
wire [5:0] \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.b ;
wire [5:0] \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.bin_s0 ;
wire \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.ce ;
wire \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.clk ;
wire \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.facout_s1 ;
wire \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.facout_s2 ;
wire [2:0] \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.fas_s1 ;
wire [2:0] \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.fas_s2 ;
wire \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.reset ;
wire [5:0] \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.s ;
wire [2:0] \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.u1.a ;
wire [2:0] \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.u1.b ;
wire \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.u1.cin ;
wire \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.u1.cout ;
wire [2:0] \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.u1.s ;
wire [2:0] \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.u2.a ;
wire [2:0] \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.u2.b ;
wire \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.u2.cin ;
wire \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.u2.cout ;
wire [2:0] \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.u2.s ;
wire \add_6s_6ns_6_2_1_U12.ce ;
wire \add_6s_6ns_6_2_1_U12.clk ;
wire [5:0] \add_6s_6ns_6_2_1_U12.din0 ;
wire [5:0] \add_6s_6ns_6_2_1_U12.din1 ;
wire [5:0] \add_6s_6ns_6_2_1_U12.dout ;
wire \add_6s_6ns_6_2_1_U12.reset ;
wire [5:0] \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.a ;
wire [5:0] \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.ain_s0 ;
wire [5:0] \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.b ;
wire [5:0] \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.bin_s0 ;
wire \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.ce ;
wire \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.clk ;
wire \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.facout_s1 ;
wire \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.facout_s2 ;
wire [2:0] \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.fas_s1 ;
wire [2:0] \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.fas_s2 ;
wire \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.reset ;
wire [5:0] \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.s ;
wire [2:0] \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.u1.a ;
wire [2:0] \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.u1.b ;
wire \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.u1.cin ;
wire \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.u1.cout ;
wire [2:0] \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.u1.s ;
wire [2:0] \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.u2.a ;
wire [2:0] \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.u2.b ;
wire \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.u2.cin ;
wire \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.u2.cout ;
wire [2:0] \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.u2.s ;
wire and_ln384_fu_881_p2;
wire and_ln414_fu_339_p2;
wire and_ln780_fu_409_p2;
wire and_ln781_fu_498_p2;
wire and_ln785_1_fu_534_p2;
wire and_ln785_fu_525_p2;
wire and_ln786_fu_420_p2;
wire and_ln850_fu_774_p2;
wire ap_CS_fsm_state1;
wire ap_CS_fsm_state10;
wire ap_CS_fsm_state11;
wire ap_CS_fsm_state12;
wire ap_CS_fsm_state13;
wire ap_CS_fsm_state14;
wire ap_CS_fsm_state15;
wire ap_CS_fsm_state16;
wire ap_CS_fsm_state17;
wire ap_CS_fsm_state18;
wire ap_CS_fsm_state19;
wire ap_CS_fsm_state2;
wire ap_CS_fsm_state20;
wire ap_CS_fsm_state21;
wire ap_CS_fsm_state22;
wire ap_CS_fsm_state23;
wire ap_CS_fsm_state24;
wire ap_CS_fsm_state25;
wire ap_CS_fsm_state26;
wire ap_CS_fsm_state27;
wire ap_CS_fsm_state28;
wire ap_CS_fsm_state29;
wire ap_CS_fsm_state3;
wire ap_CS_fsm_state30;
wire ap_CS_fsm_state4;
wire ap_CS_fsm_state5;
wire ap_CS_fsm_state6;
wire ap_CS_fsm_state7;
wire ap_CS_fsm_state8;
wire ap_CS_fsm_state9;
wire [29:0] ap_NS_fsm;
wire ap_clk;
wire ap_done;
wire ap_idle;
wire ap_ready;
wire ap_rst;
wire ap_start;
wire carry_1_fu_383_p2;
wire deleted_ones_fu_414_p3;
wire deleted_zeros_fu_391_p3;
wire [15:0] empty_fu_387_p0;
wire [14:0] empty_fu_387_p1;
wire [8:0] grp_fu_221_p0;
wire [8:0] grp_fu_221_p1;
wire [8:0] grp_fu_221_p2;
wire [1:0] grp_fu_314_p2;
wire [1:0] grp_fu_365_p1;
wire [1:0] grp_fu_365_p2;
wire [2:0] grp_fu_493_p2;
wire [2:0] grp_fu_578_p0;
wire [2:0] grp_fu_578_p1;
wire [2:0] grp_fu_578_p2;
wire [14:0] grp_fu_591_p0;
wire [14:0] grp_fu_591_p2;
wire [3:0] grp_fu_600_p0;
wire [3:0] grp_fu_600_p1;
wire [3:0] grp_fu_600_p2;
wire [16:0] grp_fu_633_p0;
wire [16:0] grp_fu_633_p1;
wire [16:0] grp_fu_633_p2;
wire [1:0] grp_fu_639_p2;
wire [4:0] grp_fu_647_p0;
wire [4:0] grp_fu_647_p1;
wire [4:0] grp_fu_647_p2;
wire [9:0] grp_fu_692_p0;
wire [9:0] grp_fu_692_p1;
wire [9:0] grp_fu_692_p2;
wire [5:0] grp_fu_721_p0;
wire [5:0] grp_fu_721_p2;
wire [5:0] grp_fu_749_p1;
wire [5:0] grp_fu_749_p2;
wire [4:0] grp_fu_793_p0;
wire [4:0] grp_fu_793_p1;
wire [4:0] grp_fu_793_p2;
wire [5:0] grp_fu_829_p2;
wire [5:0] grp_fu_862_p2;
wire [5:0] grp_fu_935_p2;
wire icmp_ln414_fu_319_p2;
wire icmp_ln768_fu_833_p2;
wire icmp_ln786_fu_838_p2;
wire icmp_ln851_1_fu_309_p2;
wire icmp_ln851_2_fu_456_p2;
wire icmp_ln851_3_fu_702_p2;
wire icmp_ln851_fu_488_p2;
wire [15:0] lhs_1_fu_425_p3;
wire lhs_V_1_fu_676_p2;
wire [4:0] lhs_fu_205_p3;
wire neg_src_fu_508_p2;
wire newsignbit_fu_815_p1;
wire [1:0] op_0;
wire [3:0] op_1;
wire [3:0] op_10;
wire [1:0] op_12;
wire [3:0] op_13;
wire [7:0] op_14;
wire op_19_V_fu_902_p3;
wire [7:0] op_2;
wire [31:0] op_28;
wire op_28_ap_vld;
wire [15:0] op_3;
wire [1:0] op_5_V_fu_539_p3;
wire [1:0] op_7;
wire [1:0] op_8;
wire or_ln340_1_fu_897_p2;
wire or_ln340_2_fu_513_p2;
wire or_ln340_fu_483_p2;
wire or_ln384_fu_876_p2;
wire or_ln388_fu_867_p2;
wire or_ln785_1_fu_843_p2;
wire or_ln785_2_fu_529_p2;
wire or_ln785_fu_467_p2;
wire or_ln786_fu_852_p2;
wire overflow_1_fu_892_p2;
wire overflow_fu_477_p2;
wire p_Result_2_fu_343_p3;
wire p_Result_3_fu_762_p3;
wire p_Result_5_fu_653_p3;
wire p_Result_8_fu_727_p3;
wire p_Result_9_fu_908_p3;
wire p_Result_s_16_fu_545_p3;
wire [15:0] ret_V_18_fu_432_p1;
wire [15:0] ret_V_18_fu_432_p2;
wire [2:0] ret_V_19_fu_557_p3;
wire [7:0] ret_V_20_fu_239_p1;
wire [7:0] ret_V_20_fu_239_p2;
wire [1:0] ret_V_21_fu_355_p3;
wire ret_V_22_fu_780_p2;
wire [1:0] ret_V_25_fu_665_p3;
wire [5:0] ret_V_27_fu_739_p3;
wire [5:0] ret_V_28_fu_920_p3;
wire ret_V_8_fu_754_p3;
wire [15:0] rhs_3_fu_622_p3;
wire [3:0] rhs_fu_227_p3;
wire [5:0] select_ln1192_fu_927_p3;
wire [1:0] select_ln340_fu_518_p3;
wire [1:0] select_ln69_fu_799_p3;
wire [1:0] select_ln850_1_fu_350_p3;
wire [1:0] select_ln850_2_fu_660_p3;
wire [5:0] select_ln850_3_fu_734_p3;
wire [5:0] select_ln850_4_fu_915_p3;
wire [2:0] select_ln850_fu_552_p3;
wire [7:0] sext_ln1192_2_fu_681_p0;
wire [15:0] sext_ln1192_fu_619_p0;
wire [7:0] sext_ln1195_fu_235_p1;
wire [7:0] sext_ln703_fu_217_p0;
wire [5:0] sext_ln850_fu_718_p1;
wire \sub_5s_5s_5_2_1_U14.ce ;
wire \sub_5s_5s_5_2_1_U14.clk ;
wire [4:0] \sub_5s_5s_5_2_1_U14.din0 ;
wire [4:0] \sub_5s_5s_5_2_1_U14.din1 ;
wire [4:0] \sub_5s_5s_5_2_1_U14.dout ;
wire \sub_5s_5s_5_2_1_U14.reset ;
wire [4:0] \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.a ;
wire [4:0] \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.ain_s0 ;
wire [4:0] \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.b ;
wire [4:0] \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.bin_s0 ;
wire \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.ce ;
wire \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.clk ;
wire \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.facout_s1 ;
wire \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.facout_s2 ;
wire [1:0] \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.fas_s1 ;
wire [2:0] \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.fas_s2 ;
wire \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.reset ;
wire [4:0] \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.s ;
wire [1:0] \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.u1.a ;
wire [1:0] \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.u1.b ;
wire \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.u1.cin ;
wire \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.u1.cout ;
wire [1:0] \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.u1.s ;
wire [2:0] \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.u2.a ;
wire [2:0] \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.u2.b ;
wire \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.u2.cin ;
wire \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.u2.cout ;
wire [2:0] \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.u2.s ;
wire \sub_9s_9s_9_2_1_U1.ce ;
wire \sub_9s_9s_9_2_1_U1.clk ;
wire [8:0] \sub_9s_9s_9_2_1_U1.din0 ;
wire [8:0] \sub_9s_9s_9_2_1_U1.din1 ;
wire [8:0] \sub_9s_9s_9_2_1_U1.dout ;
wire \sub_9s_9s_9_2_1_U1.reset ;
wire [8:0] \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.a ;
wire [8:0] \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.ain_s0 ;
wire [8:0] \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.b ;
wire [8:0] \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.bin_s0 ;
wire \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.ce ;
wire \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.clk ;
wire \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.facout_s1 ;
wire \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.facout_s2 ;
wire [3:0] \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.fas_s1 ;
wire [4:0] \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.fas_s2 ;
wire \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.reset ;
wire [8:0] \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.s ;
wire [3:0] \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.u1.a ;
wire [3:0] \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.u1.b ;
wire \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.u1.cin ;
wire \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.u1.cout ;
wire [3:0] \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.u1.s ;
wire [4:0] \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.u2.a ;
wire [4:0] \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.u2.b ;
wire \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.u2.cin ;
wire \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.u2.cout ;
wire [4:0] \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.u2.s ;
wire tmp_fu_396_p3;
wire [1:0] trunc_ln414_fu_285_p1;
wire [1:0] trunc_ln728_fu_564_p1;
wire [1:0] trunc_ln851_1_fu_255_p1;
wire trunc_ln851_2_fu_770_p1;
wire [15:0] trunc_ln851_3_fu_452_p0;
wire [12:0] trunc_ln851_3_fu_452_p1;
wire [7:0] trunc_ln851_4_fu_698_p0;
wire [4:0] trunc_ln851_4_fu_698_p1;
wire [12:0] trunc_ln851_fu_448_p1;
wire underflow_1_fu_857_p2;
wire xor_ln384_fu_871_p2;
wire xor_ln416_fu_378_p2;
wire xor_ln780_fu_403_p2;
wire xor_ln781_fu_502_p2;
wire xor_ln785_1_fu_472_p2;
wire xor_ln785_2_fu_887_p2;
wire xor_ln785_fu_462_p2;
wire xor_ln786_fu_847_p2;
wire [2:0] zext_ln886_fu_672_p1;


assign _065_ = icmp_ln851_3_reg_1262 & ap_CS_fsm[19];
assign _066_ = lhs_V_1_reg_1247 & ap_CS_fsm[26];
assign _067_ = ap_CS_fsm[15] & icmp_ln851_2_reg_1127;
assign _068_ = _070_ & ap_CS_fsm[0];
assign _069_ = ap_start & ap_CS_fsm[0];
assign and_ln384_fu_881_p2 = or_ln388_fu_867_p2 & or_ln384_fu_876_p2;
assign and_ln414_fu_339_p2 = p_Result_10_reg_981 & icmp_ln414_reg_1020;
assign and_ln780_fu_409_p2 = xor_ln780_fu_403_p2 & Range2_all_ones_reg_1025;
assign and_ln781_fu_498_p2 = carry_1_reg_1081 & Range1_all_ones_reg_1030;
assign and_ln785_1_fu_534_p2 = or_ln785_2_fu_529_p2 & and_ln786_reg_1104;
assign and_ln785_fu_525_p2 = xor_ln416_reg_1075 & deleted_zeros_reg_1098;
assign and_ln786_fu_420_p2 = p_Result_12_reg_1068 & deleted_ones_fu_414_p3;
assign and_ln850_fu_774_p2 = op_8[0] & op_8[1];
assign carry_1_fu_383_p2 = xor_ln416_reg_1075 & p_Result_11_reg_994;
assign neg_src_fu_508_p2 = xor_ln781_fu_502_p2 & p_Result_10_reg_981;
assign overflow_1_fu_892_p2 = xor_ln785_2_fu_887_p2 & or_ln785_1_reg_1358;
assign overflow_fu_477_p2 = xor_ln785_1_fu_472_p2 & or_ln785_fu_467_p2;
assign underflow_1_fu_857_p2 = p_Result_13_reg_1319 & or_ln786_fu_852_p2;
assign xor_ln384_fu_871_p2 = ~ or_ln785_1_reg_1358;
assign xor_ln780_fu_403_p2 = ~ ret_V_17_reg_976[4];
assign xor_ln781_fu_502_p2 = ~ and_ln781_fu_498_p2;
assign xor_ln785_2_fu_887_p2 = ~ p_Result_13_reg_1319;
assign xor_ln785_fu_462_p2 = ~ deleted_zeros_reg_1098;
assign xor_ln785_1_fu_472_p2 = ~ p_Result_10_reg_981;
assign xor_ln786_fu_847_p2 = ~ newsignbit_reg_1326;
assign xor_ln416_fu_378_p2 = ~ p_Result_12_reg_1068;
assign _070_ = ~ ap_start;
assign _071_ = p_Result_1_reg_1009 == 5'h1f;
assign _072_ = ! p_Result_1_reg_1009;
assign _073_ = p_Result_s_reg_1004 == 4'hf;
assign _074_ = ! trunc_ln851_1_reg_971;
assign _075_ = ! trunc_ln851_reg_1122;
always @(posedge \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.clk )
\add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.bin_s1  <= _077_;
always @(posedge \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.clk )
\add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.ain_s1  <= _076_;
always @(posedge \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.clk )
\add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.sum_s1  <= _079_;
always @(posedge \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.clk )
\add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.carry_s1  <= _078_;
assign _077_ = \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.ce  ? \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.b [9:5] : \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.bin_s1 ;
assign _076_ = \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.ce  ? \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.a [9:5] : \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.ain_s1 ;
assign _078_ = \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.ce  ? \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.facout_s1  : \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.carry_s1 ;
assign _079_ = \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.ce  ? \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.fas_s1  : \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.sum_s1 ;
assign _080_ = \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.u1.a  + \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.u1.b ;
assign { \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.u1.cout , \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.u1.s  } = _080_ + \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.u1.cin ;
assign _081_ = \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.u2.a  + \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.u2.b ;
assign { \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.u2.cout , \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.u2.s  } = _081_ + \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.u2.cin ;
always @(posedge \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.clk )
\add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.bin_s1  <= _083_;
always @(posedge \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.clk )
\add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.ain_s1  <= _082_;
always @(posedge \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.clk )
\add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.sum_s1  <= _085_;
always @(posedge \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.clk )
\add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.carry_s1  <= _084_;
assign _083_ = \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.ce  ? \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.b [14:7] : \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.bin_s1 ;
assign _082_ = \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.ce  ? \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.a [14:7] : \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.ain_s1 ;
assign _084_ = \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.ce  ? \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.facout_s1  : \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.carry_s1 ;
assign _085_ = \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.ce  ? \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.fas_s1  : \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.sum_s1 ;
assign _086_ = \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.u1.a  + \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.u1.b ;
assign { \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.u1.cout , \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.u1.s  } = _086_ + \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.u1.cin ;
assign _087_ = \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.u2.a  + \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.u2.b ;
assign { \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.u2.cout , \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.u2.s  } = _087_ + \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.u2.cin ;
always @(posedge \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.clk )
\add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.bin_s1  <= _089_;
always @(posedge \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.clk )
\add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.ain_s1  <= _088_;
always @(posedge \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.clk )
\add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.sum_s1  <= _091_;
always @(posedge \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.clk )
\add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.carry_s1  <= _090_;
assign _089_ = \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.ce  ? \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.b [16:8] : \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.bin_s1 ;
assign _088_ = \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.ce  ? \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.a [16:8] : \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.ain_s1 ;
assign _090_ = \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.ce  ? \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.facout_s1  : \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.carry_s1 ;
assign _091_ = \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.ce  ? \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.fas_s1  : \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.sum_s1 ;
assign _092_ = \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.u1.a  + \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.u1.b ;
assign { \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.u1.cout , \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.u1.s  } = _092_ + \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.u1.cin ;
assign _093_ = \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.u2.a  + \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.u2.b ;
assign { \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.u2.cout , \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.u2.s  } = _093_ + \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.u2.cin ;
always @(posedge \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.clk )
\add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.bin_s1  <= _095_;
always @(posedge \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.clk )
\add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.ain_s1  <= _094_;
always @(posedge \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.clk )
\add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.sum_s1  <= _097_;
always @(posedge \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.clk )
\add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.carry_s1  <= _096_;
assign _095_ = \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.ce  ? \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.b [1] : \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.bin_s1 ;
assign _094_ = \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.ce  ? \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.a [1] : \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.ain_s1 ;
assign _096_ = \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.ce  ? \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.facout_s1  : \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.carry_s1 ;
assign _097_ = \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.ce  ? \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.fas_s1  : \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.sum_s1 ;
assign _098_ = \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.a  + \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.b ;
assign { \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.cout , \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.s  } = _098_ + \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.cin ;
assign _099_ = \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.a  + \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.b ;
assign { \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.cout , \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.s  } = _099_ + \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.cin ;
always @(posedge \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.clk )
\add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.bin_s1  <= _101_;
always @(posedge \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.clk )
\add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.ain_s1  <= _100_;
always @(posedge \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.clk )
\add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.sum_s1  <= _103_;
always @(posedge \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.clk )
\add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.carry_s1  <= _102_;
assign _101_ = \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.ce  ? \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.b [1] : \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.bin_s1 ;
assign _100_ = \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.ce  ? \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.a [1] : \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.ain_s1 ;
assign _102_ = \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.ce  ? \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.facout_s1  : \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.carry_s1 ;
assign _103_ = \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.ce  ? \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.fas_s1  : \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.sum_s1 ;
assign _104_ = \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.a  + \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.b ;
assign { \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.cout , \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.s  } = _104_ + \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.cin ;
assign _105_ = \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.a  + \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.b ;
assign { \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.cout , \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.s  } = _105_ + \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.cin ;
always @(posedge \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.clk )
\add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.bin_s1  <= _107_;
always @(posedge \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.clk )
\add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.ain_s1  <= _106_;
always @(posedge \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.clk )
\add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.sum_s1  <= _109_;
always @(posedge \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.clk )
\add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.carry_s1  <= _108_;
assign _107_ = \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.ce  ? \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.b [1] : \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.bin_s1 ;
assign _106_ = \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.ce  ? \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.a [1] : \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.ain_s1 ;
assign _108_ = \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.ce  ? \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.facout_s1  : \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.carry_s1 ;
assign _109_ = \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.ce  ? \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.fas_s1  : \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.sum_s1 ;
assign _110_ = \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.a  + \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.b ;
assign { \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.cout , \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.s  } = _110_ + \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.cin ;
assign _111_ = \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.a  + \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.b ;
assign { \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.cout , \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.s  } = _111_ + \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.cin ;
always @(posedge \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.clk )
\add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.bin_s1  <= _113_;
always @(posedge \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.clk )
\add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.ain_s1  <= _112_;
always @(posedge \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.clk )
\add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.sum_s1  <= _115_;
always @(posedge \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.clk )
\add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.carry_s1  <= _114_;
assign _113_ = \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.ce  ? \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.b [2:1] : \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.bin_s1 ;
assign _112_ = \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.ce  ? \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.a [2:1] : \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.ain_s1 ;
assign _114_ = \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.ce  ? \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.facout_s1  : \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.carry_s1 ;
assign _115_ = \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.ce  ? \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.fas_s1  : \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.sum_s1 ;
assign _116_ = \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.u1.a  + \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.u1.b ;
assign { \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.u1.cout , \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.u1.s  } = _116_ + \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.u1.cin ;
assign _117_ = \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.u2.a  + \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.u2.b ;
assign { \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.u2.cout , \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.u2.s  } = _117_ + \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.u2.cin ;
always @(posedge \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.clk )
\add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.bin_s1  <= _119_;
always @(posedge \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.clk )
\add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.ain_s1  <= _118_;
always @(posedge \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.clk )
\add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.sum_s1  <= _121_;
always @(posedge \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.clk )
\add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.carry_s1  <= _120_;
assign _119_ = \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.ce  ? \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.b [2:1] : \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.bin_s1 ;
assign _118_ = \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.ce  ? \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.a [2:1] : \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.ain_s1 ;
assign _120_ = \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.ce  ? \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.facout_s1  : \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.carry_s1 ;
assign _121_ = \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.ce  ? \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.fas_s1  : \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.sum_s1 ;
assign _122_ = \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.u1.a  + \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.u1.b ;
assign { \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.u1.cout , \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.u1.s  } = _122_ + \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.u1.cin ;
assign _123_ = \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.u2.a  + \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.u2.b ;
assign { \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.u2.cout , \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.u2.s  } = _123_ + \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.u2.cin ;
always @(posedge \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.clk )
\add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.bin_s1  <= _125_;
always @(posedge \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.clk )
\add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.ain_s1  <= _124_;
always @(posedge \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.clk )
\add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.sum_s1  <= _127_;
always @(posedge \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.clk )
\add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.carry_s1  <= _126_;
assign _125_ = \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.ce  ? \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.b [3:2] : \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.bin_s1 ;
assign _124_ = \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.ce  ? \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.a [3:2] : \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.ain_s1 ;
assign _126_ = \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.ce  ? \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.facout_s1  : \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.carry_s1 ;
assign _127_ = \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.ce  ? \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.fas_s1  : \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.sum_s1 ;
assign _128_ = \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.u1.a  + \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.u1.b ;
assign { \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.u1.cout , \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.u1.s  } = _128_ + \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.u1.cin ;
assign _129_ = \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.u2.a  + \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.u2.b ;
assign { \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.u2.cout , \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.u2.s  } = _129_ + \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.u2.cin ;
always @(posedge \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.clk )
\add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.bin_s1  <= _131_;
always @(posedge \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.clk )
\add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.ain_s1  <= _130_;
always @(posedge \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.clk )
\add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.sum_s1  <= _133_;
always @(posedge \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.clk )
\add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.carry_s1  <= _132_;
assign _131_ = \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.ce  ? \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.b [4:2] : \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.bin_s1 ;
assign _130_ = \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.ce  ? \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.a [4:2] : \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.ain_s1 ;
assign _132_ = \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.ce  ? \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.facout_s1  : \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.carry_s1 ;
assign _133_ = \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.ce  ? \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.fas_s1  : \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.sum_s1 ;
assign _134_ = \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.u1.a  + \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.u1.b ;
assign { \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.u1.cout , \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.u1.s  } = _134_ + \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.u1.cin ;
assign _135_ = \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.u2.a  + \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.u2.b ;
assign { \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.u2.cout , \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.u2.s  } = _135_ + \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.u2.cin ;
always @(posedge \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.clk )
\add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.bin_s1  <= _137_;
always @(posedge \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.clk )
\add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.ain_s1  <= _136_;
always @(posedge \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.clk )
\add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.sum_s1  <= _139_;
always @(posedge \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.clk )
\add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.carry_s1  <= _138_;
assign _137_ = \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.ce  ? \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.b [5:3] : \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.bin_s1 ;
assign _136_ = \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.ce  ? \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.a [5:3] : \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.ain_s1 ;
assign _138_ = \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.ce  ? \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.facout_s1  : \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.carry_s1 ;
assign _139_ = \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.ce  ? \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.fas_s1  : \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.sum_s1 ;
assign _140_ = \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.u1.a  + \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.u1.b ;
assign { \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.u1.cout , \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.u1.s  } = _140_ + \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.u1.cin ;
assign _141_ = \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.u2.a  + \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.u2.b ;
assign { \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.u2.cout , \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.u2.s  } = _141_ + \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.u2.cin ;
always @(posedge \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.clk )
\add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.bin_s1  <= _143_;
always @(posedge \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.clk )
\add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.ain_s1  <= _142_;
always @(posedge \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.clk )
\add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.sum_s1  <= _145_;
always @(posedge \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.clk )
\add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.carry_s1  <= _144_;
assign _143_ = \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.ce  ? \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.b [5:3] : \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.bin_s1 ;
assign _142_ = \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.ce  ? \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.a [5:3] : \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.ain_s1 ;
assign _144_ = \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.ce  ? \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.facout_s1  : \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.carry_s1 ;
assign _145_ = \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.ce  ? \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.fas_s1  : \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.sum_s1 ;
assign _146_ = \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.u1.a  + \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.u1.b ;
assign { \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.u1.cout , \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.u1.s  } = _146_ + \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.u1.cin ;
assign _147_ = \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.u2.a  + \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.u2.b ;
assign { \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.u2.cout , \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.u2.s  } = _147_ + \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.u2.cin ;
always @(posedge \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.clk )
\add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.bin_s1  <= _149_;
always @(posedge \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.clk )
\add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.ain_s1  <= _148_;
always @(posedge \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.clk )
\add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.sum_s1  <= _151_;
always @(posedge \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.clk )
\add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.carry_s1  <= _150_;
assign _149_ = \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.ce  ? \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.b [5:3] : \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.bin_s1 ;
assign _148_ = \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.ce  ? \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.a [5:3] : \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.ain_s1 ;
assign _150_ = \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.ce  ? \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.facout_s1  : \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.carry_s1 ;
assign _151_ = \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.ce  ? \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.fas_s1  : \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.sum_s1 ;
assign _152_ = \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.u1.a  + \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.u1.b ;
assign { \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.u1.cout , \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.u1.s  } = _152_ + \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.u1.cin ;
assign _153_ = \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.u2.a  + \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.u2.b ;
assign { \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.u2.cout , \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.u2.s  } = _153_ + \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.u2.cin ;
always @(posedge \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.clk )
\add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.bin_s1  <= _155_;
always @(posedge \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.clk )
\add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.ain_s1  <= _154_;
always @(posedge \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.clk )
\add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.sum_s1  <= _157_;
always @(posedge \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.clk )
\add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.carry_s1  <= _156_;
assign _155_ = \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.ce  ? \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.b [5:3] : \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.bin_s1 ;
assign _154_ = \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.ce  ? \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.a [5:3] : \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.ain_s1 ;
assign _156_ = \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.ce  ? \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.facout_s1  : \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.carry_s1 ;
assign _157_ = \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.ce  ? \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.fas_s1  : \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.sum_s1 ;
assign _158_ = \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.u1.a  + \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.u1.b ;
assign { \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.u1.cout , \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.u1.s  } = _158_ + \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.u1.cin ;
assign _159_ = \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.u2.a  + \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.u2.b ;
assign { \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.u2.cout , \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.u2.s  } = _159_ + \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.u2.cin ;
always @(posedge \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.clk )
\add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.bin_s1  <= _161_;
always @(posedge \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.clk )
\add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.ain_s1  <= _160_;
always @(posedge \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.clk )
\add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.sum_s1  <= _163_;
always @(posedge \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.clk )
\add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.carry_s1  <= _162_;
assign _161_ = \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.ce  ? \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.b [5:3] : \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.bin_s1 ;
assign _160_ = \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.ce  ? \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.a [5:3] : \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.ain_s1 ;
assign _162_ = \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.ce  ? \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.facout_s1  : \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.carry_s1 ;
assign _163_ = \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.ce  ? \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.fas_s1  : \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.sum_s1 ;
assign _164_ = \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.u1.a  + \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.u1.b ;
assign { \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.u1.cout , \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.u1.s  } = _164_ + \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.u1.cin ;
assign _165_ = \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.u2.a  + \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.u2.b ;
assign { \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.u2.cout , \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.u2.s  } = _165_ + \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.u2.cin ;
assign \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.bin_s0  = ~ \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.b ;
always @(posedge \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.clk )
\sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.bin_s1  <= _167_;
always @(posedge \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.clk )
\sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.ain_s1  <= _166_;
always @(posedge \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.clk )
\sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.sum_s1  <= _169_;
always @(posedge \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.clk )
\sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.carry_s1  <= _168_;
assign _167_ = \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.ce  ? \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.bin_s0 [4:2] : \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.bin_s1 ;
assign _166_ = \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.ce  ? \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.a [4:2] : \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.ain_s1 ;
assign _168_ = \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.ce  ? \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.facout_s1  : \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.carry_s1 ;
assign _169_ = \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.ce  ? \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.fas_s1  : \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.sum_s1 ;
assign _170_ = \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.u1.a  + \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.u1.b ;
assign { \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.u1.cout , \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.u1.s  } = _170_ + \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.u1.cin ;
assign _171_ = \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.u2.a  + \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.u2.b ;
assign { \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.u2.cout , \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.u2.s  } = _171_ + \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.u2.cin ;
assign \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.bin_s0  = ~ \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.b ;
always @(posedge \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.clk )
\sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.bin_s1  <= _173_;
always @(posedge \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.clk )
\sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.ain_s1  <= _172_;
always @(posedge \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.clk )
\sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.sum_s1  <= _175_;
always @(posedge \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.clk )
\sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.carry_s1  <= _174_;
assign _173_ = \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.ce  ? \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.bin_s0 [8:4] : \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.bin_s1 ;
assign _172_ = \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.ce  ? \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.a [8:4] : \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.ain_s1 ;
assign _174_ = \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.ce  ? \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.facout_s1  : \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.carry_s1 ;
assign _175_ = \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.ce  ? \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.fas_s1  : \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.sum_s1 ;
assign _176_ = \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.u1.a  + \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.u1.b ;
assign { \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.u1.cout , \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.u1.s  } = _176_ + \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.u1.cin ;
assign _177_ = \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.u2.a  + \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.u2.b ;
assign { \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.u2.cout , \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.u2.s  } = _177_ + \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.u2.cin ;
assign _178_ = $signed(ret_V_19_reg_1157) > $signed({ 1'h0, ret_V_25_fu_665_p3 });
assign _179_ = | trunc_ln414_reg_999;
assign _180_ = | tmp_2_reg_1334;
assign _181_ = tmp_2_reg_1334 != 4'hf;
assign _182_ = | op_3[12:0];
assign _183_ = | op_14[4:0];
assign or_ln340_1_fu_897_p2 = underflow_1_reg_1364 | overflow_1_fu_892_p2;
assign or_ln340_2_fu_513_p2 = or_ln340_reg_1132 | neg_src_fu_508_p2;
assign or_ln340_fu_483_p2 = overflow_fu_477_p2 | and_ln786_reg_1104;
assign or_ln384_fu_876_p2 = xor_ln384_fu_871_p2 | p_Result_13_reg_1319;
assign or_ln388_fu_867_p2 = underflow_1_reg_1364 | newsignbit_reg_1326;
assign or_ln785_1_fu_843_p2 = newsignbit_reg_1326 | icmp_ln768_reg_1340;
assign or_ln785_2_fu_529_p2 = p_Result_10_reg_981 | and_ln785_fu_525_p2;
assign or_ln785_fu_467_p2 = xor_ln785_fu_462_p2 | p_Result_12_reg_1068;
assign or_ln786_fu_852_p2 = xor_ln786_fu_847_p2 | icmp_ln786_reg_1345;
assign ret_V_18_fu_432_p2 = op_3 | { op_1, 12'h000 };
assign ret_V_20_fu_239_p2 = $signed({ op_7, 2'h0 }) | $signed(op_2);
always @(posedge ap_clk)
select_ln69_reg_1309[5:2] <= 4'h0;
always @(posedge ap_clk)
xor_ln416_reg_1075 <= _063_;
always @(posedge ap_clk)
sext_ln850_reg_1277 <= _055_;
always @(posedge ap_clk)
select_ln340_reg_1142 <= _053_;
always @(posedge ap_clk)
ret_V_3_reg_1147 <= _048_;
always @(posedge ap_clk)
ret_V_28_reg_1380 <= _047_;
always @(posedge ap_clk)
select_ln1192_reg_1385 <= _052_;
always @(posedge ap_clk)
ret_V_27_reg_1289 <= _046_;
always @(posedge ap_clk)
ret_V_26_reg_1267 <= _045_;
always @(posedge ap_clk)
tmp_3_reg_1272 <= _057_;
always @(posedge ap_clk)
ret_V_20_reg_959 <= _040_;
always @(posedge ap_clk)
ret_V_4_cast_reg_964 <= _049_;
always @(posedge ap_clk)
trunc_ln851_1_reg_971 <= _060_;
always @(posedge ap_clk)
p_Val2_2_reg_1062 <= _036_;
always @(posedge ap_clk)
p_Result_12_reg_1068 <= _031_;
always @(posedge ap_clk)
or_ln785_1_reg_1358 <= _028_;
always @(posedge ap_clk)
underflow_1_reg_1364 <= _062_;
always @(posedge ap_clk)
op_5_V_reg_1152 <= _026_;
always @(posedge ap_clk)
ret_V_19_reg_1157 <= _039_;
always @(posedge ap_clk)
trunc_ln728_reg_1165 <= _059_;
always @(posedge ap_clk)
ret_V_24_reg_1232 <= _044_;
always @(posedge ap_clk)
op_22_V_reg_1242 <= _024_;
always @(posedge ap_clk)
p_Result_13_reg_1319 <= _032_;
always @(posedge ap_clk)
newsignbit_reg_1326 <= _023_;
always @(posedge ap_clk)
tmp_2_reg_1334 <= _056_;
always @(posedge ap_clk)
or_ln340_reg_1132 <= _027_;
always @(posedge ap_clk)
icmp_ln851_reg_1137 <= _021_;
always @(posedge ap_clk)
lhs_V_1_reg_1247 <= _022_;
always @(posedge ap_clk)
icmp_ln851_3_reg_1262 <= _020_;
always @(posedge ap_clk)
ret_V_17_reg_976 <= _037_;
always @(posedge ap_clk)
p_Result_10_reg_981 <= _029_;
always @(posedge ap_clk)
p_Val2_1_reg_989 <= _035_;
always @(posedge ap_clk)
p_Result_11_reg_994 <= _030_;
always @(posedge ap_clk)
trunc_ln414_reg_999 <= _058_;
always @(posedge ap_clk)
p_Result_s_reg_1004 <= _034_;
always @(posedge ap_clk)
p_Result_1_reg_1009 <= _033_;
always @(posedge ap_clk)
icmp_ln851_1_reg_1015 <= _018_;
always @(posedge ap_clk)
icmp_ln768_reg_1340 <= _016_;
always @(posedge ap_clk)
icmp_ln786_reg_1345 <= _017_;
always @(posedge ap_clk)
op_25_V_reg_1350 <= _025_;
always @(posedge ap_clk)
carry_1_reg_1081 <= _012_;
always @(posedge ap_clk)
empty_reg_1093 <= _014_;
always @(posedge ap_clk)
deleted_zeros_reg_1098 <= _013_;
always @(posedge ap_clk)
and_ln786_reg_1104 <= _010_;
always @(posedge ap_clk)
ret_V_18_reg_1110 <= _038_;
always @(posedge ap_clk)
ret_V_reg_1115 <= _051_;
always @(posedge ap_clk)
trunc_ln851_reg_1122 <= _061_;
always @(posedge ap_clk)
icmp_ln851_2_reg_1127 <= _019_;
always @(posedge ap_clk)
and_ln414_reg_1047 <= _009_;
always @(posedge ap_clk)
ret_V_21_reg_1052 <= _042_;
always @(posedge ap_clk)
and_ln384_reg_1370 <= _008_;
always @(posedge ap_clk)
ret_V_23_reg_1195 <= _043_;
always @(posedge ap_clk)
ret_V_21_cast_reg_1200 <= _041_;
always @(posedge ap_clk)
add_ln69_reg_1207 <= _007_;
always @(posedge ap_clk)
select_ln69_reg_1309[1:0] <= _054_;
always @(posedge ap_clk)
add_ln69_2_reg_1314 <= _006_;
always @(posedge ap_clk)
add_ln691_reg_1237 <= _005_;
always @(posedge ap_clk)
add_ln691_2_reg_1375 <= _004_;
always @(posedge ap_clk)
add_ln691_1_reg_1284 <= _003_;
always @(posedge ap_clk)
icmp_ln414_reg_1020 <= _015_;
always @(posedge ap_clk)
Range2_all_ones_reg_1025 <= _002_;
always @(posedge ap_clk)
Range1_all_ones_reg_1030 <= _000_;
always @(posedge ap_clk)
Range1_all_zeros_reg_1037 <= _001_;
always @(posedge ap_clk)
ret_V_6_reg_1042 <= _050_;
always @(posedge ap_clk)
ap_CS_fsm <= _011_;
assign _064_ = _069_ ? 2'h2 : 2'h1;
assign _184_ = ap_CS_fsm == 1'h1;
function [29:0] _536_;
input [29:0] a;
input [899:0] b;
input [29:0] s;
case (s)
30'b000000000000000000000000000001:
_536_ = b[29:0];
30'b000000000000000000000000000010:
_536_ = b[59:30];
30'b000000000000000000000000000100:
_536_ = b[89:60];
30'b000000000000000000000000001000:
_536_ = b[119:90];
30'b000000000000000000000000010000:
_536_ = b[149:120];
30'b000000000000000000000000100000:
_536_ = b[179:150];
30'b000000000000000000000001000000:
_536_ = b[209:180];
30'b000000000000000000000010000000:
_536_ = b[239:210];
30'b000000000000000000000100000000:
_536_ = b[269:240];
30'b000000000000000000001000000000:
_536_ = b[299:270];
30'b000000000000000000010000000000:
_536_ = b[329:300];
30'b000000000000000000100000000000:
_536_ = b[359:330];
30'b000000000000000001000000000000:
_536_ = b[389:360];
30'b000000000000000010000000000000:
_536_ = b[419:390];
30'b000000000000000100000000000000:
_536_ = b[449:420];
30'b000000000000001000000000000000:
_536_ = b[479:450];
30'b000000000000010000000000000000:
_536_ = b[509:480];
30'b000000000000100000000000000000:
_536_ = b[539:510];
30'b000000000001000000000000000000:
_536_ = b[569:540];
30'b000000000010000000000000000000:
_536_ = b[599:570];
30'b000000000100000000000000000000:
_536_ = b[629:600];
30'b000000001000000000000000000000:
_536_ = b[659:630];
30'b000000010000000000000000000000:
_536_ = b[689:660];
30'b000000100000000000000000000000:
_536_ = b[719:690];
30'b000001000000000000000000000000:
_536_ = b[749:720];
30'b000010000000000000000000000000:
_536_ = b[779:750];
30'b000100000000000000000000000000:
_536_ = b[809:780];
30'b001000000000000000000000000000:
_536_ = b[839:810];
30'b010000000000000000000000000000:
_536_ = b[869:840];
30'b100000000000000000000000000000:
_536_ = b[899:870];
30'b000000000000000000000000000000:
_536_ = a;
default:
_536_ = 30'bx;
endcase
endfunction
assign ap_NS_fsm = _536_(30'hxxxxxxxx, { 28'h0000000, _064_, 870'h00000004000000200000010000000800000040000002000000100000008000000400000020000001000000080000004000000200000010000000800000040000002000000100000008000000400000020000001000000080000004000000200000010000000800000000000001 }, { _184_, _213_, _212_, _211_, _210_, _209_, _208_, _207_, _206_, _205_, _204_, _203_, _202_, _201_, _200_, _199_, _198_, _197_, _196_, _195_, _194_, _193_, _192_, _191_, _190_, _189_, _188_, _187_, _186_, _185_ });
assign _185_ = ap_CS_fsm == 30'h20000000;
assign _186_ = ap_CS_fsm == 29'h10000000;
assign _187_ = ap_CS_fsm == 28'h8000000;
assign _188_ = ap_CS_fsm == 27'h4000000;
assign _189_ = ap_CS_fsm == 26'h2000000;
assign _190_ = ap_CS_fsm == 25'h1000000;
assign _191_ = ap_CS_fsm == 24'h800000;
assign _192_ = ap_CS_fsm == 23'h400000;
assign _193_ = ap_CS_fsm == 22'h200000;
assign _194_ = ap_CS_fsm == 21'h100000;
assign _195_ = ap_CS_fsm == 20'h80000;
assign _196_ = ap_CS_fsm == 19'h40000;
assign _197_ = ap_CS_fsm == 18'h20000;
assign _198_ = ap_CS_fsm == 17'h10000;
assign _199_ = ap_CS_fsm == 16'h8000;
assign _200_ = ap_CS_fsm == 15'h4000;
assign _201_ = ap_CS_fsm == 14'h2000;
assign _202_ = ap_CS_fsm == 13'h1000;
assign _203_ = ap_CS_fsm == 12'h800;
assign _204_ = ap_CS_fsm == 11'h400;
assign _205_ = ap_CS_fsm == 10'h200;
assign _206_ = ap_CS_fsm == 9'h100;
assign _207_ = ap_CS_fsm == 8'h80;
assign _208_ = ap_CS_fsm == 7'h40;
assign _209_ = ap_CS_fsm == 6'h20;
assign _210_ = ap_CS_fsm == 5'h10;
assign _211_ = ap_CS_fsm == 4'h8;
assign _212_ = ap_CS_fsm == 3'h4;
assign _213_ = ap_CS_fsm == 2'h2;
assign op_28_ap_vld = ap_CS_fsm[29] ? 1'h1 : 1'h0;
assign ap_idle = _068_ ? 1'h1 : 1'h0;
assign _063_ = ap_CS_fsm[6] ? xor_ln416_fu_378_p2 : xor_ln416_reg_1075;
assign _055_ = ap_CS_fsm[18] ? { tmp_3_reg_1272[4], tmp_3_reg_1272 } : sext_ln850_reg_1277;
assign _048_ = ap_CS_fsm[10] ? grp_fu_493_p2 : ret_V_3_reg_1147;
assign _053_ = ap_CS_fsm[10] ? select_ln340_fu_518_p3 : select_ln340_reg_1142;
assign _052_ = ap_CS_fsm[27] ? select_ln1192_fu_927_p3 : select_ln1192_reg_1385;
assign _047_ = ap_CS_fsm[27] ? ret_V_28_fu_920_p3 : ret_V_28_reg_1380;
assign _046_ = ap_CS_fsm[20] ? ret_V_27_fu_739_p3 : ret_V_27_reg_1289;
assign _057_ = ap_CS_fsm[17] ? grp_fu_692_p2[9:5] : tmp_3_reg_1272;
assign _045_ = ap_CS_fsm[17] ? grp_fu_692_p2 : ret_V_26_reg_1267;
assign _060_ = ap_CS_fsm[0] ? ret_V_20_fu_239_p2[1:0] : trunc_ln851_1_reg_971;
assign _049_ = ap_CS_fsm[0] ? ret_V_20_fu_239_p2[3:2] : ret_V_4_cast_reg_964;
assign _040_ = ap_CS_fsm[0] ? ret_V_20_fu_239_p2 : ret_V_20_reg_959;
assign _031_ = ap_CS_fsm[5] ? grp_fu_365_p2[1] : p_Result_12_reg_1068;
assign _036_ = ap_CS_fsm[5] ? grp_fu_365_p2 : p_Val2_2_reg_1062;
assign _062_ = ap_CS_fsm[25] ? underflow_1_fu_857_p2 : underflow_1_reg_1364;
assign _028_ = ap_CS_fsm[25] ? or_ln785_1_fu_843_p2 : or_ln785_1_reg_1358;
assign _059_ = ap_CS_fsm[11] ? ret_V_19_fu_557_p3[1:0] : trunc_ln728_reg_1165;
assign _039_ = ap_CS_fsm[11] ? ret_V_19_fu_557_p3 : ret_V_19_reg_1157;
assign _026_ = ap_CS_fsm[11] ? op_5_V_fu_539_p3 : op_5_V_reg_1152;
assign _024_ = ap_CS_fsm[15] ? grp_fu_647_p2 : op_22_V_reg_1242;
assign _044_ = ap_CS_fsm[15] ? grp_fu_633_p2 : ret_V_24_reg_1232;
assign _056_ = ap_CS_fsm[23] ? grp_fu_793_p2[4:1] : tmp_2_reg_1334;
assign _023_ = ap_CS_fsm[23] ? grp_fu_793_p2[0] : newsignbit_reg_1326;
assign _032_ = ap_CS_fsm[23] ? grp_fu_793_p2[4] : p_Result_13_reg_1319;
assign _021_ = ap_CS_fsm[9] ? icmp_ln851_fu_488_p2 : icmp_ln851_reg_1137;
assign _027_ = ap_CS_fsm[9] ? or_ln340_fu_483_p2 : or_ln340_reg_1132;
assign _020_ = ap_CS_fsm[16] ? icmp_ln851_3_fu_702_p2 : icmp_ln851_3_reg_1262;
assign _022_ = ap_CS_fsm[16] ? lhs_V_1_fu_676_p2 : lhs_V_1_reg_1247;
assign _018_ = ap_CS_fsm[1] ? icmp_ln851_1_fu_309_p2 : icmp_ln851_1_reg_1015;
assign _033_ = ap_CS_fsm[1] ? grp_fu_221_p2[8:4] : p_Result_1_reg_1009;
assign _034_ = ap_CS_fsm[1] ? grp_fu_221_p2[8:5] : p_Result_s_reg_1004;
assign _058_ = ap_CS_fsm[1] ? grp_fu_221_p2[1:0] : trunc_ln414_reg_999;
assign _030_ = ap_CS_fsm[1] ? grp_fu_221_p2[3] : p_Result_11_reg_994;
assign _035_ = ap_CS_fsm[1] ? grp_fu_221_p2[3:2] : p_Val2_1_reg_989;
assign _029_ = ap_CS_fsm[1] ? grp_fu_221_p2[8] : p_Result_10_reg_981;
assign _037_ = ap_CS_fsm[1] ? grp_fu_221_p2 : ret_V_17_reg_976;
assign _025_ = ap_CS_fsm[24] ? grp_fu_829_p2 : op_25_V_reg_1350;
assign _017_ = ap_CS_fsm[24] ? icmp_ln786_fu_838_p2 : icmp_ln786_reg_1345;
assign _016_ = ap_CS_fsm[24] ? icmp_ln768_fu_833_p2 : icmp_ln768_reg_1340;
assign _012_ = ap_CS_fsm[7] ? carry_1_fu_383_p2 : carry_1_reg_1081;
assign _019_ = ap_CS_fsm[8] ? icmp_ln851_2_fu_456_p2 : icmp_ln851_2_reg_1127;
assign _061_ = ap_CS_fsm[8] ? ret_V_18_fu_432_p2[12:0] : trunc_ln851_reg_1122;
assign _051_ = ap_CS_fsm[8] ? ret_V_18_fu_432_p2[15:13] : ret_V_reg_1115;
assign _038_ = ap_CS_fsm[8] ? ret_V_18_fu_432_p2 : ret_V_18_reg_1110;
assign _010_ = ap_CS_fsm[8] ? and_ln786_fu_420_p2 : and_ln786_reg_1104;
assign _013_ = ap_CS_fsm[8] ? deleted_zeros_fu_391_p3 : deleted_zeros_reg_1098;
assign _014_ = ap_CS_fsm[8] ? op_3[14:0] : empty_reg_1093;
assign _042_ = ap_CS_fsm[3] ? ret_V_21_fu_355_p3 : ret_V_21_reg_1052;
assign _009_ = ap_CS_fsm[3] ? and_ln414_fu_339_p2 : and_ln414_reg_1047;
assign _008_ = ap_CS_fsm[26] ? and_ln384_fu_881_p2 : and_ln384_reg_1370;
assign _007_ = ap_CS_fsm[13] ? grp_fu_600_p2 : add_ln69_reg_1207;
assign _041_ = ap_CS_fsm[13] ? grp_fu_591_p2[14:13] : ret_V_21_cast_reg_1200;
assign _043_ = ap_CS_fsm[13] ? grp_fu_578_p2 : ret_V_23_reg_1195;
assign _006_ = ap_CS_fsm[22] ? grp_fu_749_p2 : add_ln69_2_reg_1314;
assign _054_ = ap_CS_fsm[22] ? select_ln69_fu_799_p3 : select_ln69_reg_1309[1:0];
assign _005_ = _067_ ? grp_fu_639_p2 : add_ln691_reg_1237;
assign _004_ = _066_ ? grp_fu_862_p2 : add_ln691_2_reg_1375;
assign _003_ = _065_ ? grp_fu_721_p2 : add_ln691_1_reg_1284;
assign _050_ = ap_CS_fsm[2] ? grp_fu_314_p2 : ret_V_6_reg_1042;
assign _001_ = ap_CS_fsm[2] ? Range1_all_zeros_fu_334_p2 : Range1_all_zeros_reg_1037;
assign _000_ = ap_CS_fsm[2] ? Range1_all_ones_fu_329_p2 : Range1_all_ones_reg_1030;
assign _002_ = ap_CS_fsm[2] ? Range2_all_ones_fu_324_p2 : Range2_all_ones_reg_1025;
assign _015_ = ap_CS_fsm[2] ? icmp_ln414_fu_319_p2 : icmp_ln414_reg_1020;
assign _011_ = ap_rst ? 30'h00000001 : ap_NS_fsm;
assign Range1_all_ones_fu_329_p2 = _071_ ? 1'h1 : 1'h0;
assign Range1_all_zeros_fu_334_p2 = _072_ ? 1'h1 : 1'h0;
assign Range2_all_ones_fu_324_p2 = _073_ ? 1'h1 : 1'h0;
assign deleted_ones_fu_414_p3 = carry_1_reg_1081 ? and_ln780_fu_409_p2 : Range1_all_ones_reg_1030;
assign deleted_zeros_fu_391_p3 = carry_1_reg_1081 ? Range1_all_ones_reg_1030 : Range1_all_zeros_reg_1037;
assign icmp_ln414_fu_319_p2 = _179_ ? 1'h1 : 1'h0;
assign icmp_ln768_fu_833_p2 = _180_ ? 1'h1 : 1'h0;
assign icmp_ln786_fu_838_p2 = _181_ ? 1'h1 : 1'h0;
assign icmp_ln851_1_fu_309_p2 = _074_ ? 1'h1 : 1'h0;
assign icmp_ln851_2_fu_456_p2 = _182_ ? 1'h1 : 1'h0;
assign icmp_ln851_3_fu_702_p2 = _183_ ? 1'h1 : 1'h0;
assign icmp_ln851_fu_488_p2 = _075_ ? 1'h1 : 1'h0;
assign lhs_V_1_fu_676_p2 = _178_ ? 1'h1 : 1'h0;
assign op_19_V_fu_902_p3 = or_ln340_1_fu_897_p2 ? and_ln384_reg_1370 : newsignbit_reg_1326;
assign op_5_V_fu_539_p3 = and_ln785_1_fu_534_p2 ? p_Val2_2_reg_1062 : select_ln340_reg_1142;
assign ret_V_19_fu_557_p3 = ret_V_18_reg_1110[15] ? select_ln850_fu_552_p3 : ret_V_reg_1115;
assign ret_V_21_fu_355_p3 = ret_V_20_reg_959[7] ? select_ln850_1_fu_350_p3 : ret_V_4_cast_reg_964;
assign ret_V_25_fu_665_p3 = ret_V_24_reg_1232[16] ? select_ln850_2_fu_660_p3 : ret_V_21_cast_reg_1200;
assign ret_V_27_fu_739_p3 = ret_V_26_reg_1267[9] ? select_ln850_3_fu_734_p3 : sext_ln850_reg_1277;
assign ret_V_28_fu_920_p3 = op_25_V_reg_1350[5] ? select_ln850_4_fu_915_p3 : { 1'h0, op_25_V_reg_1350[4:0] };
assign select_ln1192_fu_927_p3 = op_19_V_fu_902_p3 ? 6'h3f : 6'h00;
assign select_ln340_fu_518_p3 = or_ln340_2_fu_513_p2 ? 2'h0 : p_Val2_2_reg_1062;
assign select_ln69_fu_799_p3 = ret_V_22_fu_780_p2 ? 2'h2 : 2'h1;
assign select_ln850_1_fu_350_p3 = icmp_ln851_1_reg_1015 ? ret_V_4_cast_reg_964 : ret_V_6_reg_1042;
assign select_ln850_2_fu_660_p3 = icmp_ln851_2_reg_1127 ? add_ln691_reg_1237 : ret_V_21_cast_reg_1200;
assign select_ln850_3_fu_734_p3 = icmp_ln851_3_reg_1262 ? add_ln691_1_reg_1284 : sext_ln850_reg_1277;
assign select_ln850_4_fu_915_p3 = lhs_V_1_reg_1247 ? add_ln691_2_reg_1375 : { 1'h1, op_25_V_reg_1350[4:0] };
assign select_ln850_fu_552_p3 = icmp_ln851_reg_1137 ? ret_V_reg_1115 : ret_V_3_reg_1147;
assign ret_V_22_fu_780_p2 = op_8[1] ^ and_ln850_fu_774_p2;
assign ap_CS_fsm_state1 = ap_CS_fsm[0];
assign ap_CS_fsm_state10 = ap_CS_fsm[9];
assign ap_CS_fsm_state11 = ap_CS_fsm[10];
assign ap_CS_fsm_state12 = ap_CS_fsm[11];
assign ap_CS_fsm_state13 = ap_CS_fsm[12];
assign ap_CS_fsm_state14 = ap_CS_fsm[13];
assign ap_CS_fsm_state15 = ap_CS_fsm[14];
assign ap_CS_fsm_state16 = ap_CS_fsm[15];
assign ap_CS_fsm_state17 = ap_CS_fsm[16];
assign ap_CS_fsm_state18 = ap_CS_fsm[17];
assign ap_CS_fsm_state19 = ap_CS_fsm[18];
assign ap_CS_fsm_state2 = ap_CS_fsm[1];
assign ap_CS_fsm_state20 = ap_CS_fsm[19];
assign ap_CS_fsm_state21 = ap_CS_fsm[20];
assign ap_CS_fsm_state22 = ap_CS_fsm[21];
assign ap_CS_fsm_state23 = ap_CS_fsm[22];
assign ap_CS_fsm_state24 = ap_CS_fsm[23];
assign ap_CS_fsm_state25 = ap_CS_fsm[24];
assign ap_CS_fsm_state26 = ap_CS_fsm[25];
assign ap_CS_fsm_state27 = ap_CS_fsm[26];
assign ap_CS_fsm_state28 = ap_CS_fsm[27];
assign ap_CS_fsm_state29 = ap_CS_fsm[28];
assign ap_CS_fsm_state3 = ap_CS_fsm[2];
assign ap_CS_fsm_state30 = ap_CS_fsm[29];
assign ap_CS_fsm_state4 = ap_CS_fsm[3];
assign ap_CS_fsm_state5 = ap_CS_fsm[4];
assign ap_CS_fsm_state6 = ap_CS_fsm[5];
assign ap_CS_fsm_state7 = ap_CS_fsm[6];
assign ap_CS_fsm_state8 = ap_CS_fsm[7];
assign ap_CS_fsm_state9 = ap_CS_fsm[8];
assign ap_done = op_28_ap_vld;
assign ap_ready = op_28_ap_vld;
assign empty_fu_387_p0 = op_3;
assign empty_fu_387_p1 = op_3[14:0];
assign grp_fu_221_p0 = { op_1[3], op_1[3], op_1[3], op_1[3], op_1, 1'h0 };
assign grp_fu_221_p1 = { op_2[7], op_2 };
assign grp_fu_365_p1 = { 1'h0, and_ln414_reg_1047 };
assign grp_fu_578_p0 = { op_5_V_reg_1152[1], op_5_V_reg_1152 };
assign grp_fu_578_p1 = { op_0[1], op_0 };
assign grp_fu_591_p0 = { trunc_ln728_reg_1165, 13'h0000 };
assign grp_fu_600_p0 = { ret_V_19_reg_1157[2], ret_V_19_reg_1157 };
assign grp_fu_600_p1 = { 2'h0, op_12 };
assign grp_fu_633_p0 = { ret_V_19_reg_1157[2], ret_V_19_reg_1157, 13'h0000 };
assign grp_fu_633_p1 = { op_3[15], op_3 };
assign grp_fu_647_p0 = { add_ln69_reg_1207[3], add_ln69_reg_1207 };
assign grp_fu_647_p1 = { ret_V_23_reg_1195[2], ret_V_23_reg_1195[2], ret_V_23_reg_1195 };
assign grp_fu_692_p0 = { op_22_V_reg_1242, 5'h00 };
assign grp_fu_692_p1 = { op_14[7], op_14[7], op_14 };
assign grp_fu_721_p0 = { tmp_3_reg_1272[4], tmp_3_reg_1272 };
assign grp_fu_749_p1 = { ret_V_21_reg_1052[1], ret_V_21_reg_1052[1], ret_V_21_reg_1052[1], ret_V_21_reg_1052[1], ret_V_21_reg_1052 };
assign grp_fu_793_p0 = { ret_V_19_reg_1157[2], ret_V_19_reg_1157[2], ret_V_19_reg_1157 };
assign grp_fu_793_p1 = { op_13[3], op_13 };
assign lhs_1_fu_425_p3 = { op_1, 12'h000 };
assign lhs_fu_205_p3 = { op_1, 1'h0 };
assign newsignbit_fu_815_p1 = grp_fu_793_p2[0];
assign op_28 = { grp_fu_935_p2[5], grp_fu_935_p2[5], grp_fu_935_p2[5], grp_fu_935_p2[5], grp_fu_935_p2[5], grp_fu_935_p2[5], grp_fu_935_p2[5], grp_fu_935_p2[5], grp_fu_935_p2[5], grp_fu_935_p2[5], grp_fu_935_p2[5], grp_fu_935_p2[5], grp_fu_935_p2[5], grp_fu_935_p2[5], grp_fu_935_p2[5], grp_fu_935_p2[5], grp_fu_935_p2[5], grp_fu_935_p2[5], grp_fu_935_p2[5], grp_fu_935_p2[5], grp_fu_935_p2[5], grp_fu_935_p2[5], grp_fu_935_p2[5], grp_fu_935_p2[5], grp_fu_935_p2[5], grp_fu_935_p2[5], grp_fu_935_p2 };
assign p_Result_2_fu_343_p3 = ret_V_20_reg_959[7];
assign p_Result_3_fu_762_p3 = op_8[1];
assign p_Result_5_fu_653_p3 = ret_V_24_reg_1232[16];
assign p_Result_8_fu_727_p3 = ret_V_26_reg_1267[9];
assign p_Result_9_fu_908_p3 = op_25_V_reg_1350[5];
assign p_Result_s_16_fu_545_p3 = ret_V_18_reg_1110[15];
assign ret_V_18_fu_432_p1 = op_3;
assign ret_V_20_fu_239_p1 = op_2;
assign ret_V_8_fu_754_p3 = op_8[1];
assign rhs_3_fu_622_p3 = { ret_V_19_reg_1157, 13'h0000 };
assign rhs_fu_227_p3 = { op_7, 2'h0 };
assign sext_ln1192_2_fu_681_p0 = op_14;
assign sext_ln1192_fu_619_p0 = op_3;
assign sext_ln1195_fu_235_p1 = { op_7[1], op_7[1], op_7[1], op_7[1], op_7, 2'h0 };
assign sext_ln703_fu_217_p0 = op_2;
assign sext_ln850_fu_718_p1 = { tmp_3_reg_1272[4], tmp_3_reg_1272 };
assign tmp_fu_396_p3 = ret_V_17_reg_976[4];
assign trunc_ln414_fu_285_p1 = grp_fu_221_p2[1:0];
assign trunc_ln728_fu_564_p1 = ret_V_19_fu_557_p3[1:0];
assign trunc_ln851_1_fu_255_p1 = ret_V_20_fu_239_p2[1:0];
assign trunc_ln851_2_fu_770_p1 = op_8[0];
assign trunc_ln851_3_fu_452_p0 = op_3;
assign trunc_ln851_3_fu_452_p1 = op_3[12:0];
assign trunc_ln851_4_fu_698_p0 = op_14;
assign trunc_ln851_4_fu_698_p1 = op_14[4:0];
assign trunc_ln851_fu_448_p1 = ret_V_18_fu_432_p2[12:0];
assign zext_ln886_fu_672_p1 = { 1'h0, ret_V_25_fu_665_p3 };
assign \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.ain_s0  = \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.a ;
assign \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.s  = { \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.fas_s2 , \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.sum_s1  };
assign \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.u2.a  = \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.ain_s1 ;
assign \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.u2.b  = \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.bin_s1 ;
assign \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.u2.cin  = \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.carry_s1 ;
assign \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.facout_s2  = \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.u2.cout ;
assign \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.fas_s2  = \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.u2.s ;
assign \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.u1.a  = \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.a [3:0];
assign \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.u1.b  = \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.bin_s0 [3:0];
assign \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.u1.cin  = 1'h1;
assign \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.facout_s1  = \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.u1.cout ;
assign \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.fas_s1  = \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.u1.s ;
assign \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.a  = \sub_9s_9s_9_2_1_U1.din0 ;
assign \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.b  = \sub_9s_9s_9_2_1_U1.din1 ;
assign \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.ce  = \sub_9s_9s_9_2_1_U1.ce ;
assign \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.clk  = \sub_9s_9s_9_2_1_U1.clk ;
assign \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.reset  = \sub_9s_9s_9_2_1_U1.reset ;
assign \sub_9s_9s_9_2_1_U1.dout  = \sub_9s_9s_9_2_1_U1.top_sub_9s_9s_9_2_1_Adder_0_U.s ;
assign \sub_9s_9s_9_2_1_U1.ce  = 1'h1;
assign \sub_9s_9s_9_2_1_U1.clk  = ap_clk;
assign \sub_9s_9s_9_2_1_U1.din0  = { op_1[3], op_1[3], op_1[3], op_1[3], op_1, 1'h0 };
assign \sub_9s_9s_9_2_1_U1.din1  = { op_2[7], op_2 };
assign grp_fu_221_p2 = \sub_9s_9s_9_2_1_U1.dout ;
assign \sub_9s_9s_9_2_1_U1.reset  = ap_rst;
assign \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.ain_s0  = \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.a ;
assign \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.s  = { \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.fas_s2 , \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.sum_s1  };
assign \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.u2.a  = \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.ain_s1 ;
assign \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.u2.b  = \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.bin_s1 ;
assign \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.u2.cin  = \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.carry_s1 ;
assign \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.facout_s2  = \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.u2.cout ;
assign \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.fas_s2  = \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.u2.s ;
assign \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.u1.a  = \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.a [1:0];
assign \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.u1.b  = \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.bin_s0 [1:0];
assign \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.u1.cin  = 1'h1;
assign \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.facout_s1  = \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.u1.cout ;
assign \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.fas_s1  = \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.u1.s ;
assign \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.a  = \sub_5s_5s_5_2_1_U14.din0 ;
assign \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.b  = \sub_5s_5s_5_2_1_U14.din1 ;
assign \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.ce  = \sub_5s_5s_5_2_1_U14.ce ;
assign \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.clk  = \sub_5s_5s_5_2_1_U14.clk ;
assign \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.reset  = \sub_5s_5s_5_2_1_U14.reset ;
assign \sub_5s_5s_5_2_1_U14.dout  = \sub_5s_5s_5_2_1_U14.top_sub_5s_5s_5_2_1_Adder_11_U.s ;
assign \sub_5s_5s_5_2_1_U14.ce  = 1'h1;
assign \sub_5s_5s_5_2_1_U14.clk  = ap_clk;
assign \sub_5s_5s_5_2_1_U14.din0  = { ret_V_19_reg_1157[2], ret_V_19_reg_1157[2], ret_V_19_reg_1157 };
assign \sub_5s_5s_5_2_1_U14.din1  = { op_13[3], op_13 };
assign grp_fu_793_p2 = \sub_5s_5s_5_2_1_U14.dout ;
assign \sub_5s_5s_5_2_1_U14.reset  = ap_rst;
assign \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.ain_s0  = \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.a ;
assign \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.bin_s0  = \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.b ;
assign \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.s  = { \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.fas_s2 , \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.sum_s1  };
assign \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.u2.a  = \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.ain_s1 ;
assign \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.u2.b  = \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.bin_s1 ;
assign \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.u2.cin  = \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.carry_s1 ;
assign \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.facout_s2  = \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.u2.cout ;
assign \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.fas_s2  = \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.u2.s ;
assign \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.u1.a  = \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.a [2:0];
assign \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.u1.b  = \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.b [2:0];
assign \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.u1.cin  = 1'h0;
assign \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.facout_s1  = \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.u1.cout ;
assign \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.fas_s1  = \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.u1.s ;
assign \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.a  = \add_6s_6ns_6_2_1_U12.din0 ;
assign \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.b  = \add_6s_6ns_6_2_1_U12.din1 ;
assign \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.ce  = \add_6s_6ns_6_2_1_U12.ce ;
assign \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.clk  = \add_6s_6ns_6_2_1_U12.clk ;
assign \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.reset  = \add_6s_6ns_6_2_1_U12.reset ;
assign \add_6s_6ns_6_2_1_U12.dout  = \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_9_U.s ;
assign \add_6s_6ns_6_2_1_U12.ce  = 1'h1;
assign \add_6s_6ns_6_2_1_U12.clk  = ap_clk;
assign \add_6s_6ns_6_2_1_U12.din0  = { tmp_3_reg_1272[4], tmp_3_reg_1272 };
assign \add_6s_6ns_6_2_1_U12.din1  = 6'h01;
assign grp_fu_721_p2 = \add_6s_6ns_6_2_1_U12.dout ;
assign \add_6s_6ns_6_2_1_U12.reset  = ap_rst;
assign \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.ain_s0  = \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.a ;
assign \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.bin_s0  = \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.b ;
assign \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.s  = { \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.fas_s2 , \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.sum_s1  };
assign \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.u2.a  = \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.ain_s1 ;
assign \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.u2.b  = \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.bin_s1 ;
assign \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.u2.cin  = \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.carry_s1 ;
assign \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.facout_s2  = \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.u2.cout ;
assign \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.fas_s2  = \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.u2.s ;
assign \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.u1.a  = \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.a [2:0];
assign \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.u1.b  = \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.b [2:0];
assign \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.u1.cin  = 1'h0;
assign \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.facout_s1  = \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.u1.cout ;
assign \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.fas_s1  = \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.u1.s ;
assign \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.a  = \add_6ns_6s_6_2_1_U13.din0 ;
assign \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.b  = \add_6ns_6s_6_2_1_U13.din1 ;
assign \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.ce  = \add_6ns_6s_6_2_1_U13.ce ;
assign \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.clk  = \add_6ns_6s_6_2_1_U13.clk ;
assign \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.reset  = \add_6ns_6s_6_2_1_U13.reset ;
assign \add_6ns_6s_6_2_1_U13.dout  = \add_6ns_6s_6_2_1_U13.top_add_6ns_6s_6_2_1_Adder_10_U.s ;
assign \add_6ns_6s_6_2_1_U13.ce  = 1'h1;
assign \add_6ns_6s_6_2_1_U13.clk  = ap_clk;
assign \add_6ns_6s_6_2_1_U13.din0  = ret_V_27_reg_1289;
assign \add_6ns_6s_6_2_1_U13.din1  = { ret_V_21_reg_1052[1], ret_V_21_reg_1052[1], ret_V_21_reg_1052[1], ret_V_21_reg_1052[1], ret_V_21_reg_1052 };
assign grp_fu_749_p2 = \add_6ns_6s_6_2_1_U13.dout ;
assign \add_6ns_6s_6_2_1_U13.reset  = ap_rst;
assign \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.ain_s0  = \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.a ;
assign \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.bin_s0  = \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.b ;
assign \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.s  = { \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.fas_s2 , \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.sum_s1  };
assign \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.u2.a  = \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.ain_s1 ;
assign \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.u2.b  = \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.bin_s1 ;
assign \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.u2.cin  = \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.carry_s1 ;
assign \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.facout_s2  = \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.u2.cout ;
assign \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.fas_s2  = \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.u2.s ;
assign \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.u1.a  = \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.a [2:0];
assign \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.u1.b  = \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.b [2:0];
assign \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.u1.cin  = 1'h0;
assign \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.facout_s1  = \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.u1.cout ;
assign \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.fas_s1  = \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.u1.s ;
assign \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.a  = \add_6ns_6ns_6_2_1_U17.din0 ;
assign \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.b  = \add_6ns_6ns_6_2_1_U17.din1 ;
assign \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.ce  = \add_6ns_6ns_6_2_1_U17.ce ;
assign \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.clk  = \add_6ns_6ns_6_2_1_U17.clk ;
assign \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.reset  = \add_6ns_6ns_6_2_1_U17.reset ;
assign \add_6ns_6ns_6_2_1_U17.dout  = \add_6ns_6ns_6_2_1_U17.top_add_6ns_6ns_6_2_1_Adder_12_U.s ;
assign \add_6ns_6ns_6_2_1_U17.ce  = 1'h1;
assign \add_6ns_6ns_6_2_1_U17.clk  = ap_clk;
assign \add_6ns_6ns_6_2_1_U17.din0  = ret_V_28_reg_1380;
assign \add_6ns_6ns_6_2_1_U17.din1  = select_ln1192_reg_1385;
assign grp_fu_935_p2 = \add_6ns_6ns_6_2_1_U17.dout ;
assign \add_6ns_6ns_6_2_1_U17.reset  = ap_rst;
assign \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.ain_s0  = \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.a ;
assign \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.bin_s0  = \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.b ;
assign \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.s  = { \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.fas_s2 , \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.sum_s1  };
assign \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.u2.a  = \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.ain_s1 ;
assign \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.u2.b  = \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.bin_s1 ;
assign \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.u2.cin  = \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.carry_s1 ;
assign \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.facout_s2  = \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.u2.cout ;
assign \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.fas_s2  = \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.u2.s ;
assign \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.u1.a  = \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.a [2:0];
assign \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.u1.b  = \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.b [2:0];
assign \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.u1.cin  = 1'h0;
assign \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.facout_s1  = \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.u1.cout ;
assign \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.fas_s1  = \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.u1.s ;
assign \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.a  = \add_6ns_6ns_6_2_1_U16.din0 ;
assign \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.b  = \add_6ns_6ns_6_2_1_U16.din1 ;
assign \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.ce  = \add_6ns_6ns_6_2_1_U16.ce ;
assign \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.clk  = \add_6ns_6ns_6_2_1_U16.clk ;
assign \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.reset  = \add_6ns_6ns_6_2_1_U16.reset ;
assign \add_6ns_6ns_6_2_1_U16.dout  = \add_6ns_6ns_6_2_1_U16.top_add_6ns_6ns_6_2_1_Adder_12_U.s ;
assign \add_6ns_6ns_6_2_1_U16.ce  = 1'h1;
assign \add_6ns_6ns_6_2_1_U16.clk  = ap_clk;
assign \add_6ns_6ns_6_2_1_U16.din0  = op_25_V_reg_1350;
assign \add_6ns_6ns_6_2_1_U16.din1  = 6'h01;
assign grp_fu_862_p2 = \add_6ns_6ns_6_2_1_U16.dout ;
assign \add_6ns_6ns_6_2_1_U16.reset  = ap_rst;
assign \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.ain_s0  = \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.a ;
assign \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.bin_s0  = \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.b ;
assign \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.s  = { \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.fas_s2 , \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.sum_s1  };
assign \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.u2.a  = \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.ain_s1 ;
assign \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.u2.b  = \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.bin_s1 ;
assign \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.u2.cin  = \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.carry_s1 ;
assign \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.facout_s2  = \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.u2.cout ;
assign \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.fas_s2  = \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.u2.s ;
assign \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.u1.a  = \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.a [2:0];
assign \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.u1.b  = \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.b [2:0];
assign \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.u1.cin  = 1'h0;
assign \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.facout_s1  = \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.u1.cout ;
assign \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.fas_s1  = \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.u1.s ;
assign \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.a  = \add_6ns_6ns_6_2_1_U15.din0 ;
assign \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.b  = \add_6ns_6ns_6_2_1_U15.din1 ;
assign \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.ce  = \add_6ns_6ns_6_2_1_U15.ce ;
assign \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.clk  = \add_6ns_6ns_6_2_1_U15.clk ;
assign \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.reset  = \add_6ns_6ns_6_2_1_U15.reset ;
assign \add_6ns_6ns_6_2_1_U15.dout  = \add_6ns_6ns_6_2_1_U15.top_add_6ns_6ns_6_2_1_Adder_12_U.s ;
assign \add_6ns_6ns_6_2_1_U15.ce  = 1'h1;
assign \add_6ns_6ns_6_2_1_U15.clk  = ap_clk;
assign \add_6ns_6ns_6_2_1_U15.din0  = add_ln69_2_reg_1314;
assign \add_6ns_6ns_6_2_1_U15.din1  = select_ln69_reg_1309;
assign grp_fu_829_p2 = \add_6ns_6ns_6_2_1_U15.dout ;
assign \add_6ns_6ns_6_2_1_U15.reset  = ap_rst;
assign \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.ain_s0  = \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.a ;
assign \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.bin_s0  = \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.b ;
assign \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.s  = { \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.fas_s2 , \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.sum_s1  };
assign \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.u2.a  = \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.ain_s1 ;
assign \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.u2.b  = \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.bin_s1 ;
assign \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.u2.cin  = \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.carry_s1 ;
assign \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.facout_s2  = \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.u2.cout ;
assign \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.fas_s2  = \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.u2.s ;
assign \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.u1.a  = \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.a [1:0];
assign \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.u1.b  = \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.b [1:0];
assign \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.u1.cin  = 1'h0;
assign \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.facout_s1  = \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.u1.cout ;
assign \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.fas_s1  = \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.u1.s ;
assign \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.a  = \add_5s_5s_5_2_1_U10.din0 ;
assign \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.b  = \add_5s_5s_5_2_1_U10.din1 ;
assign \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.ce  = \add_5s_5s_5_2_1_U10.ce ;
assign \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.clk  = \add_5s_5s_5_2_1_U10.clk ;
assign \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.reset  = \add_5s_5s_5_2_1_U10.reset ;
assign \add_5s_5s_5_2_1_U10.dout  = \add_5s_5s_5_2_1_U10.top_add_5s_5s_5_2_1_Adder_7_U.s ;
assign \add_5s_5s_5_2_1_U10.ce  = 1'h1;
assign \add_5s_5s_5_2_1_U10.clk  = ap_clk;
assign \add_5s_5s_5_2_1_U10.din0  = { add_ln69_reg_1207[3], add_ln69_reg_1207 };
assign \add_5s_5s_5_2_1_U10.din1  = { ret_V_23_reg_1195[2], ret_V_23_reg_1195[2], ret_V_23_reg_1195 };
assign grp_fu_647_p2 = \add_5s_5s_5_2_1_U10.dout ;
assign \add_5s_5s_5_2_1_U10.reset  = ap_rst;
assign \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.ain_s0  = \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.a ;
assign \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.bin_s0  = \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.b ;
assign \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.s  = { \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.fas_s2 , \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.sum_s1  };
assign \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.u2.a  = \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.ain_s1 ;
assign \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.u2.b  = \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.bin_s1 ;
assign \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.u2.cin  = \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.carry_s1 ;
assign \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.facout_s2  = \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.u2.cout ;
assign \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.fas_s2  = \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.u2.s ;
assign \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.u1.a  = \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.a [1:0];
assign \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.u1.b  = \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.b [1:0];
assign \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.u1.cin  = 1'h0;
assign \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.facout_s1  = \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.u1.cout ;
assign \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.fas_s1  = \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.u1.s ;
assign \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.a  = \add_4s_4ns_4_2_1_U7.din0 ;
assign \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.b  = \add_4s_4ns_4_2_1_U7.din1 ;
assign \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.ce  = \add_4s_4ns_4_2_1_U7.ce ;
assign \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.clk  = \add_4s_4ns_4_2_1_U7.clk ;
assign \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.reset  = \add_4s_4ns_4_2_1_U7.reset ;
assign \add_4s_4ns_4_2_1_U7.dout  = \add_4s_4ns_4_2_1_U7.top_add_4s_4ns_4_2_1_Adder_5_U.s ;
assign \add_4s_4ns_4_2_1_U7.ce  = 1'h1;
assign \add_4s_4ns_4_2_1_U7.clk  = ap_clk;
assign \add_4s_4ns_4_2_1_U7.din0  = { ret_V_19_reg_1157[2], ret_V_19_reg_1157 };
assign \add_4s_4ns_4_2_1_U7.din1  = { 2'h0, op_12 };
assign grp_fu_600_p2 = \add_4s_4ns_4_2_1_U7.dout ;
assign \add_4s_4ns_4_2_1_U7.reset  = ap_rst;
assign \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.ain_s0  = \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.a ;
assign \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.bin_s0  = \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.b ;
assign \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.s  = { \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.fas_s2 , \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.sum_s1  };
assign \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.u2.a  = \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.ain_s1 ;
assign \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.u2.b  = \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.bin_s1 ;
assign \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.u2.cin  = \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.carry_s1 ;
assign \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.facout_s2  = \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.u2.cout ;
assign \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.fas_s2  = \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.u2.s ;
assign \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.u1.a  = \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.a [0];
assign \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.u1.b  = \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.b [0];
assign \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.u1.cin  = 1'h0;
assign \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.facout_s1  = \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.u1.cout ;
assign \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.fas_s1  = \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.u1.s ;
assign \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.a  = \add_3s_3s_3_2_1_U5.din0 ;
assign \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.b  = \add_3s_3s_3_2_1_U5.din1 ;
assign \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.ce  = \add_3s_3s_3_2_1_U5.ce ;
assign \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.clk  = \add_3s_3s_3_2_1_U5.clk ;
assign \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.reset  = \add_3s_3s_3_2_1_U5.reset ;
assign \add_3s_3s_3_2_1_U5.dout  = \add_3s_3s_3_2_1_U5.top_add_3s_3s_3_2_1_Adder_3_U.s ;
assign \add_3s_3s_3_2_1_U5.ce  = 1'h1;
assign \add_3s_3s_3_2_1_U5.clk  = ap_clk;
assign \add_3s_3s_3_2_1_U5.din0  = { op_5_V_reg_1152[1], op_5_V_reg_1152 };
assign \add_3s_3s_3_2_1_U5.din1  = { op_0[1], op_0 };
assign grp_fu_578_p2 = \add_3s_3s_3_2_1_U5.dout ;
assign \add_3s_3s_3_2_1_U5.reset  = ap_rst;
assign \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.ain_s0  = \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.a ;
assign \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.bin_s0  = \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.b ;
assign \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.s  = { \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.fas_s2 , \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.sum_s1  };
assign \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.u2.a  = \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.ain_s1 ;
assign \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.u2.b  = \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.bin_s1 ;
assign \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.u2.cin  = \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.carry_s1 ;
assign \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.facout_s2  = \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.u2.cout ;
assign \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.fas_s2  = \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.u2.s ;
assign \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.u1.a  = \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.a [0];
assign \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.u1.b  = \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.b [0];
assign \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.u1.cin  = 1'h0;
assign \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.facout_s1  = \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.u1.cout ;
assign \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.fas_s1  = \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.u1.s ;
assign \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.a  = \add_3ns_3ns_3_2_1_U4.din0 ;
assign \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.b  = \add_3ns_3ns_3_2_1_U4.din1 ;
assign \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.ce  = \add_3ns_3ns_3_2_1_U4.ce ;
assign \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.clk  = \add_3ns_3ns_3_2_1_U4.clk ;
assign \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.reset  = \add_3ns_3ns_3_2_1_U4.reset ;
assign \add_3ns_3ns_3_2_1_U4.dout  = \add_3ns_3ns_3_2_1_U4.top_add_3ns_3ns_3_2_1_Adder_2_U.s ;
assign \add_3ns_3ns_3_2_1_U4.ce  = 1'h1;
assign \add_3ns_3ns_3_2_1_U4.clk  = ap_clk;
assign \add_3ns_3ns_3_2_1_U4.din0  = ret_V_reg_1115;
assign \add_3ns_3ns_3_2_1_U4.din1  = 3'h1;
assign grp_fu_493_p2 = \add_3ns_3ns_3_2_1_U4.dout ;
assign \add_3ns_3ns_3_2_1_U4.reset  = ap_rst;
assign \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.ain_s0  = \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.a ;
assign \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.bin_s0  = \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.b ;
assign \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.s  = { \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.fas_s2 , \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.sum_s1  };
assign \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.a  = \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.ain_s1 ;
assign \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.b  = \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.bin_s1 ;
assign \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.cin  = \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.carry_s1 ;
assign \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.facout_s2  = \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.cout ;
assign \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.fas_s2  = \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.s ;
assign \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.a  = \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.a [0];
assign \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.b  = \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.b [0];
assign \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.cin  = 1'h0;
assign \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.facout_s1  = \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.cout ;
assign \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.fas_s1  = \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.s ;
assign \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.a  = \add_2ns_2ns_2_2_1_U9.din0 ;
assign \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.b  = \add_2ns_2ns_2_2_1_U9.din1 ;
assign \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.ce  = \add_2ns_2ns_2_2_1_U9.ce ;
assign \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.clk  = \add_2ns_2ns_2_2_1_U9.clk ;
assign \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.reset  = \add_2ns_2ns_2_2_1_U9.reset ;
assign \add_2ns_2ns_2_2_1_U9.dout  = \add_2ns_2ns_2_2_1_U9.top_add_2ns_2ns_2_2_1_Adder_1_U.s ;
assign \add_2ns_2ns_2_2_1_U9.ce  = 1'h1;
assign \add_2ns_2ns_2_2_1_U9.clk  = ap_clk;
assign \add_2ns_2ns_2_2_1_U9.din0  = ret_V_21_cast_reg_1200;
assign \add_2ns_2ns_2_2_1_U9.din1  = 2'h1;
assign grp_fu_639_p2 = \add_2ns_2ns_2_2_1_U9.dout ;
assign \add_2ns_2ns_2_2_1_U9.reset  = ap_rst;
assign \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.ain_s0  = \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.a ;
assign \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.bin_s0  = \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.b ;
assign \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.s  = { \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.fas_s2 , \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.sum_s1  };
assign \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.a  = \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.ain_s1 ;
assign \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.b  = \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.bin_s1 ;
assign \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.cin  = \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.carry_s1 ;
assign \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.facout_s2  = \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.cout ;
assign \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.fas_s2  = \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.s ;
assign \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.a  = \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.a [0];
assign \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.b  = \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.b [0];
assign \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.cin  = 1'h0;
assign \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.facout_s1  = \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.cout ;
assign \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.fas_s1  = \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.s ;
assign \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.a  = \add_2ns_2ns_2_2_1_U3.din0 ;
assign \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.b  = \add_2ns_2ns_2_2_1_U3.din1 ;
assign \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.ce  = \add_2ns_2ns_2_2_1_U3.ce ;
assign \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.clk  = \add_2ns_2ns_2_2_1_U3.clk ;
assign \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.reset  = \add_2ns_2ns_2_2_1_U3.reset ;
assign \add_2ns_2ns_2_2_1_U3.dout  = \add_2ns_2ns_2_2_1_U3.top_add_2ns_2ns_2_2_1_Adder_1_U.s ;
assign \add_2ns_2ns_2_2_1_U3.ce  = 1'h1;
assign \add_2ns_2ns_2_2_1_U3.clk  = ap_clk;
assign \add_2ns_2ns_2_2_1_U3.din0  = p_Val2_1_reg_989;
assign \add_2ns_2ns_2_2_1_U3.din1  = { 1'h0, and_ln414_reg_1047 };
assign grp_fu_365_p2 = \add_2ns_2ns_2_2_1_U3.dout ;
assign \add_2ns_2ns_2_2_1_U3.reset  = ap_rst;
assign \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.ain_s0  = \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.a ;
assign \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.bin_s0  = \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.b ;
assign \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.s  = { \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.fas_s2 , \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.sum_s1  };
assign \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.a  = \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.ain_s1 ;
assign \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.b  = \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.bin_s1 ;
assign \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.cin  = \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.carry_s1 ;
assign \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.facout_s2  = \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.cout ;
assign \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.fas_s2  = \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u2.s ;
assign \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.a  = \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.a [0];
assign \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.b  = \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.b [0];
assign \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.cin  = 1'h0;
assign \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.facout_s1  = \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.cout ;
assign \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.fas_s1  = \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.u1.s ;
assign \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.a  = \add_2ns_2ns_2_2_1_U2.din0 ;
assign \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.b  = \add_2ns_2ns_2_2_1_U2.din1 ;
assign \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.ce  = \add_2ns_2ns_2_2_1_U2.ce ;
assign \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.clk  = \add_2ns_2ns_2_2_1_U2.clk ;
assign \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.reset  = \add_2ns_2ns_2_2_1_U2.reset ;
assign \add_2ns_2ns_2_2_1_U2.dout  = \add_2ns_2ns_2_2_1_U2.top_add_2ns_2ns_2_2_1_Adder_1_U.s ;
assign \add_2ns_2ns_2_2_1_U2.ce  = 1'h1;
assign \add_2ns_2ns_2_2_1_U2.clk  = ap_clk;
assign \add_2ns_2ns_2_2_1_U2.din0  = ret_V_4_cast_reg_964;
assign \add_2ns_2ns_2_2_1_U2.din1  = 2'h1;
assign grp_fu_314_p2 = \add_2ns_2ns_2_2_1_U2.dout ;
assign \add_2ns_2ns_2_2_1_U2.reset  = ap_rst;
assign \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.ain_s0  = \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.a ;
assign \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.bin_s0  = \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.b ;
assign \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.s  = { \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.fas_s2 , \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.sum_s1  };
assign \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.u2.a  = \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.ain_s1 ;
assign \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.u2.b  = \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.bin_s1 ;
assign \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.u2.cin  = \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.carry_s1 ;
assign \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.facout_s2  = \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.u2.cout ;
assign \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.fas_s2  = \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.u2.s ;
assign \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.u1.a  = \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.a [7:0];
assign \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.u1.b  = \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.b [7:0];
assign \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.u1.cin  = 1'h0;
assign \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.facout_s1  = \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.u1.cout ;
assign \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.fas_s1  = \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.u1.s ;
assign \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.a  = \add_17s_17s_17_2_1_U8.din0 ;
assign \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.b  = \add_17s_17s_17_2_1_U8.din1 ;
assign \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.ce  = \add_17s_17s_17_2_1_U8.ce ;
assign \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.clk  = \add_17s_17s_17_2_1_U8.clk ;
assign \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.reset  = \add_17s_17s_17_2_1_U8.reset ;
assign \add_17s_17s_17_2_1_U8.dout  = \add_17s_17s_17_2_1_U8.top_add_17s_17s_17_2_1_Adder_6_U.s ;
assign \add_17s_17s_17_2_1_U8.ce  = 1'h1;
assign \add_17s_17s_17_2_1_U8.clk  = ap_clk;
assign \add_17s_17s_17_2_1_U8.din0  = { ret_V_19_reg_1157[2], ret_V_19_reg_1157, 13'h0000 };
assign \add_17s_17s_17_2_1_U8.din1  = { op_3[15], op_3 };
assign grp_fu_633_p2 = \add_17s_17s_17_2_1_U8.dout ;
assign \add_17s_17s_17_2_1_U8.reset  = ap_rst;
assign \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.ain_s0  = \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.a ;
assign \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.bin_s0  = \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.b ;
assign \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.s  = { \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.fas_s2 , \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.sum_s1  };
assign \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.u2.a  = \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.ain_s1 ;
assign \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.u2.b  = \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.bin_s1 ;
assign \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.u2.cin  = \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.carry_s1 ;
assign \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.facout_s2  = \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.u2.cout ;
assign \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.fas_s2  = \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.u2.s ;
assign \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.u1.a  = \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.a [6:0];
assign \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.u1.b  = \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.b [6:0];
assign \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.u1.cin  = 1'h0;
assign \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.facout_s1  = \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.u1.cout ;
assign \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.fas_s1  = \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.u1.s ;
assign \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.a  = \add_15ns_15ns_15_2_1_U6.din0 ;
assign \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.b  = \add_15ns_15ns_15_2_1_U6.din1 ;
assign \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.ce  = \add_15ns_15ns_15_2_1_U6.ce ;
assign \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.clk  = \add_15ns_15ns_15_2_1_U6.clk ;
assign \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.reset  = \add_15ns_15ns_15_2_1_U6.reset ;
assign \add_15ns_15ns_15_2_1_U6.dout  = \add_15ns_15ns_15_2_1_U6.top_add_15ns_15ns_15_2_1_Adder_4_U.s ;
assign \add_15ns_15ns_15_2_1_U6.ce  = 1'h1;
assign \add_15ns_15ns_15_2_1_U6.clk  = ap_clk;
assign \add_15ns_15ns_15_2_1_U6.din0  = { trunc_ln728_reg_1165, 13'h0000 };
assign \add_15ns_15ns_15_2_1_U6.din1  = empty_reg_1093;
assign grp_fu_591_p2 = \add_15ns_15ns_15_2_1_U6.dout ;
assign \add_15ns_15ns_15_2_1_U6.reset  = ap_rst;
assign \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.ain_s0  = \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.a ;
assign \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.bin_s0  = \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.b ;
assign \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.s  = { \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.fas_s2 , \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.sum_s1  };
assign \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.u2.a  = \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.ain_s1 ;
assign \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.u2.b  = \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.bin_s1 ;
assign \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.u2.cin  = \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.carry_s1 ;
assign \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.facout_s2  = \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.u2.cout ;
assign \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.fas_s2  = \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.u2.s ;
assign \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.u1.a  = \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.a [4:0];
assign \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.u1.b  = \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.b [4:0];
assign \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.u1.cin  = 1'h0;
assign \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.facout_s1  = \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.u1.cout ;
assign \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.fas_s1  = \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.u1.s ;
assign \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.a  = \add_10ns_10s_10_2_1_U11.din0 ;
assign \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.b  = \add_10ns_10s_10_2_1_U11.din1 ;
assign \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.ce  = \add_10ns_10s_10_2_1_U11.ce ;
assign \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.clk  = \add_10ns_10s_10_2_1_U11.clk ;
assign \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.reset  = \add_10ns_10s_10_2_1_U11.reset ;
assign \add_10ns_10s_10_2_1_U11.dout  = \add_10ns_10s_10_2_1_U11.top_add_10ns_10s_10_2_1_Adder_8_U.s ;
assign \add_10ns_10s_10_2_1_U11.ce  = 1'h1;
assign \add_10ns_10s_10_2_1_U11.clk  = ap_clk;
assign \add_10ns_10s_10_2_1_U11.din0  = { op_22_V_reg_1242, 5'h00 };
assign \add_10ns_10s_10_2_1_U11.din1  = { op_14[7], op_14[7], op_14 };
assign grp_fu_692_p2 = \add_10ns_10s_10_2_1_U11.dout ;
assign \add_10ns_10s_10_2_1_U11.reset  = ap_rst;
endmodule


// Product machine:
module top_A_times_top_B (ap_start, op_0, op_1, op_10, op_12, op_13, op_14, op_2, op_3, op_7, op_8, ap_clk, unsafe_signal);
input ap_start;
input [1:0] op_0;
input [3:0] op_1;
input [3:0] op_10;
input [1:0] op_12;
input [3:0] op_13;
input [7:0] op_14;
input [7:0] op_2;
input [15:0] op_3;
input [1:0] op_7;
input [1:0] op_8;
input ap_clk;
output unsafe_signal;
reg _setup;
initial _setup = 1'b0;
always @ (posedge ap_clk) _setup <= 1'b1;
reg ap_start_internal;
always @ (posedge ap_clk) if (!_setup) ap_start_internal <= ap_start;
reg [1:0] op_0_internal;
always @ (posedge ap_clk) if (!_setup) op_0_internal <= op_0;
reg [3:0] op_1_internal;
always @ (posedge ap_clk) if (!_setup) op_1_internal <= op_1;
reg [3:0] op_10_internal;
always @ (posedge ap_clk) if (!_setup) op_10_internal <= op_10;
reg [1:0] op_12_internal;
always @ (posedge ap_clk) if (!_setup) op_12_internal <= op_12;
reg [3:0] op_13_internal;
always @ (posedge ap_clk) if (!_setup) op_13_internal <= op_13;
reg [7:0] op_14_internal;
always @ (posedge ap_clk) if (!_setup) op_14_internal <= op_14;
reg [7:0] op_2_internal;
always @ (posedge ap_clk) if (!_setup) op_2_internal <= op_2;
reg [15:0] op_3_internal;
always @ (posedge ap_clk) if (!_setup) op_3_internal <= op_3;
reg [1:0] op_7_internal;
always @ (posedge ap_clk) if (!_setup) op_7_internal <= op_7;
reg [1:0] op_8_internal;
always @ (posedge ap_clk) if (!_setup) op_8_internal <= op_8;
wire ap_done_A;
wire ap_done_B;
wire ap_done_eq;
assign ap_done_eq = ap_done_A == ap_done_B;
wire ap_idle_A;
wire ap_idle_B;
wire ap_idle_eq;
assign ap_idle_eq = ap_idle_A == ap_idle_B;
wire ap_ready_A;
wire ap_ready_B;
wire ap_ready_eq;
assign ap_ready_eq = ap_ready_A == ap_ready_B;
wire [31:0] op_28_A;
wire [31:0] op_28_B;
wire op_28_eq;
assign op_28_eq = op_28_A == op_28_B;
wire op_28_ap_vld_A;
wire op_28_ap_vld_B;
wire clk_enable_A;
wire clk_enable_B;
assign clk_enable_A = _setup & (~op_28_ap_vld_A | op_28_ap_vld_B);
assign clk_enable_B = _setup;
wire divergent;
assign divergent = ~(ap_done_eq & ap_idle_eq & ap_ready_eq & op_28_eq);
assign unsafe_signal = op_28_ap_vld_A & op_28_ap_vld_B & divergent;
top_A instance_A (
    .ap_clk(ap_clk),
    .clk_enable(clk_enable_A),
    .ap_start(ap_start_internal),
    .op_0(op_0_internal),
    .op_1(op_1_internal),
    .op_10(op_10_internal),
    .op_12(op_12_internal),
    .op_13(op_13_internal),
    .op_14(op_14_internal),
    .op_2(op_2_internal),
    .op_3(op_3_internal),
    .op_7(op_7_internal),
    .op_8(op_8_internal),
    .ap_done(ap_done_A),
    .ap_idle(ap_idle_A),
    .ap_ready(ap_ready_A),
    .op_28(op_28_A),
    .op_28_ap_vld(op_28_ap_vld_A)
);
top_B instance_B (
    .ap_clk(ap_clk),
    .clk_enable(clk_enable_B),
    .ap_start(ap_start_internal),
    .op_0(op_0_internal),
    .op_1(op_1_internal),
    .op_10(op_10_internal),
    .op_12(op_12_internal),
    .op_13(op_13_internal),
    .op_14(op_14_internal),
    .op_2(op_2_internal),
    .op_3(op_3_internal),
    .op_7(op_7_internal),
    .op_8(op_8_internal),
    .ap_done(ap_done_B),
    .ap_idle(ap_idle_B),
    .ap_ready(ap_ready_B),
    .op_28(op_28_B),
    .op_28_ap_vld(op_28_ap_vld_B)
);
endmodule
