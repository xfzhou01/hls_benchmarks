// Processed by function `construct_kairos` in `verilog_tricks.py`.
// Machine A:
// Processed by function `add_clk_enable_signal` in `verilog_tricks.py`.
// Processed by function `remove_reset_signal` in `verilog_tricks.py`.
module top_A (
  ap_clk,
  ap_start,
  ap_done,
  ap_idle,
  ap_ready,
  op_0,
  op_1,
  op_2,
  op_5,
  op_7,
  op_12,
  op_13,
  op_15,
  op_16,
  op_18,
  op_19,
  op_30,
  op_30_ap_vld,
clk_enable
);
input clk_enable;


input ap_clk;
wire ap_rst;
assign ap_rst = op_30_ap_vld;
input ap_start;
input [7:0] op_0;
input [31:0] op_1;
input [1:0] op_12;
input [31:0] op_13;
input [31:0] op_15;
input [31:0] op_16;
input [1:0] op_18;
input op_19;
input [15:0] op_2;
input [1:0] op_5;
input [31:0] op_7;
output ap_done;
output ap_idle;
output ap_ready;
output [31:0] op_30;
output op_30_ap_vld;


reg [31:0] add_ln691_1_reg_1274;
reg [8:0] ap_CS_fsm = 9'h001;
reg icmp_ln1499_reg_1248;
reg icmp_ln768_reg_1163;
reg icmp_ln786_reg_1168;
reg icmp_ln851_1_reg_1243;
reg icmp_ln851_2_reg_1207;
reg icmp_ln851_reg_1228;
reg [3:0] op_14_V_reg_1202;
reg [31:0] op_24_V_reg_1258;
reg [31:0] op_28_V_reg_1284;
reg p_Result_14_reg_1151;
reg p_Result_15_reg_1157;
reg p_Result_17_reg_1183;
reg p_Result_18_reg_1189;
reg [7:0] ret_V_15_reg_1212;
reg [32:0] ret_V_16_reg_1217;
reg [17:0] ret_V_18_reg_1253;
reg [31:0] ret_V_22_reg_1279;
reg [31:0] ret_V_23_cast_reg_1268;
reg [33:0] ret_V_23_reg_1294;
reg [31:0] ret_V_27_cast_reg_1299;
reg [15:0] ret_V_3_reg_1222;
reg [15:0] ret_V_4_reg_1233;
reg [4:0] ret_V_5_reg_1238;
reg [32:0] ret_reg_1146;
reg [15:0] tmp_4_reg_1196;
reg [7:0] trunc_ln728_reg_1178;
reg trunc_ln790_reg_1173;
reg [34:0] _114_;
wire [31:0] _000_;
wire [8:0] _001_;
wire _002_;
wire _003_;
wire _004_;
wire _005_;
wire _006_;
wire _007_;
wire [2:0] _008_;
wire [31:0] _009_;
wire [31:0] _010_;
wire _011_;
wire _012_;
wire _013_;
wire _014_;
wire [7:0] _015_;
wire [32:0] _016_;
wire [17:0] _017_;
wire [34:0] _018_;
wire [31:0] _019_;
wire [31:0] _020_;
wire [33:0] _021_;
wire [31:0] _022_;
wire [15:0] _023_;
wire [15:0] _024_;
wire [4:0] _025_;
wire [32:0] _026_;
wire [15:0] _027_;
wire [7:0] _028_;
wire _029_;
wire [1:0] _030_;
wire _031_;
wire _032_;
wire _033_;
wire _034_;
wire _035_;
wire _036_;
wire _037_;
wire _038_;
wire _039_;
wire _040_;
wire _041_;
wire _042_;
wire _043_;
wire _044_;
wire _045_;
wire _046_;
wire _047_;
wire _048_;
wire _049_;
wire _050_;
wire _051_;
wire _052_;
wire _053_;
wire _054_;
wire _055_;
wire [31:0] add_ln691_1_fu_960_p2;
wire [31:0] add_ln691_2_fu_1035_p2;
wire [31:0] add_ln691_3_fu_1112_p2;
wire [17:0] add_ln691_fu_881_p2;
wire [31:0] add_ln69_fu_1060_p2;
wire [2:0] and_ln731_fu_449_p2;
wire ap_CS_fsm_state1;
wire ap_CS_fsm_state2;
wire ap_CS_fsm_state3;
wire ap_CS_fsm_state4;
wire ap_CS_fsm_state5;
wire ap_CS_fsm_state6;
wire ap_CS_fsm_state7;
wire ap_CS_fsm_state8;
wire ap_CS_fsm_state9;
wire [8:0] ap_NS_fsm;
wire ap_clk;
wire ap_done;
wire ap_idle;
wire ap_ready;
wire ap_rst;
wire ap_start;
wire [1:0] icmp_ln1499_fu_805_p1;
wire icmp_ln1499_fu_805_p2;
wire icmp_ln768_1_fu_371_p2;
wire icmp_ln768_2_fu_723_p2;
wire icmp_ln768_fu_307_p2;
wire icmp_ln786_1_fu_749_p2;
wire icmp_ln786_fu_313_p2;
wire icmp_ln790_fu_541_p2;
wire icmp_ln851_1_fu_799_p2;
wire icmp_ln851_2_fu_497_p2;
wire icmp_ln851_3_fu_1029_p2;
wire icmp_ln851_fu_682_p2;
wire [24:0] lhs_V_fu_646_p3;
wire [8:0] lhs_cast_fu_585_p3;
wire [7:0] op_0;
wire [31:0] op_1;
wire [22:0] op_10_V_fu_818_p3;
wire [1:0] op_12;
wire [31:0] op_13;
wire [3:0] op_14_V_fu_485_p3;
wire [31:0] op_15;
wire [31:0] op_16;
wire [1:0] op_18;
wire op_19;
wire [15:0] op_2;
wire [17:0] op_22_V_fu_905_p2;
wire [31:0] op_24_V_fu_924_p2;
wire [31:0] op_28_V_fu_1066_p2;
wire [31:0] op_30;
wire op_30_ap_vld;
wire [3:0] op_3_V_fu_577_p3;
wire [31:0] op_4_V_fu_263_p0;
wire [3:0] op_4_V_fu_263_p1;
wire [1:0] op_5;
wire [31:0] op_7;
wire [3:0] op_8_V_fu_383_p3;
wire [1:0] op_9_V_fu_779_p3;
wire [8:0] or_ln1195_fu_596_p2;
wire or_ln384_1_fu_773_p2;
wire or_ln384_fu_571_p2;
wire or_ln785_2_fu_728_p2;
wire or_ln785_fu_514_p2;
wire or_ln786_fu_754_p2;
wire or_ln788_1_fu_553_p2;
wire or_ln788_fu_547_p2;
wire overflow_1_fu_377_p2;
wire overflow_2_fu_738_p2;
wire overflow_3_fu_479_p2;
wire overflow_fu_523_p2;
wire p_Result_10_fu_873_p3;
wire p_Result_11_fu_966_p3;
wire p_Result_12_fu_1017_p3;
wire p_Result_13_fu_1102_p3;
wire [31:0] p_Result_16_fu_353_p1;
wire p_Result_16_fu_353_p3;
wire p_Result_18_fu_409_p1;
wire p_Result_19_fu_463_p3;
wire [1:0] p_Result_3_fu_612_p1;
wire p_Result_3_fu_612_p3;
wire p_Result_4_fu_811_p3;
wire [19:0] p_Result_9_fu_791_p3;
wire [2:0] p_Result_s_20_fu_534_p3;
wire [30:0] p_Result_s_fu_297_p4;
wire [3:0] p_Val2_1_fu_506_p3;
wire [3:0] p_Val2_3_fu_345_p3;
wire [1:0] p_Val2_6_fu_716_p3;
wire [3:0] p_Val2_8_fu_455_p3;
wire [3:0] r_V_fu_439_p2;
wire [16:0] ret_1_fu_395_p2;
wire [7:0] ret_V_15_fu_638_p3;
wire [32:0] ret_V_16_fu_662_p2;
wire [36:0] ret_V_17_fu_853_p2;
wire [17:0] ret_V_18_fu_894_p3;
wire [17:0] ret_V_19_fu_914_p2;
wire [35:0] ret_V_20_fu_944_p2;
wire [35:0] ret_V_20_reg_1263;
wire [53:0] ret_V_21_fu_1001_p2;
wire [31:0] ret_V_22_fu_1049_p3;
wire [31:0] ret_V_23_cast_fu_950_p4;
wire [33:0] ret_V_23_fu_1086_p2;
wire [31:0] ret_V_24_fu_1124_p3;
wire [31:0] ret_V_25_cast_fu_1007_p4;
wire [15:0] ret_V_3_fu_668_p4;
wire [15:0] ret_V_4_fu_688_p2;
wire [4:0] ret_V_5_fu_710_p2;
wire [7:0] ret_V_cast_fu_602_p4;
wire [7:0] ret_V_fu_624_p2;
wire [32:0] ret_fu_275_p2;
wire [35:0] rhs_2_fu_841_p3;
wire rhs_3_fu_335_p2;
wire [34:0] rhs_5_fu_933_p3;
wire [52:0] rhs_6_fu_989_p3;
wire [32:0] rhs_8_fu_1075_p3;
wire [1:0] rhs_fu_698_p1;
wire [2:0] rhs_fu_698_p3;
wire [2:0] select_ln1118_1_fu_431_p3;
wire [3:0] select_ln1118_fu_423_p3;
wire [31:0] select_ln1192_fu_1131_p3;
wire [31:0] select_ln353_fu_982_p3;
wire [3:0] select_ln384_1_fu_563_p3;
wire [1:0] select_ln384_fu_765_p3;
wire [15:0] select_ln850_1_fu_829_p3;
wire [17:0] select_ln850_2_fu_887_p3;
wire [15:0] select_ln850_3_fu_834_p3;
wire [31:0] select_ln850_4_fu_1041_p3;
wire [31:0] select_ln850_5_fu_1117_p3;
wire [31:0] select_ln850_6_fu_977_p3;
wire [7:0] select_ln850_fu_630_p3;
wire [36:0] sext_ln1192_1_fu_825_p1;
wire [36:0] sext_ln1192_2_fu_849_p1;
wire [17:0] sext_ln1192_3_fu_910_p1;
wire [35:0] sext_ln1192_4_fu_940_p1;
wire [53:0] sext_ln1192_5_fu_997_p1;
wire [33:0] sext_ln1192_6_fu_1082_p1;
wire [31:0] sext_ln1192_8_fu_920_p1;
wire [4:0] sext_ln1192_fu_706_p1;
wire [1:0] sext_ln1195_fu_592_p0;
wire [8:0] sext_ln1195_fu_592_p1;
wire [31:0] sext_ln215_fu_267_p0;
wire [32:0] sext_ln215_fu_267_p1;
wire [17:0] sext_ln69_fu_902_p1;
wire [4:0] sext_ln703_1_fu_694_p1;
wire [35:0] sext_ln703_2_fu_930_p1;
wire [31:0] sext_ln703_3_fu_973_p0;
wire [53:0] sext_ln703_3_fu_973_p1;
wire [1:0] sext_ln703_4_fu_1071_p0;
wire [33:0] sext_ln703_4_fu_1071_p1;
wire [31:0] sext_ln703_fu_658_p0;
wire [32:0] sext_ln703_fu_658_p1;
wire [17:0] sext_ln850_fu_869_p1;
wire [31:0] tmp_3_fu_361_p1;
wire [1:0] tmp_3_fu_361_p4;
wire [16:0] tmp_6_fu_859_p4;
wire tmp_fu_471_p3;
wire [7:0] trunc_ln728_fu_327_p1;
wire [31:0] trunc_ln731_1_fu_341_p0;
wire [1:0] trunc_ln731_1_fu_341_p1;
wire [2:0] trunc_ln731_3_fu_445_p1;
wire [1:0] trunc_ln731_fu_503_p1;
wire trunc_ln790_fu_319_p1;
wire [31:0] trunc_ln851_1_fu_678_p0;
wire [16:0] trunc_ln851_1_fu_678_p1;
wire [1:0] trunc_ln851_2_fu_787_p1;
wire [2:0] trunc_ln851_3_fu_493_p1;
wire [31:0] trunc_ln851_4_fu_1025_p0;
wire [20:0] trunc_ln851_4_fu_1025_p1;
wire [1:0] trunc_ln851_5_fu_1109_p0;
wire trunc_ln851_5_fu_1109_p1;
wire trunc_ln851_fu_620_p1;
wire underflow_1_fu_760_p2;
wire underflow_fu_558_p2;
wire xor_ln785_1_fu_733_p2;
wire xor_ln785_fu_518_p2;
wire xor_ln786_1_fu_744_p2;
wire xor_ln786_fu_529_p2;
wire [32:0] zext_ln1192_fu_654_p1;
wire [16:0] zext_ln1195_fu_323_p1;
wire [16:0] zext_ln1347_fu_391_p1;
wire [32:0] zext_ln215_fu_271_p1;
wire [31:0] zext_ln69_fu_1057_p1;
wire [15:0] zext_ln870_fu_331_p1;


assign add_ln691_1_fu_960_p2 = ret_V_20_fu_944_p2[34:3] + 1'h1;
assign add_ln691_2_fu_1035_p2 = ret_V_21_fu_1001_p2[52:21] + 1'h1;
assign add_ln691_3_fu_1112_p2 = ret_V_27_cast_reg_1299 + 1'h1;
assign add_ln691_fu_881_p2 = $signed(ret_V_17_fu_853_p2[36:20]) + $signed(2'h1);
assign add_ln69_fu_1060_p2 = icmp_ln1499_reg_1248 + op_16;
assign op_22_V_fu_905_p2 = $signed(ret_V_18_reg_1253) + $signed(ret_V_15_reg_1212);
assign op_24_V_fu_924_p2 = $signed(ret_V_19_fu_914_p2) + $signed(op_13);
assign op_28_V_fu_1066_p2 = add_ln69_fu_1060_p2 + ret_V_22_reg_1279;
assign op_30 = ret_V_24_fu_1124_p3 + select_ln1192_fu_1131_p3;
assign ret_V_16_fu_662_p2 = $signed({ 1'h0, op_0, 17'h00000 }) + $signed(op_7);
assign ret_V_17_fu_853_p2 = $signed({ select_ln850_3_fu_834_p3, 20'h00000 }) + $signed({ ret_V_5_reg_1238, 18'h00000 });
assign ret_V_19_fu_914_p2 = $signed(op_22_V_fu_905_p2) + $signed(op_12);
assign ret_V_20_fu_944_p2 = $signed({ op_24_V_reg_1258, 3'h0 }) + $signed(op_14_V_reg_1202);
assign ret_V_21_fu_1001_p2 = $signed({ select_ln353_fu_982_p3, 21'h000000 }) + $signed(op_15);
assign ret_V_23_fu_1086_p2 = $signed({ op_28_V_reg_1284, 1'h0 }) + $signed(op_18);
assign ret_V_4_fu_688_p2 = ret_V_16_fu_662_p2[32:17] + 1'h1;
assign ret_V_5_fu_710_p2 = $signed({ op_5, 1'h0 }) + $signed(op_3_V_fu_577_p3);
assign ret_V_fu_624_p2 = or_ln1195_fu_596_p2[8:1] + 1'h1;
assign _031_ = icmp_ln851_2_reg_1207 & ap_CS_fsm[4];
assign _032_ = ap_CS_fsm[0] & _034_;
assign _033_ = ap_CS_fsm[0] & ap_start;
assign and_ln731_fu_449_p2 = op_8_V_fu_383_p3[2:0] & select_ln1118_1_fu_431_p3;
assign overflow_2_fu_738_p2 = xor_ln785_1_fu_733_p2 & or_ln785_2_fu_728_p2;
assign overflow_fu_523_p2 = xor_ln785_fu_518_p2 & or_ln785_fu_514_p2;
assign r_V_fu_439_p2 = select_ln1118_fu_423_p3 & op_8_V_fu_383_p3;
assign underflow_1_fu_760_p2 = p_Result_17_reg_1183 & or_ln786_fu_754_p2;
assign underflow_fu_558_p2 = p_Result_14_reg_1151 & or_ln788_1_fu_553_p2;
assign xor_ln785_1_fu_733_p2 = ~ p_Result_17_reg_1183;
assign xor_ln786_1_fu_744_p2 = ~ p_Result_18_reg_1189;
assign xor_ln785_fu_518_p2 = ~ p_Result_14_reg_1151;
assign xor_ln786_fu_529_p2 = ~ p_Result_15_reg_1157;
assign _034_ = ~ ap_start;
assign _035_ = ! { trunc_ln790_reg_1173, 2'h0 };
assign _036_ = ! op_7[16:0];
assign _037_ = op_1[3:0] == op_2;
assign _038_ = op_9_V_fu_779_p3 != op_5;
assign _039_ = | op_1[3:2];
assign _040_ = | tmp_4_reg_1196;
assign _041_ = | ret_fu_275_p2[32:2];
assign _042_ = tmp_4_reg_1196 != 16'hffff;
assign _043_ = ret_fu_275_p2[32:2] != 31'h7fffffff;
assign _044_ = | { ret_V_5_fu_710_p2[1:0], 18'h00000 };
assign _045_ = | op_14_V_fu_485_p3[2:0];
assign _046_ = | op_15[20:0];
assign or_ln1195_fu_596_p2 = { op_5[1], op_5[1], op_5[1], op_5[1], op_5[1], op_5[1], op_5[1], op_5 } | { trunc_ln728_reg_1178, 1'h0 };
assign or_ln384_1_fu_773_p2 = underflow_1_fu_760_p2 | overflow_2_fu_738_p2;
assign or_ln384_fu_571_p2 = underflow_fu_558_p2 | overflow_fu_523_p2;
assign or_ln785_2_fu_728_p2 = p_Result_18_reg_1189 | icmp_ln768_2_fu_723_p2;
assign or_ln785_fu_514_p2 = p_Result_15_reg_1157 | icmp_ln768_reg_1163;
assign or_ln786_fu_754_p2 = xor_ln786_1_fu_744_p2 | icmp_ln786_1_fu_749_p2;
assign or_ln788_1_fu_553_p2 = or_ln788_fu_547_p2 | icmp_ln786_reg_1168;
assign or_ln788_fu_547_p2 = xor_ln786_fu_529_p2 | icmp_ln790_fu_541_p2;
assign overflow_1_fu_377_p2 = op_1[1] | icmp_ln768_1_fu_371_p2;
assign overflow_3_fu_479_p2 = r_V_fu_439_p2[3] | and_ln731_fu_449_p2[2];
always @(posedge ap_clk)
op_14_V_reg_1202[0] <= 1'h0;
always @(posedge ap_clk)
ret_V_23_reg_1294 <= _021_;
always @(posedge ap_clk)
ret_V_27_cast_reg_1299 <= _022_;
always @(posedge ap_clk)
ret_V_22_reg_1279 <= _019_;
always @(posedge ap_clk)
_114_ <= _018_;
assign ret_V_20_reg_1263[35:1] = _114_;
always @(posedge ap_clk)
ret_V_23_cast_reg_1268 <= _020_;
always @(posedge ap_clk)
ret_V_18_reg_1253 <= _017_;
always @(posedge ap_clk)
op_28_V_reg_1284 <= _010_;
always @(posedge ap_clk)
op_24_V_reg_1258 <= _009_;
always @(posedge ap_clk)
ret_reg_1146 <= _026_;
always @(posedge ap_clk)
p_Result_14_reg_1151 <= _011_;
always @(posedge ap_clk)
p_Result_15_reg_1157 <= _012_;
always @(posedge ap_clk)
icmp_ln768_reg_1163 <= _003_;
always @(posedge ap_clk)
icmp_ln786_reg_1168 <= _004_;
always @(posedge ap_clk)
trunc_ln790_reg_1173 <= _029_;
always @(posedge ap_clk)
trunc_ln728_reg_1178 <= _028_;
always @(posedge ap_clk)
p_Result_17_reg_1183 <= _013_;
always @(posedge ap_clk)
p_Result_18_reg_1189 <= _014_;
always @(posedge ap_clk)
tmp_4_reg_1196 <= _027_;
always @(posedge ap_clk)
op_14_V_reg_1202[3:1] <= _008_;
always @(posedge ap_clk)
icmp_ln851_2_reg_1207 <= _006_;
always @(posedge ap_clk)
ret_V_15_reg_1212 <= _015_;
always @(posedge ap_clk)
ret_V_16_reg_1217 <= _016_;
always @(posedge ap_clk)
ret_V_3_reg_1222 <= _023_;
always @(posedge ap_clk)
icmp_ln851_reg_1228 <= _007_;
always @(posedge ap_clk)
ret_V_4_reg_1233 <= _024_;
always @(posedge ap_clk)
ret_V_5_reg_1238 <= _025_;
always @(posedge ap_clk)
icmp_ln851_1_reg_1243 <= _005_;
always @(posedge ap_clk)
icmp_ln1499_reg_1248 <= _002_;
always @(posedge ap_clk)
add_ln691_1_reg_1274 <= _000_;
always @(posedge ap_clk)
ap_CS_fsm <= _001_;
assign _030_ = _033_ ? 2'h2 : 2'h1;
assign _047_ = ap_CS_fsm == 1'h1;
function [8:0] _143_;
input [8:0] a;
input [80:0] b;
input [8:0] s;
case (s)
9'b000000001:
_143_ = b[8:0];
9'b000000010:
_143_ = b[17:9];
9'b000000100:
_143_ = b[26:18];
9'b000001000:
_143_ = b[35:27];
9'b000010000:
_143_ = b[44:36];
9'b000100000:
_143_ = b[53:45];
9'b001000000:
_143_ = b[62:54];
9'b010000000:
_143_ = b[71:63];
9'b100000000:
_143_ = b[80:72];
9'b000000000:
_143_ = a;
default:
_143_ = 9'bx;
endcase
endfunction
assign ap_NS_fsm = _143_(9'hxxx, { 7'h00, _030_, 72'h020202020202020001 }, { _047_, _055_, _054_, _053_, _052_, _051_, _050_, _049_, _048_ });
assign _048_ = ap_CS_fsm == 9'h100;
assign _049_ = ap_CS_fsm == 8'h80;
assign _050_ = ap_CS_fsm == 7'h40;
assign _051_ = ap_CS_fsm == 6'h20;
assign _052_ = ap_CS_fsm == 5'h10;
assign _053_ = ap_CS_fsm == 4'h8;
assign _054_ = ap_CS_fsm == 3'h4;
assign _055_ = ap_CS_fsm == 2'h2;
assign op_30_ap_vld = ap_CS_fsm[8] ? 1'h1 : 1'h0;
assign ap_idle = _032_ ? 1'h1 : 1'h0;
assign _022_ = ap_CS_fsm[7] ? ret_V_23_fu_1086_p2[32:1] : ret_V_27_cast_reg_1299;
assign _021_ = ap_CS_fsm[7] ? ret_V_23_fu_1086_p2 : ret_V_23_reg_1294;
assign _019_ = ap_CS_fsm[5] ? ret_V_22_fu_1049_p3 : ret_V_22_reg_1279;
assign _020_ = ap_CS_fsm[4] ? ret_V_20_fu_944_p2[34:3] : ret_V_23_cast_reg_1268;
assign _018_ = ap_CS_fsm[4] ? ret_V_20_fu_944_p2[35:1] : ret_V_20_reg_1263[35:1];
assign _017_ = ap_CS_fsm[2] ? ret_V_18_fu_894_p3 : ret_V_18_reg_1253;
assign _010_ = ap_CS_fsm[6] ? op_28_V_fu_1066_p2 : op_28_V_reg_1284;
assign _009_ = ap_CS_fsm[3] ? op_24_V_fu_924_p2 : op_24_V_reg_1258;
assign _006_ = ap_CS_fsm[0] ? icmp_ln851_2_fu_497_p2 : icmp_ln851_2_reg_1207;
assign _008_ = ap_CS_fsm[0] ? op_14_V_fu_485_p3[3:1] : op_14_V_reg_1202[3:1];
assign _027_ = ap_CS_fsm[0] ? ret_1_fu_395_p2[16:1] : tmp_4_reg_1196;
assign _014_ = ap_CS_fsm[0] ? ret_1_fu_395_p2[0] : p_Result_18_reg_1189;
assign _013_ = ap_CS_fsm[0] ? ret_1_fu_395_p2[16] : p_Result_17_reg_1183;
assign _028_ = ap_CS_fsm[0] ? op_2[7:0] : trunc_ln728_reg_1178;
assign _029_ = ap_CS_fsm[0] ? ret_fu_275_p2[0] : trunc_ln790_reg_1173;
assign _004_ = ap_CS_fsm[0] ? icmp_ln786_fu_313_p2 : icmp_ln786_reg_1168;
assign _003_ = ap_CS_fsm[0] ? icmp_ln768_fu_307_p2 : icmp_ln768_reg_1163;
assign _012_ = ap_CS_fsm[0] ? ret_fu_275_p2[1] : p_Result_15_reg_1157;
assign _011_ = ap_CS_fsm[0] ? ret_fu_275_p2[32] : p_Result_14_reg_1151;
assign _026_ = ap_CS_fsm[0] ? ret_fu_275_p2 : ret_reg_1146;
assign _002_ = ap_CS_fsm[1] ? icmp_ln1499_fu_805_p2 : icmp_ln1499_reg_1248;
assign _005_ = ap_CS_fsm[1] ? icmp_ln851_1_fu_799_p2 : icmp_ln851_1_reg_1243;
assign _025_ = ap_CS_fsm[1] ? ret_V_5_fu_710_p2 : ret_V_5_reg_1238;
assign _024_ = ap_CS_fsm[1] ? ret_V_4_fu_688_p2 : ret_V_4_reg_1233;
assign _007_ = ap_CS_fsm[1] ? icmp_ln851_fu_682_p2 : icmp_ln851_reg_1228;
assign _023_ = ap_CS_fsm[1] ? ret_V_16_fu_662_p2[32:17] : ret_V_3_reg_1222;
assign _016_ = ap_CS_fsm[1] ? ret_V_16_fu_662_p2 : ret_V_16_reg_1217;
assign _015_ = ap_CS_fsm[1] ? ret_V_15_fu_638_p3 : ret_V_15_reg_1212;
assign _000_ = _031_ ? add_ln691_1_fu_960_p2 : add_ln691_1_reg_1274;
assign _001_ = ap_rst ? 9'h001 : ap_NS_fsm;
assign ret_1_fu_395_p2 = op_2 - rhs_3_fu_335_p2;
assign ret_fu_275_p2 = $signed(op_1) - $signed({ 1'h0, op_2 });
assign icmp_ln1499_fu_805_p2 = _038_ ? 1'h1 : 1'h0;
assign icmp_ln768_1_fu_371_p2 = _039_ ? 1'h1 : 1'h0;
assign icmp_ln768_2_fu_723_p2 = _040_ ? 1'h1 : 1'h0;
assign icmp_ln768_fu_307_p2 = _041_ ? 1'h1 : 1'h0;
assign icmp_ln786_1_fu_749_p2 = _042_ ? 1'h1 : 1'h0;
assign icmp_ln786_fu_313_p2 = _043_ ? 1'h1 : 1'h0;
assign icmp_ln790_fu_541_p2 = _035_ ? 1'h1 : 1'h0;
assign icmp_ln851_1_fu_799_p2 = _044_ ? 1'h1 : 1'h0;
assign icmp_ln851_2_fu_497_p2 = _045_ ? 1'h1 : 1'h0;
assign icmp_ln851_3_fu_1029_p2 = _046_ ? 1'h1 : 1'h0;
assign icmp_ln851_fu_682_p2 = _036_ ? 1'h1 : 1'h0;
assign op_14_V_fu_485_p3 = overflow_3_fu_479_p2 ? 4'h0 : { and_ln731_fu_449_p2, 1'h0 };
assign op_3_V_fu_577_p3 = or_ln384_fu_571_p2 ? select_ln384_1_fu_563_p3 : { ret_reg_1146[1:0], 2'h0 };
assign op_8_V_fu_383_p3 = overflow_1_fu_377_p2 ? 4'h7 : { op_1[1:0], 2'h0 };
assign op_9_V_fu_779_p3 = or_ln384_1_fu_773_p2 ? select_ln384_fu_765_p3 : { p_Result_18_reg_1189, 1'h0 };
assign ret_V_15_fu_638_p3 = op_5[1] ? select_ln850_fu_630_p3 : or_ln1195_fu_596_p2[8:1];
assign ret_V_18_fu_894_p3 = ret_V_17_fu_853_p2[36] ? select_ln850_2_fu_887_p3 : { 2'h0, ret_V_17_fu_853_p2[35:20] };
assign ret_V_22_fu_1049_p3 = ret_V_21_fu_1001_p2[53] ? select_ln850_4_fu_1041_p3 : ret_V_21_fu_1001_p2[52:21];
assign ret_V_24_fu_1124_p3 = ret_V_23_reg_1294[33] ? select_ln850_5_fu_1117_p3 : ret_V_27_cast_reg_1299;
assign rhs_3_fu_335_p2 = _037_ ? 1'h1 : 1'h0;
assign select_ln1118_1_fu_431_p3 = rhs_3_fu_335_p2 ? 3'h7 : 3'h0;
assign select_ln1118_fu_423_p3 = rhs_3_fu_335_p2 ? 4'hf : 4'h0;
assign select_ln1192_fu_1131_p3 = op_19 ? 32'd4294967295 : 32'd0;
assign select_ln353_fu_982_p3 = ret_V_20_reg_1263[35] ? select_ln850_6_fu_977_p3 : ret_V_23_cast_reg_1268;
assign select_ln384_1_fu_563_p3 = overflow_fu_523_p2 ? 4'h7 : 4'h9;
assign select_ln384_fu_765_p3 = overflow_2_fu_738_p2 ? 2'h1 : 2'h2;
assign select_ln850_1_fu_829_p3 = icmp_ln851_reg_1228 ? ret_V_3_reg_1222 : ret_V_4_reg_1233;
assign select_ln850_2_fu_887_p3 = icmp_ln851_1_reg_1243 ? add_ln691_fu_881_p2 : { 2'h3, ret_V_17_fu_853_p2[35:20] };
assign select_ln850_3_fu_834_p3 = ret_V_16_reg_1217[32] ? select_ln850_1_fu_829_p3 : ret_V_3_reg_1222;
assign select_ln850_4_fu_1041_p3 = icmp_ln851_3_fu_1029_p2 ? add_ln691_2_fu_1035_p2 : ret_V_21_fu_1001_p2[52:21];
assign select_ln850_5_fu_1117_p3 = op_18[0] ? add_ln691_3_fu_1112_p2 : ret_V_27_cast_reg_1299;
assign select_ln850_6_fu_977_p3 = icmp_ln851_2_reg_1207 ? add_ln691_1_reg_1274 : ret_V_23_cast_reg_1268;
assign select_ln850_fu_630_p3 = or_ln1195_fu_596_p2[0] ? ret_V_fu_624_p2 : or_ln1195_fu_596_p2[8:1];
assign ap_CS_fsm_state1 = ap_CS_fsm[0];
assign ap_CS_fsm_state2 = ap_CS_fsm[1];
assign ap_CS_fsm_state3 = ap_CS_fsm[2];
assign ap_CS_fsm_state4 = ap_CS_fsm[3];
assign ap_CS_fsm_state5 = ap_CS_fsm[4];
assign ap_CS_fsm_state6 = ap_CS_fsm[5];
assign ap_CS_fsm_state7 = ap_CS_fsm[6];
assign ap_CS_fsm_state8 = ap_CS_fsm[7];
assign ap_CS_fsm_state9 = ap_CS_fsm[8];
assign ap_done = op_30_ap_vld;
assign ap_ready = op_30_ap_vld;
assign icmp_ln1499_fu_805_p1 = op_5;
assign lhs_V_fu_646_p3 = { op_0, 17'h00000 };
assign lhs_cast_fu_585_p3 = { trunc_ln728_reg_1178, 1'h0 };
assign op_10_V_fu_818_p3 = { ret_V_5_reg_1238, 18'h00000 };
assign op_4_V_fu_263_p0 = op_1;
assign op_4_V_fu_263_p1 = op_1[3:0];
assign p_Result_10_fu_873_p3 = ret_V_17_fu_853_p2[36];
assign p_Result_11_fu_966_p3 = ret_V_20_reg_1263[35];
assign p_Result_12_fu_1017_p3 = ret_V_21_fu_1001_p2[53];
assign p_Result_13_fu_1102_p3 = ret_V_23_reg_1294[33];
assign p_Result_16_fu_353_p1 = op_1;
assign p_Result_16_fu_353_p3 = op_1[1];
assign p_Result_18_fu_409_p1 = ret_1_fu_395_p2[0];
assign p_Result_19_fu_463_p3 = and_ln731_fu_449_p2[2];
assign p_Result_3_fu_612_p1 = op_5;
assign p_Result_3_fu_612_p3 = op_5[1];
assign p_Result_4_fu_811_p3 = ret_V_16_reg_1217[32];
assign p_Result_9_fu_791_p3 = { ret_V_5_fu_710_p2[1:0], 18'h00000 };
assign p_Result_s_20_fu_534_p3 = { trunc_ln790_reg_1173, 2'h0 };
assign p_Result_s_fu_297_p4 = ret_fu_275_p2[32:2];
assign p_Val2_1_fu_506_p3 = { ret_reg_1146[1:0], 2'h0 };
assign p_Val2_3_fu_345_p3 = { op_1[1:0], 2'h0 };
assign p_Val2_6_fu_716_p3 = { p_Result_18_reg_1189, 1'h0 };
assign p_Val2_8_fu_455_p3 = { and_ln731_fu_449_p2, 1'h0 };
assign ret_V_23_cast_fu_950_p4 = ret_V_20_fu_944_p2[34:3];
assign ret_V_25_cast_fu_1007_p4 = ret_V_21_fu_1001_p2[52:21];
assign ret_V_3_fu_668_p4 = ret_V_16_fu_662_p2[32:17];
assign ret_V_cast_fu_602_p4 = or_ln1195_fu_596_p2[8:1];
assign rhs_2_fu_841_p3 = { select_ln850_3_fu_834_p3, 20'h00000 };
assign rhs_5_fu_933_p3 = { op_24_V_reg_1258, 3'h0 };
assign rhs_6_fu_989_p3 = { select_ln353_fu_982_p3, 21'h000000 };
assign rhs_8_fu_1075_p3 = { op_28_V_reg_1284, 1'h0 };
assign rhs_fu_698_p1 = op_5;
assign rhs_fu_698_p3 = { op_5, 1'h0 };
assign sext_ln1192_1_fu_825_p1 = { ret_V_5_reg_1238[4], ret_V_5_reg_1238[4], ret_V_5_reg_1238[4], ret_V_5_reg_1238[4], ret_V_5_reg_1238[4], ret_V_5_reg_1238[4], ret_V_5_reg_1238[4], ret_V_5_reg_1238[4], ret_V_5_reg_1238[4], ret_V_5_reg_1238[4], ret_V_5_reg_1238[4], ret_V_5_reg_1238[4], ret_V_5_reg_1238[4], ret_V_5_reg_1238[4], ret_V_5_reg_1238, 18'h00000 };
assign sext_ln1192_2_fu_849_p1 = { select_ln850_3_fu_834_p3[15], select_ln850_3_fu_834_p3, 20'h00000 };
assign sext_ln1192_3_fu_910_p1 = { op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12 };
assign sext_ln1192_4_fu_940_p1 = { op_24_V_reg_1258[31], op_24_V_reg_1258, 3'h0 };
assign sext_ln1192_5_fu_997_p1 = { select_ln353_fu_982_p3[31], select_ln353_fu_982_p3, 21'h000000 };
assign sext_ln1192_6_fu_1082_p1 = { op_28_V_reg_1284[31], op_28_V_reg_1284, 1'h0 };
assign sext_ln1192_8_fu_920_p1 = { ret_V_19_fu_914_p2[17], ret_V_19_fu_914_p2[17], ret_V_19_fu_914_p2[17], ret_V_19_fu_914_p2[17], ret_V_19_fu_914_p2[17], ret_V_19_fu_914_p2[17], ret_V_19_fu_914_p2[17], ret_V_19_fu_914_p2[17], ret_V_19_fu_914_p2[17], ret_V_19_fu_914_p2[17], ret_V_19_fu_914_p2[17], ret_V_19_fu_914_p2[17], ret_V_19_fu_914_p2[17], ret_V_19_fu_914_p2[17], ret_V_19_fu_914_p2 };
assign sext_ln1192_fu_706_p1 = { op_5[1], op_5[1], op_5, 1'h0 };
assign sext_ln1195_fu_592_p0 = op_5;
assign sext_ln1195_fu_592_p1 = { op_5[1], op_5[1], op_5[1], op_5[1], op_5[1], op_5[1], op_5[1], op_5 };
assign sext_ln215_fu_267_p0 = op_1;
assign sext_ln215_fu_267_p1 = { op_1[31], op_1 };
assign sext_ln69_fu_902_p1 = { ret_V_15_reg_1212[7], ret_V_15_reg_1212[7], ret_V_15_reg_1212[7], ret_V_15_reg_1212[7], ret_V_15_reg_1212[7], ret_V_15_reg_1212[7], ret_V_15_reg_1212[7], ret_V_15_reg_1212[7], ret_V_15_reg_1212[7], ret_V_15_reg_1212[7], ret_V_15_reg_1212 };
assign sext_ln703_1_fu_694_p1 = { op_3_V_fu_577_p3[3], op_3_V_fu_577_p3 };
assign sext_ln703_2_fu_930_p1 = { op_14_V_reg_1202[3], op_14_V_reg_1202[3], op_14_V_reg_1202[3], op_14_V_reg_1202[3], op_14_V_reg_1202[3], op_14_V_reg_1202[3], op_14_V_reg_1202[3], op_14_V_reg_1202[3], op_14_V_reg_1202[3], op_14_V_reg_1202[3], op_14_V_reg_1202[3], op_14_V_reg_1202[3], op_14_V_reg_1202[3], op_14_V_reg_1202[3], op_14_V_reg_1202[3], op_14_V_reg_1202[3], op_14_V_reg_1202[3], op_14_V_reg_1202[3], op_14_V_reg_1202[3], op_14_V_reg_1202[3], op_14_V_reg_1202[3], op_14_V_reg_1202[3], op_14_V_reg_1202[3], op_14_V_reg_1202[3], op_14_V_reg_1202[3], op_14_V_reg_1202[3], op_14_V_reg_1202[3], op_14_V_reg_1202[3], op_14_V_reg_1202[3], op_14_V_reg_1202[3], op_14_V_reg_1202[3], op_14_V_reg_1202[3], op_14_V_reg_1202 };
assign sext_ln703_3_fu_973_p0 = op_15;
assign sext_ln703_3_fu_973_p1 = { op_15[31], op_15[31], op_15[31], op_15[31], op_15[31], op_15[31], op_15[31], op_15[31], op_15[31], op_15[31], op_15[31], op_15[31], op_15[31], op_15[31], op_15[31], op_15[31], op_15[31], op_15[31], op_15[31], op_15[31], op_15[31], op_15[31], op_15 };
assign sext_ln703_4_fu_1071_p0 = op_18;
assign sext_ln703_4_fu_1071_p1 = { op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18 };
assign sext_ln703_fu_658_p0 = op_7;
assign sext_ln703_fu_658_p1 = { op_7[31], op_7 };
assign sext_ln850_fu_869_p1 = { ret_V_17_fu_853_p2[36], ret_V_17_fu_853_p2[36:20] };
assign tmp_3_fu_361_p1 = op_1;
assign tmp_3_fu_361_p4 = op_1[3:2];
assign tmp_6_fu_859_p4 = ret_V_17_fu_853_p2[36:20];
assign tmp_fu_471_p3 = r_V_fu_439_p2[3];
assign trunc_ln728_fu_327_p1 = op_2[7:0];
assign trunc_ln731_1_fu_341_p0 = op_1;
assign trunc_ln731_1_fu_341_p1 = op_1[1:0];
assign trunc_ln731_3_fu_445_p1 = op_8_V_fu_383_p3[2:0];
assign trunc_ln731_fu_503_p1 = ret_reg_1146[1:0];
assign trunc_ln790_fu_319_p1 = ret_fu_275_p2[0];
assign trunc_ln851_1_fu_678_p0 = op_7;
assign trunc_ln851_1_fu_678_p1 = op_7[16:0];
assign trunc_ln851_2_fu_787_p1 = ret_V_5_fu_710_p2[1:0];
assign trunc_ln851_3_fu_493_p1 = op_14_V_fu_485_p3[2:0];
assign trunc_ln851_4_fu_1025_p0 = op_15;
assign trunc_ln851_4_fu_1025_p1 = op_15[20:0];
assign trunc_ln851_5_fu_1109_p0 = op_18;
assign trunc_ln851_5_fu_1109_p1 = op_18[0];
assign trunc_ln851_fu_620_p1 = or_ln1195_fu_596_p2[0];
assign zext_ln1192_fu_654_p1 = { 8'h00, op_0, 17'h00000 };
assign zext_ln1195_fu_323_p1 = { 1'h0, op_2 };
assign zext_ln1347_fu_391_p1 = { 16'h0000, rhs_3_fu_335_p2 };
assign zext_ln215_fu_271_p1 = { 17'h00000, op_2 };
assign zext_ln69_fu_1057_p1 = { 31'h00000000, icmp_ln1499_reg_1248 };
assign zext_ln870_fu_331_p1 = { 12'h000, op_1[3:0] };
endmodule


// Machine B:
// Processed by function `add_clk_enable_signal` in `verilog_tricks.py`.
// Processed by function `remove_reset_signal` in `verilog_tricks.py`.
module top_B (
  ap_clk,
  ap_start,
  ap_done,
  ap_idle,
  ap_ready,
  op_0,
  op_1,
  op_2,
  op_5,
  op_7,
  op_12,
  op_13,
  op_15,
  op_16,
  op_18,
  op_19,
  op_30,
  op_30_ap_vld,
clk_enable
);
input clk_enable;


input ap_clk;
wire ap_rst;
assign ap_rst = op_30_ap_vld;
input ap_start;
input [7:0] op_0;
input [31:0] op_1;
input [1:0] op_12;
input [31:0] op_13;
input [31:0] op_15;
input [31:0] op_16;
input [1:0] op_18;
input op_19;
input [15:0] op_2;
input [1:0] op_5;
input [31:0] op_7;
output ap_done;
output ap_idle;
output ap_ready;
output [31:0] op_30;
output op_30_ap_vld;


reg [7:0] \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_3_U.ain_s1 ;
reg [7:0] \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_3_U.bin_s1 ;
reg \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_3_U.carry_s1 ;
reg [7:0] \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_3_U.sum_s1 ;
reg [8:0] \add_18ns_18s_18_2_1_U10.top_add_18ns_18s_18_2_1_Adder_8_U.ain_s1 ;
reg [8:0] \add_18ns_18s_18_2_1_U10.top_add_18ns_18s_18_2_1_Adder_8_U.bin_s1 ;
reg \add_18ns_18s_18_2_1_U10.top_add_18ns_18s_18_2_1_Adder_8_U.carry_s1 ;
reg [8:0] \add_18ns_18s_18_2_1_U10.top_add_18ns_18s_18_2_1_Adder_8_U.sum_s1 ;
reg [8:0] \add_18ns_18s_18_2_1_U9.top_add_18ns_18s_18_2_1_Adder_8_U.ain_s1 ;
reg [8:0] \add_18ns_18s_18_2_1_U9.top_add_18ns_18s_18_2_1_Adder_8_U.bin_s1 ;
reg \add_18ns_18s_18_2_1_U9.top_add_18ns_18s_18_2_1_Adder_8_U.carry_s1 ;
reg [8:0] \add_18ns_18s_18_2_1_U9.top_add_18ns_18s_18_2_1_Adder_8_U.sum_s1 ;
reg [8:0] \add_18s_18ns_18_2_1_U8.top_add_18s_18ns_18_2_1_Adder_7_U.ain_s1 ;
reg [8:0] \add_18s_18ns_18_2_1_U8.top_add_18s_18ns_18_2_1_Adder_7_U.bin_s1 ;
reg \add_18s_18ns_18_2_1_U8.top_add_18s_18ns_18_2_1_Adder_7_U.carry_s1 ;
reg [8:0] \add_18s_18ns_18_2_1_U8.top_add_18s_18ns_18_2_1_Adder_7_U.sum_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_11_U.ain_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_11_U.bin_s1 ;
reg \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_11_U.carry_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_11_U.sum_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.ain_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.bin_s1 ;
reg \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.carry_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.sum_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.ain_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.bin_s1 ;
reg \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.carry_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.sum_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.ain_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.bin_s1 ;
reg \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.carry_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.sum_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.ain_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.bin_s1 ;
reg \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.carry_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.sum_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.ain_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.bin_s1 ;
reg \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.carry_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.sum_s1 ;
reg [15:0] \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_9_U.ain_s1 ;
reg [15:0] \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_9_U.bin_s1 ;
reg \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_9_U.carry_s1 ;
reg [15:0] \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_9_U.sum_s1 ;
reg [16:0] \add_33ns_33s_33_2_1_U3.top_add_33ns_33s_33_2_1_Adder_2_U.ain_s1 ;
reg [16:0] \add_33ns_33s_33_2_1_U3.top_add_33ns_33s_33_2_1_Adder_2_U.bin_s1 ;
reg \add_33ns_33s_33_2_1_U3.top_add_33ns_33s_33_2_1_Adder_2_U.carry_s1 ;
reg [15:0] \add_33ns_33s_33_2_1_U3.top_add_33ns_33s_33_2_1_Adder_2_U.sum_s1 ;
reg [16:0] \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_13_U.ain_s1 ;
reg [16:0] \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_13_U.bin_s1 ;
reg \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_13_U.carry_s1 ;
reg [16:0] \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_13_U.sum_s1 ;
reg [17:0] \add_36s_36s_36_2_1_U12.top_add_36s_36s_36_2_1_Adder_10_U.ain_s1 ;
reg [17:0] \add_36s_36s_36_2_1_U12.top_add_36s_36s_36_2_1_Adder_10_U.bin_s1 ;
reg \add_36s_36s_36_2_1_U12.top_add_36s_36s_36_2_1_Adder_10_U.carry_s1 ;
reg [17:0] \add_36s_36s_36_2_1_U12.top_add_36s_36s_36_2_1_Adder_10_U.sum_s1 ;
reg [18:0] \add_37s_37s_37_2_1_U7.top_add_37s_37s_37_2_1_Adder_6_U.ain_s1 ;
reg [18:0] \add_37s_37s_37_2_1_U7.top_add_37s_37s_37_2_1_Adder_6_U.bin_s1 ;
reg \add_37s_37s_37_2_1_U7.top_add_37s_37s_37_2_1_Adder_6_U.carry_s1 ;
reg [17:0] \add_37s_37s_37_2_1_U7.top_add_37s_37s_37_2_1_Adder_6_U.sum_s1 ;
reg [26:0] \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_12_U.ain_s1 ;
reg [26:0] \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_12_U.bin_s1 ;
reg \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_12_U.carry_s1 ;
reg [26:0] \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_12_U.sum_s1 ;
reg [2:0] \add_5s_5s_5_2_1_U5.top_add_5s_5s_5_2_1_Adder_4_U.ain_s1 ;
reg [2:0] \add_5s_5s_5_2_1_U5.top_add_5s_5s_5_2_1_Adder_4_U.bin_s1 ;
reg \add_5s_5s_5_2_1_U5.top_add_5s_5s_5_2_1_Adder_4_U.carry_s1 ;
reg [1:0] \add_5s_5s_5_2_1_U5.top_add_5s_5s_5_2_1_Adder_4_U.sum_s1 ;
reg [3:0] \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.ain_s1 ;
reg [3:0] \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.bin_s1 ;
reg \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.carry_s1 ;
reg [3:0] \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.sum_s1 ;
reg [31:0] add_ln691_1_reg_1456;
reg [31:0] add_ln691_2_reg_1498;
reg [31:0] add_ln691_3_reg_1550;
reg [17:0] add_ln691_reg_1368;
reg [31:0] add_ln69_reg_1513;
reg [2:0] and_ln731_reg_1403;
reg [37:0] ap_CS_fsm = 38'h0000000001;
reg icmp_ln1499_reg_1306;
reg icmp_ln768_1_reg_1127;
reg icmp_ln768_2_reg_1231;
reg icmp_ln768_reg_1176;
reg icmp_ln786_1_reg_1236;
reg icmp_ln786_reg_1181;
reg icmp_ln790_reg_1211;
reg icmp_ln851_1_reg_1341;
reg icmp_ln851_2_reg_1439;
reg icmp_ln851_3_reg_1476;
reg icmp_ln851_reg_1226;
reg [3:0] op_14_V_reg_1414;
reg [17:0] op_22_V_reg_1383;
reg [31:0] op_24_V_reg_1419;
reg [31:0] op_28_V_reg_1518;
reg [3:0] op_3_V_reg_1264;
reg [3:0] op_8_V_reg_1165;
reg [1:0] op_9_V_reg_1269;
reg [8:0] or_ln1195_reg_1279;
reg or_ln384_reg_1241;
reg overflow_2_reg_1258;
reg overflow_reg_1205;
reg p_Result_14_reg_1137;
reg p_Result_15_reg_1143;
reg p_Result_17_reg_1186;
reg p_Result_18_reg_1192;
reg [30:0] p_Result_s_reg_1149;
reg [7:0] ret_V_15_reg_1346;
reg [32:0] ret_V_16_reg_1246;
reg [36:0] ret_V_17_reg_1351;
reg [17:0] ret_V_18_reg_1373;
reg [17:0] ret_V_19_reg_1393;
reg [35:0] ret_V_20_reg_1444;
reg [53:0] ret_V_21_reg_1481;
reg [31:0] ret_V_22_reg_1508;
reg [31:0] ret_V_23_cast_reg_1449;
reg [33:0] ret_V_23_reg_1538;
reg [31:0] ret_V_24_reg_1555;
reg [31:0] ret_V_25_cast_reg_1486;
reg [31:0] ret_V_27_cast_reg_1543;
reg [15:0] ret_V_3_reg_1251;
reg [15:0] ret_V_4_reg_1291;
reg [4:0] ret_V_5_reg_1311;
reg [7:0] ret_V_cast_reg_1284;
reg [7:0] ret_V_reg_1326;
reg [32:0] ret_reg_1132;
reg rhs_3_reg_1120;
reg [31:0] select_ln1192_reg_1560;
reg [31:0] select_ln353_reg_1461;
reg [15:0] select_ln850_3_reg_1316;
reg [17:0] sext_ln850_reg_1361;
reg [8:0] \sub_17ns_17ns_17_2_1_U2.top_sub_17ns_17ns_17_2_1_Adder_1_U.ain_s1 ;
reg [8:0] \sub_17ns_17ns_17_2_1_U2.top_sub_17ns_17ns_17_2_1_Adder_1_U.bin_s1 ;
reg \sub_17ns_17ns_17_2_1_U2.top_sub_17ns_17ns_17_2_1_Adder_1_U.carry_s1 ;
reg [7:0] \sub_17ns_17ns_17_2_1_U2.top_sub_17ns_17ns_17_2_1_Adder_1_U.sum_s1 ;
reg [16:0] \sub_33s_33ns_33_2_1_U1.top_sub_33s_33ns_33_2_1_Adder_0_U.ain_s1 ;
reg [16:0] \sub_33s_33ns_33_2_1_U1.top_sub_33s_33ns_33_2_1_Adder_0_U.bin_s1 ;
reg \sub_33s_33ns_33_2_1_U1.top_sub_33s_33ns_33_2_1_Adder_0_U.carry_s1 ;
reg [15:0] \sub_33s_33ns_33_2_1_U1.top_sub_33s_33ns_33_2_1_Adder_0_U.sum_s1 ;
reg [15:0] tmp_4_reg_1199;
reg [16:0] tmp_6_reg_1356;
reg [7:0] trunc_ln728_reg_1115;
reg trunc_ln790_reg_1155;
reg [1:0] trunc_ln851_2_reg_1321;
reg [2:0] trunc_ln851_3_reg_1424;
wire [31:0] _000_;
wire [31:0] _001_;
wire [31:0] _002_;
wire [17:0] _003_;
wire [31:0] _004_;
wire [2:0] _005_;
wire [37:0] _006_;
wire _007_;
wire _008_;
wire _009_;
wire _010_;
wire _011_;
wire _012_;
wire _013_;
wire _014_;
wire _015_;
wire _016_;
wire _017_;
wire [2:0] _018_;
wire [17:0] _019_;
wire [31:0] _020_;
wire [31:0] _021_;
wire [3:0] _022_;
wire [3:0] _023_;
wire [1:0] _024_;
wire [8:0] _025_;
wire _026_;
wire _027_;
wire _028_;
wire _029_;
wire _030_;
wire _031_;
wire _032_;
wire [30:0] _033_;
wire [7:0] _034_;
wire [32:0] _035_;
wire [36:0] _036_;
wire [17:0] _037_;
wire [17:0] _038_;
wire [35:0] _039_;
wire [53:0] _040_;
wire [31:0] _041_;
wire [31:0] _042_;
wire [33:0] _043_;
wire [31:0] _044_;
wire [31:0] _045_;
wire [31:0] _046_;
wire [15:0] _047_;
wire [15:0] _048_;
wire [4:0] _049_;
wire [7:0] _050_;
wire [7:0] _051_;
wire [32:0] _052_;
wire _053_;
wire [31:0] _054_;
wire [31:0] _055_;
wire [15:0] _056_;
wire [17:0] _057_;
wire [15:0] _058_;
wire [16:0] _059_;
wire [7:0] _060_;
wire _061_;
wire [1:0] _062_;
wire [1:0] _063_;
wire [1:0] _064_;
wire _065_;
wire _066_;
wire _067_;
wire _068_;
wire _069_;
wire _070_;
wire _071_;
wire _072_;
wire _073_;
wire _074_;
wire _075_;
wire [7:0] _076_;
wire [7:0] _077_;
wire _078_;
wire [7:0] _079_;
wire [8:0] _080_;
wire [8:0] _081_;
wire [8:0] _082_;
wire [8:0] _083_;
wire _084_;
wire [8:0] _085_;
wire [9:0] _086_;
wire [9:0] _087_;
wire [8:0] _088_;
wire [8:0] _089_;
wire _090_;
wire [8:0] _091_;
wire [9:0] _092_;
wire [9:0] _093_;
wire [8:0] _094_;
wire [8:0] _095_;
wire _096_;
wire [8:0] _097_;
wire [9:0] _098_;
wire [9:0] _099_;
wire [15:0] _100_;
wire [15:0] _101_;
wire _102_;
wire [15:0] _103_;
wire [16:0] _104_;
wire [16:0] _105_;
wire [15:0] _106_;
wire [15:0] _107_;
wire _108_;
wire [15:0] _109_;
wire [16:0] _110_;
wire [16:0] _111_;
wire [15:0] _112_;
wire [15:0] _113_;
wire _114_;
wire [15:0] _115_;
wire [16:0] _116_;
wire [16:0] _117_;
wire [15:0] _118_;
wire [15:0] _119_;
wire _120_;
wire [15:0] _121_;
wire [16:0] _122_;
wire [16:0] _123_;
wire [15:0] _124_;
wire [15:0] _125_;
wire _126_;
wire [15:0] _127_;
wire [16:0] _128_;
wire [16:0] _129_;
wire [15:0] _130_;
wire [15:0] _131_;
wire _132_;
wire [15:0] _133_;
wire [16:0] _134_;
wire [16:0] _135_;
wire [15:0] _136_;
wire [15:0] _137_;
wire _138_;
wire [15:0] _139_;
wire [16:0] _140_;
wire [16:0] _141_;
wire [16:0] _142_;
wire [16:0] _143_;
wire _144_;
wire [15:0] _145_;
wire [16:0] _146_;
wire [17:0] _147_;
wire [16:0] _148_;
wire [16:0] _149_;
wire _150_;
wire [16:0] _151_;
wire [17:0] _152_;
wire [17:0] _153_;
wire [17:0] _154_;
wire [17:0] _155_;
wire _156_;
wire [17:0] _157_;
wire [18:0] _158_;
wire [18:0] _159_;
wire [18:0] _160_;
wire [18:0] _161_;
wire _162_;
wire [17:0] _163_;
wire [18:0] _164_;
wire [19:0] _165_;
wire [26:0] _166_;
wire [26:0] _167_;
wire _168_;
wire [26:0] _169_;
wire [27:0] _170_;
wire [27:0] _171_;
wire [2:0] _172_;
wire [2:0] _173_;
wire _174_;
wire [1:0] _175_;
wire [2:0] _176_;
wire [3:0] _177_;
wire [3:0] _178_;
wire [3:0] _179_;
wire _180_;
wire [3:0] _181_;
wire [4:0] _182_;
wire [4:0] _183_;
wire [8:0] _184_;
wire [8:0] _185_;
wire _186_;
wire [7:0] _187_;
wire [8:0] _188_;
wire [9:0] _189_;
wire [16:0] _190_;
wire [16:0] _191_;
wire _192_;
wire [15:0] _193_;
wire [16:0] _194_;
wire [17:0] _195_;
wire _196_;
wire _197_;
wire _198_;
wire _199_;
wire _200_;
wire _201_;
wire _202_;
wire _203_;
wire _204_;
wire _205_;
wire _206_;
wire _207_;
wire _208_;
wire _209_;
wire _210_;
wire _211_;
wire _212_;
wire _213_;
wire _214_;
wire _215_;
wire _216_;
wire _217_;
wire _218_;
wire _219_;
wire _220_;
wire _221_;
wire _222_;
wire _223_;
wire _224_;
wire _225_;
wire _226_;
wire _227_;
wire _228_;
wire _229_;
wire _230_;
wire _231_;
wire _232_;
wire _233_;
wire _234_;
wire _235_;
wire _236_;
wire _237_;
wire _238_;
wire _239_;
wire _240_;
wire _241_;
wire _242_;
wire \add_16ns_16ns_16_2_1_U4.ce ;
wire \add_16ns_16ns_16_2_1_U4.clk ;
wire [15:0] \add_16ns_16ns_16_2_1_U4.din0 ;
wire [15:0] \add_16ns_16ns_16_2_1_U4.din1 ;
wire [15:0] \add_16ns_16ns_16_2_1_U4.dout ;
wire \add_16ns_16ns_16_2_1_U4.reset ;
wire [15:0] \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_3_U.a ;
wire [15:0] \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_3_U.ain_s0 ;
wire [15:0] \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_3_U.b ;
wire [15:0] \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_3_U.bin_s0 ;
wire \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_3_U.ce ;
wire \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_3_U.clk ;
wire \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_3_U.facout_s1 ;
wire \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_3_U.facout_s2 ;
wire [7:0] \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_3_U.fas_s1 ;
wire [7:0] \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_3_U.fas_s2 ;
wire \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_3_U.reset ;
wire [15:0] \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_3_U.s ;
wire [7:0] \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_3_U.u1.a ;
wire [7:0] \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_3_U.u1.b ;
wire \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_3_U.u1.cin ;
wire \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_3_U.u1.cout ;
wire [7:0] \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_3_U.u1.s ;
wire [7:0] \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_3_U.u2.a ;
wire [7:0] \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_3_U.u2.b ;
wire \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_3_U.u2.cin ;
wire \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_3_U.u2.cout ;
wire [7:0] \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_3_U.u2.s ;
wire \add_18ns_18s_18_2_1_U10.ce ;
wire \add_18ns_18s_18_2_1_U10.clk ;
wire [17:0] \add_18ns_18s_18_2_1_U10.din0 ;
wire [17:0] \add_18ns_18s_18_2_1_U10.din1 ;
wire [17:0] \add_18ns_18s_18_2_1_U10.dout ;
wire \add_18ns_18s_18_2_1_U10.reset ;
wire [17:0] \add_18ns_18s_18_2_1_U10.top_add_18ns_18s_18_2_1_Adder_8_U.a ;
wire [17:0] \add_18ns_18s_18_2_1_U10.top_add_18ns_18s_18_2_1_Adder_8_U.ain_s0 ;
wire [17:0] \add_18ns_18s_18_2_1_U10.top_add_18ns_18s_18_2_1_Adder_8_U.b ;
wire [17:0] \add_18ns_18s_18_2_1_U10.top_add_18ns_18s_18_2_1_Adder_8_U.bin_s0 ;
wire \add_18ns_18s_18_2_1_U10.top_add_18ns_18s_18_2_1_Adder_8_U.ce ;
wire \add_18ns_18s_18_2_1_U10.top_add_18ns_18s_18_2_1_Adder_8_U.clk ;
wire \add_18ns_18s_18_2_1_U10.top_add_18ns_18s_18_2_1_Adder_8_U.facout_s1 ;
wire \add_18ns_18s_18_2_1_U10.top_add_18ns_18s_18_2_1_Adder_8_U.facout_s2 ;
wire [8:0] \add_18ns_18s_18_2_1_U10.top_add_18ns_18s_18_2_1_Adder_8_U.fas_s1 ;
wire [8:0] \add_18ns_18s_18_2_1_U10.top_add_18ns_18s_18_2_1_Adder_8_U.fas_s2 ;
wire \add_18ns_18s_18_2_1_U10.top_add_18ns_18s_18_2_1_Adder_8_U.reset ;
wire [17:0] \add_18ns_18s_18_2_1_U10.top_add_18ns_18s_18_2_1_Adder_8_U.s ;
wire [8:0] \add_18ns_18s_18_2_1_U10.top_add_18ns_18s_18_2_1_Adder_8_U.u1.a ;
wire [8:0] \add_18ns_18s_18_2_1_U10.top_add_18ns_18s_18_2_1_Adder_8_U.u1.b ;
wire \add_18ns_18s_18_2_1_U10.top_add_18ns_18s_18_2_1_Adder_8_U.u1.cin ;
wire \add_18ns_18s_18_2_1_U10.top_add_18ns_18s_18_2_1_Adder_8_U.u1.cout ;
wire [8:0] \add_18ns_18s_18_2_1_U10.top_add_18ns_18s_18_2_1_Adder_8_U.u1.s ;
wire [8:0] \add_18ns_18s_18_2_1_U10.top_add_18ns_18s_18_2_1_Adder_8_U.u2.a ;
wire [8:0] \add_18ns_18s_18_2_1_U10.top_add_18ns_18s_18_2_1_Adder_8_U.u2.b ;
wire \add_18ns_18s_18_2_1_U10.top_add_18ns_18s_18_2_1_Adder_8_U.u2.cin ;
wire \add_18ns_18s_18_2_1_U10.top_add_18ns_18s_18_2_1_Adder_8_U.u2.cout ;
wire [8:0] \add_18ns_18s_18_2_1_U10.top_add_18ns_18s_18_2_1_Adder_8_U.u2.s ;
wire \add_18ns_18s_18_2_1_U9.ce ;
wire \add_18ns_18s_18_2_1_U9.clk ;
wire [17:0] \add_18ns_18s_18_2_1_U9.din0 ;
wire [17:0] \add_18ns_18s_18_2_1_U9.din1 ;
wire [17:0] \add_18ns_18s_18_2_1_U9.dout ;
wire \add_18ns_18s_18_2_1_U9.reset ;
wire [17:0] \add_18ns_18s_18_2_1_U9.top_add_18ns_18s_18_2_1_Adder_8_U.a ;
wire [17:0] \add_18ns_18s_18_2_1_U9.top_add_18ns_18s_18_2_1_Adder_8_U.ain_s0 ;
wire [17:0] \add_18ns_18s_18_2_1_U9.top_add_18ns_18s_18_2_1_Adder_8_U.b ;
wire [17:0] \add_18ns_18s_18_2_1_U9.top_add_18ns_18s_18_2_1_Adder_8_U.bin_s0 ;
wire \add_18ns_18s_18_2_1_U9.top_add_18ns_18s_18_2_1_Adder_8_U.ce ;
wire \add_18ns_18s_18_2_1_U9.top_add_18ns_18s_18_2_1_Adder_8_U.clk ;
wire \add_18ns_18s_18_2_1_U9.top_add_18ns_18s_18_2_1_Adder_8_U.facout_s1 ;
wire \add_18ns_18s_18_2_1_U9.top_add_18ns_18s_18_2_1_Adder_8_U.facout_s2 ;
wire [8:0] \add_18ns_18s_18_2_1_U9.top_add_18ns_18s_18_2_1_Adder_8_U.fas_s1 ;
wire [8:0] \add_18ns_18s_18_2_1_U9.top_add_18ns_18s_18_2_1_Adder_8_U.fas_s2 ;
wire \add_18ns_18s_18_2_1_U9.top_add_18ns_18s_18_2_1_Adder_8_U.reset ;
wire [17:0] \add_18ns_18s_18_2_1_U9.top_add_18ns_18s_18_2_1_Adder_8_U.s ;
wire [8:0] \add_18ns_18s_18_2_1_U9.top_add_18ns_18s_18_2_1_Adder_8_U.u1.a ;
wire [8:0] \add_18ns_18s_18_2_1_U9.top_add_18ns_18s_18_2_1_Adder_8_U.u1.b ;
wire \add_18ns_18s_18_2_1_U9.top_add_18ns_18s_18_2_1_Adder_8_U.u1.cin ;
wire \add_18ns_18s_18_2_1_U9.top_add_18ns_18s_18_2_1_Adder_8_U.u1.cout ;
wire [8:0] \add_18ns_18s_18_2_1_U9.top_add_18ns_18s_18_2_1_Adder_8_U.u1.s ;
wire [8:0] \add_18ns_18s_18_2_1_U9.top_add_18ns_18s_18_2_1_Adder_8_U.u2.a ;
wire [8:0] \add_18ns_18s_18_2_1_U9.top_add_18ns_18s_18_2_1_Adder_8_U.u2.b ;
wire \add_18ns_18s_18_2_1_U9.top_add_18ns_18s_18_2_1_Adder_8_U.u2.cin ;
wire \add_18ns_18s_18_2_1_U9.top_add_18ns_18s_18_2_1_Adder_8_U.u2.cout ;
wire [8:0] \add_18ns_18s_18_2_1_U9.top_add_18ns_18s_18_2_1_Adder_8_U.u2.s ;
wire \add_18s_18ns_18_2_1_U8.ce ;
wire \add_18s_18ns_18_2_1_U8.clk ;
wire [17:0] \add_18s_18ns_18_2_1_U8.din0 ;
wire [17:0] \add_18s_18ns_18_2_1_U8.din1 ;
wire [17:0] \add_18s_18ns_18_2_1_U8.dout ;
wire \add_18s_18ns_18_2_1_U8.reset ;
wire [17:0] \add_18s_18ns_18_2_1_U8.top_add_18s_18ns_18_2_1_Adder_7_U.a ;
wire [17:0] \add_18s_18ns_18_2_1_U8.top_add_18s_18ns_18_2_1_Adder_7_U.ain_s0 ;
wire [17:0] \add_18s_18ns_18_2_1_U8.top_add_18s_18ns_18_2_1_Adder_7_U.b ;
wire [17:0] \add_18s_18ns_18_2_1_U8.top_add_18s_18ns_18_2_1_Adder_7_U.bin_s0 ;
wire \add_18s_18ns_18_2_1_U8.top_add_18s_18ns_18_2_1_Adder_7_U.ce ;
wire \add_18s_18ns_18_2_1_U8.top_add_18s_18ns_18_2_1_Adder_7_U.clk ;
wire \add_18s_18ns_18_2_1_U8.top_add_18s_18ns_18_2_1_Adder_7_U.facout_s1 ;
wire \add_18s_18ns_18_2_1_U8.top_add_18s_18ns_18_2_1_Adder_7_U.facout_s2 ;
wire [8:0] \add_18s_18ns_18_2_1_U8.top_add_18s_18ns_18_2_1_Adder_7_U.fas_s1 ;
wire [8:0] \add_18s_18ns_18_2_1_U8.top_add_18s_18ns_18_2_1_Adder_7_U.fas_s2 ;
wire \add_18s_18ns_18_2_1_U8.top_add_18s_18ns_18_2_1_Adder_7_U.reset ;
wire [17:0] \add_18s_18ns_18_2_1_U8.top_add_18s_18ns_18_2_1_Adder_7_U.s ;
wire [8:0] \add_18s_18ns_18_2_1_U8.top_add_18s_18ns_18_2_1_Adder_7_U.u1.a ;
wire [8:0] \add_18s_18ns_18_2_1_U8.top_add_18s_18ns_18_2_1_Adder_7_U.u1.b ;
wire \add_18s_18ns_18_2_1_U8.top_add_18s_18ns_18_2_1_Adder_7_U.u1.cin ;
wire \add_18s_18ns_18_2_1_U8.top_add_18s_18ns_18_2_1_Adder_7_U.u1.cout ;
wire [8:0] \add_18s_18ns_18_2_1_U8.top_add_18s_18ns_18_2_1_Adder_7_U.u1.s ;
wire [8:0] \add_18s_18ns_18_2_1_U8.top_add_18s_18ns_18_2_1_Adder_7_U.u2.a ;
wire [8:0] \add_18s_18ns_18_2_1_U8.top_add_18s_18ns_18_2_1_Adder_7_U.u2.b ;
wire \add_18s_18ns_18_2_1_U8.top_add_18s_18ns_18_2_1_Adder_7_U.u2.cin ;
wire \add_18s_18ns_18_2_1_U8.top_add_18s_18ns_18_2_1_Adder_7_U.u2.cout ;
wire [8:0] \add_18s_18ns_18_2_1_U8.top_add_18s_18ns_18_2_1_Adder_7_U.u2.s ;
wire \add_32ns_32ns_32_2_1_U13.ce ;
wire \add_32ns_32ns_32_2_1_U13.clk ;
wire [31:0] \add_32ns_32ns_32_2_1_U13.din0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U13.din1 ;
wire [31:0] \add_32ns_32ns_32_2_1_U13.dout ;
wire \add_32ns_32ns_32_2_1_U13.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_11_U.a ;
wire [31:0] \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_11_U.ain_s0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_11_U.b ;
wire [31:0] \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_11_U.bin_s0 ;
wire \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_11_U.ce ;
wire \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_11_U.clk ;
wire \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_11_U.facout_s1 ;
wire \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_11_U.facout_s2 ;
wire [15:0] \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_11_U.fas_s1 ;
wire [15:0] \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_11_U.fas_s2 ;
wire \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_11_U.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_11_U.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.b ;
wire \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.cin ;
wire \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.b ;
wire \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.cin ;
wire \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.s ;
wire \add_32ns_32ns_32_2_1_U15.ce ;
wire \add_32ns_32ns_32_2_1_U15.clk ;
wire [31:0] \add_32ns_32ns_32_2_1_U15.din0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U15.din1 ;
wire [31:0] \add_32ns_32ns_32_2_1_U15.dout ;
wire \add_32ns_32ns_32_2_1_U15.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.a ;
wire [31:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.ain_s0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.b ;
wire [31:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.bin_s0 ;
wire \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.ce ;
wire \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.clk ;
wire \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.facout_s1 ;
wire \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.facout_s2 ;
wire [15:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.fas_s1 ;
wire [15:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.fas_s2 ;
wire \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.b ;
wire \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.cin ;
wire \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.b ;
wire \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.cin ;
wire \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.s ;
wire \add_32ns_32ns_32_2_1_U16.ce ;
wire \add_32ns_32ns_32_2_1_U16.clk ;
wire [31:0] \add_32ns_32ns_32_2_1_U16.din0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U16.din1 ;
wire [31:0] \add_32ns_32ns_32_2_1_U16.dout ;
wire \add_32ns_32ns_32_2_1_U16.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.a ;
wire [31:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.ain_s0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.b ;
wire [31:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.bin_s0 ;
wire \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.ce ;
wire \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.clk ;
wire \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.facout_s1 ;
wire \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.facout_s2 ;
wire [15:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.fas_s1 ;
wire [15:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.fas_s2 ;
wire \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.b ;
wire \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.cin ;
wire \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.b ;
wire \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.cin ;
wire \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.s ;
wire \add_32ns_32ns_32_2_1_U17.ce ;
wire \add_32ns_32ns_32_2_1_U17.clk ;
wire [31:0] \add_32ns_32ns_32_2_1_U17.din0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U17.din1 ;
wire [31:0] \add_32ns_32ns_32_2_1_U17.dout ;
wire \add_32ns_32ns_32_2_1_U17.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.a ;
wire [31:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.ain_s0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.b ;
wire [31:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.bin_s0 ;
wire \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.ce ;
wire \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.clk ;
wire \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.facout_s1 ;
wire \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.facout_s2 ;
wire [15:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.fas_s1 ;
wire [15:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.fas_s2 ;
wire \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.b ;
wire \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.cin ;
wire \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.b ;
wire \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.cin ;
wire \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.s ;
wire \add_32ns_32ns_32_2_1_U19.ce ;
wire \add_32ns_32ns_32_2_1_U19.clk ;
wire [31:0] \add_32ns_32ns_32_2_1_U19.din0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U19.din1 ;
wire [31:0] \add_32ns_32ns_32_2_1_U19.dout ;
wire \add_32ns_32ns_32_2_1_U19.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.a ;
wire [31:0] \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.ain_s0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.b ;
wire [31:0] \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.bin_s0 ;
wire \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.ce ;
wire \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.clk ;
wire \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.facout_s1 ;
wire \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.facout_s2 ;
wire [15:0] \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.fas_s1 ;
wire [15:0] \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.fas_s2 ;
wire \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.b ;
wire \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.cin ;
wire \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.b ;
wire \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.cin ;
wire \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.s ;
wire \add_32ns_32ns_32_2_1_U20.ce ;
wire \add_32ns_32ns_32_2_1_U20.clk ;
wire [31:0] \add_32ns_32ns_32_2_1_U20.din0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U20.din1 ;
wire [31:0] \add_32ns_32ns_32_2_1_U20.dout ;
wire \add_32ns_32ns_32_2_1_U20.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.a ;
wire [31:0] \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.ain_s0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.b ;
wire [31:0] \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.bin_s0 ;
wire \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.ce ;
wire \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.clk ;
wire \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.facout_s1 ;
wire \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.facout_s2 ;
wire [15:0] \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.fas_s1 ;
wire [15:0] \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.fas_s2 ;
wire \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.b ;
wire \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.cin ;
wire \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.b ;
wire \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.cin ;
wire \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.s ;
wire \add_32s_32ns_32_2_1_U11.ce ;
wire \add_32s_32ns_32_2_1_U11.clk ;
wire [31:0] \add_32s_32ns_32_2_1_U11.din0 ;
wire [31:0] \add_32s_32ns_32_2_1_U11.din1 ;
wire [31:0] \add_32s_32ns_32_2_1_U11.dout ;
wire \add_32s_32ns_32_2_1_U11.reset ;
wire [31:0] \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_9_U.a ;
wire [31:0] \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_9_U.ain_s0 ;
wire [31:0] \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_9_U.b ;
wire [31:0] \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_9_U.bin_s0 ;
wire \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_9_U.ce ;
wire \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_9_U.clk ;
wire \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_9_U.facout_s1 ;
wire \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_9_U.facout_s2 ;
wire [15:0] \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_9_U.fas_s1 ;
wire [15:0] \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_9_U.fas_s2 ;
wire \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_9_U.reset ;
wire [31:0] \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_9_U.s ;
wire [15:0] \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_9_U.u1.a ;
wire [15:0] \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_9_U.u1.b ;
wire \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_9_U.u1.cin ;
wire \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_9_U.u1.cout ;
wire [15:0] \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_9_U.u1.s ;
wire [15:0] \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_9_U.u2.a ;
wire [15:0] \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_9_U.u2.b ;
wire \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_9_U.u2.cin ;
wire \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_9_U.u2.cout ;
wire [15:0] \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_9_U.u2.s ;
wire \add_33ns_33s_33_2_1_U3.ce ;
wire \add_33ns_33s_33_2_1_U3.clk ;
wire [32:0] \add_33ns_33s_33_2_1_U3.din0 ;
wire [32:0] \add_33ns_33s_33_2_1_U3.din1 ;
wire [32:0] \add_33ns_33s_33_2_1_U3.dout ;
wire \add_33ns_33s_33_2_1_U3.reset ;
wire [32:0] \add_33ns_33s_33_2_1_U3.top_add_33ns_33s_33_2_1_Adder_2_U.a ;
wire [32:0] \add_33ns_33s_33_2_1_U3.top_add_33ns_33s_33_2_1_Adder_2_U.ain_s0 ;
wire [32:0] \add_33ns_33s_33_2_1_U3.top_add_33ns_33s_33_2_1_Adder_2_U.b ;
wire [32:0] \add_33ns_33s_33_2_1_U3.top_add_33ns_33s_33_2_1_Adder_2_U.bin_s0 ;
wire \add_33ns_33s_33_2_1_U3.top_add_33ns_33s_33_2_1_Adder_2_U.ce ;
wire \add_33ns_33s_33_2_1_U3.top_add_33ns_33s_33_2_1_Adder_2_U.clk ;
wire \add_33ns_33s_33_2_1_U3.top_add_33ns_33s_33_2_1_Adder_2_U.facout_s1 ;
wire \add_33ns_33s_33_2_1_U3.top_add_33ns_33s_33_2_1_Adder_2_U.facout_s2 ;
wire [15:0] \add_33ns_33s_33_2_1_U3.top_add_33ns_33s_33_2_1_Adder_2_U.fas_s1 ;
wire [16:0] \add_33ns_33s_33_2_1_U3.top_add_33ns_33s_33_2_1_Adder_2_U.fas_s2 ;
wire \add_33ns_33s_33_2_1_U3.top_add_33ns_33s_33_2_1_Adder_2_U.reset ;
wire [32:0] \add_33ns_33s_33_2_1_U3.top_add_33ns_33s_33_2_1_Adder_2_U.s ;
wire [15:0] \add_33ns_33s_33_2_1_U3.top_add_33ns_33s_33_2_1_Adder_2_U.u1.a ;
wire [15:0] \add_33ns_33s_33_2_1_U3.top_add_33ns_33s_33_2_1_Adder_2_U.u1.b ;
wire \add_33ns_33s_33_2_1_U3.top_add_33ns_33s_33_2_1_Adder_2_U.u1.cin ;
wire \add_33ns_33s_33_2_1_U3.top_add_33ns_33s_33_2_1_Adder_2_U.u1.cout ;
wire [15:0] \add_33ns_33s_33_2_1_U3.top_add_33ns_33s_33_2_1_Adder_2_U.u1.s ;
wire [16:0] \add_33ns_33s_33_2_1_U3.top_add_33ns_33s_33_2_1_Adder_2_U.u2.a ;
wire [16:0] \add_33ns_33s_33_2_1_U3.top_add_33ns_33s_33_2_1_Adder_2_U.u2.b ;
wire \add_33ns_33s_33_2_1_U3.top_add_33ns_33s_33_2_1_Adder_2_U.u2.cin ;
wire \add_33ns_33s_33_2_1_U3.top_add_33ns_33s_33_2_1_Adder_2_U.u2.cout ;
wire [16:0] \add_33ns_33s_33_2_1_U3.top_add_33ns_33s_33_2_1_Adder_2_U.u2.s ;
wire \add_34s_34s_34_2_1_U18.ce ;
wire \add_34s_34s_34_2_1_U18.clk ;
wire [33:0] \add_34s_34s_34_2_1_U18.din0 ;
wire [33:0] \add_34s_34s_34_2_1_U18.din1 ;
wire [33:0] \add_34s_34s_34_2_1_U18.dout ;
wire \add_34s_34s_34_2_1_U18.reset ;
wire [33:0] \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_13_U.a ;
wire [33:0] \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_13_U.ain_s0 ;
wire [33:0] \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_13_U.b ;
wire [33:0] \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_13_U.bin_s0 ;
wire \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_13_U.ce ;
wire \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_13_U.clk ;
wire \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_13_U.facout_s1 ;
wire \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_13_U.facout_s2 ;
wire [16:0] \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_13_U.fas_s1 ;
wire [16:0] \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_13_U.fas_s2 ;
wire \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_13_U.reset ;
wire [33:0] \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_13_U.s ;
wire [16:0] \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_13_U.u1.a ;
wire [16:0] \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_13_U.u1.b ;
wire \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_13_U.u1.cin ;
wire \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_13_U.u1.cout ;
wire [16:0] \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_13_U.u1.s ;
wire [16:0] \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_13_U.u2.a ;
wire [16:0] \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_13_U.u2.b ;
wire \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_13_U.u2.cin ;
wire \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_13_U.u2.cout ;
wire [16:0] \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_13_U.u2.s ;
wire \add_36s_36s_36_2_1_U12.ce ;
wire \add_36s_36s_36_2_1_U12.clk ;
wire [35:0] \add_36s_36s_36_2_1_U12.din0 ;
wire [35:0] \add_36s_36s_36_2_1_U12.din1 ;
wire [35:0] \add_36s_36s_36_2_1_U12.dout ;
wire \add_36s_36s_36_2_1_U12.reset ;
wire [35:0] \add_36s_36s_36_2_1_U12.top_add_36s_36s_36_2_1_Adder_10_U.a ;
wire [35:0] \add_36s_36s_36_2_1_U12.top_add_36s_36s_36_2_1_Adder_10_U.ain_s0 ;
wire [35:0] \add_36s_36s_36_2_1_U12.top_add_36s_36s_36_2_1_Adder_10_U.b ;
wire [35:0] \add_36s_36s_36_2_1_U12.top_add_36s_36s_36_2_1_Adder_10_U.bin_s0 ;
wire \add_36s_36s_36_2_1_U12.top_add_36s_36s_36_2_1_Adder_10_U.ce ;
wire \add_36s_36s_36_2_1_U12.top_add_36s_36s_36_2_1_Adder_10_U.clk ;
wire \add_36s_36s_36_2_1_U12.top_add_36s_36s_36_2_1_Adder_10_U.facout_s1 ;
wire \add_36s_36s_36_2_1_U12.top_add_36s_36s_36_2_1_Adder_10_U.facout_s2 ;
wire [17:0] \add_36s_36s_36_2_1_U12.top_add_36s_36s_36_2_1_Adder_10_U.fas_s1 ;
wire [17:0] \add_36s_36s_36_2_1_U12.top_add_36s_36s_36_2_1_Adder_10_U.fas_s2 ;
wire \add_36s_36s_36_2_1_U12.top_add_36s_36s_36_2_1_Adder_10_U.reset ;
wire [35:0] \add_36s_36s_36_2_1_U12.top_add_36s_36s_36_2_1_Adder_10_U.s ;
wire [17:0] \add_36s_36s_36_2_1_U12.top_add_36s_36s_36_2_1_Adder_10_U.u1.a ;
wire [17:0] \add_36s_36s_36_2_1_U12.top_add_36s_36s_36_2_1_Adder_10_U.u1.b ;
wire \add_36s_36s_36_2_1_U12.top_add_36s_36s_36_2_1_Adder_10_U.u1.cin ;
wire \add_36s_36s_36_2_1_U12.top_add_36s_36s_36_2_1_Adder_10_U.u1.cout ;
wire [17:0] \add_36s_36s_36_2_1_U12.top_add_36s_36s_36_2_1_Adder_10_U.u1.s ;
wire [17:0] \add_36s_36s_36_2_1_U12.top_add_36s_36s_36_2_1_Adder_10_U.u2.a ;
wire [17:0] \add_36s_36s_36_2_1_U12.top_add_36s_36s_36_2_1_Adder_10_U.u2.b ;
wire \add_36s_36s_36_2_1_U12.top_add_36s_36s_36_2_1_Adder_10_U.u2.cin ;
wire \add_36s_36s_36_2_1_U12.top_add_36s_36s_36_2_1_Adder_10_U.u2.cout ;
wire [17:0] \add_36s_36s_36_2_1_U12.top_add_36s_36s_36_2_1_Adder_10_U.u2.s ;
wire \add_37s_37s_37_2_1_U7.ce ;
wire \add_37s_37s_37_2_1_U7.clk ;
wire [36:0] \add_37s_37s_37_2_1_U7.din0 ;
wire [36:0] \add_37s_37s_37_2_1_U7.din1 ;
wire [36:0] \add_37s_37s_37_2_1_U7.dout ;
wire \add_37s_37s_37_2_1_U7.reset ;
wire [36:0] \add_37s_37s_37_2_1_U7.top_add_37s_37s_37_2_1_Adder_6_U.a ;
wire [36:0] \add_37s_37s_37_2_1_U7.top_add_37s_37s_37_2_1_Adder_6_U.ain_s0 ;
wire [36:0] \add_37s_37s_37_2_1_U7.top_add_37s_37s_37_2_1_Adder_6_U.b ;
wire [36:0] \add_37s_37s_37_2_1_U7.top_add_37s_37s_37_2_1_Adder_6_U.bin_s0 ;
wire \add_37s_37s_37_2_1_U7.top_add_37s_37s_37_2_1_Adder_6_U.ce ;
wire \add_37s_37s_37_2_1_U7.top_add_37s_37s_37_2_1_Adder_6_U.clk ;
wire \add_37s_37s_37_2_1_U7.top_add_37s_37s_37_2_1_Adder_6_U.facout_s1 ;
wire \add_37s_37s_37_2_1_U7.top_add_37s_37s_37_2_1_Adder_6_U.facout_s2 ;
wire [17:0] \add_37s_37s_37_2_1_U7.top_add_37s_37s_37_2_1_Adder_6_U.fas_s1 ;
wire [18:0] \add_37s_37s_37_2_1_U7.top_add_37s_37s_37_2_1_Adder_6_U.fas_s2 ;
wire \add_37s_37s_37_2_1_U7.top_add_37s_37s_37_2_1_Adder_6_U.reset ;
wire [36:0] \add_37s_37s_37_2_1_U7.top_add_37s_37s_37_2_1_Adder_6_U.s ;
wire [17:0] \add_37s_37s_37_2_1_U7.top_add_37s_37s_37_2_1_Adder_6_U.u1.a ;
wire [17:0] \add_37s_37s_37_2_1_U7.top_add_37s_37s_37_2_1_Adder_6_U.u1.b ;
wire \add_37s_37s_37_2_1_U7.top_add_37s_37s_37_2_1_Adder_6_U.u1.cin ;
wire \add_37s_37s_37_2_1_U7.top_add_37s_37s_37_2_1_Adder_6_U.u1.cout ;
wire [17:0] \add_37s_37s_37_2_1_U7.top_add_37s_37s_37_2_1_Adder_6_U.u1.s ;
wire [18:0] \add_37s_37s_37_2_1_U7.top_add_37s_37s_37_2_1_Adder_6_U.u2.a ;
wire [18:0] \add_37s_37s_37_2_1_U7.top_add_37s_37s_37_2_1_Adder_6_U.u2.b ;
wire \add_37s_37s_37_2_1_U7.top_add_37s_37s_37_2_1_Adder_6_U.u2.cin ;
wire \add_37s_37s_37_2_1_U7.top_add_37s_37s_37_2_1_Adder_6_U.u2.cout ;
wire [18:0] \add_37s_37s_37_2_1_U7.top_add_37s_37s_37_2_1_Adder_6_U.u2.s ;
wire \add_54s_54s_54_2_1_U14.ce ;
wire \add_54s_54s_54_2_1_U14.clk ;
wire [53:0] \add_54s_54s_54_2_1_U14.din0 ;
wire [53:0] \add_54s_54s_54_2_1_U14.din1 ;
wire [53:0] \add_54s_54s_54_2_1_U14.dout ;
wire \add_54s_54s_54_2_1_U14.reset ;
wire [53:0] \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_12_U.a ;
wire [53:0] \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_12_U.ain_s0 ;
wire [53:0] \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_12_U.b ;
wire [53:0] \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_12_U.bin_s0 ;
wire \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_12_U.ce ;
wire \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_12_U.clk ;
wire \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_12_U.facout_s1 ;
wire \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_12_U.facout_s2 ;
wire [26:0] \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_12_U.fas_s1 ;
wire [26:0] \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_12_U.fas_s2 ;
wire \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_12_U.reset ;
wire [53:0] \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_12_U.s ;
wire [26:0] \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_12_U.u1.a ;
wire [26:0] \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_12_U.u1.b ;
wire \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_12_U.u1.cin ;
wire \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_12_U.u1.cout ;
wire [26:0] \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_12_U.u1.s ;
wire [26:0] \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_12_U.u2.a ;
wire [26:0] \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_12_U.u2.b ;
wire \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_12_U.u2.cin ;
wire \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_12_U.u2.cout ;
wire [26:0] \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_12_U.u2.s ;
wire \add_5s_5s_5_2_1_U5.ce ;
wire \add_5s_5s_5_2_1_U5.clk ;
wire [4:0] \add_5s_5s_5_2_1_U5.din0 ;
wire [4:0] \add_5s_5s_5_2_1_U5.din1 ;
wire [4:0] \add_5s_5s_5_2_1_U5.dout ;
wire \add_5s_5s_5_2_1_U5.reset ;
wire [4:0] \add_5s_5s_5_2_1_U5.top_add_5s_5s_5_2_1_Adder_4_U.a ;
wire [4:0] \add_5s_5s_5_2_1_U5.top_add_5s_5s_5_2_1_Adder_4_U.ain_s0 ;
wire [4:0] \add_5s_5s_5_2_1_U5.top_add_5s_5s_5_2_1_Adder_4_U.b ;
wire [4:0] \add_5s_5s_5_2_1_U5.top_add_5s_5s_5_2_1_Adder_4_U.bin_s0 ;
wire \add_5s_5s_5_2_1_U5.top_add_5s_5s_5_2_1_Adder_4_U.ce ;
wire \add_5s_5s_5_2_1_U5.top_add_5s_5s_5_2_1_Adder_4_U.clk ;
wire \add_5s_5s_5_2_1_U5.top_add_5s_5s_5_2_1_Adder_4_U.facout_s1 ;
wire \add_5s_5s_5_2_1_U5.top_add_5s_5s_5_2_1_Adder_4_U.facout_s2 ;
wire [1:0] \add_5s_5s_5_2_1_U5.top_add_5s_5s_5_2_1_Adder_4_U.fas_s1 ;
wire [2:0] \add_5s_5s_5_2_1_U5.top_add_5s_5s_5_2_1_Adder_4_U.fas_s2 ;
wire \add_5s_5s_5_2_1_U5.top_add_5s_5s_5_2_1_Adder_4_U.reset ;
wire [4:0] \add_5s_5s_5_2_1_U5.top_add_5s_5s_5_2_1_Adder_4_U.s ;
wire [1:0] \add_5s_5s_5_2_1_U5.top_add_5s_5s_5_2_1_Adder_4_U.u1.a ;
wire [1:0] \add_5s_5s_5_2_1_U5.top_add_5s_5s_5_2_1_Adder_4_U.u1.b ;
wire \add_5s_5s_5_2_1_U5.top_add_5s_5s_5_2_1_Adder_4_U.u1.cin ;
wire \add_5s_5s_5_2_1_U5.top_add_5s_5s_5_2_1_Adder_4_U.u1.cout ;
wire [1:0] \add_5s_5s_5_2_1_U5.top_add_5s_5s_5_2_1_Adder_4_U.u1.s ;
wire [2:0] \add_5s_5s_5_2_1_U5.top_add_5s_5s_5_2_1_Adder_4_U.u2.a ;
wire [2:0] \add_5s_5s_5_2_1_U5.top_add_5s_5s_5_2_1_Adder_4_U.u2.b ;
wire \add_5s_5s_5_2_1_U5.top_add_5s_5s_5_2_1_Adder_4_U.u2.cin ;
wire \add_5s_5s_5_2_1_U5.top_add_5s_5s_5_2_1_Adder_4_U.u2.cout ;
wire [2:0] \add_5s_5s_5_2_1_U5.top_add_5s_5s_5_2_1_Adder_4_U.u2.s ;
wire \add_8ns_8ns_8_2_1_U6.ce ;
wire \add_8ns_8ns_8_2_1_U6.clk ;
wire [7:0] \add_8ns_8ns_8_2_1_U6.din0 ;
wire [7:0] \add_8ns_8ns_8_2_1_U6.din1 ;
wire [7:0] \add_8ns_8ns_8_2_1_U6.dout ;
wire \add_8ns_8ns_8_2_1_U6.reset ;
wire [7:0] \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.a ;
wire [7:0] \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.ain_s0 ;
wire [7:0] \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.b ;
wire [7:0] \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.bin_s0 ;
wire \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.ce ;
wire \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.clk ;
wire \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.facout_s1 ;
wire \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.facout_s2 ;
wire [3:0] \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.fas_s1 ;
wire [3:0] \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.fas_s2 ;
wire \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.reset ;
wire [7:0] \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.s ;
wire [3:0] \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.u1.a ;
wire [3:0] \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.u1.b ;
wire \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.u1.cin ;
wire \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.u1.cout ;
wire [3:0] \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.u1.s ;
wire [3:0] \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.u2.a ;
wire [3:0] \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.u2.b ;
wire \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.u2.cin ;
wire \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.u2.cout ;
wire [3:0] \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.u2.s ;
wire [2:0] and_ln731_fu_818_p2;
wire ap_CS_fsm_state1;
wire ap_CS_fsm_state10;
wire ap_CS_fsm_state11;
wire ap_CS_fsm_state12;
wire ap_CS_fsm_state13;
wire ap_CS_fsm_state14;
wire ap_CS_fsm_state15;
wire ap_CS_fsm_state16;
wire ap_CS_fsm_state17;
wire ap_CS_fsm_state18;
wire ap_CS_fsm_state19;
wire ap_CS_fsm_state2;
wire ap_CS_fsm_state20;
wire ap_CS_fsm_state21;
wire ap_CS_fsm_state22;
wire ap_CS_fsm_state23;
wire ap_CS_fsm_state24;
wire ap_CS_fsm_state25;
wire ap_CS_fsm_state26;
wire ap_CS_fsm_state27;
wire ap_CS_fsm_state28;
wire ap_CS_fsm_state29;
wire ap_CS_fsm_state3;
wire ap_CS_fsm_state30;
wire ap_CS_fsm_state31;
wire ap_CS_fsm_state32;
wire ap_CS_fsm_state33;
wire ap_CS_fsm_state34;
wire ap_CS_fsm_state35;
wire ap_CS_fsm_state36;
wire ap_CS_fsm_state37;
wire ap_CS_fsm_state38;
wire ap_CS_fsm_state4;
wire ap_CS_fsm_state5;
wire ap_CS_fsm_state6;
wire ap_CS_fsm_state7;
wire ap_CS_fsm_state8;
wire ap_CS_fsm_state9;
wire [37:0] ap_NS_fsm;
wire ap_clk;
wire ap_done;
wire ap_idle;
wire ap_ready;
wire ap_rst;
wire ap_start;
wire [31:0] grp_fu_1018_p2;
wire [33:0] grp_fu_1037_p0;
wire [33:0] grp_fu_1037_p1;
wire [33:0] grp_fu_1037_p2;
wire [31:0] grp_fu_1053_p2;
wire [31:0] grp_fu_1089_p2;
wire [32:0] grp_fu_275_p0;
wire [32:0] grp_fu_275_p1;
wire [32:0] grp_fu_275_p2;
wire [16:0] grp_fu_378_p0;
wire [16:0] grp_fu_378_p1;
wire [16:0] grp_fu_378_p2;
wire [32:0] grp_fu_460_p0;
wire [32:0] grp_fu_460_p1;
wire [32:0] grp_fu_460_p2;
wire [15:0] grp_fu_561_p2;
wire [4:0] grp_fu_650_p0;
wire [4:0] grp_fu_650_p1;
wire [4:0] grp_fu_650_p2;
wire [7:0] grp_fu_661_p2;
wire [36:0] grp_fu_711_p0;
wire [36:0] grp_fu_711_p1;
wire [36:0] grp_fu_711_p2;
wire [17:0] grp_fu_766_p0;
wire [17:0] grp_fu_766_p2;
wire [17:0] grp_fu_794_p1;
wire [17:0] grp_fu_794_p2;
wire [17:0] grp_fu_803_p1;
wire [17:0] grp_fu_803_p2;
wire [31:0] grp_fu_827_p0;
wire [31:0] grp_fu_827_p2;
wire [35:0] grp_fu_899_p0;
wire [35:0] grp_fu_899_p1;
wire [35:0] grp_fu_899_p2;
wire [31:0] grp_fu_920_p2;
wire [53:0] grp_fu_959_p0;
wire [53:0] grp_fu_959_p1;
wire [53:0] grp_fu_959_p2;
wire [31:0] grp_fu_985_p2;
wire [31:0] grp_fu_993_p0;
wire [31:0] grp_fu_993_p2;
wire [1:0] icmp_ln1499_fu_656_p1;
wire icmp_ln1499_fu_656_p2;
wire icmp_ln768_1_fu_305_p2;
wire icmp_ln768_2_fu_476_p2;
wire icmp_ln768_fu_384_p2;
wire icmp_ln786_1_fu_481_p2;
wire icmp_ln786_fu_389_p2;
wire icmp_ln790_fu_438_p2;
wire icmp_ln851_1_fu_724_p2;
wire icmp_ln851_2_fu_905_p2;
wire icmp_ln851_3_fu_969_p2;
wire icmp_ln851_fu_470_p2;
wire [24:0] lhs_V_fu_444_p3;
wire [8:0] lhs_cast_fu_608_p3;
wire [7:0] op_0;
wire [31:0] op_1;
wire [22:0] op_10_V_fu_689_p3;
wire [1:0] op_12;
wire [31:0] op_13;
wire [3:0] op_14_V_fu_873_p3;
wire [31:0] op_15;
wire [31:0] op_16;
wire [1:0] op_18;
wire op_19;
wire [15:0] op_2;
wire [31:0] op_30;
wire op_30_ap_vld;
wire [3:0] op_3_V_fu_554_p3;
wire [31:0] op_4_V_fu_263_p0;
wire [3:0] op_4_V_fu_263_p1;
wire [1:0] op_5;
wire [31:0] op_7;
wire [3:0] op_8_V_fu_367_p3;
wire [1:0] op_9_V_fu_600_p3;
wire [8:0] or_ln1195_fu_619_p2;
wire or_ln384_1_fu_595_p2;
wire or_ln384_fu_506_p2;
wire or_ln785_2_fu_521_p2;
wire or_ln785_fu_416_p2;
wire or_ln786_fu_578_p2;
wire or_ln788_1_fu_496_p2;
wire or_ln788_fu_491_p2;
wire overflow_1_fu_362_p2;
wire overflow_2_fu_530_p2;
wire overflow_3_fu_867_p2;
wire overflow_fu_425_p2;
wire p_Result_10_fu_772_p3;
wire p_Result_11_fu_925_p3;
wire p_Result_12_fu_999_p3;
wire p_Result_13_fu_1058_p3;
wire [31:0] p_Result_16_fu_355_p1;
wire p_Result_16_fu_355_p3;
wire p_Result_18_fu_402_p1;
wire p_Result_19_fu_852_p3;
wire [1:0] p_Result_3_fu_730_p1;
wire p_Result_3_fu_730_p3;
wire p_Result_4_fu_666_p3;
wire [19:0] p_Result_9_fu_717_p3;
wire [2:0] p_Result_s_20_fu_431_p3;
wire [3:0] p_Val2_1_fu_539_p3;
wire [3:0] p_Val2_3_fu_347_p3;
wire [1:0] p_Val2_6_fu_566_p3;
wire [3:0] p_Val2_8_fu_845_p3;
wire [3:0] r_V_fu_840_p2;
wire [7:0] ret_V_15_fu_746_p3;
wire [17:0] ret_V_18_fu_784_p3;
wire [31:0] ret_V_22_fu_1011_p3;
wire [31:0] ret_V_24_fu_1074_p3;
wire [35:0] rhs_2_fu_700_p3;
wire rhs_3_fu_289_p2;
wire [34:0] rhs_5_fu_888_p3;
wire [52:0] rhs_6_fu_948_p3;
wire [32:0] rhs_8_fu_1026_p3;
wire [1:0] rhs_fu_638_p1;
wire [2:0] rhs_fu_638_p3;
wire [2:0] select_ln1118_1_fu_808_p3;
wire [3:0] select_ln1118_fu_833_p3;
wire [31:0] select_ln1192_fu_1081_p3;
wire [31:0] select_ln353_fu_937_p3;
wire [3:0] select_ln384_1_fu_547_p3;
wire [1:0] select_ln384_fu_588_p3;
wire [15:0] select_ln850_1_fu_673_p3;
wire [17:0] select_ln850_2_fu_779_p3;
wire [15:0] select_ln850_3_fu_678_p3;
wire [31:0] select_ln850_4_fu_1006_p3;
wire [31:0] select_ln850_5_fu_1068_p3;
wire [31:0] select_ln850_6_fu_932_p3;
wire [7:0] select_ln850_fu_740_p3;
wire [1:0] sext_ln1195_fu_615_p0;
wire [8:0] sext_ln1195_fu_615_p1;
wire [31:0] sext_ln215_fu_267_p0;
wire [31:0] sext_ln703_3_fu_944_p0;
wire [1:0] sext_ln703_4_fu_1022_p0;
wire [31:0] sext_ln703_fu_456_p0;
wire [17:0] sext_ln850_fu_763_p1;
wire \sub_17ns_17ns_17_2_1_U2.ce ;
wire \sub_17ns_17ns_17_2_1_U2.clk ;
wire [16:0] \sub_17ns_17ns_17_2_1_U2.din0 ;
wire [16:0] \sub_17ns_17ns_17_2_1_U2.din1 ;
wire [16:0] \sub_17ns_17ns_17_2_1_U2.dout ;
wire \sub_17ns_17ns_17_2_1_U2.reset ;
wire [16:0] \sub_17ns_17ns_17_2_1_U2.top_sub_17ns_17ns_17_2_1_Adder_1_U.a ;
wire [16:0] \sub_17ns_17ns_17_2_1_U2.top_sub_17ns_17ns_17_2_1_Adder_1_U.ain_s0 ;
wire [16:0] \sub_17ns_17ns_17_2_1_U2.top_sub_17ns_17ns_17_2_1_Adder_1_U.b ;
wire [16:0] \sub_17ns_17ns_17_2_1_U2.top_sub_17ns_17ns_17_2_1_Adder_1_U.bin_s0 ;
wire \sub_17ns_17ns_17_2_1_U2.top_sub_17ns_17ns_17_2_1_Adder_1_U.ce ;
wire \sub_17ns_17ns_17_2_1_U2.top_sub_17ns_17ns_17_2_1_Adder_1_U.clk ;
wire \sub_17ns_17ns_17_2_1_U2.top_sub_17ns_17ns_17_2_1_Adder_1_U.facout_s1 ;
wire \sub_17ns_17ns_17_2_1_U2.top_sub_17ns_17ns_17_2_1_Adder_1_U.facout_s2 ;
wire [7:0] \sub_17ns_17ns_17_2_1_U2.top_sub_17ns_17ns_17_2_1_Adder_1_U.fas_s1 ;
wire [8:0] \sub_17ns_17ns_17_2_1_U2.top_sub_17ns_17ns_17_2_1_Adder_1_U.fas_s2 ;
wire \sub_17ns_17ns_17_2_1_U2.top_sub_17ns_17ns_17_2_1_Adder_1_U.reset ;
wire [16:0] \sub_17ns_17ns_17_2_1_U2.top_sub_17ns_17ns_17_2_1_Adder_1_U.s ;
wire [7:0] \sub_17ns_17ns_17_2_1_U2.top_sub_17ns_17ns_17_2_1_Adder_1_U.u1.a ;
wire [7:0] \sub_17ns_17ns_17_2_1_U2.top_sub_17ns_17ns_17_2_1_Adder_1_U.u1.b ;
wire \sub_17ns_17ns_17_2_1_U2.top_sub_17ns_17ns_17_2_1_Adder_1_U.u1.cin ;
wire \sub_17ns_17ns_17_2_1_U2.top_sub_17ns_17ns_17_2_1_Adder_1_U.u1.cout ;
wire [7:0] \sub_17ns_17ns_17_2_1_U2.top_sub_17ns_17ns_17_2_1_Adder_1_U.u1.s ;
wire [8:0] \sub_17ns_17ns_17_2_1_U2.top_sub_17ns_17ns_17_2_1_Adder_1_U.u2.a ;
wire [8:0] \sub_17ns_17ns_17_2_1_U2.top_sub_17ns_17ns_17_2_1_Adder_1_U.u2.b ;
wire \sub_17ns_17ns_17_2_1_U2.top_sub_17ns_17ns_17_2_1_Adder_1_U.u2.cin ;
wire \sub_17ns_17ns_17_2_1_U2.top_sub_17ns_17ns_17_2_1_Adder_1_U.u2.cout ;
wire [8:0] \sub_17ns_17ns_17_2_1_U2.top_sub_17ns_17ns_17_2_1_Adder_1_U.u2.s ;
wire \sub_33s_33ns_33_2_1_U1.ce ;
wire \sub_33s_33ns_33_2_1_U1.clk ;
wire [32:0] \sub_33s_33ns_33_2_1_U1.din0 ;
wire [32:0] \sub_33s_33ns_33_2_1_U1.din1 ;
wire [32:0] \sub_33s_33ns_33_2_1_U1.dout ;
wire \sub_33s_33ns_33_2_1_U1.reset ;
wire [32:0] \sub_33s_33ns_33_2_1_U1.top_sub_33s_33ns_33_2_1_Adder_0_U.a ;
wire [32:0] \sub_33s_33ns_33_2_1_U1.top_sub_33s_33ns_33_2_1_Adder_0_U.ain_s0 ;
wire [32:0] \sub_33s_33ns_33_2_1_U1.top_sub_33s_33ns_33_2_1_Adder_0_U.b ;
wire [32:0] \sub_33s_33ns_33_2_1_U1.top_sub_33s_33ns_33_2_1_Adder_0_U.bin_s0 ;
wire \sub_33s_33ns_33_2_1_U1.top_sub_33s_33ns_33_2_1_Adder_0_U.ce ;
wire \sub_33s_33ns_33_2_1_U1.top_sub_33s_33ns_33_2_1_Adder_0_U.clk ;
wire \sub_33s_33ns_33_2_1_U1.top_sub_33s_33ns_33_2_1_Adder_0_U.facout_s1 ;
wire \sub_33s_33ns_33_2_1_U1.top_sub_33s_33ns_33_2_1_Adder_0_U.facout_s2 ;
wire [15:0] \sub_33s_33ns_33_2_1_U1.top_sub_33s_33ns_33_2_1_Adder_0_U.fas_s1 ;
wire [16:0] \sub_33s_33ns_33_2_1_U1.top_sub_33s_33ns_33_2_1_Adder_0_U.fas_s2 ;
wire \sub_33s_33ns_33_2_1_U1.top_sub_33s_33ns_33_2_1_Adder_0_U.reset ;
wire [32:0] \sub_33s_33ns_33_2_1_U1.top_sub_33s_33ns_33_2_1_Adder_0_U.s ;
wire [15:0] \sub_33s_33ns_33_2_1_U1.top_sub_33s_33ns_33_2_1_Adder_0_U.u1.a ;
wire [15:0] \sub_33s_33ns_33_2_1_U1.top_sub_33s_33ns_33_2_1_Adder_0_U.u1.b ;
wire \sub_33s_33ns_33_2_1_U1.top_sub_33s_33ns_33_2_1_Adder_0_U.u1.cin ;
wire \sub_33s_33ns_33_2_1_U1.top_sub_33s_33ns_33_2_1_Adder_0_U.u1.cout ;
wire [15:0] \sub_33s_33ns_33_2_1_U1.top_sub_33s_33ns_33_2_1_Adder_0_U.u1.s ;
wire [16:0] \sub_33s_33ns_33_2_1_U1.top_sub_33s_33ns_33_2_1_Adder_0_U.u2.a ;
wire [16:0] \sub_33s_33ns_33_2_1_U1.top_sub_33s_33ns_33_2_1_Adder_0_U.u2.b ;
wire \sub_33s_33ns_33_2_1_U1.top_sub_33s_33ns_33_2_1_Adder_0_U.u2.cin ;
wire \sub_33s_33ns_33_2_1_U1.top_sub_33s_33ns_33_2_1_Adder_0_U.u2.cout ;
wire [16:0] \sub_33s_33ns_33_2_1_U1.top_sub_33s_33ns_33_2_1_Adder_0_U.u2.s ;
wire [31:0] tmp_3_fu_295_p1;
wire [1:0] tmp_3_fu_295_p4;
wire tmp_fu_859_p3;
wire [7:0] trunc_ln728_fu_281_p1;
wire [31:0] trunc_ln731_1_fu_344_p0;
wire [1:0] trunc_ln731_1_fu_344_p1;
wire [2:0] trunc_ln731_3_fu_815_p1;
wire [1:0] trunc_ln731_fu_536_p1;
wire trunc_ln790_fu_337_p1;
wire [31:0] trunc_ln851_1_fu_466_p0;
wire [16:0] trunc_ln851_1_fu_466_p1;
wire [1:0] trunc_ln851_2_fu_685_p1;
wire [2:0] trunc_ln851_3_fu_881_p1;
wire [31:0] trunc_ln851_4_fu_965_p0;
wire [20:0] trunc_ln851_4_fu_965_p1;
wire [1:0] trunc_ln851_5_fu_1065_p0;
wire trunc_ln851_5_fu_1065_p1;
wire trunc_ln851_fu_737_p1;
wire underflow_1_fu_583_p2;
wire underflow_fu_501_p2;
wire xor_ln785_1_fu_525_p2;
wire xor_ln785_fu_420_p2;
wire xor_ln786_1_fu_573_p2;
wire xor_ln786_fu_486_p2;
wire [15:0] zext_ln870_fu_285_p1;


assign _065_ = icmp_ln851_2_reg_1439 & ap_CS_fsm[22];
assign _066_ = icmp_ln851_3_reg_1476 & ap_CS_fsm[27];
assign _067_ = icmp_ln851_1_reg_1341 & ap_CS_fsm[11];
assign _068_ = ap_CS_fsm[6] & _071_;
assign _069_ = _072_ & ap_CS_fsm[0];
assign _070_ = ap_start & ap_CS_fsm[0];
assign and_ln731_fu_818_p2 = op_8_V_reg_1165[2:0] & select_ln1118_1_fu_808_p3;
assign overflow_2_fu_530_p2 = xor_ln785_1_fu_525_p2 & or_ln785_2_fu_521_p2;
assign overflow_fu_425_p2 = xor_ln785_fu_420_p2 & or_ln785_fu_416_p2;
assign r_V_fu_840_p2 = select_ln1118_fu_833_p3 & op_8_V_reg_1165;
assign underflow_1_fu_583_p2 = p_Result_17_reg_1186 & or_ln786_fu_578_p2;
assign underflow_fu_501_p2 = p_Result_14_reg_1137 & or_ln788_1_fu_496_p2;
assign xor_ln786_1_fu_573_p2 = ~ p_Result_18_reg_1192;
assign xor_ln786_fu_486_p2 = ~ p_Result_15_reg_1143;
assign xor_ln785_1_fu_525_p2 = ~ p_Result_17_reg_1186;
assign xor_ln785_fu_420_p2 = ~ p_Result_14_reg_1137;
assign _071_ = ~ icmp_ln851_reg_1226;
assign _072_ = ~ ap_start;
assign _073_ = ! { trunc_ln790_reg_1155, 2'h0 };
assign _074_ = ! op_7[16:0];
assign _075_ = op_1[3:0] == op_2;
always @(posedge \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_3_U.clk )
\add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_3_U.bin_s1  <= _077_;
always @(posedge \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_3_U.clk )
\add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_3_U.ain_s1  <= _076_;
always @(posedge \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_3_U.clk )
\add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_3_U.sum_s1  <= _079_;
always @(posedge \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_3_U.clk )
\add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_3_U.carry_s1  <= _078_;
assign _077_ = \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_3_U.ce  ? \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_3_U.b [15:8] : \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_3_U.bin_s1 ;
assign _076_ = \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_3_U.ce  ? \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_3_U.a [15:8] : \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_3_U.ain_s1 ;
assign _078_ = \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_3_U.ce  ? \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_3_U.facout_s1  : \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_3_U.carry_s1 ;
assign _079_ = \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_3_U.ce  ? \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_3_U.fas_s1  : \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_3_U.sum_s1 ;
assign _080_ = \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_3_U.u1.a  + \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_3_U.u1.b ;
assign { \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_3_U.u1.cout , \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_3_U.u1.s  } = _080_ + \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_3_U.u1.cin ;
assign _081_ = \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_3_U.u2.a  + \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_3_U.u2.b ;
assign { \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_3_U.u2.cout , \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_3_U.u2.s  } = _081_ + \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_3_U.u2.cin ;
always @(posedge \add_18ns_18s_18_2_1_U10.top_add_18ns_18s_18_2_1_Adder_8_U.clk )
\add_18ns_18s_18_2_1_U10.top_add_18ns_18s_18_2_1_Adder_8_U.bin_s1  <= _083_;
always @(posedge \add_18ns_18s_18_2_1_U10.top_add_18ns_18s_18_2_1_Adder_8_U.clk )
\add_18ns_18s_18_2_1_U10.top_add_18ns_18s_18_2_1_Adder_8_U.ain_s1  <= _082_;
always @(posedge \add_18ns_18s_18_2_1_U10.top_add_18ns_18s_18_2_1_Adder_8_U.clk )
\add_18ns_18s_18_2_1_U10.top_add_18ns_18s_18_2_1_Adder_8_U.sum_s1  <= _085_;
always @(posedge \add_18ns_18s_18_2_1_U10.top_add_18ns_18s_18_2_1_Adder_8_U.clk )
\add_18ns_18s_18_2_1_U10.top_add_18ns_18s_18_2_1_Adder_8_U.carry_s1  <= _084_;
assign _083_ = \add_18ns_18s_18_2_1_U10.top_add_18ns_18s_18_2_1_Adder_8_U.ce  ? \add_18ns_18s_18_2_1_U10.top_add_18ns_18s_18_2_1_Adder_8_U.b [17:9] : \add_18ns_18s_18_2_1_U10.top_add_18ns_18s_18_2_1_Adder_8_U.bin_s1 ;
assign _082_ = \add_18ns_18s_18_2_1_U10.top_add_18ns_18s_18_2_1_Adder_8_U.ce  ? \add_18ns_18s_18_2_1_U10.top_add_18ns_18s_18_2_1_Adder_8_U.a [17:9] : \add_18ns_18s_18_2_1_U10.top_add_18ns_18s_18_2_1_Adder_8_U.ain_s1 ;
assign _084_ = \add_18ns_18s_18_2_1_U10.top_add_18ns_18s_18_2_1_Adder_8_U.ce  ? \add_18ns_18s_18_2_1_U10.top_add_18ns_18s_18_2_1_Adder_8_U.facout_s1  : \add_18ns_18s_18_2_1_U10.top_add_18ns_18s_18_2_1_Adder_8_U.carry_s1 ;
assign _085_ = \add_18ns_18s_18_2_1_U10.top_add_18ns_18s_18_2_1_Adder_8_U.ce  ? \add_18ns_18s_18_2_1_U10.top_add_18ns_18s_18_2_1_Adder_8_U.fas_s1  : \add_18ns_18s_18_2_1_U10.top_add_18ns_18s_18_2_1_Adder_8_U.sum_s1 ;
assign _086_ = \add_18ns_18s_18_2_1_U10.top_add_18ns_18s_18_2_1_Adder_8_U.u1.a  + \add_18ns_18s_18_2_1_U10.top_add_18ns_18s_18_2_1_Adder_8_U.u1.b ;
assign { \add_18ns_18s_18_2_1_U10.top_add_18ns_18s_18_2_1_Adder_8_U.u1.cout , \add_18ns_18s_18_2_1_U10.top_add_18ns_18s_18_2_1_Adder_8_U.u1.s  } = _086_ + \add_18ns_18s_18_2_1_U10.top_add_18ns_18s_18_2_1_Adder_8_U.u1.cin ;
assign _087_ = \add_18ns_18s_18_2_1_U10.top_add_18ns_18s_18_2_1_Adder_8_U.u2.a  + \add_18ns_18s_18_2_1_U10.top_add_18ns_18s_18_2_1_Adder_8_U.u2.b ;
assign { \add_18ns_18s_18_2_1_U10.top_add_18ns_18s_18_2_1_Adder_8_U.u2.cout , \add_18ns_18s_18_2_1_U10.top_add_18ns_18s_18_2_1_Adder_8_U.u2.s  } = _087_ + \add_18ns_18s_18_2_1_U10.top_add_18ns_18s_18_2_1_Adder_8_U.u2.cin ;
always @(posedge \add_18ns_18s_18_2_1_U9.top_add_18ns_18s_18_2_1_Adder_8_U.clk )
\add_18ns_18s_18_2_1_U9.top_add_18ns_18s_18_2_1_Adder_8_U.bin_s1  <= _089_;
always @(posedge \add_18ns_18s_18_2_1_U9.top_add_18ns_18s_18_2_1_Adder_8_U.clk )
\add_18ns_18s_18_2_1_U9.top_add_18ns_18s_18_2_1_Adder_8_U.ain_s1  <= _088_;
always @(posedge \add_18ns_18s_18_2_1_U9.top_add_18ns_18s_18_2_1_Adder_8_U.clk )
\add_18ns_18s_18_2_1_U9.top_add_18ns_18s_18_2_1_Adder_8_U.sum_s1  <= _091_;
always @(posedge \add_18ns_18s_18_2_1_U9.top_add_18ns_18s_18_2_1_Adder_8_U.clk )
\add_18ns_18s_18_2_1_U9.top_add_18ns_18s_18_2_1_Adder_8_U.carry_s1  <= _090_;
assign _089_ = \add_18ns_18s_18_2_1_U9.top_add_18ns_18s_18_2_1_Adder_8_U.ce  ? \add_18ns_18s_18_2_1_U9.top_add_18ns_18s_18_2_1_Adder_8_U.b [17:9] : \add_18ns_18s_18_2_1_U9.top_add_18ns_18s_18_2_1_Adder_8_U.bin_s1 ;
assign _088_ = \add_18ns_18s_18_2_1_U9.top_add_18ns_18s_18_2_1_Adder_8_U.ce  ? \add_18ns_18s_18_2_1_U9.top_add_18ns_18s_18_2_1_Adder_8_U.a [17:9] : \add_18ns_18s_18_2_1_U9.top_add_18ns_18s_18_2_1_Adder_8_U.ain_s1 ;
assign _090_ = \add_18ns_18s_18_2_1_U9.top_add_18ns_18s_18_2_1_Adder_8_U.ce  ? \add_18ns_18s_18_2_1_U9.top_add_18ns_18s_18_2_1_Adder_8_U.facout_s1  : \add_18ns_18s_18_2_1_U9.top_add_18ns_18s_18_2_1_Adder_8_U.carry_s1 ;
assign _091_ = \add_18ns_18s_18_2_1_U9.top_add_18ns_18s_18_2_1_Adder_8_U.ce  ? \add_18ns_18s_18_2_1_U9.top_add_18ns_18s_18_2_1_Adder_8_U.fas_s1  : \add_18ns_18s_18_2_1_U9.top_add_18ns_18s_18_2_1_Adder_8_U.sum_s1 ;
assign _092_ = \add_18ns_18s_18_2_1_U9.top_add_18ns_18s_18_2_1_Adder_8_U.u1.a  + \add_18ns_18s_18_2_1_U9.top_add_18ns_18s_18_2_1_Adder_8_U.u1.b ;
assign { \add_18ns_18s_18_2_1_U9.top_add_18ns_18s_18_2_1_Adder_8_U.u1.cout , \add_18ns_18s_18_2_1_U9.top_add_18ns_18s_18_2_1_Adder_8_U.u1.s  } = _092_ + \add_18ns_18s_18_2_1_U9.top_add_18ns_18s_18_2_1_Adder_8_U.u1.cin ;
assign _093_ = \add_18ns_18s_18_2_1_U9.top_add_18ns_18s_18_2_1_Adder_8_U.u2.a  + \add_18ns_18s_18_2_1_U9.top_add_18ns_18s_18_2_1_Adder_8_U.u2.b ;
assign { \add_18ns_18s_18_2_1_U9.top_add_18ns_18s_18_2_1_Adder_8_U.u2.cout , \add_18ns_18s_18_2_1_U9.top_add_18ns_18s_18_2_1_Adder_8_U.u2.s  } = _093_ + \add_18ns_18s_18_2_1_U9.top_add_18ns_18s_18_2_1_Adder_8_U.u2.cin ;
always @(posedge \add_18s_18ns_18_2_1_U8.top_add_18s_18ns_18_2_1_Adder_7_U.clk )
\add_18s_18ns_18_2_1_U8.top_add_18s_18ns_18_2_1_Adder_7_U.bin_s1  <= _095_;
always @(posedge \add_18s_18ns_18_2_1_U8.top_add_18s_18ns_18_2_1_Adder_7_U.clk )
\add_18s_18ns_18_2_1_U8.top_add_18s_18ns_18_2_1_Adder_7_U.ain_s1  <= _094_;
always @(posedge \add_18s_18ns_18_2_1_U8.top_add_18s_18ns_18_2_1_Adder_7_U.clk )
\add_18s_18ns_18_2_1_U8.top_add_18s_18ns_18_2_1_Adder_7_U.sum_s1  <= _097_;
always @(posedge \add_18s_18ns_18_2_1_U8.top_add_18s_18ns_18_2_1_Adder_7_U.clk )
\add_18s_18ns_18_2_1_U8.top_add_18s_18ns_18_2_1_Adder_7_U.carry_s1  <= _096_;
assign _095_ = \add_18s_18ns_18_2_1_U8.top_add_18s_18ns_18_2_1_Adder_7_U.ce  ? \add_18s_18ns_18_2_1_U8.top_add_18s_18ns_18_2_1_Adder_7_U.b [17:9] : \add_18s_18ns_18_2_1_U8.top_add_18s_18ns_18_2_1_Adder_7_U.bin_s1 ;
assign _094_ = \add_18s_18ns_18_2_1_U8.top_add_18s_18ns_18_2_1_Adder_7_U.ce  ? \add_18s_18ns_18_2_1_U8.top_add_18s_18ns_18_2_1_Adder_7_U.a [17:9] : \add_18s_18ns_18_2_1_U8.top_add_18s_18ns_18_2_1_Adder_7_U.ain_s1 ;
assign _096_ = \add_18s_18ns_18_2_1_U8.top_add_18s_18ns_18_2_1_Adder_7_U.ce  ? \add_18s_18ns_18_2_1_U8.top_add_18s_18ns_18_2_1_Adder_7_U.facout_s1  : \add_18s_18ns_18_2_1_U8.top_add_18s_18ns_18_2_1_Adder_7_U.carry_s1 ;
assign _097_ = \add_18s_18ns_18_2_1_U8.top_add_18s_18ns_18_2_1_Adder_7_U.ce  ? \add_18s_18ns_18_2_1_U8.top_add_18s_18ns_18_2_1_Adder_7_U.fas_s1  : \add_18s_18ns_18_2_1_U8.top_add_18s_18ns_18_2_1_Adder_7_U.sum_s1 ;
assign _098_ = \add_18s_18ns_18_2_1_U8.top_add_18s_18ns_18_2_1_Adder_7_U.u1.a  + \add_18s_18ns_18_2_1_U8.top_add_18s_18ns_18_2_1_Adder_7_U.u1.b ;
assign { \add_18s_18ns_18_2_1_U8.top_add_18s_18ns_18_2_1_Adder_7_U.u1.cout , \add_18s_18ns_18_2_1_U8.top_add_18s_18ns_18_2_1_Adder_7_U.u1.s  } = _098_ + \add_18s_18ns_18_2_1_U8.top_add_18s_18ns_18_2_1_Adder_7_U.u1.cin ;
assign _099_ = \add_18s_18ns_18_2_1_U8.top_add_18s_18ns_18_2_1_Adder_7_U.u2.a  + \add_18s_18ns_18_2_1_U8.top_add_18s_18ns_18_2_1_Adder_7_U.u2.b ;
assign { \add_18s_18ns_18_2_1_U8.top_add_18s_18ns_18_2_1_Adder_7_U.u2.cout , \add_18s_18ns_18_2_1_U8.top_add_18s_18ns_18_2_1_Adder_7_U.u2.s  } = _099_ + \add_18s_18ns_18_2_1_U8.top_add_18s_18ns_18_2_1_Adder_7_U.u2.cin ;
always @(posedge \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_11_U.clk )
\add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_11_U.bin_s1  <= _101_;
always @(posedge \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_11_U.clk )
\add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_11_U.ain_s1  <= _100_;
always @(posedge \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_11_U.clk )
\add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_11_U.sum_s1  <= _103_;
always @(posedge \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_11_U.clk )
\add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_11_U.carry_s1  <= _102_;
assign _101_ = \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_11_U.ce  ? \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_11_U.b [31:16] : \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_11_U.bin_s1 ;
assign _100_ = \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_11_U.ce  ? \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_11_U.a [31:16] : \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_11_U.ain_s1 ;
assign _102_ = \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_11_U.ce  ? \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_11_U.facout_s1  : \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_11_U.carry_s1 ;
assign _103_ = \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_11_U.ce  ? \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_11_U.fas_s1  : \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_11_U.sum_s1 ;
assign _104_ = \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.a  + \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.b ;
assign { \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.cout , \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.s  } = _104_ + \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.cin ;
assign _105_ = \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.a  + \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.b ;
assign { \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.cout , \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.s  } = _105_ + \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.cin ;
always @(posedge \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.clk )
\add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.bin_s1  <= _107_;
always @(posedge \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.clk )
\add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.ain_s1  <= _106_;
always @(posedge \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.clk )
\add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.sum_s1  <= _109_;
always @(posedge \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.clk )
\add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.carry_s1  <= _108_;
assign _107_ = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.ce  ? \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.b [31:16] : \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.bin_s1 ;
assign _106_ = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.ce  ? \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.a [31:16] : \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.ain_s1 ;
assign _108_ = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.ce  ? \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.facout_s1  : \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.carry_s1 ;
assign _109_ = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.ce  ? \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.fas_s1  : \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.sum_s1 ;
assign _110_ = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.a  + \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.b ;
assign { \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.cout , \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.s  } = _110_ + \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.cin ;
assign _111_ = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.a  + \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.b ;
assign { \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.cout , \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.s  } = _111_ + \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.cin ;
always @(posedge \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.clk )
\add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.bin_s1  <= _113_;
always @(posedge \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.clk )
\add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.ain_s1  <= _112_;
always @(posedge \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.clk )
\add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.sum_s1  <= _115_;
always @(posedge \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.clk )
\add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.carry_s1  <= _114_;
assign _113_ = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.ce  ? \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.b [31:16] : \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.bin_s1 ;
assign _112_ = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.ce  ? \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.a [31:16] : \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.ain_s1 ;
assign _114_ = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.ce  ? \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.facout_s1  : \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.carry_s1 ;
assign _115_ = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.ce  ? \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.fas_s1  : \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.sum_s1 ;
assign _116_ = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.a  + \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.b ;
assign { \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.cout , \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.s  } = _116_ + \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.cin ;
assign _117_ = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.a  + \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.b ;
assign { \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.cout , \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.s  } = _117_ + \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.cin ;
always @(posedge \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.clk )
\add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.bin_s1  <= _119_;
always @(posedge \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.clk )
\add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.ain_s1  <= _118_;
always @(posedge \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.clk )
\add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.sum_s1  <= _121_;
always @(posedge \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.clk )
\add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.carry_s1  <= _120_;
assign _119_ = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.ce  ? \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.b [31:16] : \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.bin_s1 ;
assign _118_ = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.ce  ? \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.a [31:16] : \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.ain_s1 ;
assign _120_ = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.ce  ? \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.facout_s1  : \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.carry_s1 ;
assign _121_ = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.ce  ? \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.fas_s1  : \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.sum_s1 ;
assign _122_ = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.a  + \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.b ;
assign { \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.cout , \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.s  } = _122_ + \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.cin ;
assign _123_ = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.a  + \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.b ;
assign { \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.cout , \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.s  } = _123_ + \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.cin ;
always @(posedge \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.clk )
\add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.bin_s1  <= _125_;
always @(posedge \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.clk )
\add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.ain_s1  <= _124_;
always @(posedge \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.clk )
\add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.sum_s1  <= _127_;
always @(posedge \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.clk )
\add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.carry_s1  <= _126_;
assign _125_ = \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.ce  ? \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.b [31:16] : \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.bin_s1 ;
assign _124_ = \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.ce  ? \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.a [31:16] : \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.ain_s1 ;
assign _126_ = \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.ce  ? \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.facout_s1  : \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.carry_s1 ;
assign _127_ = \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.ce  ? \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.fas_s1  : \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.sum_s1 ;
assign _128_ = \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.a  + \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.b ;
assign { \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.cout , \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.s  } = _128_ + \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.cin ;
assign _129_ = \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.a  + \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.b ;
assign { \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.cout , \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.s  } = _129_ + \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.cin ;
always @(posedge \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.clk )
\add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.bin_s1  <= _131_;
always @(posedge \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.clk )
\add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.ain_s1  <= _130_;
always @(posedge \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.clk )
\add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.sum_s1  <= _133_;
always @(posedge \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.clk )
\add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.carry_s1  <= _132_;
assign _131_ = \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.ce  ? \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.b [31:16] : \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.bin_s1 ;
assign _130_ = \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.ce  ? \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.a [31:16] : \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.ain_s1 ;
assign _132_ = \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.ce  ? \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.facout_s1  : \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.carry_s1 ;
assign _133_ = \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.ce  ? \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.fas_s1  : \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.sum_s1 ;
assign _134_ = \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.a  + \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.b ;
assign { \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.cout , \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.s  } = _134_ + \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.cin ;
assign _135_ = \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.a  + \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.b ;
assign { \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.cout , \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.s  } = _135_ + \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.cin ;
always @(posedge \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_9_U.clk )
\add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_9_U.bin_s1  <= _137_;
always @(posedge \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_9_U.clk )
\add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_9_U.ain_s1  <= _136_;
always @(posedge \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_9_U.clk )
\add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_9_U.sum_s1  <= _139_;
always @(posedge \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_9_U.clk )
\add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_9_U.carry_s1  <= _138_;
assign _137_ = \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_9_U.ce  ? \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_9_U.b [31:16] : \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_9_U.bin_s1 ;
assign _136_ = \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_9_U.ce  ? \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_9_U.a [31:16] : \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_9_U.ain_s1 ;
assign _138_ = \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_9_U.ce  ? \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_9_U.facout_s1  : \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_9_U.carry_s1 ;
assign _139_ = \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_9_U.ce  ? \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_9_U.fas_s1  : \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_9_U.sum_s1 ;
assign _140_ = \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_9_U.u1.a  + \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_9_U.u1.b ;
assign { \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_9_U.u1.cout , \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_9_U.u1.s  } = _140_ + \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_9_U.u1.cin ;
assign _141_ = \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_9_U.u2.a  + \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_9_U.u2.b ;
assign { \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_9_U.u2.cout , \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_9_U.u2.s  } = _141_ + \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_9_U.u2.cin ;
always @(posedge \add_33ns_33s_33_2_1_U3.top_add_33ns_33s_33_2_1_Adder_2_U.clk )
\add_33ns_33s_33_2_1_U3.top_add_33ns_33s_33_2_1_Adder_2_U.bin_s1  <= _143_;
always @(posedge \add_33ns_33s_33_2_1_U3.top_add_33ns_33s_33_2_1_Adder_2_U.clk )
\add_33ns_33s_33_2_1_U3.top_add_33ns_33s_33_2_1_Adder_2_U.ain_s1  <= _142_;
always @(posedge \add_33ns_33s_33_2_1_U3.top_add_33ns_33s_33_2_1_Adder_2_U.clk )
\add_33ns_33s_33_2_1_U3.top_add_33ns_33s_33_2_1_Adder_2_U.sum_s1  <= _145_;
always @(posedge \add_33ns_33s_33_2_1_U3.top_add_33ns_33s_33_2_1_Adder_2_U.clk )
\add_33ns_33s_33_2_1_U3.top_add_33ns_33s_33_2_1_Adder_2_U.carry_s1  <= _144_;
assign _143_ = \add_33ns_33s_33_2_1_U3.top_add_33ns_33s_33_2_1_Adder_2_U.ce  ? \add_33ns_33s_33_2_1_U3.top_add_33ns_33s_33_2_1_Adder_2_U.b [32:16] : \add_33ns_33s_33_2_1_U3.top_add_33ns_33s_33_2_1_Adder_2_U.bin_s1 ;
assign _142_ = \add_33ns_33s_33_2_1_U3.top_add_33ns_33s_33_2_1_Adder_2_U.ce  ? \add_33ns_33s_33_2_1_U3.top_add_33ns_33s_33_2_1_Adder_2_U.a [32:16] : \add_33ns_33s_33_2_1_U3.top_add_33ns_33s_33_2_1_Adder_2_U.ain_s1 ;
assign _144_ = \add_33ns_33s_33_2_1_U3.top_add_33ns_33s_33_2_1_Adder_2_U.ce  ? \add_33ns_33s_33_2_1_U3.top_add_33ns_33s_33_2_1_Adder_2_U.facout_s1  : \add_33ns_33s_33_2_1_U3.top_add_33ns_33s_33_2_1_Adder_2_U.carry_s1 ;
assign _145_ = \add_33ns_33s_33_2_1_U3.top_add_33ns_33s_33_2_1_Adder_2_U.ce  ? \add_33ns_33s_33_2_1_U3.top_add_33ns_33s_33_2_1_Adder_2_U.fas_s1  : \add_33ns_33s_33_2_1_U3.top_add_33ns_33s_33_2_1_Adder_2_U.sum_s1 ;
assign _146_ = \add_33ns_33s_33_2_1_U3.top_add_33ns_33s_33_2_1_Adder_2_U.u1.a  + \add_33ns_33s_33_2_1_U3.top_add_33ns_33s_33_2_1_Adder_2_U.u1.b ;
assign { \add_33ns_33s_33_2_1_U3.top_add_33ns_33s_33_2_1_Adder_2_U.u1.cout , \add_33ns_33s_33_2_1_U3.top_add_33ns_33s_33_2_1_Adder_2_U.u1.s  } = _146_ + \add_33ns_33s_33_2_1_U3.top_add_33ns_33s_33_2_1_Adder_2_U.u1.cin ;
assign _147_ = \add_33ns_33s_33_2_1_U3.top_add_33ns_33s_33_2_1_Adder_2_U.u2.a  + \add_33ns_33s_33_2_1_U3.top_add_33ns_33s_33_2_1_Adder_2_U.u2.b ;
assign { \add_33ns_33s_33_2_1_U3.top_add_33ns_33s_33_2_1_Adder_2_U.u2.cout , \add_33ns_33s_33_2_1_U3.top_add_33ns_33s_33_2_1_Adder_2_U.u2.s  } = _147_ + \add_33ns_33s_33_2_1_U3.top_add_33ns_33s_33_2_1_Adder_2_U.u2.cin ;
always @(posedge \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_13_U.clk )
\add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_13_U.bin_s1  <= _149_;
always @(posedge \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_13_U.clk )
\add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_13_U.ain_s1  <= _148_;
always @(posedge \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_13_U.clk )
\add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_13_U.sum_s1  <= _151_;
always @(posedge \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_13_U.clk )
\add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_13_U.carry_s1  <= _150_;
assign _149_ = \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_13_U.ce  ? \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_13_U.b [33:17] : \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_13_U.bin_s1 ;
assign _148_ = \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_13_U.ce  ? \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_13_U.a [33:17] : \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_13_U.ain_s1 ;
assign _150_ = \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_13_U.ce  ? \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_13_U.facout_s1  : \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_13_U.carry_s1 ;
assign _151_ = \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_13_U.ce  ? \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_13_U.fas_s1  : \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_13_U.sum_s1 ;
assign _152_ = \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_13_U.u1.a  + \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_13_U.u1.b ;
assign { \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_13_U.u1.cout , \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_13_U.u1.s  } = _152_ + \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_13_U.u1.cin ;
assign _153_ = \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_13_U.u2.a  + \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_13_U.u2.b ;
assign { \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_13_U.u2.cout , \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_13_U.u2.s  } = _153_ + \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_13_U.u2.cin ;
always @(posedge \add_36s_36s_36_2_1_U12.top_add_36s_36s_36_2_1_Adder_10_U.clk )
\add_36s_36s_36_2_1_U12.top_add_36s_36s_36_2_1_Adder_10_U.bin_s1  <= _155_;
always @(posedge \add_36s_36s_36_2_1_U12.top_add_36s_36s_36_2_1_Adder_10_U.clk )
\add_36s_36s_36_2_1_U12.top_add_36s_36s_36_2_1_Adder_10_U.ain_s1  <= _154_;
always @(posedge \add_36s_36s_36_2_1_U12.top_add_36s_36s_36_2_1_Adder_10_U.clk )
\add_36s_36s_36_2_1_U12.top_add_36s_36s_36_2_1_Adder_10_U.sum_s1  <= _157_;
always @(posedge \add_36s_36s_36_2_1_U12.top_add_36s_36s_36_2_1_Adder_10_U.clk )
\add_36s_36s_36_2_1_U12.top_add_36s_36s_36_2_1_Adder_10_U.carry_s1  <= _156_;
assign _155_ = \add_36s_36s_36_2_1_U12.top_add_36s_36s_36_2_1_Adder_10_U.ce  ? \add_36s_36s_36_2_1_U12.top_add_36s_36s_36_2_1_Adder_10_U.b [35:18] : \add_36s_36s_36_2_1_U12.top_add_36s_36s_36_2_1_Adder_10_U.bin_s1 ;
assign _154_ = \add_36s_36s_36_2_1_U12.top_add_36s_36s_36_2_1_Adder_10_U.ce  ? \add_36s_36s_36_2_1_U12.top_add_36s_36s_36_2_1_Adder_10_U.a [35:18] : \add_36s_36s_36_2_1_U12.top_add_36s_36s_36_2_1_Adder_10_U.ain_s1 ;
assign _156_ = \add_36s_36s_36_2_1_U12.top_add_36s_36s_36_2_1_Adder_10_U.ce  ? \add_36s_36s_36_2_1_U12.top_add_36s_36s_36_2_1_Adder_10_U.facout_s1  : \add_36s_36s_36_2_1_U12.top_add_36s_36s_36_2_1_Adder_10_U.carry_s1 ;
assign _157_ = \add_36s_36s_36_2_1_U12.top_add_36s_36s_36_2_1_Adder_10_U.ce  ? \add_36s_36s_36_2_1_U12.top_add_36s_36s_36_2_1_Adder_10_U.fas_s1  : \add_36s_36s_36_2_1_U12.top_add_36s_36s_36_2_1_Adder_10_U.sum_s1 ;
assign _158_ = \add_36s_36s_36_2_1_U12.top_add_36s_36s_36_2_1_Adder_10_U.u1.a  + \add_36s_36s_36_2_1_U12.top_add_36s_36s_36_2_1_Adder_10_U.u1.b ;
assign { \add_36s_36s_36_2_1_U12.top_add_36s_36s_36_2_1_Adder_10_U.u1.cout , \add_36s_36s_36_2_1_U12.top_add_36s_36s_36_2_1_Adder_10_U.u1.s  } = _158_ + \add_36s_36s_36_2_1_U12.top_add_36s_36s_36_2_1_Adder_10_U.u1.cin ;
assign _159_ = \add_36s_36s_36_2_1_U12.top_add_36s_36s_36_2_1_Adder_10_U.u2.a  + \add_36s_36s_36_2_1_U12.top_add_36s_36s_36_2_1_Adder_10_U.u2.b ;
assign { \add_36s_36s_36_2_1_U12.top_add_36s_36s_36_2_1_Adder_10_U.u2.cout , \add_36s_36s_36_2_1_U12.top_add_36s_36s_36_2_1_Adder_10_U.u2.s  } = _159_ + \add_36s_36s_36_2_1_U12.top_add_36s_36s_36_2_1_Adder_10_U.u2.cin ;
always @(posedge \add_37s_37s_37_2_1_U7.top_add_37s_37s_37_2_1_Adder_6_U.clk )
\add_37s_37s_37_2_1_U7.top_add_37s_37s_37_2_1_Adder_6_U.bin_s1  <= _161_;
always @(posedge \add_37s_37s_37_2_1_U7.top_add_37s_37s_37_2_1_Adder_6_U.clk )
\add_37s_37s_37_2_1_U7.top_add_37s_37s_37_2_1_Adder_6_U.ain_s1  <= _160_;
always @(posedge \add_37s_37s_37_2_1_U7.top_add_37s_37s_37_2_1_Adder_6_U.clk )
\add_37s_37s_37_2_1_U7.top_add_37s_37s_37_2_1_Adder_6_U.sum_s1  <= _163_;
always @(posedge \add_37s_37s_37_2_1_U7.top_add_37s_37s_37_2_1_Adder_6_U.clk )
\add_37s_37s_37_2_1_U7.top_add_37s_37s_37_2_1_Adder_6_U.carry_s1  <= _162_;
assign _161_ = \add_37s_37s_37_2_1_U7.top_add_37s_37s_37_2_1_Adder_6_U.ce  ? \add_37s_37s_37_2_1_U7.top_add_37s_37s_37_2_1_Adder_6_U.b [36:18] : \add_37s_37s_37_2_1_U7.top_add_37s_37s_37_2_1_Adder_6_U.bin_s1 ;
assign _160_ = \add_37s_37s_37_2_1_U7.top_add_37s_37s_37_2_1_Adder_6_U.ce  ? \add_37s_37s_37_2_1_U7.top_add_37s_37s_37_2_1_Adder_6_U.a [36:18] : \add_37s_37s_37_2_1_U7.top_add_37s_37s_37_2_1_Adder_6_U.ain_s1 ;
assign _162_ = \add_37s_37s_37_2_1_U7.top_add_37s_37s_37_2_1_Adder_6_U.ce  ? \add_37s_37s_37_2_1_U7.top_add_37s_37s_37_2_1_Adder_6_U.facout_s1  : \add_37s_37s_37_2_1_U7.top_add_37s_37s_37_2_1_Adder_6_U.carry_s1 ;
assign _163_ = \add_37s_37s_37_2_1_U7.top_add_37s_37s_37_2_1_Adder_6_U.ce  ? \add_37s_37s_37_2_1_U7.top_add_37s_37s_37_2_1_Adder_6_U.fas_s1  : \add_37s_37s_37_2_1_U7.top_add_37s_37s_37_2_1_Adder_6_U.sum_s1 ;
assign _164_ = \add_37s_37s_37_2_1_U7.top_add_37s_37s_37_2_1_Adder_6_U.u1.a  + \add_37s_37s_37_2_1_U7.top_add_37s_37s_37_2_1_Adder_6_U.u1.b ;
assign { \add_37s_37s_37_2_1_U7.top_add_37s_37s_37_2_1_Adder_6_U.u1.cout , \add_37s_37s_37_2_1_U7.top_add_37s_37s_37_2_1_Adder_6_U.u1.s  } = _164_ + \add_37s_37s_37_2_1_U7.top_add_37s_37s_37_2_1_Adder_6_U.u1.cin ;
assign _165_ = \add_37s_37s_37_2_1_U7.top_add_37s_37s_37_2_1_Adder_6_U.u2.a  + \add_37s_37s_37_2_1_U7.top_add_37s_37s_37_2_1_Adder_6_U.u2.b ;
assign { \add_37s_37s_37_2_1_U7.top_add_37s_37s_37_2_1_Adder_6_U.u2.cout , \add_37s_37s_37_2_1_U7.top_add_37s_37s_37_2_1_Adder_6_U.u2.s  } = _165_ + \add_37s_37s_37_2_1_U7.top_add_37s_37s_37_2_1_Adder_6_U.u2.cin ;
always @(posedge \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_12_U.clk )
\add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_12_U.bin_s1  <= _167_;
always @(posedge \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_12_U.clk )
\add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_12_U.ain_s1  <= _166_;
always @(posedge \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_12_U.clk )
\add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_12_U.sum_s1  <= _169_;
always @(posedge \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_12_U.clk )
\add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_12_U.carry_s1  <= _168_;
assign _167_ = \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_12_U.ce  ? \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_12_U.b [53:27] : \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_12_U.bin_s1 ;
assign _166_ = \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_12_U.ce  ? \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_12_U.a [53:27] : \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_12_U.ain_s1 ;
assign _168_ = \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_12_U.ce  ? \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_12_U.facout_s1  : \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_12_U.carry_s1 ;
assign _169_ = \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_12_U.ce  ? \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_12_U.fas_s1  : \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_12_U.sum_s1 ;
assign _170_ = \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_12_U.u1.a  + \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_12_U.u1.b ;
assign { \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_12_U.u1.cout , \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_12_U.u1.s  } = _170_ + \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_12_U.u1.cin ;
assign _171_ = \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_12_U.u2.a  + \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_12_U.u2.b ;
assign { \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_12_U.u2.cout , \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_12_U.u2.s  } = _171_ + \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_12_U.u2.cin ;
always @(posedge \add_5s_5s_5_2_1_U5.top_add_5s_5s_5_2_1_Adder_4_U.clk )
\add_5s_5s_5_2_1_U5.top_add_5s_5s_5_2_1_Adder_4_U.bin_s1  <= _173_;
always @(posedge \add_5s_5s_5_2_1_U5.top_add_5s_5s_5_2_1_Adder_4_U.clk )
\add_5s_5s_5_2_1_U5.top_add_5s_5s_5_2_1_Adder_4_U.ain_s1  <= _172_;
always @(posedge \add_5s_5s_5_2_1_U5.top_add_5s_5s_5_2_1_Adder_4_U.clk )
\add_5s_5s_5_2_1_U5.top_add_5s_5s_5_2_1_Adder_4_U.sum_s1  <= _175_;
always @(posedge \add_5s_5s_5_2_1_U5.top_add_5s_5s_5_2_1_Adder_4_U.clk )
\add_5s_5s_5_2_1_U5.top_add_5s_5s_5_2_1_Adder_4_U.carry_s1  <= _174_;
assign _173_ = \add_5s_5s_5_2_1_U5.top_add_5s_5s_5_2_1_Adder_4_U.ce  ? \add_5s_5s_5_2_1_U5.top_add_5s_5s_5_2_1_Adder_4_U.b [4:2] : \add_5s_5s_5_2_1_U5.top_add_5s_5s_5_2_1_Adder_4_U.bin_s1 ;
assign _172_ = \add_5s_5s_5_2_1_U5.top_add_5s_5s_5_2_1_Adder_4_U.ce  ? \add_5s_5s_5_2_1_U5.top_add_5s_5s_5_2_1_Adder_4_U.a [4:2] : \add_5s_5s_5_2_1_U5.top_add_5s_5s_5_2_1_Adder_4_U.ain_s1 ;
assign _174_ = \add_5s_5s_5_2_1_U5.top_add_5s_5s_5_2_1_Adder_4_U.ce  ? \add_5s_5s_5_2_1_U5.top_add_5s_5s_5_2_1_Adder_4_U.facout_s1  : \add_5s_5s_5_2_1_U5.top_add_5s_5s_5_2_1_Adder_4_U.carry_s1 ;
assign _175_ = \add_5s_5s_5_2_1_U5.top_add_5s_5s_5_2_1_Adder_4_U.ce  ? \add_5s_5s_5_2_1_U5.top_add_5s_5s_5_2_1_Adder_4_U.fas_s1  : \add_5s_5s_5_2_1_U5.top_add_5s_5s_5_2_1_Adder_4_U.sum_s1 ;
assign _176_ = \add_5s_5s_5_2_1_U5.top_add_5s_5s_5_2_1_Adder_4_U.u1.a  + \add_5s_5s_5_2_1_U5.top_add_5s_5s_5_2_1_Adder_4_U.u1.b ;
assign { \add_5s_5s_5_2_1_U5.top_add_5s_5s_5_2_1_Adder_4_U.u1.cout , \add_5s_5s_5_2_1_U5.top_add_5s_5s_5_2_1_Adder_4_U.u1.s  } = _176_ + \add_5s_5s_5_2_1_U5.top_add_5s_5s_5_2_1_Adder_4_U.u1.cin ;
assign _177_ = \add_5s_5s_5_2_1_U5.top_add_5s_5s_5_2_1_Adder_4_U.u2.a  + \add_5s_5s_5_2_1_U5.top_add_5s_5s_5_2_1_Adder_4_U.u2.b ;
assign { \add_5s_5s_5_2_1_U5.top_add_5s_5s_5_2_1_Adder_4_U.u2.cout , \add_5s_5s_5_2_1_U5.top_add_5s_5s_5_2_1_Adder_4_U.u2.s  } = _177_ + \add_5s_5s_5_2_1_U5.top_add_5s_5s_5_2_1_Adder_4_U.u2.cin ;
always @(posedge \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.clk )
\add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.bin_s1  <= _179_;
always @(posedge \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.clk )
\add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.ain_s1  <= _178_;
always @(posedge \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.clk )
\add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.sum_s1  <= _181_;
always @(posedge \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.clk )
\add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.carry_s1  <= _180_;
assign _179_ = \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.ce  ? \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.b [7:4] : \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.bin_s1 ;
assign _178_ = \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.ce  ? \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.a [7:4] : \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.ain_s1 ;
assign _180_ = \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.ce  ? \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.facout_s1  : \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.carry_s1 ;
assign _181_ = \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.ce  ? \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.fas_s1  : \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.sum_s1 ;
assign _182_ = \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.u1.a  + \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.u1.b ;
assign { \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.u1.cout , \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.u1.s  } = _182_ + \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.u1.cin ;
assign _183_ = \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.u2.a  + \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.u2.b ;
assign { \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.u2.cout , \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.u2.s  } = _183_ + \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.u2.cin ;
assign \sub_17ns_17ns_17_2_1_U2.top_sub_17ns_17ns_17_2_1_Adder_1_U.bin_s0  = ~ \sub_17ns_17ns_17_2_1_U2.top_sub_17ns_17ns_17_2_1_Adder_1_U.b ;
always @(posedge \sub_17ns_17ns_17_2_1_U2.top_sub_17ns_17ns_17_2_1_Adder_1_U.clk )
\sub_17ns_17ns_17_2_1_U2.top_sub_17ns_17ns_17_2_1_Adder_1_U.bin_s1  <= _185_;
always @(posedge \sub_17ns_17ns_17_2_1_U2.top_sub_17ns_17ns_17_2_1_Adder_1_U.clk )
\sub_17ns_17ns_17_2_1_U2.top_sub_17ns_17ns_17_2_1_Adder_1_U.ain_s1  <= _184_;
always @(posedge \sub_17ns_17ns_17_2_1_U2.top_sub_17ns_17ns_17_2_1_Adder_1_U.clk )
\sub_17ns_17ns_17_2_1_U2.top_sub_17ns_17ns_17_2_1_Adder_1_U.sum_s1  <= _187_;
always @(posedge \sub_17ns_17ns_17_2_1_U2.top_sub_17ns_17ns_17_2_1_Adder_1_U.clk )
\sub_17ns_17ns_17_2_1_U2.top_sub_17ns_17ns_17_2_1_Adder_1_U.carry_s1  <= _186_;
assign _185_ = \sub_17ns_17ns_17_2_1_U2.top_sub_17ns_17ns_17_2_1_Adder_1_U.ce  ? \sub_17ns_17ns_17_2_1_U2.top_sub_17ns_17ns_17_2_1_Adder_1_U.bin_s0 [16:8] : \sub_17ns_17ns_17_2_1_U2.top_sub_17ns_17ns_17_2_1_Adder_1_U.bin_s1 ;
assign _184_ = \sub_17ns_17ns_17_2_1_U2.top_sub_17ns_17ns_17_2_1_Adder_1_U.ce  ? \sub_17ns_17ns_17_2_1_U2.top_sub_17ns_17ns_17_2_1_Adder_1_U.a [16:8] : \sub_17ns_17ns_17_2_1_U2.top_sub_17ns_17ns_17_2_1_Adder_1_U.ain_s1 ;
assign _186_ = \sub_17ns_17ns_17_2_1_U2.top_sub_17ns_17ns_17_2_1_Adder_1_U.ce  ? \sub_17ns_17ns_17_2_1_U2.top_sub_17ns_17ns_17_2_1_Adder_1_U.facout_s1  : \sub_17ns_17ns_17_2_1_U2.top_sub_17ns_17ns_17_2_1_Adder_1_U.carry_s1 ;
assign _187_ = \sub_17ns_17ns_17_2_1_U2.top_sub_17ns_17ns_17_2_1_Adder_1_U.ce  ? \sub_17ns_17ns_17_2_1_U2.top_sub_17ns_17ns_17_2_1_Adder_1_U.fas_s1  : \sub_17ns_17ns_17_2_1_U2.top_sub_17ns_17ns_17_2_1_Adder_1_U.sum_s1 ;
assign _188_ = \sub_17ns_17ns_17_2_1_U2.top_sub_17ns_17ns_17_2_1_Adder_1_U.u1.a  + \sub_17ns_17ns_17_2_1_U2.top_sub_17ns_17ns_17_2_1_Adder_1_U.u1.b ;
assign { \sub_17ns_17ns_17_2_1_U2.top_sub_17ns_17ns_17_2_1_Adder_1_U.u1.cout , \sub_17ns_17ns_17_2_1_U2.top_sub_17ns_17ns_17_2_1_Adder_1_U.u1.s  } = _188_ + \sub_17ns_17ns_17_2_1_U2.top_sub_17ns_17ns_17_2_1_Adder_1_U.u1.cin ;
assign _189_ = \sub_17ns_17ns_17_2_1_U2.top_sub_17ns_17ns_17_2_1_Adder_1_U.u2.a  + \sub_17ns_17ns_17_2_1_U2.top_sub_17ns_17ns_17_2_1_Adder_1_U.u2.b ;
assign { \sub_17ns_17ns_17_2_1_U2.top_sub_17ns_17ns_17_2_1_Adder_1_U.u2.cout , \sub_17ns_17ns_17_2_1_U2.top_sub_17ns_17ns_17_2_1_Adder_1_U.u2.s  } = _189_ + \sub_17ns_17ns_17_2_1_U2.top_sub_17ns_17ns_17_2_1_Adder_1_U.u2.cin ;
assign \sub_33s_33ns_33_2_1_U1.top_sub_33s_33ns_33_2_1_Adder_0_U.bin_s0  = ~ \sub_33s_33ns_33_2_1_U1.top_sub_33s_33ns_33_2_1_Adder_0_U.b ;
always @(posedge \sub_33s_33ns_33_2_1_U1.top_sub_33s_33ns_33_2_1_Adder_0_U.clk )
\sub_33s_33ns_33_2_1_U1.top_sub_33s_33ns_33_2_1_Adder_0_U.bin_s1  <= _191_;
always @(posedge \sub_33s_33ns_33_2_1_U1.top_sub_33s_33ns_33_2_1_Adder_0_U.clk )
\sub_33s_33ns_33_2_1_U1.top_sub_33s_33ns_33_2_1_Adder_0_U.ain_s1  <= _190_;
always @(posedge \sub_33s_33ns_33_2_1_U1.top_sub_33s_33ns_33_2_1_Adder_0_U.clk )
\sub_33s_33ns_33_2_1_U1.top_sub_33s_33ns_33_2_1_Adder_0_U.sum_s1  <= _193_;
always @(posedge \sub_33s_33ns_33_2_1_U1.top_sub_33s_33ns_33_2_1_Adder_0_U.clk )
\sub_33s_33ns_33_2_1_U1.top_sub_33s_33ns_33_2_1_Adder_0_U.carry_s1  <= _192_;
assign _191_ = \sub_33s_33ns_33_2_1_U1.top_sub_33s_33ns_33_2_1_Adder_0_U.ce  ? \sub_33s_33ns_33_2_1_U1.top_sub_33s_33ns_33_2_1_Adder_0_U.bin_s0 [32:16] : \sub_33s_33ns_33_2_1_U1.top_sub_33s_33ns_33_2_1_Adder_0_U.bin_s1 ;
assign _190_ = \sub_33s_33ns_33_2_1_U1.top_sub_33s_33ns_33_2_1_Adder_0_U.ce  ? \sub_33s_33ns_33_2_1_U1.top_sub_33s_33ns_33_2_1_Adder_0_U.a [32:16] : \sub_33s_33ns_33_2_1_U1.top_sub_33s_33ns_33_2_1_Adder_0_U.ain_s1 ;
assign _192_ = \sub_33s_33ns_33_2_1_U1.top_sub_33s_33ns_33_2_1_Adder_0_U.ce  ? \sub_33s_33ns_33_2_1_U1.top_sub_33s_33ns_33_2_1_Adder_0_U.facout_s1  : \sub_33s_33ns_33_2_1_U1.top_sub_33s_33ns_33_2_1_Adder_0_U.carry_s1 ;
assign _193_ = \sub_33s_33ns_33_2_1_U1.top_sub_33s_33ns_33_2_1_Adder_0_U.ce  ? \sub_33s_33ns_33_2_1_U1.top_sub_33s_33ns_33_2_1_Adder_0_U.fas_s1  : \sub_33s_33ns_33_2_1_U1.top_sub_33s_33ns_33_2_1_Adder_0_U.sum_s1 ;
assign _194_ = \sub_33s_33ns_33_2_1_U1.top_sub_33s_33ns_33_2_1_Adder_0_U.u1.a  + \sub_33s_33ns_33_2_1_U1.top_sub_33s_33ns_33_2_1_Adder_0_U.u1.b ;
assign { \sub_33s_33ns_33_2_1_U1.top_sub_33s_33ns_33_2_1_Adder_0_U.u1.cout , \sub_33s_33ns_33_2_1_U1.top_sub_33s_33ns_33_2_1_Adder_0_U.u1.s  } = _194_ + \sub_33s_33ns_33_2_1_U1.top_sub_33s_33ns_33_2_1_Adder_0_U.u1.cin ;
assign _195_ = \sub_33s_33ns_33_2_1_U1.top_sub_33s_33ns_33_2_1_Adder_0_U.u2.a  + \sub_33s_33ns_33_2_1_U1.top_sub_33s_33ns_33_2_1_Adder_0_U.u2.b ;
assign { \sub_33s_33ns_33_2_1_U1.top_sub_33s_33ns_33_2_1_Adder_0_U.u2.cout , \sub_33s_33ns_33_2_1_U1.top_sub_33s_33ns_33_2_1_Adder_0_U.u2.s  } = _195_ + \sub_33s_33ns_33_2_1_U1.top_sub_33s_33ns_33_2_1_Adder_0_U.u2.cin ;
assign _196_ = op_9_V_reg_1269 != op_5;
assign _197_ = | op_1[3:2];
assign _198_ = | tmp_4_reg_1199;
assign _199_ = | p_Result_s_reg_1149;
assign _200_ = tmp_4_reg_1199 != 16'hffff;
assign _201_ = p_Result_s_reg_1149 != 31'h7fffffff;
assign _202_ = | { trunc_ln851_2_reg_1321, 18'h00000 };
assign _203_ = | trunc_ln851_3_reg_1424;
assign _204_ = | op_15[20:0];
assign or_ln1195_fu_619_p2 = { op_5[1], op_5[1], op_5[1], op_5[1], op_5[1], op_5[1], op_5[1], op_5 } | { trunc_ln728_reg_1115, 1'h0 };
assign or_ln384_1_fu_595_p2 = underflow_1_fu_583_p2 | overflow_2_reg_1258;
assign or_ln384_fu_506_p2 = underflow_fu_501_p2 | overflow_reg_1205;
assign or_ln785_2_fu_521_p2 = p_Result_18_reg_1192 | icmp_ln768_2_reg_1231;
assign or_ln785_fu_416_p2 = p_Result_15_reg_1143 | icmp_ln768_reg_1176;
assign or_ln786_fu_578_p2 = xor_ln786_1_fu_573_p2 | icmp_ln786_1_reg_1236;
assign or_ln788_1_fu_496_p2 = or_ln788_fu_491_p2 | icmp_ln786_reg_1181;
assign or_ln788_fu_491_p2 = xor_ln786_fu_486_p2 | icmp_ln790_reg_1211;
assign overflow_1_fu_362_p2 = op_1[1] | icmp_ln768_1_reg_1127;
assign overflow_3_fu_867_p2 = r_V_fu_840_p2[3] | and_ln731_reg_1403[2];
always @(posedge ap_clk)
op_14_V_reg_1414[0] <= 1'h0;
always @(posedge ap_clk)
trunc_ln851_3_reg_1424[0] <= 1'h0;
always @(posedge ap_clk)
sext_ln850_reg_1361 <= _057_;
always @(posedge ap_clk)
select_ln353_reg_1461 <= _055_;
always @(posedge ap_clk)
ret_V_5_reg_1311 <= _049_;
always @(posedge ap_clk)
select_ln850_3_reg_1316 <= _056_;
always @(posedge ap_clk)
trunc_ln851_2_reg_1321 <= _062_;
always @(posedge ap_clk)
ret_V_4_reg_1291 <= _048_;
always @(posedge ap_clk)
ret_V_24_reg_1555 <= _044_;
always @(posedge ap_clk)
select_ln1192_reg_1560 <= _054_;
always @(posedge ap_clk)
ret_V_23_reg_1538 <= _043_;
always @(posedge ap_clk)
ret_V_27_cast_reg_1543 <= _046_;
always @(posedge ap_clk)
ret_V_21_reg_1481 <= _040_;
always @(posedge ap_clk)
ret_V_25_cast_reg_1486 <= _045_;
always @(posedge ap_clk)
ret_V_20_reg_1444 <= _039_;
always @(posedge ap_clk)
ret_V_23_cast_reg_1449 <= _042_;
always @(posedge ap_clk)
ret_V_19_reg_1393 <= _038_;
always @(posedge ap_clk)
ret_V_18_reg_1373 <= _037_;
always @(posedge ap_clk)
ret_V_15_reg_1346 <= _034_;
always @(posedge ap_clk)
ret_V_17_reg_1351 <= _036_;
always @(posedge ap_clk)
tmp_6_reg_1356 <= _059_;
always @(posedge ap_clk)
or_ln384_reg_1241 <= _026_;
always @(posedge ap_clk)
ret_V_16_reg_1246 <= _035_;
always @(posedge ap_clk)
ret_V_3_reg_1251 <= _047_;
always @(posedge ap_clk)
overflow_2_reg_1258 <= _027_;
always @(posedge ap_clk)
ret_reg_1132 <= _052_;
always @(posedge ap_clk)
p_Result_14_reg_1137 <= _029_;
always @(posedge ap_clk)
p_Result_15_reg_1143 <= _030_;
always @(posedge ap_clk)
p_Result_s_reg_1149 <= _033_;
always @(posedge ap_clk)
trunc_ln790_reg_1155 <= _061_;
always @(posedge ap_clk)
op_8_V_reg_1165 <= _023_;
always @(posedge ap_clk)
op_3_V_reg_1264 <= _022_;
always @(posedge ap_clk)
op_9_V_reg_1269 <= _024_;
always @(posedge ap_clk)
op_28_V_reg_1518 <= _021_;
always @(posedge ap_clk)
op_22_V_reg_1383 <= _019_;
always @(posedge ap_clk)
op_14_V_reg_1414[3:1] <= _018_;
always @(posedge ap_clk)
op_24_V_reg_1419 <= _020_;
always @(posedge ap_clk)
trunc_ln851_3_reg_1424[2:1] <= _063_;
always @(posedge ap_clk)
icmp_ln851_3_reg_1476 <= _016_;
always @(posedge ap_clk)
icmp_ln851_2_reg_1439 <= _015_;
always @(posedge ap_clk)
ret_V_reg_1326 <= _051_;
always @(posedge ap_clk)
icmp_ln851_1_reg_1341 <= _014_;
always @(posedge ap_clk)
icmp_ln768_reg_1176 <= _010_;
always @(posedge ap_clk)
icmp_ln786_reg_1181 <= _012_;
always @(posedge ap_clk)
p_Result_17_reg_1186 <= _031_;
always @(posedge ap_clk)
p_Result_18_reg_1192 <= _032_;
always @(posedge ap_clk)
tmp_4_reg_1199 <= _058_;
always @(posedge ap_clk)
overflow_reg_1205 <= _028_;
always @(posedge ap_clk)
icmp_ln790_reg_1211 <= _013_;
always @(posedge ap_clk)
icmp_ln851_reg_1226 <= _017_;
always @(posedge ap_clk)
icmp_ln768_2_reg_1231 <= _009_;
always @(posedge ap_clk)
icmp_ln786_1_reg_1236 <= _011_;
always @(posedge ap_clk)
trunc_ln728_reg_1115 <= _060_;
always @(posedge ap_clk)
rhs_3_reg_1120 <= _053_;
always @(posedge ap_clk)
icmp_ln768_1_reg_1127 <= _008_;
always @(posedge ap_clk)
or_ln1195_reg_1279 <= _025_;
always @(posedge ap_clk)
ret_V_cast_reg_1284 <= _050_;
always @(posedge ap_clk)
icmp_ln1499_reg_1306 <= _007_;
always @(posedge ap_clk)
and_ln731_reg_1403 <= _005_;
always @(posedge ap_clk)
ret_V_22_reg_1508 <= _041_;
always @(posedge ap_clk)
add_ln69_reg_1513 <= _004_;
always @(posedge ap_clk)
add_ln691_reg_1368 <= _003_;
always @(posedge ap_clk)
add_ln691_3_reg_1550 <= _002_;
always @(posedge ap_clk)
add_ln691_2_reg_1498 <= _001_;
always @(posedge ap_clk)
add_ln691_1_reg_1456 <= _000_;
always @(posedge ap_clk)
ap_CS_fsm <= _006_;
assign _064_ = _070_ ? 2'h2 : 2'h1;
assign _205_ = ap_CS_fsm == 1'h1;
function [37:0] _593_;
input [37:0] a;
input [1443:0] b;
input [37:0] s;
case (s)
38'b00000000000000000000000000000000000001:
_593_ = b[37:0];
38'b00000000000000000000000000000000000010:
_593_ = b[75:38];
38'b00000000000000000000000000000000000100:
_593_ = b[113:76];
38'b00000000000000000000000000000000001000:
_593_ = b[151:114];
38'b00000000000000000000000000000000010000:
_593_ = b[189:152];
38'b00000000000000000000000000000000100000:
_593_ = b[227:190];
38'b00000000000000000000000000000001000000:
_593_ = b[265:228];
38'b00000000000000000000000000000010000000:
_593_ = b[303:266];
38'b00000000000000000000000000000100000000:
_593_ = b[341:304];
38'b00000000000000000000000000001000000000:
_593_ = b[379:342];
38'b00000000000000000000000000010000000000:
_593_ = b[417:380];
38'b00000000000000000000000000100000000000:
_593_ = b[455:418];
38'b00000000000000000000000001000000000000:
_593_ = b[493:456];
38'b00000000000000000000000010000000000000:
_593_ = b[531:494];
38'b00000000000000000000000100000000000000:
_593_ = b[569:532];
38'b00000000000000000000001000000000000000:
_593_ = b[607:570];
38'b00000000000000000000010000000000000000:
_593_ = b[645:608];
38'b00000000000000000000100000000000000000:
_593_ = b[683:646];
38'b00000000000000000001000000000000000000:
_593_ = b[721:684];
38'b00000000000000000010000000000000000000:
_593_ = b[759:722];
38'b00000000000000000100000000000000000000:
_593_ = b[797:760];
38'b00000000000000001000000000000000000000:
_593_ = b[835:798];
38'b00000000000000010000000000000000000000:
_593_ = b[873:836];
38'b00000000000000100000000000000000000000:
_593_ = b[911:874];
38'b00000000000001000000000000000000000000:
_593_ = b[949:912];
38'b00000000000010000000000000000000000000:
_593_ = b[987:950];
38'b00000000000100000000000000000000000000:
_593_ = b[1025:988];
38'b00000000001000000000000000000000000000:
_593_ = b[1063:1026];
38'b00000000010000000000000000000000000000:
_593_ = b[1101:1064];
38'b00000000100000000000000000000000000000:
_593_ = b[1139:1102];
38'b00000001000000000000000000000000000000:
_593_ = b[1177:1140];
38'b00000010000000000000000000000000000000:
_593_ = b[1215:1178];
38'b00000100000000000000000000000000000000:
_593_ = b[1253:1216];
38'b00001000000000000000000000000000000000:
_593_ = b[1291:1254];
38'b00010000000000000000000000000000000000:
_593_ = b[1329:1292];
38'b00100000000000000000000000000000000000:
_593_ = b[1367:1330];
38'b01000000000000000000000000000000000000:
_593_ = b[1405:1368];
38'b10000000000000000000000000000000000000:
_593_ = b[1443:1406];
38'b00000000000000000000000000000000000000:
_593_ = a;
default:
_593_ = 38'bx;
endcase
endfunction
assign ap_NS_fsm = _593_(38'hxxxxxxxxxx, { 36'h000000000, _064_, 1406'h0000000004000000002000000001000000000800000000400000000200000000100000000080000000040000000020000000010000000008000000004000000002000000001000000000800000000400000000200000000100000000080000000040000000020000000010000000008000000004000000002000000001000000000800000000400000000200000000100000000080000000040000000020000000010000000008000000000000000001 }, { _205_, _242_, _241_, _240_, _239_, _238_, _237_, _236_, _235_, _234_, _233_, _232_, _231_, _230_, _229_, _228_, _227_, _226_, _225_, _224_, _223_, _222_, _221_, _220_, _219_, _218_, _217_, _216_, _215_, _214_, _213_, _212_, _211_, _210_, _209_, _208_, _207_, _206_ });
assign _206_ = ap_CS_fsm == 38'h2000000000;
assign _207_ = ap_CS_fsm == 37'h1000000000;
assign _208_ = ap_CS_fsm == 36'h800000000;
assign _209_ = ap_CS_fsm == 35'h400000000;
assign _210_ = ap_CS_fsm == 34'h200000000;
assign _211_ = ap_CS_fsm == 33'h100000000;
assign _212_ = ap_CS_fsm == 32'd2147483648;
assign _213_ = ap_CS_fsm == 31'h40000000;
assign _214_ = ap_CS_fsm == 30'h20000000;
assign _215_ = ap_CS_fsm == 29'h10000000;
assign _216_ = ap_CS_fsm == 28'h8000000;
assign _217_ = ap_CS_fsm == 27'h4000000;
assign _218_ = ap_CS_fsm == 26'h2000000;
assign _219_ = ap_CS_fsm == 25'h1000000;
assign _220_ = ap_CS_fsm == 24'h800000;
assign _221_ = ap_CS_fsm == 23'h400000;
assign _222_ = ap_CS_fsm == 22'h200000;
assign _223_ = ap_CS_fsm == 21'h100000;
assign _224_ = ap_CS_fsm == 20'h80000;
assign _225_ = ap_CS_fsm == 19'h40000;
assign _226_ = ap_CS_fsm == 18'h20000;
assign _227_ = ap_CS_fsm == 17'h10000;
assign _228_ = ap_CS_fsm == 16'h8000;
assign _229_ = ap_CS_fsm == 15'h4000;
assign _230_ = ap_CS_fsm == 14'h2000;
assign _231_ = ap_CS_fsm == 13'h1000;
assign _232_ = ap_CS_fsm == 12'h800;
assign _233_ = ap_CS_fsm == 11'h400;
assign _234_ = ap_CS_fsm == 10'h200;
assign _235_ = ap_CS_fsm == 9'h100;
assign _236_ = ap_CS_fsm == 8'h80;
assign _237_ = ap_CS_fsm == 7'h40;
assign _238_ = ap_CS_fsm == 6'h20;
assign _239_ = ap_CS_fsm == 5'h10;
assign _240_ = ap_CS_fsm == 4'h8;
assign _241_ = ap_CS_fsm == 3'h4;
assign _242_ = ap_CS_fsm == 2'h2;
assign op_30_ap_vld = ap_CS_fsm[37] ? 1'h1 : 1'h0;
assign ap_idle = _069_ ? 1'h1 : 1'h0;
assign _057_ = ap_CS_fsm[10] ? { tmp_6_reg_1356[16], tmp_6_reg_1356 } : sext_ln850_reg_1361;
assign _055_ = ap_CS_fsm[23] ? select_ln353_fu_937_p3 : select_ln353_reg_1461;
assign _062_ = ap_CS_fsm[7] ? grp_fu_650_p2[1:0] : trunc_ln851_2_reg_1321;
assign _056_ = ap_CS_fsm[7] ? select_ln850_3_fu_678_p3 : select_ln850_3_reg_1316;
assign _049_ = ap_CS_fsm[7] ? grp_fu_650_p2 : ret_V_5_reg_1311;
assign _048_ = _068_ ? grp_fu_561_p2 : ret_V_4_reg_1291;
assign _054_ = ap_CS_fsm[35] ? select_ln1192_fu_1081_p3 : select_ln1192_reg_1560;
assign _044_ = ap_CS_fsm[35] ? ret_V_24_fu_1074_p3 : ret_V_24_reg_1555;
assign _046_ = ap_CS_fsm[32] ? grp_fu_1037_p2[32:1] : ret_V_27_cast_reg_1543;
assign _043_ = ap_CS_fsm[32] ? grp_fu_1037_p2 : ret_V_23_reg_1538;
assign _045_ = ap_CS_fsm[25] ? grp_fu_959_p2[52:21] : ret_V_25_cast_reg_1486;
assign _040_ = ap_CS_fsm[25] ? grp_fu_959_p2 : ret_V_21_reg_1481;
assign _042_ = ap_CS_fsm[20] ? grp_fu_899_p2[34:3] : ret_V_23_cast_reg_1449;
assign _039_ = ap_CS_fsm[20] ? grp_fu_899_p2 : ret_V_20_reg_1444;
assign _038_ = ap_CS_fsm[16] ? grp_fu_803_p2 : ret_V_19_reg_1393;
assign _037_ = ap_CS_fsm[12] ? ret_V_18_fu_784_p3 : ret_V_18_reg_1373;
assign _059_ = ap_CS_fsm[9] ? grp_fu_711_p2[36:20] : tmp_6_reg_1356;
assign _036_ = ap_CS_fsm[9] ? grp_fu_711_p2 : ret_V_17_reg_1351;
assign _034_ = ap_CS_fsm[9] ? ret_V_15_fu_746_p3 : ret_V_15_reg_1346;
assign _027_ = ap_CS_fsm[4] ? overflow_2_fu_530_p2 : overflow_2_reg_1258;
assign _047_ = ap_CS_fsm[4] ? grp_fu_460_p2[32:17] : ret_V_3_reg_1251;
assign _035_ = ap_CS_fsm[4] ? grp_fu_460_p2 : ret_V_16_reg_1246;
assign _026_ = ap_CS_fsm[4] ? or_ln384_fu_506_p2 : or_ln384_reg_1241;
assign _023_ = ap_CS_fsm[1] ? op_8_V_fu_367_p3 : op_8_V_reg_1165;
assign _061_ = ap_CS_fsm[1] ? grp_fu_275_p2[0] : trunc_ln790_reg_1155;
assign _033_ = ap_CS_fsm[1] ? grp_fu_275_p2[32:2] : p_Result_s_reg_1149;
assign _030_ = ap_CS_fsm[1] ? grp_fu_275_p2[1] : p_Result_15_reg_1143;
assign _029_ = ap_CS_fsm[1] ? grp_fu_275_p2[32] : p_Result_14_reg_1137;
assign _052_ = ap_CS_fsm[1] ? grp_fu_275_p2 : ret_reg_1132;
assign _024_ = ap_CS_fsm[5] ? op_9_V_fu_600_p3 : op_9_V_reg_1269;
assign _022_ = ap_CS_fsm[5] ? op_3_V_fu_554_p3 : op_3_V_reg_1264;
assign _021_ = ap_CS_fsm[30] ? grp_fu_1018_p2 : op_28_V_reg_1518;
assign _019_ = ap_CS_fsm[14] ? grp_fu_794_p2 : op_22_V_reg_1383;
assign _063_ = ap_CS_fsm[18] ? op_14_V_fu_873_p3[2:1] : trunc_ln851_3_reg_1424[2:1];
assign _020_ = ap_CS_fsm[18] ? grp_fu_827_p2 : op_24_V_reg_1419;
assign _018_ = ap_CS_fsm[18] ? op_14_V_fu_873_p3[3:1] : op_14_V_reg_1414[3:1];
assign _016_ = ap_CS_fsm[24] ? icmp_ln851_3_fu_969_p2 : icmp_ln851_3_reg_1476;
assign _015_ = ap_CS_fsm[19] ? icmp_ln851_2_fu_905_p2 : icmp_ln851_2_reg_1439;
assign _014_ = ap_CS_fsm[8] ? icmp_ln851_1_fu_724_p2 : icmp_ln851_1_reg_1341;
assign _051_ = ap_CS_fsm[8] ? grp_fu_661_p2 : ret_V_reg_1326;
assign _058_ = ap_CS_fsm[2] ? grp_fu_378_p2[16:1] : tmp_4_reg_1199;
assign _032_ = ap_CS_fsm[2] ? grp_fu_378_p2[0] : p_Result_18_reg_1192;
assign _031_ = ap_CS_fsm[2] ? grp_fu_378_p2[16] : p_Result_17_reg_1186;
assign _012_ = ap_CS_fsm[2] ? icmp_ln786_fu_389_p2 : icmp_ln786_reg_1181;
assign _010_ = ap_CS_fsm[2] ? icmp_ln768_fu_384_p2 : icmp_ln768_reg_1176;
assign _011_ = ap_CS_fsm[3] ? icmp_ln786_1_fu_481_p2 : icmp_ln786_1_reg_1236;
assign _009_ = ap_CS_fsm[3] ? icmp_ln768_2_fu_476_p2 : icmp_ln768_2_reg_1231;
assign _017_ = ap_CS_fsm[3] ? icmp_ln851_fu_470_p2 : icmp_ln851_reg_1226;
assign _013_ = ap_CS_fsm[3] ? icmp_ln790_fu_438_p2 : icmp_ln790_reg_1211;
assign _028_ = ap_CS_fsm[3] ? overflow_fu_425_p2 : overflow_reg_1205;
assign _008_ = ap_CS_fsm[0] ? icmp_ln768_1_fu_305_p2 : icmp_ln768_1_reg_1127;
assign _053_ = ap_CS_fsm[0] ? rhs_3_fu_289_p2 : rhs_3_reg_1120;
assign _060_ = ap_CS_fsm[0] ? op_2[7:0] : trunc_ln728_reg_1115;
assign _007_ = ap_CS_fsm[6] ? icmp_ln1499_fu_656_p2 : icmp_ln1499_reg_1306;
assign _050_ = ap_CS_fsm[6] ? or_ln1195_fu_619_p2[8:1] : ret_V_cast_reg_1284;
assign _025_ = ap_CS_fsm[6] ? or_ln1195_fu_619_p2 : or_ln1195_reg_1279;
assign _005_ = ap_CS_fsm[17] ? and_ln731_fu_818_p2 : and_ln731_reg_1403;
assign _004_ = ap_CS_fsm[28] ? grp_fu_993_p2 : add_ln69_reg_1513;
assign _041_ = ap_CS_fsm[28] ? ret_V_22_fu_1011_p3 : ret_V_22_reg_1508;
assign _003_ = _067_ ? grp_fu_766_p2 : add_ln691_reg_1368;
assign _002_ = ap_CS_fsm[34] ? grp_fu_1053_p2 : add_ln691_3_reg_1550;
assign _001_ = _066_ ? grp_fu_985_p2 : add_ln691_2_reg_1498;
assign _000_ = _065_ ? grp_fu_920_p2 : add_ln691_1_reg_1456;
assign _006_ = ap_rst ? 38'h0000000001 : ap_NS_fsm;
assign icmp_ln1499_fu_656_p2 = _196_ ? 1'h1 : 1'h0;
assign icmp_ln768_1_fu_305_p2 = _197_ ? 1'h1 : 1'h0;
assign icmp_ln768_2_fu_476_p2 = _198_ ? 1'h1 : 1'h0;
assign icmp_ln768_fu_384_p2 = _199_ ? 1'h1 : 1'h0;
assign icmp_ln786_1_fu_481_p2 = _200_ ? 1'h1 : 1'h0;
assign icmp_ln786_fu_389_p2 = _201_ ? 1'h1 : 1'h0;
assign icmp_ln790_fu_438_p2 = _073_ ? 1'h1 : 1'h0;
assign icmp_ln851_1_fu_724_p2 = _202_ ? 1'h1 : 1'h0;
assign icmp_ln851_2_fu_905_p2 = _203_ ? 1'h1 : 1'h0;
assign icmp_ln851_3_fu_969_p2 = _204_ ? 1'h1 : 1'h0;
assign icmp_ln851_fu_470_p2 = _074_ ? 1'h1 : 1'h0;
assign op_14_V_fu_873_p3 = overflow_3_fu_867_p2 ? 4'h0 : { and_ln731_reg_1403, 1'h0 };
assign op_3_V_fu_554_p3 = or_ln384_reg_1241 ? select_ln384_1_fu_547_p3 : { ret_reg_1132[1:0], 2'h0 };
assign op_8_V_fu_367_p3 = overflow_1_fu_362_p2 ? 4'h7 : { op_1[1:0], 2'h0 };
assign op_9_V_fu_600_p3 = or_ln384_1_fu_595_p2 ? select_ln384_fu_588_p3 : { p_Result_18_reg_1192, 1'h0 };
assign ret_V_15_fu_746_p3 = op_5[1] ? select_ln850_fu_740_p3 : ret_V_cast_reg_1284;
assign ret_V_18_fu_784_p3 = ret_V_17_reg_1351[36] ? select_ln850_2_fu_779_p3 : sext_ln850_reg_1361;
assign ret_V_22_fu_1011_p3 = ret_V_21_reg_1481[53] ? select_ln850_4_fu_1006_p3 : ret_V_25_cast_reg_1486;
assign ret_V_24_fu_1074_p3 = ret_V_23_reg_1538[33] ? select_ln850_5_fu_1068_p3 : ret_V_27_cast_reg_1543;
assign rhs_3_fu_289_p2 = _075_ ? 1'h1 : 1'h0;
assign select_ln1118_1_fu_808_p3 = rhs_3_reg_1120 ? 3'h7 : 3'h0;
assign select_ln1118_fu_833_p3 = rhs_3_reg_1120 ? 4'hf : 4'h0;
assign select_ln1192_fu_1081_p3 = op_19 ? 32'd4294967295 : 32'd0;
assign select_ln353_fu_937_p3 = ret_V_20_reg_1444[35] ? select_ln850_6_fu_932_p3 : ret_V_23_cast_reg_1449;
assign select_ln384_1_fu_547_p3 = overflow_reg_1205 ? 4'h7 : 4'h9;
assign select_ln384_fu_588_p3 = overflow_2_reg_1258 ? 2'h1 : 2'h2;
assign select_ln850_1_fu_673_p3 = icmp_ln851_reg_1226 ? ret_V_3_reg_1251 : ret_V_4_reg_1291;
assign select_ln850_2_fu_779_p3 = icmp_ln851_1_reg_1341 ? add_ln691_reg_1368 : sext_ln850_reg_1361;
assign select_ln850_3_fu_678_p3 = ret_V_16_reg_1246[32] ? select_ln850_1_fu_673_p3 : ret_V_3_reg_1251;
assign select_ln850_4_fu_1006_p3 = icmp_ln851_3_reg_1476 ? add_ln691_2_reg_1498 : ret_V_25_cast_reg_1486;
assign select_ln850_5_fu_1068_p3 = op_18[0] ? add_ln691_3_reg_1550 : ret_V_27_cast_reg_1543;
assign select_ln850_6_fu_932_p3 = icmp_ln851_2_reg_1439 ? add_ln691_1_reg_1456 : ret_V_23_cast_reg_1449;
assign select_ln850_fu_740_p3 = or_ln1195_reg_1279[0] ? ret_V_reg_1326 : ret_V_cast_reg_1284;
assign ap_CS_fsm_state1 = ap_CS_fsm[0];
assign ap_CS_fsm_state10 = ap_CS_fsm[9];
assign ap_CS_fsm_state11 = ap_CS_fsm[10];
assign ap_CS_fsm_state12 = ap_CS_fsm[11];
assign ap_CS_fsm_state13 = ap_CS_fsm[12];
assign ap_CS_fsm_state14 = ap_CS_fsm[13];
assign ap_CS_fsm_state15 = ap_CS_fsm[14];
assign ap_CS_fsm_state16 = ap_CS_fsm[15];
assign ap_CS_fsm_state17 = ap_CS_fsm[16];
assign ap_CS_fsm_state18 = ap_CS_fsm[17];
assign ap_CS_fsm_state19 = ap_CS_fsm[18];
assign ap_CS_fsm_state2 = ap_CS_fsm[1];
assign ap_CS_fsm_state20 = ap_CS_fsm[19];
assign ap_CS_fsm_state21 = ap_CS_fsm[20];
assign ap_CS_fsm_state22 = ap_CS_fsm[21];
assign ap_CS_fsm_state23 = ap_CS_fsm[22];
assign ap_CS_fsm_state24 = ap_CS_fsm[23];
assign ap_CS_fsm_state25 = ap_CS_fsm[24];
assign ap_CS_fsm_state26 = ap_CS_fsm[25];
assign ap_CS_fsm_state27 = ap_CS_fsm[26];
assign ap_CS_fsm_state28 = ap_CS_fsm[27];
assign ap_CS_fsm_state29 = ap_CS_fsm[28];
assign ap_CS_fsm_state3 = ap_CS_fsm[2];
assign ap_CS_fsm_state30 = ap_CS_fsm[29];
assign ap_CS_fsm_state31 = ap_CS_fsm[30];
assign ap_CS_fsm_state32 = ap_CS_fsm[31];
assign ap_CS_fsm_state33 = ap_CS_fsm[32];
assign ap_CS_fsm_state34 = ap_CS_fsm[33];
assign ap_CS_fsm_state35 = ap_CS_fsm[34];
assign ap_CS_fsm_state36 = ap_CS_fsm[35];
assign ap_CS_fsm_state37 = ap_CS_fsm[36];
assign ap_CS_fsm_state38 = ap_CS_fsm[37];
assign ap_CS_fsm_state4 = ap_CS_fsm[3];
assign ap_CS_fsm_state5 = ap_CS_fsm[4];
assign ap_CS_fsm_state6 = ap_CS_fsm[5];
assign ap_CS_fsm_state7 = ap_CS_fsm[6];
assign ap_CS_fsm_state8 = ap_CS_fsm[7];
assign ap_CS_fsm_state9 = ap_CS_fsm[8];
assign ap_done = op_30_ap_vld;
assign ap_ready = op_30_ap_vld;
assign grp_fu_1037_p0 = { op_28_V_reg_1518[31], op_28_V_reg_1518, 1'h0 };
assign grp_fu_1037_p1 = { op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18 };
assign grp_fu_275_p0 = { op_1[31], op_1 };
assign grp_fu_275_p1 = { 17'h00000, op_2 };
assign grp_fu_378_p0 = { 1'h0, op_2 };
assign grp_fu_378_p1 = { 16'h0000, rhs_3_reg_1120 };
assign grp_fu_460_p0 = { 8'h00, op_0, 17'h00000 };
assign grp_fu_460_p1 = { op_7[31], op_7 };
assign grp_fu_650_p0 = { op_5[1], op_5[1], op_5, 1'h0 };
assign grp_fu_650_p1 = { op_3_V_reg_1264[3], op_3_V_reg_1264 };
assign grp_fu_711_p0 = { select_ln850_3_reg_1316[15], select_ln850_3_reg_1316, 20'h00000 };
assign grp_fu_711_p1 = { ret_V_5_reg_1311[4], ret_V_5_reg_1311[4], ret_V_5_reg_1311[4], ret_V_5_reg_1311[4], ret_V_5_reg_1311[4], ret_V_5_reg_1311[4], ret_V_5_reg_1311[4], ret_V_5_reg_1311[4], ret_V_5_reg_1311[4], ret_V_5_reg_1311[4], ret_V_5_reg_1311[4], ret_V_5_reg_1311[4], ret_V_5_reg_1311[4], ret_V_5_reg_1311[4], ret_V_5_reg_1311, 18'h00000 };
assign grp_fu_766_p0 = { tmp_6_reg_1356[16], tmp_6_reg_1356 };
assign grp_fu_794_p1 = { ret_V_15_reg_1346[7], ret_V_15_reg_1346[7], ret_V_15_reg_1346[7], ret_V_15_reg_1346[7], ret_V_15_reg_1346[7], ret_V_15_reg_1346[7], ret_V_15_reg_1346[7], ret_V_15_reg_1346[7], ret_V_15_reg_1346[7], ret_V_15_reg_1346[7], ret_V_15_reg_1346 };
assign grp_fu_803_p1 = { op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12 };
assign grp_fu_827_p0 = { ret_V_19_reg_1393[17], ret_V_19_reg_1393[17], ret_V_19_reg_1393[17], ret_V_19_reg_1393[17], ret_V_19_reg_1393[17], ret_V_19_reg_1393[17], ret_V_19_reg_1393[17], ret_V_19_reg_1393[17], ret_V_19_reg_1393[17], ret_V_19_reg_1393[17], ret_V_19_reg_1393[17], ret_V_19_reg_1393[17], ret_V_19_reg_1393[17], ret_V_19_reg_1393[17], ret_V_19_reg_1393 };
assign grp_fu_899_p0 = { op_24_V_reg_1419[31], op_24_V_reg_1419, 3'h0 };
assign grp_fu_899_p1 = { op_14_V_reg_1414[3], op_14_V_reg_1414[3], op_14_V_reg_1414[3], op_14_V_reg_1414[3], op_14_V_reg_1414[3], op_14_V_reg_1414[3], op_14_V_reg_1414[3], op_14_V_reg_1414[3], op_14_V_reg_1414[3], op_14_V_reg_1414[3], op_14_V_reg_1414[3], op_14_V_reg_1414[3], op_14_V_reg_1414[3], op_14_V_reg_1414[3], op_14_V_reg_1414[3], op_14_V_reg_1414[3], op_14_V_reg_1414[3], op_14_V_reg_1414[3], op_14_V_reg_1414[3], op_14_V_reg_1414[3], op_14_V_reg_1414[3], op_14_V_reg_1414[3], op_14_V_reg_1414[3], op_14_V_reg_1414[3], op_14_V_reg_1414[3], op_14_V_reg_1414[3], op_14_V_reg_1414[3], op_14_V_reg_1414[3], op_14_V_reg_1414[3], op_14_V_reg_1414[3], op_14_V_reg_1414[3], op_14_V_reg_1414[3], op_14_V_reg_1414 };
assign grp_fu_959_p0 = { select_ln353_reg_1461[31], select_ln353_reg_1461, 21'h000000 };
assign grp_fu_959_p1 = { op_15[31], op_15[31], op_15[31], op_15[31], op_15[31], op_15[31], op_15[31], op_15[31], op_15[31], op_15[31], op_15[31], op_15[31], op_15[31], op_15[31], op_15[31], op_15[31], op_15[31], op_15[31], op_15[31], op_15[31], op_15[31], op_15[31], op_15 };
assign grp_fu_993_p0 = { 31'h00000000, icmp_ln1499_reg_1306 };
assign icmp_ln1499_fu_656_p1 = op_5;
assign lhs_V_fu_444_p3 = { op_0, 17'h00000 };
assign lhs_cast_fu_608_p3 = { trunc_ln728_reg_1115, 1'h0 };
assign op_10_V_fu_689_p3 = { ret_V_5_reg_1311, 18'h00000 };
assign op_30 = grp_fu_1089_p2;
assign op_4_V_fu_263_p0 = op_1;
assign op_4_V_fu_263_p1 = op_1[3:0];
assign p_Result_10_fu_772_p3 = ret_V_17_reg_1351[36];
assign p_Result_11_fu_925_p3 = ret_V_20_reg_1444[35];
assign p_Result_12_fu_999_p3 = ret_V_21_reg_1481[53];
assign p_Result_13_fu_1058_p3 = ret_V_23_reg_1538[33];
assign p_Result_16_fu_355_p1 = op_1;
assign p_Result_16_fu_355_p3 = op_1[1];
assign p_Result_18_fu_402_p1 = grp_fu_378_p2[0];
assign p_Result_19_fu_852_p3 = and_ln731_reg_1403[2];
assign p_Result_3_fu_730_p1 = op_5;
assign p_Result_3_fu_730_p3 = op_5[1];
assign p_Result_4_fu_666_p3 = ret_V_16_reg_1246[32];
assign p_Result_9_fu_717_p3 = { trunc_ln851_2_reg_1321, 18'h00000 };
assign p_Result_s_20_fu_431_p3 = { trunc_ln790_reg_1155, 2'h0 };
assign p_Val2_1_fu_539_p3 = { ret_reg_1132[1:0], 2'h0 };
assign p_Val2_3_fu_347_p3 = { op_1[1:0], 2'h0 };
assign p_Val2_6_fu_566_p3 = { p_Result_18_reg_1192, 1'h0 };
assign p_Val2_8_fu_845_p3 = { and_ln731_reg_1403, 1'h0 };
assign rhs_2_fu_700_p3 = { select_ln850_3_reg_1316, 20'h00000 };
assign rhs_5_fu_888_p3 = { op_24_V_reg_1419, 3'h0 };
assign rhs_6_fu_948_p3 = { select_ln353_reg_1461, 21'h000000 };
assign rhs_8_fu_1026_p3 = { op_28_V_reg_1518, 1'h0 };
assign rhs_fu_638_p1 = op_5;
assign rhs_fu_638_p3 = { op_5, 1'h0 };
assign sext_ln1195_fu_615_p0 = op_5;
assign sext_ln1195_fu_615_p1 = { op_5[1], op_5[1], op_5[1], op_5[1], op_5[1], op_5[1], op_5[1], op_5 };
assign sext_ln215_fu_267_p0 = op_1;
assign sext_ln703_3_fu_944_p0 = op_15;
assign sext_ln703_4_fu_1022_p0 = op_18;
assign sext_ln703_fu_456_p0 = op_7;
assign sext_ln850_fu_763_p1 = { tmp_6_reg_1356[16], tmp_6_reg_1356 };
assign tmp_3_fu_295_p1 = op_1;
assign tmp_3_fu_295_p4 = op_1[3:2];
assign tmp_fu_859_p3 = r_V_fu_840_p2[3];
assign trunc_ln728_fu_281_p1 = op_2[7:0];
assign trunc_ln731_1_fu_344_p0 = op_1;
assign trunc_ln731_1_fu_344_p1 = op_1[1:0];
assign trunc_ln731_3_fu_815_p1 = op_8_V_reg_1165[2:0];
assign trunc_ln731_fu_536_p1 = ret_reg_1132[1:0];
assign trunc_ln790_fu_337_p1 = grp_fu_275_p2[0];
assign trunc_ln851_1_fu_466_p0 = op_7;
assign trunc_ln851_1_fu_466_p1 = op_7[16:0];
assign trunc_ln851_2_fu_685_p1 = grp_fu_650_p2[1:0];
assign trunc_ln851_3_fu_881_p1 = op_14_V_fu_873_p3[2:0];
assign trunc_ln851_4_fu_965_p0 = op_15;
assign trunc_ln851_4_fu_965_p1 = op_15[20:0];
assign trunc_ln851_5_fu_1065_p0 = op_18;
assign trunc_ln851_5_fu_1065_p1 = op_18[0];
assign trunc_ln851_fu_737_p1 = or_ln1195_reg_1279[0];
assign zext_ln870_fu_285_p1 = { 12'h000, op_1[3:0] };
assign \sub_33s_33ns_33_2_1_U1.top_sub_33s_33ns_33_2_1_Adder_0_U.ain_s0  = \sub_33s_33ns_33_2_1_U1.top_sub_33s_33ns_33_2_1_Adder_0_U.a ;
assign \sub_33s_33ns_33_2_1_U1.top_sub_33s_33ns_33_2_1_Adder_0_U.s  = { \sub_33s_33ns_33_2_1_U1.top_sub_33s_33ns_33_2_1_Adder_0_U.fas_s2 , \sub_33s_33ns_33_2_1_U1.top_sub_33s_33ns_33_2_1_Adder_0_U.sum_s1  };
assign \sub_33s_33ns_33_2_1_U1.top_sub_33s_33ns_33_2_1_Adder_0_U.u2.a  = \sub_33s_33ns_33_2_1_U1.top_sub_33s_33ns_33_2_1_Adder_0_U.ain_s1 ;
assign \sub_33s_33ns_33_2_1_U1.top_sub_33s_33ns_33_2_1_Adder_0_U.u2.b  = \sub_33s_33ns_33_2_1_U1.top_sub_33s_33ns_33_2_1_Adder_0_U.bin_s1 ;
assign \sub_33s_33ns_33_2_1_U1.top_sub_33s_33ns_33_2_1_Adder_0_U.u2.cin  = \sub_33s_33ns_33_2_1_U1.top_sub_33s_33ns_33_2_1_Adder_0_U.carry_s1 ;
assign \sub_33s_33ns_33_2_1_U1.top_sub_33s_33ns_33_2_1_Adder_0_U.facout_s2  = \sub_33s_33ns_33_2_1_U1.top_sub_33s_33ns_33_2_1_Adder_0_U.u2.cout ;
assign \sub_33s_33ns_33_2_1_U1.top_sub_33s_33ns_33_2_1_Adder_0_U.fas_s2  = \sub_33s_33ns_33_2_1_U1.top_sub_33s_33ns_33_2_1_Adder_0_U.u2.s ;
assign \sub_33s_33ns_33_2_1_U1.top_sub_33s_33ns_33_2_1_Adder_0_U.u1.a  = \sub_33s_33ns_33_2_1_U1.top_sub_33s_33ns_33_2_1_Adder_0_U.a [15:0];
assign \sub_33s_33ns_33_2_1_U1.top_sub_33s_33ns_33_2_1_Adder_0_U.u1.b  = \sub_33s_33ns_33_2_1_U1.top_sub_33s_33ns_33_2_1_Adder_0_U.bin_s0 [15:0];
assign \sub_33s_33ns_33_2_1_U1.top_sub_33s_33ns_33_2_1_Adder_0_U.u1.cin  = 1'h1;
assign \sub_33s_33ns_33_2_1_U1.top_sub_33s_33ns_33_2_1_Adder_0_U.facout_s1  = \sub_33s_33ns_33_2_1_U1.top_sub_33s_33ns_33_2_1_Adder_0_U.u1.cout ;
assign \sub_33s_33ns_33_2_1_U1.top_sub_33s_33ns_33_2_1_Adder_0_U.fas_s1  = \sub_33s_33ns_33_2_1_U1.top_sub_33s_33ns_33_2_1_Adder_0_U.u1.s ;
assign \sub_33s_33ns_33_2_1_U1.top_sub_33s_33ns_33_2_1_Adder_0_U.a  = \sub_33s_33ns_33_2_1_U1.din0 ;
assign \sub_33s_33ns_33_2_1_U1.top_sub_33s_33ns_33_2_1_Adder_0_U.b  = \sub_33s_33ns_33_2_1_U1.din1 ;
assign \sub_33s_33ns_33_2_1_U1.top_sub_33s_33ns_33_2_1_Adder_0_U.ce  = \sub_33s_33ns_33_2_1_U1.ce ;
assign \sub_33s_33ns_33_2_1_U1.top_sub_33s_33ns_33_2_1_Adder_0_U.clk  = \sub_33s_33ns_33_2_1_U1.clk ;
assign \sub_33s_33ns_33_2_1_U1.top_sub_33s_33ns_33_2_1_Adder_0_U.reset  = \sub_33s_33ns_33_2_1_U1.reset ;
assign \sub_33s_33ns_33_2_1_U1.dout  = \sub_33s_33ns_33_2_1_U1.top_sub_33s_33ns_33_2_1_Adder_0_U.s ;
assign \sub_33s_33ns_33_2_1_U1.ce  = 1'h1;
assign \sub_33s_33ns_33_2_1_U1.clk  = ap_clk;
assign \sub_33s_33ns_33_2_1_U1.din0  = { op_1[31], op_1 };
assign \sub_33s_33ns_33_2_1_U1.din1  = { 17'h00000, op_2 };
assign grp_fu_275_p2 = \sub_33s_33ns_33_2_1_U1.dout ;
assign \sub_33s_33ns_33_2_1_U1.reset  = ap_rst;
assign \sub_17ns_17ns_17_2_1_U2.top_sub_17ns_17ns_17_2_1_Adder_1_U.ain_s0  = \sub_17ns_17ns_17_2_1_U2.top_sub_17ns_17ns_17_2_1_Adder_1_U.a ;
assign \sub_17ns_17ns_17_2_1_U2.top_sub_17ns_17ns_17_2_1_Adder_1_U.s  = { \sub_17ns_17ns_17_2_1_U2.top_sub_17ns_17ns_17_2_1_Adder_1_U.fas_s2 , \sub_17ns_17ns_17_2_1_U2.top_sub_17ns_17ns_17_2_1_Adder_1_U.sum_s1  };
assign \sub_17ns_17ns_17_2_1_U2.top_sub_17ns_17ns_17_2_1_Adder_1_U.u2.a  = \sub_17ns_17ns_17_2_1_U2.top_sub_17ns_17ns_17_2_1_Adder_1_U.ain_s1 ;
assign \sub_17ns_17ns_17_2_1_U2.top_sub_17ns_17ns_17_2_1_Adder_1_U.u2.b  = \sub_17ns_17ns_17_2_1_U2.top_sub_17ns_17ns_17_2_1_Adder_1_U.bin_s1 ;
assign \sub_17ns_17ns_17_2_1_U2.top_sub_17ns_17ns_17_2_1_Adder_1_U.u2.cin  = \sub_17ns_17ns_17_2_1_U2.top_sub_17ns_17ns_17_2_1_Adder_1_U.carry_s1 ;
assign \sub_17ns_17ns_17_2_1_U2.top_sub_17ns_17ns_17_2_1_Adder_1_U.facout_s2  = \sub_17ns_17ns_17_2_1_U2.top_sub_17ns_17ns_17_2_1_Adder_1_U.u2.cout ;
assign \sub_17ns_17ns_17_2_1_U2.top_sub_17ns_17ns_17_2_1_Adder_1_U.fas_s2  = \sub_17ns_17ns_17_2_1_U2.top_sub_17ns_17ns_17_2_1_Adder_1_U.u2.s ;
assign \sub_17ns_17ns_17_2_1_U2.top_sub_17ns_17ns_17_2_1_Adder_1_U.u1.a  = \sub_17ns_17ns_17_2_1_U2.top_sub_17ns_17ns_17_2_1_Adder_1_U.a [7:0];
assign \sub_17ns_17ns_17_2_1_U2.top_sub_17ns_17ns_17_2_1_Adder_1_U.u1.b  = \sub_17ns_17ns_17_2_1_U2.top_sub_17ns_17ns_17_2_1_Adder_1_U.bin_s0 [7:0];
assign \sub_17ns_17ns_17_2_1_U2.top_sub_17ns_17ns_17_2_1_Adder_1_U.u1.cin  = 1'h1;
assign \sub_17ns_17ns_17_2_1_U2.top_sub_17ns_17ns_17_2_1_Adder_1_U.facout_s1  = \sub_17ns_17ns_17_2_1_U2.top_sub_17ns_17ns_17_2_1_Adder_1_U.u1.cout ;
assign \sub_17ns_17ns_17_2_1_U2.top_sub_17ns_17ns_17_2_1_Adder_1_U.fas_s1  = \sub_17ns_17ns_17_2_1_U2.top_sub_17ns_17ns_17_2_1_Adder_1_U.u1.s ;
assign \sub_17ns_17ns_17_2_1_U2.top_sub_17ns_17ns_17_2_1_Adder_1_U.a  = \sub_17ns_17ns_17_2_1_U2.din0 ;
assign \sub_17ns_17ns_17_2_1_U2.top_sub_17ns_17ns_17_2_1_Adder_1_U.b  = \sub_17ns_17ns_17_2_1_U2.din1 ;
assign \sub_17ns_17ns_17_2_1_U2.top_sub_17ns_17ns_17_2_1_Adder_1_U.ce  = \sub_17ns_17ns_17_2_1_U2.ce ;
assign \sub_17ns_17ns_17_2_1_U2.top_sub_17ns_17ns_17_2_1_Adder_1_U.clk  = \sub_17ns_17ns_17_2_1_U2.clk ;
assign \sub_17ns_17ns_17_2_1_U2.top_sub_17ns_17ns_17_2_1_Adder_1_U.reset  = \sub_17ns_17ns_17_2_1_U2.reset ;
assign \sub_17ns_17ns_17_2_1_U2.dout  = \sub_17ns_17ns_17_2_1_U2.top_sub_17ns_17ns_17_2_1_Adder_1_U.s ;
assign \sub_17ns_17ns_17_2_1_U2.ce  = 1'h1;
assign \sub_17ns_17ns_17_2_1_U2.clk  = ap_clk;
assign \sub_17ns_17ns_17_2_1_U2.din0  = { 1'h0, op_2 };
assign \sub_17ns_17ns_17_2_1_U2.din1  = { 16'h0000, rhs_3_reg_1120 };
assign grp_fu_378_p2 = \sub_17ns_17ns_17_2_1_U2.dout ;
assign \sub_17ns_17ns_17_2_1_U2.reset  = ap_rst;
assign \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.ain_s0  = \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.a ;
assign \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.bin_s0  = \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.b ;
assign \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.s  = { \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.fas_s2 , \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.sum_s1  };
assign \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.u2.a  = \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.ain_s1 ;
assign \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.u2.b  = \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.bin_s1 ;
assign \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.u2.cin  = \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.carry_s1 ;
assign \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.facout_s2  = \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.u2.cout ;
assign \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.fas_s2  = \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.u2.s ;
assign \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.u1.a  = \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.a [3:0];
assign \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.u1.b  = \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.b [3:0];
assign \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.u1.cin  = 1'h0;
assign \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.facout_s1  = \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.u1.cout ;
assign \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.fas_s1  = \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.u1.s ;
assign \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.a  = \add_8ns_8ns_8_2_1_U6.din0 ;
assign \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.b  = \add_8ns_8ns_8_2_1_U6.din1 ;
assign \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.ce  = \add_8ns_8ns_8_2_1_U6.ce ;
assign \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.clk  = \add_8ns_8ns_8_2_1_U6.clk ;
assign \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.reset  = \add_8ns_8ns_8_2_1_U6.reset ;
assign \add_8ns_8ns_8_2_1_U6.dout  = \add_8ns_8ns_8_2_1_U6.top_add_8ns_8ns_8_2_1_Adder_5_U.s ;
assign \add_8ns_8ns_8_2_1_U6.ce  = 1'h1;
assign \add_8ns_8ns_8_2_1_U6.clk  = ap_clk;
assign \add_8ns_8ns_8_2_1_U6.din0  = ret_V_cast_reg_1284;
assign \add_8ns_8ns_8_2_1_U6.din1  = 8'h01;
assign grp_fu_661_p2 = \add_8ns_8ns_8_2_1_U6.dout ;
assign \add_8ns_8ns_8_2_1_U6.reset  = ap_rst;
assign \add_5s_5s_5_2_1_U5.top_add_5s_5s_5_2_1_Adder_4_U.ain_s0  = \add_5s_5s_5_2_1_U5.top_add_5s_5s_5_2_1_Adder_4_U.a ;
assign \add_5s_5s_5_2_1_U5.top_add_5s_5s_5_2_1_Adder_4_U.bin_s0  = \add_5s_5s_5_2_1_U5.top_add_5s_5s_5_2_1_Adder_4_U.b ;
assign \add_5s_5s_5_2_1_U5.top_add_5s_5s_5_2_1_Adder_4_U.s  = { \add_5s_5s_5_2_1_U5.top_add_5s_5s_5_2_1_Adder_4_U.fas_s2 , \add_5s_5s_5_2_1_U5.top_add_5s_5s_5_2_1_Adder_4_U.sum_s1  };
assign \add_5s_5s_5_2_1_U5.top_add_5s_5s_5_2_1_Adder_4_U.u2.a  = \add_5s_5s_5_2_1_U5.top_add_5s_5s_5_2_1_Adder_4_U.ain_s1 ;
assign \add_5s_5s_5_2_1_U5.top_add_5s_5s_5_2_1_Adder_4_U.u2.b  = \add_5s_5s_5_2_1_U5.top_add_5s_5s_5_2_1_Adder_4_U.bin_s1 ;
assign \add_5s_5s_5_2_1_U5.top_add_5s_5s_5_2_1_Adder_4_U.u2.cin  = \add_5s_5s_5_2_1_U5.top_add_5s_5s_5_2_1_Adder_4_U.carry_s1 ;
assign \add_5s_5s_5_2_1_U5.top_add_5s_5s_5_2_1_Adder_4_U.facout_s2  = \add_5s_5s_5_2_1_U5.top_add_5s_5s_5_2_1_Adder_4_U.u2.cout ;
assign \add_5s_5s_5_2_1_U5.top_add_5s_5s_5_2_1_Adder_4_U.fas_s2  = \add_5s_5s_5_2_1_U5.top_add_5s_5s_5_2_1_Adder_4_U.u2.s ;
assign \add_5s_5s_5_2_1_U5.top_add_5s_5s_5_2_1_Adder_4_U.u1.a  = \add_5s_5s_5_2_1_U5.top_add_5s_5s_5_2_1_Adder_4_U.a [1:0];
assign \add_5s_5s_5_2_1_U5.top_add_5s_5s_5_2_1_Adder_4_U.u1.b  = \add_5s_5s_5_2_1_U5.top_add_5s_5s_5_2_1_Adder_4_U.b [1:0];
assign \add_5s_5s_5_2_1_U5.top_add_5s_5s_5_2_1_Adder_4_U.u1.cin  = 1'h0;
assign \add_5s_5s_5_2_1_U5.top_add_5s_5s_5_2_1_Adder_4_U.facout_s1  = \add_5s_5s_5_2_1_U5.top_add_5s_5s_5_2_1_Adder_4_U.u1.cout ;
assign \add_5s_5s_5_2_1_U5.top_add_5s_5s_5_2_1_Adder_4_U.fas_s1  = \add_5s_5s_5_2_1_U5.top_add_5s_5s_5_2_1_Adder_4_U.u1.s ;
assign \add_5s_5s_5_2_1_U5.top_add_5s_5s_5_2_1_Adder_4_U.a  = \add_5s_5s_5_2_1_U5.din0 ;
assign \add_5s_5s_5_2_1_U5.top_add_5s_5s_5_2_1_Adder_4_U.b  = \add_5s_5s_5_2_1_U5.din1 ;
assign \add_5s_5s_5_2_1_U5.top_add_5s_5s_5_2_1_Adder_4_U.ce  = \add_5s_5s_5_2_1_U5.ce ;
assign \add_5s_5s_5_2_1_U5.top_add_5s_5s_5_2_1_Adder_4_U.clk  = \add_5s_5s_5_2_1_U5.clk ;
assign \add_5s_5s_5_2_1_U5.top_add_5s_5s_5_2_1_Adder_4_U.reset  = \add_5s_5s_5_2_1_U5.reset ;
assign \add_5s_5s_5_2_1_U5.dout  = \add_5s_5s_5_2_1_U5.top_add_5s_5s_5_2_1_Adder_4_U.s ;
assign \add_5s_5s_5_2_1_U5.ce  = 1'h1;
assign \add_5s_5s_5_2_1_U5.clk  = ap_clk;
assign \add_5s_5s_5_2_1_U5.din0  = { op_5[1], op_5[1], op_5, 1'h0 };
assign \add_5s_5s_5_2_1_U5.din1  = { op_3_V_reg_1264[3], op_3_V_reg_1264 };
assign grp_fu_650_p2 = \add_5s_5s_5_2_1_U5.dout ;
assign \add_5s_5s_5_2_1_U5.reset  = ap_rst;
assign \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_12_U.ain_s0  = \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_12_U.a ;
assign \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_12_U.bin_s0  = \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_12_U.b ;
assign \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_12_U.s  = { \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_12_U.fas_s2 , \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_12_U.sum_s1  };
assign \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_12_U.u2.a  = \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_12_U.ain_s1 ;
assign \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_12_U.u2.b  = \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_12_U.bin_s1 ;
assign \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_12_U.u2.cin  = \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_12_U.carry_s1 ;
assign \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_12_U.facout_s2  = \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_12_U.u2.cout ;
assign \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_12_U.fas_s2  = \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_12_U.u2.s ;
assign \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_12_U.u1.a  = \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_12_U.a [26:0];
assign \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_12_U.u1.b  = \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_12_U.b [26:0];
assign \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_12_U.u1.cin  = 1'h0;
assign \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_12_U.facout_s1  = \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_12_U.u1.cout ;
assign \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_12_U.fas_s1  = \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_12_U.u1.s ;
assign \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_12_U.a  = \add_54s_54s_54_2_1_U14.din0 ;
assign \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_12_U.b  = \add_54s_54s_54_2_1_U14.din1 ;
assign \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_12_U.ce  = \add_54s_54s_54_2_1_U14.ce ;
assign \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_12_U.clk  = \add_54s_54s_54_2_1_U14.clk ;
assign \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_12_U.reset  = \add_54s_54s_54_2_1_U14.reset ;
assign \add_54s_54s_54_2_1_U14.dout  = \add_54s_54s_54_2_1_U14.top_add_54s_54s_54_2_1_Adder_12_U.s ;
assign \add_54s_54s_54_2_1_U14.ce  = 1'h1;
assign \add_54s_54s_54_2_1_U14.clk  = ap_clk;
assign \add_54s_54s_54_2_1_U14.din0  = { select_ln353_reg_1461[31], select_ln353_reg_1461, 21'h000000 };
assign \add_54s_54s_54_2_1_U14.din1  = { op_15[31], op_15[31], op_15[31], op_15[31], op_15[31], op_15[31], op_15[31], op_15[31], op_15[31], op_15[31], op_15[31], op_15[31], op_15[31], op_15[31], op_15[31], op_15[31], op_15[31], op_15[31], op_15[31], op_15[31], op_15[31], op_15[31], op_15 };
assign grp_fu_959_p2 = \add_54s_54s_54_2_1_U14.dout ;
assign \add_54s_54s_54_2_1_U14.reset  = ap_rst;
assign \add_37s_37s_37_2_1_U7.top_add_37s_37s_37_2_1_Adder_6_U.ain_s0  = \add_37s_37s_37_2_1_U7.top_add_37s_37s_37_2_1_Adder_6_U.a ;
assign \add_37s_37s_37_2_1_U7.top_add_37s_37s_37_2_1_Adder_6_U.bin_s0  = \add_37s_37s_37_2_1_U7.top_add_37s_37s_37_2_1_Adder_6_U.b ;
assign \add_37s_37s_37_2_1_U7.top_add_37s_37s_37_2_1_Adder_6_U.s  = { \add_37s_37s_37_2_1_U7.top_add_37s_37s_37_2_1_Adder_6_U.fas_s2 , \add_37s_37s_37_2_1_U7.top_add_37s_37s_37_2_1_Adder_6_U.sum_s1  };
assign \add_37s_37s_37_2_1_U7.top_add_37s_37s_37_2_1_Adder_6_U.u2.a  = \add_37s_37s_37_2_1_U7.top_add_37s_37s_37_2_1_Adder_6_U.ain_s1 ;
assign \add_37s_37s_37_2_1_U7.top_add_37s_37s_37_2_1_Adder_6_U.u2.b  = \add_37s_37s_37_2_1_U7.top_add_37s_37s_37_2_1_Adder_6_U.bin_s1 ;
assign \add_37s_37s_37_2_1_U7.top_add_37s_37s_37_2_1_Adder_6_U.u2.cin  = \add_37s_37s_37_2_1_U7.top_add_37s_37s_37_2_1_Adder_6_U.carry_s1 ;
assign \add_37s_37s_37_2_1_U7.top_add_37s_37s_37_2_1_Adder_6_U.facout_s2  = \add_37s_37s_37_2_1_U7.top_add_37s_37s_37_2_1_Adder_6_U.u2.cout ;
assign \add_37s_37s_37_2_1_U7.top_add_37s_37s_37_2_1_Adder_6_U.fas_s2  = \add_37s_37s_37_2_1_U7.top_add_37s_37s_37_2_1_Adder_6_U.u2.s ;
assign \add_37s_37s_37_2_1_U7.top_add_37s_37s_37_2_1_Adder_6_U.u1.a  = \add_37s_37s_37_2_1_U7.top_add_37s_37s_37_2_1_Adder_6_U.a [17:0];
assign \add_37s_37s_37_2_1_U7.top_add_37s_37s_37_2_1_Adder_6_U.u1.b  = \add_37s_37s_37_2_1_U7.top_add_37s_37s_37_2_1_Adder_6_U.b [17:0];
assign \add_37s_37s_37_2_1_U7.top_add_37s_37s_37_2_1_Adder_6_U.u1.cin  = 1'h0;
assign \add_37s_37s_37_2_1_U7.top_add_37s_37s_37_2_1_Adder_6_U.facout_s1  = \add_37s_37s_37_2_1_U7.top_add_37s_37s_37_2_1_Adder_6_U.u1.cout ;
assign \add_37s_37s_37_2_1_U7.top_add_37s_37s_37_2_1_Adder_6_U.fas_s1  = \add_37s_37s_37_2_1_U7.top_add_37s_37s_37_2_1_Adder_6_U.u1.s ;
assign \add_37s_37s_37_2_1_U7.top_add_37s_37s_37_2_1_Adder_6_U.a  = \add_37s_37s_37_2_1_U7.din0 ;
assign \add_37s_37s_37_2_1_U7.top_add_37s_37s_37_2_1_Adder_6_U.b  = \add_37s_37s_37_2_1_U7.din1 ;
assign \add_37s_37s_37_2_1_U7.top_add_37s_37s_37_2_1_Adder_6_U.ce  = \add_37s_37s_37_2_1_U7.ce ;
assign \add_37s_37s_37_2_1_U7.top_add_37s_37s_37_2_1_Adder_6_U.clk  = \add_37s_37s_37_2_1_U7.clk ;
assign \add_37s_37s_37_2_1_U7.top_add_37s_37s_37_2_1_Adder_6_U.reset  = \add_37s_37s_37_2_1_U7.reset ;
assign \add_37s_37s_37_2_1_U7.dout  = \add_37s_37s_37_2_1_U7.top_add_37s_37s_37_2_1_Adder_6_U.s ;
assign \add_37s_37s_37_2_1_U7.ce  = 1'h1;
assign \add_37s_37s_37_2_1_U7.clk  = ap_clk;
assign \add_37s_37s_37_2_1_U7.din0  = { select_ln850_3_reg_1316[15], select_ln850_3_reg_1316, 20'h00000 };
assign \add_37s_37s_37_2_1_U7.din1  = { ret_V_5_reg_1311[4], ret_V_5_reg_1311[4], ret_V_5_reg_1311[4], ret_V_5_reg_1311[4], ret_V_5_reg_1311[4], ret_V_5_reg_1311[4], ret_V_5_reg_1311[4], ret_V_5_reg_1311[4], ret_V_5_reg_1311[4], ret_V_5_reg_1311[4], ret_V_5_reg_1311[4], ret_V_5_reg_1311[4], ret_V_5_reg_1311[4], ret_V_5_reg_1311[4], ret_V_5_reg_1311, 18'h00000 };
assign grp_fu_711_p2 = \add_37s_37s_37_2_1_U7.dout ;
assign \add_37s_37s_37_2_1_U7.reset  = ap_rst;
assign \add_36s_36s_36_2_1_U12.top_add_36s_36s_36_2_1_Adder_10_U.ain_s0  = \add_36s_36s_36_2_1_U12.top_add_36s_36s_36_2_1_Adder_10_U.a ;
assign \add_36s_36s_36_2_1_U12.top_add_36s_36s_36_2_1_Adder_10_U.bin_s0  = \add_36s_36s_36_2_1_U12.top_add_36s_36s_36_2_1_Adder_10_U.b ;
assign \add_36s_36s_36_2_1_U12.top_add_36s_36s_36_2_1_Adder_10_U.s  = { \add_36s_36s_36_2_1_U12.top_add_36s_36s_36_2_1_Adder_10_U.fas_s2 , \add_36s_36s_36_2_1_U12.top_add_36s_36s_36_2_1_Adder_10_U.sum_s1  };
assign \add_36s_36s_36_2_1_U12.top_add_36s_36s_36_2_1_Adder_10_U.u2.a  = \add_36s_36s_36_2_1_U12.top_add_36s_36s_36_2_1_Adder_10_U.ain_s1 ;
assign \add_36s_36s_36_2_1_U12.top_add_36s_36s_36_2_1_Adder_10_U.u2.b  = \add_36s_36s_36_2_1_U12.top_add_36s_36s_36_2_1_Adder_10_U.bin_s1 ;
assign \add_36s_36s_36_2_1_U12.top_add_36s_36s_36_2_1_Adder_10_U.u2.cin  = \add_36s_36s_36_2_1_U12.top_add_36s_36s_36_2_1_Adder_10_U.carry_s1 ;
assign \add_36s_36s_36_2_1_U12.top_add_36s_36s_36_2_1_Adder_10_U.facout_s2  = \add_36s_36s_36_2_1_U12.top_add_36s_36s_36_2_1_Adder_10_U.u2.cout ;
assign \add_36s_36s_36_2_1_U12.top_add_36s_36s_36_2_1_Adder_10_U.fas_s2  = \add_36s_36s_36_2_1_U12.top_add_36s_36s_36_2_1_Adder_10_U.u2.s ;
assign \add_36s_36s_36_2_1_U12.top_add_36s_36s_36_2_1_Adder_10_U.u1.a  = \add_36s_36s_36_2_1_U12.top_add_36s_36s_36_2_1_Adder_10_U.a [17:0];
assign \add_36s_36s_36_2_1_U12.top_add_36s_36s_36_2_1_Adder_10_U.u1.b  = \add_36s_36s_36_2_1_U12.top_add_36s_36s_36_2_1_Adder_10_U.b [17:0];
assign \add_36s_36s_36_2_1_U12.top_add_36s_36s_36_2_1_Adder_10_U.u1.cin  = 1'h0;
assign \add_36s_36s_36_2_1_U12.top_add_36s_36s_36_2_1_Adder_10_U.facout_s1  = \add_36s_36s_36_2_1_U12.top_add_36s_36s_36_2_1_Adder_10_U.u1.cout ;
assign \add_36s_36s_36_2_1_U12.top_add_36s_36s_36_2_1_Adder_10_U.fas_s1  = \add_36s_36s_36_2_1_U12.top_add_36s_36s_36_2_1_Adder_10_U.u1.s ;
assign \add_36s_36s_36_2_1_U12.top_add_36s_36s_36_2_1_Adder_10_U.a  = \add_36s_36s_36_2_1_U12.din0 ;
assign \add_36s_36s_36_2_1_U12.top_add_36s_36s_36_2_1_Adder_10_U.b  = \add_36s_36s_36_2_1_U12.din1 ;
assign \add_36s_36s_36_2_1_U12.top_add_36s_36s_36_2_1_Adder_10_U.ce  = \add_36s_36s_36_2_1_U12.ce ;
assign \add_36s_36s_36_2_1_U12.top_add_36s_36s_36_2_1_Adder_10_U.clk  = \add_36s_36s_36_2_1_U12.clk ;
assign \add_36s_36s_36_2_1_U12.top_add_36s_36s_36_2_1_Adder_10_U.reset  = \add_36s_36s_36_2_1_U12.reset ;
assign \add_36s_36s_36_2_1_U12.dout  = \add_36s_36s_36_2_1_U12.top_add_36s_36s_36_2_1_Adder_10_U.s ;
assign \add_36s_36s_36_2_1_U12.ce  = 1'h1;
assign \add_36s_36s_36_2_1_U12.clk  = ap_clk;
assign \add_36s_36s_36_2_1_U12.din0  = { op_24_V_reg_1419[31], op_24_V_reg_1419, 3'h0 };
assign \add_36s_36s_36_2_1_U12.din1  = { op_14_V_reg_1414[3], op_14_V_reg_1414[3], op_14_V_reg_1414[3], op_14_V_reg_1414[3], op_14_V_reg_1414[3], op_14_V_reg_1414[3], op_14_V_reg_1414[3], op_14_V_reg_1414[3], op_14_V_reg_1414[3], op_14_V_reg_1414[3], op_14_V_reg_1414[3], op_14_V_reg_1414[3], op_14_V_reg_1414[3], op_14_V_reg_1414[3], op_14_V_reg_1414[3], op_14_V_reg_1414[3], op_14_V_reg_1414[3], op_14_V_reg_1414[3], op_14_V_reg_1414[3], op_14_V_reg_1414[3], op_14_V_reg_1414[3], op_14_V_reg_1414[3], op_14_V_reg_1414[3], op_14_V_reg_1414[3], op_14_V_reg_1414[3], op_14_V_reg_1414[3], op_14_V_reg_1414[3], op_14_V_reg_1414[3], op_14_V_reg_1414[3], op_14_V_reg_1414[3], op_14_V_reg_1414[3], op_14_V_reg_1414[3], op_14_V_reg_1414 };
assign grp_fu_899_p2 = \add_36s_36s_36_2_1_U12.dout ;
assign \add_36s_36s_36_2_1_U12.reset  = ap_rst;
assign \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_13_U.ain_s0  = \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_13_U.a ;
assign \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_13_U.bin_s0  = \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_13_U.b ;
assign \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_13_U.s  = { \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_13_U.fas_s2 , \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_13_U.sum_s1  };
assign \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_13_U.u2.a  = \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_13_U.ain_s1 ;
assign \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_13_U.u2.b  = \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_13_U.bin_s1 ;
assign \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_13_U.u2.cin  = \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_13_U.carry_s1 ;
assign \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_13_U.facout_s2  = \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_13_U.u2.cout ;
assign \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_13_U.fas_s2  = \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_13_U.u2.s ;
assign \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_13_U.u1.a  = \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_13_U.a [16:0];
assign \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_13_U.u1.b  = \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_13_U.b [16:0];
assign \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_13_U.u1.cin  = 1'h0;
assign \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_13_U.facout_s1  = \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_13_U.u1.cout ;
assign \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_13_U.fas_s1  = \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_13_U.u1.s ;
assign \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_13_U.a  = \add_34s_34s_34_2_1_U18.din0 ;
assign \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_13_U.b  = \add_34s_34s_34_2_1_U18.din1 ;
assign \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_13_U.ce  = \add_34s_34s_34_2_1_U18.ce ;
assign \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_13_U.clk  = \add_34s_34s_34_2_1_U18.clk ;
assign \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_13_U.reset  = \add_34s_34s_34_2_1_U18.reset ;
assign \add_34s_34s_34_2_1_U18.dout  = \add_34s_34s_34_2_1_U18.top_add_34s_34s_34_2_1_Adder_13_U.s ;
assign \add_34s_34s_34_2_1_U18.ce  = 1'h1;
assign \add_34s_34s_34_2_1_U18.clk  = ap_clk;
assign \add_34s_34s_34_2_1_U18.din0  = { op_28_V_reg_1518[31], op_28_V_reg_1518, 1'h0 };
assign \add_34s_34s_34_2_1_U18.din1  = { op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18[1], op_18 };
assign grp_fu_1037_p2 = \add_34s_34s_34_2_1_U18.dout ;
assign \add_34s_34s_34_2_1_U18.reset  = ap_rst;
assign \add_33ns_33s_33_2_1_U3.top_add_33ns_33s_33_2_1_Adder_2_U.ain_s0  = \add_33ns_33s_33_2_1_U3.top_add_33ns_33s_33_2_1_Adder_2_U.a ;
assign \add_33ns_33s_33_2_1_U3.top_add_33ns_33s_33_2_1_Adder_2_U.bin_s0  = \add_33ns_33s_33_2_1_U3.top_add_33ns_33s_33_2_1_Adder_2_U.b ;
assign \add_33ns_33s_33_2_1_U3.top_add_33ns_33s_33_2_1_Adder_2_U.s  = { \add_33ns_33s_33_2_1_U3.top_add_33ns_33s_33_2_1_Adder_2_U.fas_s2 , \add_33ns_33s_33_2_1_U3.top_add_33ns_33s_33_2_1_Adder_2_U.sum_s1  };
assign \add_33ns_33s_33_2_1_U3.top_add_33ns_33s_33_2_1_Adder_2_U.u2.a  = \add_33ns_33s_33_2_1_U3.top_add_33ns_33s_33_2_1_Adder_2_U.ain_s1 ;
assign \add_33ns_33s_33_2_1_U3.top_add_33ns_33s_33_2_1_Adder_2_U.u2.b  = \add_33ns_33s_33_2_1_U3.top_add_33ns_33s_33_2_1_Adder_2_U.bin_s1 ;
assign \add_33ns_33s_33_2_1_U3.top_add_33ns_33s_33_2_1_Adder_2_U.u2.cin  = \add_33ns_33s_33_2_1_U3.top_add_33ns_33s_33_2_1_Adder_2_U.carry_s1 ;
assign \add_33ns_33s_33_2_1_U3.top_add_33ns_33s_33_2_1_Adder_2_U.facout_s2  = \add_33ns_33s_33_2_1_U3.top_add_33ns_33s_33_2_1_Adder_2_U.u2.cout ;
assign \add_33ns_33s_33_2_1_U3.top_add_33ns_33s_33_2_1_Adder_2_U.fas_s2  = \add_33ns_33s_33_2_1_U3.top_add_33ns_33s_33_2_1_Adder_2_U.u2.s ;
assign \add_33ns_33s_33_2_1_U3.top_add_33ns_33s_33_2_1_Adder_2_U.u1.a  = \add_33ns_33s_33_2_1_U3.top_add_33ns_33s_33_2_1_Adder_2_U.a [15:0];
assign \add_33ns_33s_33_2_1_U3.top_add_33ns_33s_33_2_1_Adder_2_U.u1.b  = \add_33ns_33s_33_2_1_U3.top_add_33ns_33s_33_2_1_Adder_2_U.b [15:0];
assign \add_33ns_33s_33_2_1_U3.top_add_33ns_33s_33_2_1_Adder_2_U.u1.cin  = 1'h0;
assign \add_33ns_33s_33_2_1_U3.top_add_33ns_33s_33_2_1_Adder_2_U.facout_s1  = \add_33ns_33s_33_2_1_U3.top_add_33ns_33s_33_2_1_Adder_2_U.u1.cout ;
assign \add_33ns_33s_33_2_1_U3.top_add_33ns_33s_33_2_1_Adder_2_U.fas_s1  = \add_33ns_33s_33_2_1_U3.top_add_33ns_33s_33_2_1_Adder_2_U.u1.s ;
assign \add_33ns_33s_33_2_1_U3.top_add_33ns_33s_33_2_1_Adder_2_U.a  = \add_33ns_33s_33_2_1_U3.din0 ;
assign \add_33ns_33s_33_2_1_U3.top_add_33ns_33s_33_2_1_Adder_2_U.b  = \add_33ns_33s_33_2_1_U3.din1 ;
assign \add_33ns_33s_33_2_1_U3.top_add_33ns_33s_33_2_1_Adder_2_U.ce  = \add_33ns_33s_33_2_1_U3.ce ;
assign \add_33ns_33s_33_2_1_U3.top_add_33ns_33s_33_2_1_Adder_2_U.clk  = \add_33ns_33s_33_2_1_U3.clk ;
assign \add_33ns_33s_33_2_1_U3.top_add_33ns_33s_33_2_1_Adder_2_U.reset  = \add_33ns_33s_33_2_1_U3.reset ;
assign \add_33ns_33s_33_2_1_U3.dout  = \add_33ns_33s_33_2_1_U3.top_add_33ns_33s_33_2_1_Adder_2_U.s ;
assign \add_33ns_33s_33_2_1_U3.ce  = 1'h1;
assign \add_33ns_33s_33_2_1_U3.clk  = ap_clk;
assign \add_33ns_33s_33_2_1_U3.din0  = { 8'h00, op_0, 17'h00000 };
assign \add_33ns_33s_33_2_1_U3.din1  = { op_7[31], op_7 };
assign grp_fu_460_p2 = \add_33ns_33s_33_2_1_U3.dout ;
assign \add_33ns_33s_33_2_1_U3.reset  = ap_rst;
assign \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_9_U.ain_s0  = \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_9_U.a ;
assign \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_9_U.bin_s0  = \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_9_U.b ;
assign \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_9_U.s  = { \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_9_U.fas_s2 , \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_9_U.sum_s1  };
assign \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_9_U.u2.a  = \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_9_U.ain_s1 ;
assign \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_9_U.u2.b  = \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_9_U.bin_s1 ;
assign \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_9_U.u2.cin  = \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_9_U.carry_s1 ;
assign \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_9_U.facout_s2  = \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_9_U.u2.cout ;
assign \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_9_U.fas_s2  = \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_9_U.u2.s ;
assign \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_9_U.u1.a  = \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_9_U.a [15:0];
assign \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_9_U.u1.b  = \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_9_U.b [15:0];
assign \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_9_U.u1.cin  = 1'h0;
assign \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_9_U.facout_s1  = \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_9_U.u1.cout ;
assign \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_9_U.fas_s1  = \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_9_U.u1.s ;
assign \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_9_U.a  = \add_32s_32ns_32_2_1_U11.din0 ;
assign \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_9_U.b  = \add_32s_32ns_32_2_1_U11.din1 ;
assign \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_9_U.ce  = \add_32s_32ns_32_2_1_U11.ce ;
assign \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_9_U.clk  = \add_32s_32ns_32_2_1_U11.clk ;
assign \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_9_U.reset  = \add_32s_32ns_32_2_1_U11.reset ;
assign \add_32s_32ns_32_2_1_U11.dout  = \add_32s_32ns_32_2_1_U11.top_add_32s_32ns_32_2_1_Adder_9_U.s ;
assign \add_32s_32ns_32_2_1_U11.ce  = 1'h1;
assign \add_32s_32ns_32_2_1_U11.clk  = ap_clk;
assign \add_32s_32ns_32_2_1_U11.din0  = { ret_V_19_reg_1393[17], ret_V_19_reg_1393[17], ret_V_19_reg_1393[17], ret_V_19_reg_1393[17], ret_V_19_reg_1393[17], ret_V_19_reg_1393[17], ret_V_19_reg_1393[17], ret_V_19_reg_1393[17], ret_V_19_reg_1393[17], ret_V_19_reg_1393[17], ret_V_19_reg_1393[17], ret_V_19_reg_1393[17], ret_V_19_reg_1393[17], ret_V_19_reg_1393[17], ret_V_19_reg_1393 };
assign \add_32s_32ns_32_2_1_U11.din1  = op_13;
assign grp_fu_827_p2 = \add_32s_32ns_32_2_1_U11.dout ;
assign \add_32s_32ns_32_2_1_U11.reset  = ap_rst;
assign \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.ain_s0  = \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.a ;
assign \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.bin_s0  = \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.b ;
assign \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.s  = { \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.fas_s2 , \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.sum_s1  };
assign \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.a  = \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.ain_s1 ;
assign \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.b  = \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.bin_s1 ;
assign \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.cin  = \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.carry_s1 ;
assign \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.facout_s2  = \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.cout ;
assign \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.fas_s2  = \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.s ;
assign \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.a  = \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.a [15:0];
assign \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.b  = \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.b [15:0];
assign \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.cin  = 1'h0;
assign \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.facout_s1  = \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.cout ;
assign \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.fas_s1  = \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.s ;
assign \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.a  = \add_32ns_32ns_32_2_1_U20.din0 ;
assign \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.b  = \add_32ns_32ns_32_2_1_U20.din1 ;
assign \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.ce  = \add_32ns_32ns_32_2_1_U20.ce ;
assign \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.clk  = \add_32ns_32ns_32_2_1_U20.clk ;
assign \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.reset  = \add_32ns_32ns_32_2_1_U20.reset ;
assign \add_32ns_32ns_32_2_1_U20.dout  = \add_32ns_32ns_32_2_1_U20.top_add_32ns_32ns_32_2_1_Adder_11_U.s ;
assign \add_32ns_32ns_32_2_1_U20.ce  = 1'h1;
assign \add_32ns_32ns_32_2_1_U20.clk  = ap_clk;
assign \add_32ns_32ns_32_2_1_U20.din0  = ret_V_24_reg_1555;
assign \add_32ns_32ns_32_2_1_U20.din1  = select_ln1192_reg_1560;
assign grp_fu_1089_p2 = \add_32ns_32ns_32_2_1_U20.dout ;
assign \add_32ns_32ns_32_2_1_U20.reset  = ap_rst;
assign \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.ain_s0  = \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.a ;
assign \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.bin_s0  = \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.b ;
assign \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.s  = { \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.fas_s2 , \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.sum_s1  };
assign \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.a  = \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.ain_s1 ;
assign \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.b  = \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.bin_s1 ;
assign \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.cin  = \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.carry_s1 ;
assign \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.facout_s2  = \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.cout ;
assign \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.fas_s2  = \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.s ;
assign \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.a  = \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.a [15:0];
assign \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.b  = \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.b [15:0];
assign \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.cin  = 1'h0;
assign \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.facout_s1  = \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.cout ;
assign \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.fas_s1  = \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.s ;
assign \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.a  = \add_32ns_32ns_32_2_1_U19.din0 ;
assign \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.b  = \add_32ns_32ns_32_2_1_U19.din1 ;
assign \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.ce  = \add_32ns_32ns_32_2_1_U19.ce ;
assign \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.clk  = \add_32ns_32ns_32_2_1_U19.clk ;
assign \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.reset  = \add_32ns_32ns_32_2_1_U19.reset ;
assign \add_32ns_32ns_32_2_1_U19.dout  = \add_32ns_32ns_32_2_1_U19.top_add_32ns_32ns_32_2_1_Adder_11_U.s ;
assign \add_32ns_32ns_32_2_1_U19.ce  = 1'h1;
assign \add_32ns_32ns_32_2_1_U19.clk  = ap_clk;
assign \add_32ns_32ns_32_2_1_U19.din0  = ret_V_27_cast_reg_1543;
assign \add_32ns_32ns_32_2_1_U19.din1  = 32'd1;
assign grp_fu_1053_p2 = \add_32ns_32ns_32_2_1_U19.dout ;
assign \add_32ns_32ns_32_2_1_U19.reset  = ap_rst;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.ain_s0  = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.a ;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.bin_s0  = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.b ;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.s  = { \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.fas_s2 , \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.sum_s1  };
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.a  = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.ain_s1 ;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.b  = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.bin_s1 ;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.cin  = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.carry_s1 ;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.facout_s2  = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.cout ;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.fas_s2  = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.s ;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.a  = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.a [15:0];
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.b  = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.b [15:0];
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.cin  = 1'h0;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.facout_s1  = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.cout ;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.fas_s1  = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.s ;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.a  = \add_32ns_32ns_32_2_1_U17.din0 ;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.b  = \add_32ns_32ns_32_2_1_U17.din1 ;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.ce  = \add_32ns_32ns_32_2_1_U17.ce ;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.clk  = \add_32ns_32ns_32_2_1_U17.clk ;
assign \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.reset  = \add_32ns_32ns_32_2_1_U17.reset ;
assign \add_32ns_32ns_32_2_1_U17.dout  = \add_32ns_32ns_32_2_1_U17.top_add_32ns_32ns_32_2_1_Adder_11_U.s ;
assign \add_32ns_32ns_32_2_1_U17.ce  = 1'h1;
assign \add_32ns_32ns_32_2_1_U17.clk  = ap_clk;
assign \add_32ns_32ns_32_2_1_U17.din0  = add_ln69_reg_1513;
assign \add_32ns_32ns_32_2_1_U17.din1  = ret_V_22_reg_1508;
assign grp_fu_1018_p2 = \add_32ns_32ns_32_2_1_U17.dout ;
assign \add_32ns_32ns_32_2_1_U17.reset  = ap_rst;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.ain_s0  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.a ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.bin_s0  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.b ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.s  = { \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.fas_s2 , \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.sum_s1  };
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.a  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.ain_s1 ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.b  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.bin_s1 ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.cin  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.carry_s1 ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.facout_s2  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.cout ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.fas_s2  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.s ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.a  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.a [15:0];
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.b  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.b [15:0];
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.cin  = 1'h0;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.facout_s1  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.cout ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.fas_s1  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.s ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.a  = \add_32ns_32ns_32_2_1_U16.din0 ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.b  = \add_32ns_32ns_32_2_1_U16.din1 ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.ce  = \add_32ns_32ns_32_2_1_U16.ce ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.clk  = \add_32ns_32ns_32_2_1_U16.clk ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.reset  = \add_32ns_32ns_32_2_1_U16.reset ;
assign \add_32ns_32ns_32_2_1_U16.dout  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.s ;
assign \add_32ns_32ns_32_2_1_U16.ce  = 1'h1;
assign \add_32ns_32ns_32_2_1_U16.clk  = ap_clk;
assign \add_32ns_32ns_32_2_1_U16.din0  = { 31'h00000000, icmp_ln1499_reg_1306 };
assign \add_32ns_32ns_32_2_1_U16.din1  = op_16;
assign grp_fu_993_p2 = \add_32ns_32ns_32_2_1_U16.dout ;
assign \add_32ns_32ns_32_2_1_U16.reset  = ap_rst;
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.ain_s0  = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.a ;
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.bin_s0  = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.b ;
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.s  = { \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.fas_s2 , \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.sum_s1  };
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.a  = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.ain_s1 ;
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.b  = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.bin_s1 ;
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.cin  = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.carry_s1 ;
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.facout_s2  = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.cout ;
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.fas_s2  = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.s ;
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.a  = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.a [15:0];
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.b  = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.b [15:0];
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.cin  = 1'h0;
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.facout_s1  = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.cout ;
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.fas_s1  = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.s ;
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.a  = \add_32ns_32ns_32_2_1_U15.din0 ;
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.b  = \add_32ns_32ns_32_2_1_U15.din1 ;
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.ce  = \add_32ns_32ns_32_2_1_U15.ce ;
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.clk  = \add_32ns_32ns_32_2_1_U15.clk ;
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.reset  = \add_32ns_32ns_32_2_1_U15.reset ;
assign \add_32ns_32ns_32_2_1_U15.dout  = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.s ;
assign \add_32ns_32ns_32_2_1_U15.ce  = 1'h1;
assign \add_32ns_32ns_32_2_1_U15.clk  = ap_clk;
assign \add_32ns_32ns_32_2_1_U15.din0  = ret_V_25_cast_reg_1486;
assign \add_32ns_32ns_32_2_1_U15.din1  = 32'd1;
assign grp_fu_985_p2 = \add_32ns_32ns_32_2_1_U15.dout ;
assign \add_32ns_32ns_32_2_1_U15.reset  = ap_rst;
assign \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_11_U.ain_s0  = \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_11_U.a ;
assign \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_11_U.bin_s0  = \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_11_U.b ;
assign \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_11_U.s  = { \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_11_U.fas_s2 , \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_11_U.sum_s1  };
assign \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.a  = \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_11_U.ain_s1 ;
assign \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.b  = \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_11_U.bin_s1 ;
assign \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.cin  = \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_11_U.carry_s1 ;
assign \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_11_U.facout_s2  = \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.cout ;
assign \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_11_U.fas_s2  = \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.s ;
assign \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.a  = \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_11_U.a [15:0];
assign \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.b  = \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_11_U.b [15:0];
assign \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.cin  = 1'h0;
assign \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_11_U.facout_s1  = \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.cout ;
assign \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_11_U.fas_s1  = \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.s ;
assign \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_11_U.a  = \add_32ns_32ns_32_2_1_U13.din0 ;
assign \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_11_U.b  = \add_32ns_32ns_32_2_1_U13.din1 ;
assign \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_11_U.ce  = \add_32ns_32ns_32_2_1_U13.ce ;
assign \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_11_U.clk  = \add_32ns_32ns_32_2_1_U13.clk ;
assign \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_11_U.reset  = \add_32ns_32ns_32_2_1_U13.reset ;
assign \add_32ns_32ns_32_2_1_U13.dout  = \add_32ns_32ns_32_2_1_U13.top_add_32ns_32ns_32_2_1_Adder_11_U.s ;
assign \add_32ns_32ns_32_2_1_U13.ce  = 1'h1;
assign \add_32ns_32ns_32_2_1_U13.clk  = ap_clk;
assign \add_32ns_32ns_32_2_1_U13.din0  = ret_V_23_cast_reg_1449;
assign \add_32ns_32ns_32_2_1_U13.din1  = 32'd1;
assign grp_fu_920_p2 = \add_32ns_32ns_32_2_1_U13.dout ;
assign \add_32ns_32ns_32_2_1_U13.reset  = ap_rst;
assign \add_18s_18ns_18_2_1_U8.top_add_18s_18ns_18_2_1_Adder_7_U.ain_s0  = \add_18s_18ns_18_2_1_U8.top_add_18s_18ns_18_2_1_Adder_7_U.a ;
assign \add_18s_18ns_18_2_1_U8.top_add_18s_18ns_18_2_1_Adder_7_U.bin_s0  = \add_18s_18ns_18_2_1_U8.top_add_18s_18ns_18_2_1_Adder_7_U.b ;
assign \add_18s_18ns_18_2_1_U8.top_add_18s_18ns_18_2_1_Adder_7_U.s  = { \add_18s_18ns_18_2_1_U8.top_add_18s_18ns_18_2_1_Adder_7_U.fas_s2 , \add_18s_18ns_18_2_1_U8.top_add_18s_18ns_18_2_1_Adder_7_U.sum_s1  };
assign \add_18s_18ns_18_2_1_U8.top_add_18s_18ns_18_2_1_Adder_7_U.u2.a  = \add_18s_18ns_18_2_1_U8.top_add_18s_18ns_18_2_1_Adder_7_U.ain_s1 ;
assign \add_18s_18ns_18_2_1_U8.top_add_18s_18ns_18_2_1_Adder_7_U.u2.b  = \add_18s_18ns_18_2_1_U8.top_add_18s_18ns_18_2_1_Adder_7_U.bin_s1 ;
assign \add_18s_18ns_18_2_1_U8.top_add_18s_18ns_18_2_1_Adder_7_U.u2.cin  = \add_18s_18ns_18_2_1_U8.top_add_18s_18ns_18_2_1_Adder_7_U.carry_s1 ;
assign \add_18s_18ns_18_2_1_U8.top_add_18s_18ns_18_2_1_Adder_7_U.facout_s2  = \add_18s_18ns_18_2_1_U8.top_add_18s_18ns_18_2_1_Adder_7_U.u2.cout ;
assign \add_18s_18ns_18_2_1_U8.top_add_18s_18ns_18_2_1_Adder_7_U.fas_s2  = \add_18s_18ns_18_2_1_U8.top_add_18s_18ns_18_2_1_Adder_7_U.u2.s ;
assign \add_18s_18ns_18_2_1_U8.top_add_18s_18ns_18_2_1_Adder_7_U.u1.a  = \add_18s_18ns_18_2_1_U8.top_add_18s_18ns_18_2_1_Adder_7_U.a [8:0];
assign \add_18s_18ns_18_2_1_U8.top_add_18s_18ns_18_2_1_Adder_7_U.u1.b  = \add_18s_18ns_18_2_1_U8.top_add_18s_18ns_18_2_1_Adder_7_U.b [8:0];
assign \add_18s_18ns_18_2_1_U8.top_add_18s_18ns_18_2_1_Adder_7_U.u1.cin  = 1'h0;
assign \add_18s_18ns_18_2_1_U8.top_add_18s_18ns_18_2_1_Adder_7_U.facout_s1  = \add_18s_18ns_18_2_1_U8.top_add_18s_18ns_18_2_1_Adder_7_U.u1.cout ;
assign \add_18s_18ns_18_2_1_U8.top_add_18s_18ns_18_2_1_Adder_7_U.fas_s1  = \add_18s_18ns_18_2_1_U8.top_add_18s_18ns_18_2_1_Adder_7_U.u1.s ;
assign \add_18s_18ns_18_2_1_U8.top_add_18s_18ns_18_2_1_Adder_7_U.a  = \add_18s_18ns_18_2_1_U8.din0 ;
assign \add_18s_18ns_18_2_1_U8.top_add_18s_18ns_18_2_1_Adder_7_U.b  = \add_18s_18ns_18_2_1_U8.din1 ;
assign \add_18s_18ns_18_2_1_U8.top_add_18s_18ns_18_2_1_Adder_7_U.ce  = \add_18s_18ns_18_2_1_U8.ce ;
assign \add_18s_18ns_18_2_1_U8.top_add_18s_18ns_18_2_1_Adder_7_U.clk  = \add_18s_18ns_18_2_1_U8.clk ;
assign \add_18s_18ns_18_2_1_U8.top_add_18s_18ns_18_2_1_Adder_7_U.reset  = \add_18s_18ns_18_2_1_U8.reset ;
assign \add_18s_18ns_18_2_1_U8.dout  = \add_18s_18ns_18_2_1_U8.top_add_18s_18ns_18_2_1_Adder_7_U.s ;
assign \add_18s_18ns_18_2_1_U8.ce  = 1'h1;
assign \add_18s_18ns_18_2_1_U8.clk  = ap_clk;
assign \add_18s_18ns_18_2_1_U8.din0  = { tmp_6_reg_1356[16], tmp_6_reg_1356 };
assign \add_18s_18ns_18_2_1_U8.din1  = 18'h00001;
assign grp_fu_766_p2 = \add_18s_18ns_18_2_1_U8.dout ;
assign \add_18s_18ns_18_2_1_U8.reset  = ap_rst;
assign \add_18ns_18s_18_2_1_U9.top_add_18ns_18s_18_2_1_Adder_8_U.ain_s0  = \add_18ns_18s_18_2_1_U9.top_add_18ns_18s_18_2_1_Adder_8_U.a ;
assign \add_18ns_18s_18_2_1_U9.top_add_18ns_18s_18_2_1_Adder_8_U.bin_s0  = \add_18ns_18s_18_2_1_U9.top_add_18ns_18s_18_2_1_Adder_8_U.b ;
assign \add_18ns_18s_18_2_1_U9.top_add_18ns_18s_18_2_1_Adder_8_U.s  = { \add_18ns_18s_18_2_1_U9.top_add_18ns_18s_18_2_1_Adder_8_U.fas_s2 , \add_18ns_18s_18_2_1_U9.top_add_18ns_18s_18_2_1_Adder_8_U.sum_s1  };
assign \add_18ns_18s_18_2_1_U9.top_add_18ns_18s_18_2_1_Adder_8_U.u2.a  = \add_18ns_18s_18_2_1_U9.top_add_18ns_18s_18_2_1_Adder_8_U.ain_s1 ;
assign \add_18ns_18s_18_2_1_U9.top_add_18ns_18s_18_2_1_Adder_8_U.u2.b  = \add_18ns_18s_18_2_1_U9.top_add_18ns_18s_18_2_1_Adder_8_U.bin_s1 ;
assign \add_18ns_18s_18_2_1_U9.top_add_18ns_18s_18_2_1_Adder_8_U.u2.cin  = \add_18ns_18s_18_2_1_U9.top_add_18ns_18s_18_2_1_Adder_8_U.carry_s1 ;
assign \add_18ns_18s_18_2_1_U9.top_add_18ns_18s_18_2_1_Adder_8_U.facout_s2  = \add_18ns_18s_18_2_1_U9.top_add_18ns_18s_18_2_1_Adder_8_U.u2.cout ;
assign \add_18ns_18s_18_2_1_U9.top_add_18ns_18s_18_2_1_Adder_8_U.fas_s2  = \add_18ns_18s_18_2_1_U9.top_add_18ns_18s_18_2_1_Adder_8_U.u2.s ;
assign \add_18ns_18s_18_2_1_U9.top_add_18ns_18s_18_2_1_Adder_8_U.u1.a  = \add_18ns_18s_18_2_1_U9.top_add_18ns_18s_18_2_1_Adder_8_U.a [8:0];
assign \add_18ns_18s_18_2_1_U9.top_add_18ns_18s_18_2_1_Adder_8_U.u1.b  = \add_18ns_18s_18_2_1_U9.top_add_18ns_18s_18_2_1_Adder_8_U.b [8:0];
assign \add_18ns_18s_18_2_1_U9.top_add_18ns_18s_18_2_1_Adder_8_U.u1.cin  = 1'h0;
assign \add_18ns_18s_18_2_1_U9.top_add_18ns_18s_18_2_1_Adder_8_U.facout_s1  = \add_18ns_18s_18_2_1_U9.top_add_18ns_18s_18_2_1_Adder_8_U.u1.cout ;
assign \add_18ns_18s_18_2_1_U9.top_add_18ns_18s_18_2_1_Adder_8_U.fas_s1  = \add_18ns_18s_18_2_1_U9.top_add_18ns_18s_18_2_1_Adder_8_U.u1.s ;
assign \add_18ns_18s_18_2_1_U9.top_add_18ns_18s_18_2_1_Adder_8_U.a  = \add_18ns_18s_18_2_1_U9.din0 ;
assign \add_18ns_18s_18_2_1_U9.top_add_18ns_18s_18_2_1_Adder_8_U.b  = \add_18ns_18s_18_2_1_U9.din1 ;
assign \add_18ns_18s_18_2_1_U9.top_add_18ns_18s_18_2_1_Adder_8_U.ce  = \add_18ns_18s_18_2_1_U9.ce ;
assign \add_18ns_18s_18_2_1_U9.top_add_18ns_18s_18_2_1_Adder_8_U.clk  = \add_18ns_18s_18_2_1_U9.clk ;
assign \add_18ns_18s_18_2_1_U9.top_add_18ns_18s_18_2_1_Adder_8_U.reset  = \add_18ns_18s_18_2_1_U9.reset ;
assign \add_18ns_18s_18_2_1_U9.dout  = \add_18ns_18s_18_2_1_U9.top_add_18ns_18s_18_2_1_Adder_8_U.s ;
assign \add_18ns_18s_18_2_1_U9.ce  = 1'h1;
assign \add_18ns_18s_18_2_1_U9.clk  = ap_clk;
assign \add_18ns_18s_18_2_1_U9.din0  = ret_V_18_reg_1373;
assign \add_18ns_18s_18_2_1_U9.din1  = { ret_V_15_reg_1346[7], ret_V_15_reg_1346[7], ret_V_15_reg_1346[7], ret_V_15_reg_1346[7], ret_V_15_reg_1346[7], ret_V_15_reg_1346[7], ret_V_15_reg_1346[7], ret_V_15_reg_1346[7], ret_V_15_reg_1346[7], ret_V_15_reg_1346[7], ret_V_15_reg_1346 };
assign grp_fu_794_p2 = \add_18ns_18s_18_2_1_U9.dout ;
assign \add_18ns_18s_18_2_1_U9.reset  = ap_rst;
assign \add_18ns_18s_18_2_1_U10.top_add_18ns_18s_18_2_1_Adder_8_U.ain_s0  = \add_18ns_18s_18_2_1_U10.top_add_18ns_18s_18_2_1_Adder_8_U.a ;
assign \add_18ns_18s_18_2_1_U10.top_add_18ns_18s_18_2_1_Adder_8_U.bin_s0  = \add_18ns_18s_18_2_1_U10.top_add_18ns_18s_18_2_1_Adder_8_U.b ;
assign \add_18ns_18s_18_2_1_U10.top_add_18ns_18s_18_2_1_Adder_8_U.s  = { \add_18ns_18s_18_2_1_U10.top_add_18ns_18s_18_2_1_Adder_8_U.fas_s2 , \add_18ns_18s_18_2_1_U10.top_add_18ns_18s_18_2_1_Adder_8_U.sum_s1  };
assign \add_18ns_18s_18_2_1_U10.top_add_18ns_18s_18_2_1_Adder_8_U.u2.a  = \add_18ns_18s_18_2_1_U10.top_add_18ns_18s_18_2_1_Adder_8_U.ain_s1 ;
assign \add_18ns_18s_18_2_1_U10.top_add_18ns_18s_18_2_1_Adder_8_U.u2.b  = \add_18ns_18s_18_2_1_U10.top_add_18ns_18s_18_2_1_Adder_8_U.bin_s1 ;
assign \add_18ns_18s_18_2_1_U10.top_add_18ns_18s_18_2_1_Adder_8_U.u2.cin  = \add_18ns_18s_18_2_1_U10.top_add_18ns_18s_18_2_1_Adder_8_U.carry_s1 ;
assign \add_18ns_18s_18_2_1_U10.top_add_18ns_18s_18_2_1_Adder_8_U.facout_s2  = \add_18ns_18s_18_2_1_U10.top_add_18ns_18s_18_2_1_Adder_8_U.u2.cout ;
assign \add_18ns_18s_18_2_1_U10.top_add_18ns_18s_18_2_1_Adder_8_U.fas_s2  = \add_18ns_18s_18_2_1_U10.top_add_18ns_18s_18_2_1_Adder_8_U.u2.s ;
assign \add_18ns_18s_18_2_1_U10.top_add_18ns_18s_18_2_1_Adder_8_U.u1.a  = \add_18ns_18s_18_2_1_U10.top_add_18ns_18s_18_2_1_Adder_8_U.a [8:0];
assign \add_18ns_18s_18_2_1_U10.top_add_18ns_18s_18_2_1_Adder_8_U.u1.b  = \add_18ns_18s_18_2_1_U10.top_add_18ns_18s_18_2_1_Adder_8_U.b [8:0];
assign \add_18ns_18s_18_2_1_U10.top_add_18ns_18s_18_2_1_Adder_8_U.u1.cin  = 1'h0;
assign \add_18ns_18s_18_2_1_U10.top_add_18ns_18s_18_2_1_Adder_8_U.facout_s1  = \add_18ns_18s_18_2_1_U10.top_add_18ns_18s_18_2_1_Adder_8_U.u1.cout ;
assign \add_18ns_18s_18_2_1_U10.top_add_18ns_18s_18_2_1_Adder_8_U.fas_s1  = \add_18ns_18s_18_2_1_U10.top_add_18ns_18s_18_2_1_Adder_8_U.u1.s ;
assign \add_18ns_18s_18_2_1_U10.top_add_18ns_18s_18_2_1_Adder_8_U.a  = \add_18ns_18s_18_2_1_U10.din0 ;
assign \add_18ns_18s_18_2_1_U10.top_add_18ns_18s_18_2_1_Adder_8_U.b  = \add_18ns_18s_18_2_1_U10.din1 ;
assign \add_18ns_18s_18_2_1_U10.top_add_18ns_18s_18_2_1_Adder_8_U.ce  = \add_18ns_18s_18_2_1_U10.ce ;
assign \add_18ns_18s_18_2_1_U10.top_add_18ns_18s_18_2_1_Adder_8_U.clk  = \add_18ns_18s_18_2_1_U10.clk ;
assign \add_18ns_18s_18_2_1_U10.top_add_18ns_18s_18_2_1_Adder_8_U.reset  = \add_18ns_18s_18_2_1_U10.reset ;
assign \add_18ns_18s_18_2_1_U10.dout  = \add_18ns_18s_18_2_1_U10.top_add_18ns_18s_18_2_1_Adder_8_U.s ;
assign \add_18ns_18s_18_2_1_U10.ce  = 1'h1;
assign \add_18ns_18s_18_2_1_U10.clk  = ap_clk;
assign \add_18ns_18s_18_2_1_U10.din0  = op_22_V_reg_1383;
assign \add_18ns_18s_18_2_1_U10.din1  = { op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12[1], op_12 };
assign grp_fu_803_p2 = \add_18ns_18s_18_2_1_U10.dout ;
assign \add_18ns_18s_18_2_1_U10.reset  = ap_rst;
assign \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_3_U.ain_s0  = \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_3_U.a ;
assign \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_3_U.bin_s0  = \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_3_U.b ;
assign \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_3_U.s  = { \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_3_U.fas_s2 , \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_3_U.sum_s1  };
assign \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_3_U.u2.a  = \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_3_U.ain_s1 ;
assign \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_3_U.u2.b  = \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_3_U.bin_s1 ;
assign \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_3_U.u2.cin  = \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_3_U.carry_s1 ;
assign \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_3_U.facout_s2  = \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_3_U.u2.cout ;
assign \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_3_U.fas_s2  = \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_3_U.u2.s ;
assign \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_3_U.u1.a  = \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_3_U.a [7:0];
assign \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_3_U.u1.b  = \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_3_U.b [7:0];
assign \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_3_U.u1.cin  = 1'h0;
assign \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_3_U.facout_s1  = \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_3_U.u1.cout ;
assign \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_3_U.fas_s1  = \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_3_U.u1.s ;
assign \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_3_U.a  = \add_16ns_16ns_16_2_1_U4.din0 ;
assign \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_3_U.b  = \add_16ns_16ns_16_2_1_U4.din1 ;
assign \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_3_U.ce  = \add_16ns_16ns_16_2_1_U4.ce ;
assign \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_3_U.clk  = \add_16ns_16ns_16_2_1_U4.clk ;
assign \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_3_U.reset  = \add_16ns_16ns_16_2_1_U4.reset ;
assign \add_16ns_16ns_16_2_1_U4.dout  = \add_16ns_16ns_16_2_1_U4.top_add_16ns_16ns_16_2_1_Adder_3_U.s ;
assign \add_16ns_16ns_16_2_1_U4.ce  = 1'h1;
assign \add_16ns_16ns_16_2_1_U4.clk  = ap_clk;
assign \add_16ns_16ns_16_2_1_U4.din0  = ret_V_3_reg_1251;
assign \add_16ns_16ns_16_2_1_U4.din1  = 16'h0001;
assign grp_fu_561_p2 = \add_16ns_16ns_16_2_1_U4.dout ;
assign \add_16ns_16ns_16_2_1_U4.reset  = ap_rst;
endmodule


// Product machine:
module top_A_times_top_B (ap_start, op_0, op_1, op_12, op_13, op_15, op_16, op_18, op_19, op_2, op_5, op_7, ap_clk, unsafe_signal);
input ap_start;
input [7:0] op_0;
input [31:0] op_1;
input [1:0] op_12;
input [31:0] op_13;
input [31:0] op_15;
input [31:0] op_16;
input [1:0] op_18;
input op_19;
input [15:0] op_2;
input [1:0] op_5;
input [31:0] op_7;
input ap_clk;
output unsafe_signal;
reg _setup;
initial _setup = 1'b0;
always @ (posedge ap_clk) _setup <= 1'b1;
reg ap_start_internal;
always @ (posedge ap_clk) if (!_setup) ap_start_internal <= ap_start;
reg [7:0] op_0_internal;
always @ (posedge ap_clk) if (!_setup) op_0_internal <= op_0;
reg [31:0] op_1_internal;
always @ (posedge ap_clk) if (!_setup) op_1_internal <= op_1;
reg [1:0] op_12_internal;
always @ (posedge ap_clk) if (!_setup) op_12_internal <= op_12;
reg [31:0] op_13_internal;
always @ (posedge ap_clk) if (!_setup) op_13_internal <= op_13;
reg [31:0] op_15_internal;
always @ (posedge ap_clk) if (!_setup) op_15_internal <= op_15;
reg [31:0] op_16_internal;
always @ (posedge ap_clk) if (!_setup) op_16_internal <= op_16;
reg [1:0] op_18_internal;
always @ (posedge ap_clk) if (!_setup) op_18_internal <= op_18;
reg op_19_internal;
always @ (posedge ap_clk) if (!_setup) op_19_internal <= op_19;
reg [15:0] op_2_internal;
always @ (posedge ap_clk) if (!_setup) op_2_internal <= op_2;
reg [1:0] op_5_internal;
always @ (posedge ap_clk) if (!_setup) op_5_internal <= op_5;
reg [31:0] op_7_internal;
always @ (posedge ap_clk) if (!_setup) op_7_internal <= op_7;
wire ap_done_A;
wire ap_done_B;
wire ap_done_eq;
assign ap_done_eq = ap_done_A == ap_done_B;
wire ap_idle_A;
wire ap_idle_B;
wire ap_idle_eq;
assign ap_idle_eq = ap_idle_A == ap_idle_B;
wire ap_ready_A;
wire ap_ready_B;
wire ap_ready_eq;
assign ap_ready_eq = ap_ready_A == ap_ready_B;
wire [31:0] op_30_A;
wire [31:0] op_30_B;
wire op_30_eq;
assign op_30_eq = op_30_A == op_30_B;
wire op_30_ap_vld_A;
wire op_30_ap_vld_B;
wire clk_enable_A;
wire clk_enable_B;
assign clk_enable_A = _setup & (~op_30_ap_vld_A | op_30_ap_vld_B);
assign clk_enable_B = _setup;
wire divergent;
assign divergent = ~(ap_done_eq & ap_idle_eq & ap_ready_eq & op_30_eq);
assign unsafe_signal = op_30_ap_vld_A & op_30_ap_vld_B & divergent;
top_A instance_A (
    .ap_clk(ap_clk),
    .clk_enable(clk_enable_A),
    .ap_start(ap_start_internal),
    .op_0(op_0_internal),
    .op_1(op_1_internal),
    .op_12(op_12_internal),
    .op_13(op_13_internal),
    .op_15(op_15_internal),
    .op_16(op_16_internal),
    .op_18(op_18_internal),
    .op_19(op_19_internal),
    .op_2(op_2_internal),
    .op_5(op_5_internal),
    .op_7(op_7_internal),
    .ap_done(ap_done_A),
    .ap_idle(ap_idle_A),
    .ap_ready(ap_ready_A),
    .op_30(op_30_A),
    .op_30_ap_vld(op_30_ap_vld_A)
);
top_B instance_B (
    .ap_clk(ap_clk),
    .clk_enable(clk_enable_B),
    .ap_start(ap_start_internal),
    .op_0(op_0_internal),
    .op_1(op_1_internal),
    .op_12(op_12_internal),
    .op_13(op_13_internal),
    .op_15(op_15_internal),
    .op_16(op_16_internal),
    .op_18(op_18_internal),
    .op_19(op_19_internal),
    .op_2(op_2_internal),
    .op_5(op_5_internal),
    .op_7(op_7_internal),
    .ap_done(ap_done_B),
    .ap_idle(ap_idle_B),
    .ap_ready(ap_ready_B),
    .op_30(op_30_B),
    .op_30_ap_vld(op_30_ap_vld_B)
);
endmodule
