// Processed by function `construct_kairos` in `verilog_tricks.py`.
// Machine A:
// Processed by function `add_clk_enable_signal` in `verilog_tricks.py`.
// Processed by function `remove_reset_signal` in `verilog_tricks.py`.
module top_A (
  ap_clk,
  ap_start,
  ap_done,
  ap_idle,
  ap_ready,
  op_0,
  op_1,
  op_2,
  op_4,
  op_5,
  op_7,
  op_9,
  op_11,
  op_12,
  op_14,
  op_15,
  op_19,
  op_29,
  op_29_ap_vld,
clk_enable
);
input clk_enable;


input ap_clk;
wire ap_rst;
assign ap_rst = op_29_ap_vld;
input ap_start;
input [3:0] op_0;
input [7:0] op_1;
input [1:0] op_11;
input [1:0] op_12;
input [31:0] op_14;
input [15:0] op_15;
input [15:0] op_19;
input [15:0] op_2;
input [7:0] op_4;
input [7:0] op_5;
input [7:0] op_7;
input [1:0] op_9;
output ap_done;
output ap_idle;
output ap_ready;
output [31:0] op_29;
output op_29_ap_vld;


reg [4:0] \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.ain_s1 ;
reg [4:0] \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.bin_s1 ;
reg \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.carry_s1 ;
reg [4:0] \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.sum_s1 ;
reg [8:0] \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.ain_s1 ;
reg [8:0] \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.bin_s1 ;
reg \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.carry_s1 ;
reg [7:0] \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.sum_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.ain_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.bin_s1 ;
reg \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.carry_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.sum_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.ain_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.bin_s1 ;
reg \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.carry_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.sum_s1 ;
reg [15:0] \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.ain_s1 ;
reg [15:0] \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.bin_s1 ;
reg \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.carry_s1 ;
reg [15:0] \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.sum_s1 ;
reg [15:0] \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.ain_s1 ;
reg [15:0] \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.bin_s1 ;
reg \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.carry_s1 ;
reg [15:0] \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.sum_s1 ;
reg [15:0] \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.ain_s1 ;
reg [15:0] \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.bin_s1 ;
reg \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.carry_s1 ;
reg [15:0] \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.sum_s1 ;
reg [15:0] \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.ain_s1 ;
reg [15:0] \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.bin_s1 ;
reg \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.carry_s1 ;
reg [15:0] \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.sum_s1 ;
reg [16:0] \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.ain_s1 ;
reg [16:0] \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.bin_s1 ;
reg \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.carry_s1 ;
reg [16:0] \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.sum_s1 ;
reg [1:0] \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.ain_s1 ;
reg [1:0] \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.bin_s1 ;
reg \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.carry_s1 ;
reg \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.sum_s1 ;
reg [2:0] \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.ain_s1 ;
reg [2:0] \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.bin_s1 ;
reg \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.carry_s1 ;
reg [1:0] \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.sum_s1 ;
reg [2:0] \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.ain_s1 ;
reg [2:0] \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.bin_s1 ;
reg \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.carry_s1 ;
reg [1:0] \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.sum_s1 ;
reg [3:0] \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.ain_s1 ;
reg [3:0] \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.bin_s1 ;
reg \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.carry_s1 ;
reg [2:0] \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.sum_s1 ;
reg [31:0] add_ln691_1_reg_928;
reg [31:0] add_ln691_reg_809;
reg [2:0] add_ln69_1_reg_861;
reg [16:0] add_ln69_3_reg_963;
reg [31:0] add_ln69_reg_856;
reg [23:0] ap_CS_fsm = 24'h000001;
reg [31:0] \ashr_32s_32ns_32_7_1_U10.din1_cast_array[0] ;
reg [31:0] \ashr_32s_32ns_32_7_1_U10.din1_cast_array[1] ;
reg [31:0] \ashr_32s_32ns_32_7_1_U10.din1_cast_array[2] ;
reg [31:0] \ashr_32s_32ns_32_7_1_U10.din1_cast_array[3] ;
reg [31:0] \ashr_32s_32ns_32_7_1_U10.din1_cast_array[4] ;
reg [31:0] \ashr_32s_32ns_32_7_1_U10.din1_cast_array[5] ;
reg [31:0] \ashr_32s_32ns_32_7_1_U10.dout_array[0] ;
reg [31:0] \ashr_32s_32ns_32_7_1_U10.dout_array[1] ;
reg [31:0] \ashr_32s_32ns_32_7_1_U10.dout_array[2] ;
reg [31:0] \ashr_32s_32ns_32_7_1_U10.dout_array[3] ;
reg [31:0] \ashr_32s_32ns_32_7_1_U10.dout_array[4] ;
reg [31:0] \ashr_32s_32ns_32_7_1_U10.dout_array[5] ;
reg icmp_ln768_reg_716;
reg icmp_ln850_reg_804;
reg lhs_V_4_reg_679;
reg newsignbit_reg_673;
reg [3:0] op_16_V_reg_886;
reg [31:0] op_25_V_reg_891;
reg op_6_V_reg_699;
reg [19:0] op_8_V_reg_761;
reg p_Result_3_reg_704;
reg p_Result_4_reg_820;
reg [8:0] p_Result_s_reg_711;
reg [1:0] r_reg_933;
reg [4:0] ret_1_reg_731;
reg [4:0] ret_V_11_reg_741;
reg [6:0] ret_V_12_reg_776;
reg [31:0] ret_V_13_reg_825;
reg [33:0] ret_V_14_reg_906;
reg [31:0] ret_V_15_reg_938;
reg [31:0] ret_V_16_reg_958;
reg [31:0] ret_V_9_cast_reg_911;
reg [27:0] ret_V_9_reg_786;
reg [21:0] ret_V_reg_881;
reg [4:0] select_ln1192_reg_736;
reg [2:0] select_ln69_reg_830;
reg [31:0] sext_ln831_reg_797;
reg [31:0] sh_reg_835;
reg [31:0] \shl_32s_32ns_32_7_1_U11.din1_cast_array[0] ;
reg [31:0] \shl_32s_32ns_32_7_1_U11.din1_cast_array[1] ;
reg [31:0] \shl_32s_32ns_32_7_1_U11.din1_cast_array[2] ;
reg [31:0] \shl_32s_32ns_32_7_1_U11.din1_cast_array[3] ;
reg [31:0] \shl_32s_32ns_32_7_1_U11.din1_cast_array[4] ;
reg [31:0] \shl_32s_32ns_32_7_1_U11.din1_cast_array[5] ;
reg [31:0] \shl_32s_32ns_32_7_1_U11.dout_array[0] ;
reg [31:0] \shl_32s_32ns_32_7_1_U11.dout_array[1] ;
reg [31:0] \shl_32s_32ns_32_7_1_U11.dout_array[2] ;
reg [31:0] \shl_32s_32ns_32_7_1_U11.dout_array[3] ;
reg [31:0] \shl_32s_32ns_32_7_1_U11.dout_array[4] ;
reg [31:0] \shl_32s_32ns_32_7_1_U11.dout_array[5] ;
reg signbit_1_reg_684;
reg [10:0] \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.ain_s1 ;
reg [10:0] \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.bin_s1 ;
reg \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.carry_s1 ;
reg [10:0] \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.sum_s1 ;
reg [13:0] \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.ain_s1 ;
reg [13:0] \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.bin_s1 ;
reg \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.carry_s1 ;
reg [13:0] \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.sum_s1 ;
reg [15:0] \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.ain_s1 ;
reg [15:0] \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.bin_s1 ;
reg \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.carry_s1 ;
reg [15:0] \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.sum_s1 ;
reg [5:0] tmp_2_reg_781;
reg trunc_ln213_reg_658;
reg [2:0] trunc_ln728_reg_689;
reg [1:0] trunc_ln798_1_reg_923;
reg [1:0] trunc_ln798_reg_918;
reg [18:0] trunc_ln851_reg_792;
wire [31:0] _000_;
wire [31:0] _001_;
wire [2:0] _002_;
wire [16:0] _003_;
wire [31:0] _004_;
wire [23:0] _005_;
wire _006_;
wire _007_;
wire _008_;
wire _009_;
wire [3:0] _010_;
wire [31:0] _011_;
wire _012_;
wire _013_;
wire _014_;
wire _015_;
wire [8:0] _016_;
wire [1:0] _017_;
wire [4:0] _018_;
wire [4:0] _019_;
wire [6:0] _020_;
wire [31:0] _021_;
wire [33:0] _022_;
wire [31:0] _023_;
wire [31:0] _024_;
wire [31:0] _025_;
wire [27:0] _026_;
wire [21:0] _027_;
wire [4:0] _028_;
wire [2:0] _029_;
wire [31:0] _030_;
wire [31:0] _031_;
wire _032_;
wire [5:0] _033_;
wire _034_;
wire [2:0] _035_;
wire [1:0] _036_;
wire [1:0] _037_;
wire [18:0] _038_;
wire [1:0] _039_;
wire _040_;
wire _041_;
wire _042_;
wire _043_;
wire _044_;
wire _045_;
wire [4:0] _046_;
wire [4:0] _047_;
wire _048_;
wire [4:0] _049_;
wire [5:0] _050_;
wire [5:0] _051_;
wire [8:0] _052_;
wire [8:0] _053_;
wire _054_;
wire [7:0] _055_;
wire [8:0] _056_;
wire [9:0] _057_;
wire [15:0] _058_;
wire [15:0] _059_;
wire _060_;
wire [15:0] _061_;
wire [16:0] _062_;
wire [16:0] _063_;
wire [15:0] _064_;
wire [15:0] _065_;
wire _066_;
wire [15:0] _067_;
wire [16:0] _068_;
wire [16:0] _069_;
wire [15:0] _070_;
wire [15:0] _071_;
wire _072_;
wire [15:0] _073_;
wire [16:0] _074_;
wire [16:0] _075_;
wire [15:0] _076_;
wire [15:0] _077_;
wire _078_;
wire [15:0] _079_;
wire [16:0] _080_;
wire [16:0] _081_;
wire [15:0] _082_;
wire [15:0] _083_;
wire _084_;
wire [15:0] _085_;
wire [16:0] _086_;
wire [16:0] _087_;
wire [15:0] _088_;
wire [15:0] _089_;
wire _090_;
wire [15:0] _091_;
wire [16:0] _092_;
wire [16:0] _093_;
wire [16:0] _094_;
wire [16:0] _095_;
wire _096_;
wire [16:0] _097_;
wire [17:0] _098_;
wire [17:0] _099_;
wire [1:0] _100_;
wire [1:0] _101_;
wire _102_;
wire _103_;
wire [1:0] _104_;
wire [2:0] _105_;
wire [2:0] _106_;
wire [2:0] _107_;
wire _108_;
wire [1:0] _109_;
wire [2:0] _110_;
wire [3:0] _111_;
wire [2:0] _112_;
wire [2:0] _113_;
wire _114_;
wire [1:0] _115_;
wire [2:0] _116_;
wire [3:0] _117_;
wire [3:0] _118_;
wire [3:0] _119_;
wire _120_;
wire [2:0] _121_;
wire [3:0] _122_;
wire [4:0] _123_;
wire [31:0] _124_;
wire [31:0] _125_;
wire [31:0] _126_;
wire [31:0] _127_;
wire [31:0] _128_;
wire [31:0] _129_;
wire [31:0] _130_;
wire [31:0] _131_;
wire [31:0] _132_;
wire [31:0] _133_;
wire [31:0] _134_;
wire [31:0] _135_;
wire [31:0] _136_;
wire [31:0] _137_;
wire [31:0] _138_;
wire [31:0] _139_;
wire [31:0] _140_;
wire [31:0] _141_;
wire [31:0] _142_;
wire [31:0] _143_;
wire [31:0] _144_;
wire [31:0] _145_;
wire [31:0] _146_;
wire [31:0] _147_;
wire [31:0] _148_;
wire [31:0] _149_;
wire [31:0] _150_;
wire [31:0] _151_;
wire [31:0] _152_;
wire [31:0] _153_;
wire [31:0] _154_;
wire [31:0] _155_;
wire [31:0] _156_;
wire [31:0] _157_;
wire [31:0] _158_;
wire [31:0] _159_;
wire [31:0] _160_;
wire [31:0] _161_;
wire [31:0] _162_;
wire [31:0] _163_;
wire [31:0] _164_;
wire [31:0] _165_;
wire [31:0] _166_;
wire [31:0] _167_;
wire [31:0] _168_;
wire [31:0] _169_;
wire [31:0] _170_;
wire [31:0] _171_;
wire [31:0] _172_;
wire [31:0] _173_;
wire [31:0] _174_;
wire [31:0] _175_;
wire [31:0] _176_;
wire [31:0] _177_;
wire [31:0] _178_;
wire [31:0] _179_;
wire [31:0] _180_;
wire [31:0] _181_;
wire [31:0] _182_;
wire [31:0] _183_;
wire [10:0] _184_;
wire [10:0] _185_;
wire _186_;
wire [10:0] _187_;
wire [11:0] _188_;
wire [11:0] _189_;
wire [13:0] _190_;
wire [13:0] _191_;
wire _192_;
wire [13:0] _193_;
wire [14:0] _194_;
wire [14:0] _195_;
wire [15:0] _196_;
wire [15:0] _197_;
wire _198_;
wire [15:0] _199_;
wire [16:0] _200_;
wire [16:0] _201_;
wire _202_;
wire _203_;
wire _204_;
wire _205_;
wire _206_;
wire _207_;
wire _208_;
wire _209_;
wire _210_;
wire _211_;
wire _212_;
wire _213_;
wire _214_;
wire _215_;
wire _216_;
wire _217_;
wire _218_;
wire _219_;
wire _220_;
wire _221_;
wire _222_;
wire _223_;
wire _224_;
wire _225_;
wire _226_;
wire _227_;
wire _228_;
wire _229_;
wire \add_10ns_10s_10_2_1_U1.ce ;
wire \add_10ns_10s_10_2_1_U1.clk ;
wire [9:0] \add_10ns_10s_10_2_1_U1.din0 ;
wire [9:0] \add_10ns_10s_10_2_1_U1.din1 ;
wire [9:0] \add_10ns_10s_10_2_1_U1.dout ;
wire \add_10ns_10s_10_2_1_U1.reset ;
wire [9:0] \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.a ;
wire [9:0] \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.ain_s0 ;
wire [9:0] \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.b ;
wire [9:0] \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.bin_s0 ;
wire \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.ce ;
wire \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.clk ;
wire \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.facout_s1 ;
wire \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.facout_s2 ;
wire [4:0] \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.fas_s1 ;
wire [4:0] \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.fas_s2 ;
wire \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.reset ;
wire [9:0] \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.s ;
wire [4:0] \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.u1.a ;
wire [4:0] \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.u1.b ;
wire \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.u1.cin ;
wire \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.u1.cout ;
wire [4:0] \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.u1.s ;
wire [4:0] \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.u2.a ;
wire [4:0] \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.u2.b ;
wire \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.u2.cin ;
wire \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.u2.cout ;
wire [4:0] \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.u2.s ;
wire \add_17s_17s_17_2_1_U17.ce ;
wire \add_17s_17s_17_2_1_U17.clk ;
wire [16:0] \add_17s_17s_17_2_1_U17.din0 ;
wire [16:0] \add_17s_17s_17_2_1_U17.din1 ;
wire [16:0] \add_17s_17s_17_2_1_U17.dout ;
wire \add_17s_17s_17_2_1_U17.reset ;
wire [16:0] \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.a ;
wire [16:0] \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.ain_s0 ;
wire [16:0] \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.b ;
wire [16:0] \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.bin_s0 ;
wire \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.ce ;
wire \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.clk ;
wire \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.facout_s1 ;
wire \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.facout_s2 ;
wire [7:0] \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.fas_s1 ;
wire [8:0] \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.fas_s2 ;
wire \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.reset ;
wire [16:0] \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.s ;
wire [7:0] \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.u1.a ;
wire [7:0] \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.u1.b ;
wire \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.u1.cin ;
wire \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.u1.cout ;
wire [7:0] \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.u1.s ;
wire [8:0] \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.u2.a ;
wire [8:0] \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.u2.b ;
wire \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.u2.cin ;
wire \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.u2.cout ;
wire [8:0] \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.u2.s ;
wire \add_32ns_32ns_32_2_1_U15.ce ;
wire \add_32ns_32ns_32_2_1_U15.clk ;
wire [31:0] \add_32ns_32ns_32_2_1_U15.din0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U15.din1 ;
wire [31:0] \add_32ns_32ns_32_2_1_U15.dout ;
wire \add_32ns_32ns_32_2_1_U15.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.a ;
wire [31:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.ain_s0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.b ;
wire [31:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.bin_s0 ;
wire \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.ce ;
wire \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.clk ;
wire \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.facout_s1 ;
wire \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.facout_s2 ;
wire [15:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.fas_s1 ;
wire [15:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.fas_s2 ;
wire \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.b ;
wire \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.cin ;
wire \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.b ;
wire \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.cin ;
wire \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.s ;
wire \add_32ns_32ns_32_2_1_U16.ce ;
wire \add_32ns_32ns_32_2_1_U16.clk ;
wire [31:0] \add_32ns_32ns_32_2_1_U16.din0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U16.din1 ;
wire [31:0] \add_32ns_32ns_32_2_1_U16.dout ;
wire \add_32ns_32ns_32_2_1_U16.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.a ;
wire [31:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.ain_s0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.b ;
wire [31:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.bin_s0 ;
wire \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.ce ;
wire \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.clk ;
wire \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.facout_s1 ;
wire \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.facout_s2 ;
wire [15:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.fas_s1 ;
wire [15:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.fas_s2 ;
wire \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.b ;
wire \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.cin ;
wire \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.b ;
wire \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.cin ;
wire \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.s ;
wire \add_32ns_32s_32_2_1_U8.ce ;
wire \add_32ns_32s_32_2_1_U8.clk ;
wire [31:0] \add_32ns_32s_32_2_1_U8.din0 ;
wire [31:0] \add_32ns_32s_32_2_1_U8.din1 ;
wire [31:0] \add_32ns_32s_32_2_1_U8.dout ;
wire \add_32ns_32s_32_2_1_U8.reset ;
wire [31:0] \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.a ;
wire [31:0] \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.ain_s0 ;
wire [31:0] \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.b ;
wire [31:0] \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.bin_s0 ;
wire \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.ce ;
wire \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.clk ;
wire \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.facout_s1 ;
wire \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.facout_s2 ;
wire [15:0] \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.fas_s1 ;
wire [15:0] \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.fas_s2 ;
wire \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.reset ;
wire [31:0] \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.s ;
wire [15:0] \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.u1.a ;
wire [15:0] \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.u1.b ;
wire \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.u1.cin ;
wire \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.u1.cout ;
wire [15:0] \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.u1.s ;
wire [15:0] \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.u2.a ;
wire [15:0] \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.u2.b ;
wire \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.u2.cin ;
wire \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.u2.cout ;
wire [15:0] \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.u2.s ;
wire \add_32s_32ns_32_2_1_U13.ce ;
wire \add_32s_32ns_32_2_1_U13.clk ;
wire [31:0] \add_32s_32ns_32_2_1_U13.din0 ;
wire [31:0] \add_32s_32ns_32_2_1_U13.din1 ;
wire [31:0] \add_32s_32ns_32_2_1_U13.dout ;
wire \add_32s_32ns_32_2_1_U13.reset ;
wire [31:0] \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.a ;
wire [31:0] \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.ain_s0 ;
wire [31:0] \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.b ;
wire [31:0] \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.bin_s0 ;
wire \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.ce ;
wire \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.clk ;
wire \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.facout_s1 ;
wire \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.facout_s2 ;
wire [15:0] \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.fas_s1 ;
wire [15:0] \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.fas_s2 ;
wire \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.reset ;
wire [31:0] \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.s ;
wire [15:0] \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.u1.a ;
wire [15:0] \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.u1.b ;
wire \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.u1.cin ;
wire \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.u1.cout ;
wire [15:0] \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.u1.s ;
wire [15:0] \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.u2.a ;
wire [15:0] \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.u2.b ;
wire \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.u2.cin ;
wire \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.u2.cout ;
wire [15:0] \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.u2.s ;
wire \add_32s_32ns_32_2_1_U18.ce ;
wire \add_32s_32ns_32_2_1_U18.clk ;
wire [31:0] \add_32s_32ns_32_2_1_U18.din0 ;
wire [31:0] \add_32s_32ns_32_2_1_U18.din1 ;
wire [31:0] \add_32s_32ns_32_2_1_U18.dout ;
wire \add_32s_32ns_32_2_1_U18.reset ;
wire [31:0] \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.a ;
wire [31:0] \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.ain_s0 ;
wire [31:0] \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.b ;
wire [31:0] \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.bin_s0 ;
wire \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.ce ;
wire \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.clk ;
wire \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.facout_s1 ;
wire \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.facout_s2 ;
wire [15:0] \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.fas_s1 ;
wire [15:0] \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.fas_s2 ;
wire \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.reset ;
wire [31:0] \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.s ;
wire [15:0] \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.u1.a ;
wire [15:0] \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.u1.b ;
wire \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.u1.cin ;
wire \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.u1.cout ;
wire [15:0] \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.u1.s ;
wire [15:0] \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.u2.a ;
wire [15:0] \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.u2.b ;
wire \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.u2.cin ;
wire \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.u2.cout ;
wire [15:0] \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.u2.s ;
wire \add_32s_32ns_32_2_1_U6.ce ;
wire \add_32s_32ns_32_2_1_U6.clk ;
wire [31:0] \add_32s_32ns_32_2_1_U6.din0 ;
wire [31:0] \add_32s_32ns_32_2_1_U6.din1 ;
wire [31:0] \add_32s_32ns_32_2_1_U6.dout ;
wire \add_32s_32ns_32_2_1_U6.reset ;
wire [31:0] \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.a ;
wire [31:0] \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.ain_s0 ;
wire [31:0] \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.b ;
wire [31:0] \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.bin_s0 ;
wire \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.ce ;
wire \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.clk ;
wire \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.facout_s1 ;
wire \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.facout_s2 ;
wire [15:0] \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.fas_s1 ;
wire [15:0] \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.fas_s2 ;
wire \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.reset ;
wire [31:0] \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.s ;
wire [15:0] \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.u1.a ;
wire [15:0] \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.u1.b ;
wire \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.u1.cin ;
wire \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.u1.cout ;
wire [15:0] \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.u1.s ;
wire [15:0] \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.u2.a ;
wire [15:0] \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.u2.b ;
wire \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.u2.cin ;
wire \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.u2.cout ;
wire [15:0] \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.u2.s ;
wire \add_34s_34s_34_2_1_U14.ce ;
wire \add_34s_34s_34_2_1_U14.clk ;
wire [33:0] \add_34s_34s_34_2_1_U14.din0 ;
wire [33:0] \add_34s_34s_34_2_1_U14.din1 ;
wire [33:0] \add_34s_34s_34_2_1_U14.dout ;
wire \add_34s_34s_34_2_1_U14.reset ;
wire [33:0] \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.a ;
wire [33:0] \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.ain_s0 ;
wire [33:0] \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.b ;
wire [33:0] \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.bin_s0 ;
wire \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.ce ;
wire \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.clk ;
wire \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.facout_s1 ;
wire \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.facout_s2 ;
wire [16:0] \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.fas_s1 ;
wire [16:0] \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.fas_s2 ;
wire \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.reset ;
wire [33:0] \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.s ;
wire [16:0] \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.u1.a ;
wire [16:0] \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.u1.b ;
wire \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.u1.cin ;
wire \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.u1.cout ;
wire [16:0] \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.u1.s ;
wire [16:0] \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.u2.a ;
wire [16:0] \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.u2.b ;
wire \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.u2.cin ;
wire \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.u2.cout ;
wire [16:0] \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.u2.s ;
wire \add_3s_3ns_3_2_1_U9.ce ;
wire \add_3s_3ns_3_2_1_U9.clk ;
wire [2:0] \add_3s_3ns_3_2_1_U9.din0 ;
wire [2:0] \add_3s_3ns_3_2_1_U9.din1 ;
wire [2:0] \add_3s_3ns_3_2_1_U9.dout ;
wire \add_3s_3ns_3_2_1_U9.reset ;
wire [2:0] \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.a ;
wire [2:0] \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.ain_s0 ;
wire [2:0] \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.b ;
wire [2:0] \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.bin_s0 ;
wire \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.ce ;
wire \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.clk ;
wire \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.facout_s1 ;
wire \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.facout_s2 ;
wire \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.fas_s1 ;
wire [1:0] \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.fas_s2 ;
wire \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.reset ;
wire [2:0] \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.s ;
wire \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.u1.a ;
wire \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.u1.b ;
wire \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.u1.cin ;
wire \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.u1.cout ;
wire \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.u1.s ;
wire [1:0] \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.u2.a ;
wire [1:0] \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.u2.b ;
wire \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.u2.cin ;
wire \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.u2.cout ;
wire [1:0] \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.u2.s ;
wire \add_5ns_5ns_5_2_1_U3.ce ;
wire \add_5ns_5ns_5_2_1_U3.clk ;
wire [4:0] \add_5ns_5ns_5_2_1_U3.din0 ;
wire [4:0] \add_5ns_5ns_5_2_1_U3.din1 ;
wire [4:0] \add_5ns_5ns_5_2_1_U3.dout ;
wire \add_5ns_5ns_5_2_1_U3.reset ;
wire [4:0] \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.a ;
wire [4:0] \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.ain_s0 ;
wire [4:0] \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.b ;
wire [4:0] \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.bin_s0 ;
wire \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.ce ;
wire \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.clk ;
wire \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.facout_s1 ;
wire \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.facout_s2 ;
wire [1:0] \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.fas_s1 ;
wire [2:0] \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.fas_s2 ;
wire \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.reset ;
wire [4:0] \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.s ;
wire [1:0] \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.u1.a ;
wire [1:0] \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.u1.b ;
wire \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.u1.cin ;
wire \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.u1.cout ;
wire [1:0] \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.u1.s ;
wire [2:0] \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.u2.a ;
wire [2:0] \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.u2.b ;
wire \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.u2.cin ;
wire \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.u2.cout ;
wire [2:0] \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.u2.s ;
wire \add_5s_5ns_5_2_1_U2.ce ;
wire \add_5s_5ns_5_2_1_U2.clk ;
wire [4:0] \add_5s_5ns_5_2_1_U2.din0 ;
wire [4:0] \add_5s_5ns_5_2_1_U2.din1 ;
wire [4:0] \add_5s_5ns_5_2_1_U2.dout ;
wire \add_5s_5ns_5_2_1_U2.reset ;
wire [4:0] \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.a ;
wire [4:0] \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.ain_s0 ;
wire [4:0] \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.b ;
wire [4:0] \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.bin_s0 ;
wire \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.ce ;
wire \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.clk ;
wire \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.facout_s1 ;
wire \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.facout_s2 ;
wire [1:0] \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.fas_s1 ;
wire [2:0] \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.fas_s2 ;
wire \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.reset ;
wire [4:0] \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.s ;
wire [1:0] \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.u1.a ;
wire [1:0] \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.u1.b ;
wire \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.u1.cin ;
wire \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.u1.cout ;
wire [1:0] \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.u1.s ;
wire [2:0] \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.u2.a ;
wire [2:0] \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.u2.b ;
wire \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.u2.cin ;
wire \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.u2.cout ;
wire [2:0] \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.u2.s ;
wire \add_7s_7s_7_2_1_U4.ce ;
wire \add_7s_7s_7_2_1_U4.clk ;
wire [6:0] \add_7s_7s_7_2_1_U4.din0 ;
wire [6:0] \add_7s_7s_7_2_1_U4.din1 ;
wire [6:0] \add_7s_7s_7_2_1_U4.dout ;
wire \add_7s_7s_7_2_1_U4.reset ;
wire [6:0] \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.a ;
wire [6:0] \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.ain_s0 ;
wire [6:0] \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.b ;
wire [6:0] \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.bin_s0 ;
wire \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.ce ;
wire \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.clk ;
wire \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.facout_s1 ;
wire \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.facout_s2 ;
wire [2:0] \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.fas_s1 ;
wire [3:0] \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.fas_s2 ;
wire \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.reset ;
wire [6:0] \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.s ;
wire [2:0] \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.u1.a ;
wire [2:0] \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.u1.b ;
wire \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.u1.cin ;
wire \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.u1.cout ;
wire [2:0] \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.u1.s ;
wire [3:0] \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.u2.a ;
wire [3:0] \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.u2.b ;
wire \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.u2.cin ;
wire \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.u2.cout ;
wire [3:0] \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.u2.s ;
wire and_ln353_fu_445_p2;
wire ap_CS_fsm_state1;
wire ap_CS_fsm_state10;
wire ap_CS_fsm_state11;
wire ap_CS_fsm_state12;
wire ap_CS_fsm_state13;
wire ap_CS_fsm_state14;
wire ap_CS_fsm_state15;
wire ap_CS_fsm_state16;
wire ap_CS_fsm_state17;
wire ap_CS_fsm_state18;
wire ap_CS_fsm_state19;
wire ap_CS_fsm_state2;
wire ap_CS_fsm_state20;
wire ap_CS_fsm_state21;
wire ap_CS_fsm_state22;
wire ap_CS_fsm_state23;
wire ap_CS_fsm_state24;
wire ap_CS_fsm_state3;
wire ap_CS_fsm_state4;
wire ap_CS_fsm_state5;
wire ap_CS_fsm_state6;
wire ap_CS_fsm_state7;
wire ap_CS_fsm_state8;
wire ap_CS_fsm_state9;
wire [23:0] ap_NS_fsm;
wire ap_clk;
wire ap_done;
wire ap_idle;
wire ap_ready;
wire ap_rst;
wire ap_start;
wire \ashr_32s_32ns_32_7_1_U10.ce ;
wire \ashr_32s_32ns_32_7_1_U10.clk ;
wire [31:0] \ashr_32s_32ns_32_7_1_U10.din0 ;
wire [31:0] \ashr_32s_32ns_32_7_1_U10.din1 ;
wire [31:0] \ashr_32s_32ns_32_7_1_U10.din1_cast ;
wire [31:0] \ashr_32s_32ns_32_7_1_U10.din1_mask ;
wire [31:0] \ashr_32s_32ns_32_7_1_U10.dout ;
wire \ashr_32s_32ns_32_7_1_U10.reset ;
wire [9:0] grp_fu_221_p0;
wire [9:0] grp_fu_221_p1;
wire [9:0] grp_fu_221_p2;
wire [4:0] grp_fu_296_p0;
wire [4:0] grp_fu_296_p1;
wire [4:0] grp_fu_296_p2;
wire [4:0] grp_fu_336_p2;
wire [6:0] grp_fu_355_p0;
wire [6:0] grp_fu_355_p1;
wire [6:0] grp_fu_355_p2;
wire [27:0] grp_fu_383_p0;
wire [27:0] grp_fu_383_p1;
wire [27:0] grp_fu_383_p2;
wire [31:0] grp_fu_406_p0;
wire [31:0] grp_fu_406_p2;
wire [31:0] grp_fu_425_p2;
wire [31:0] grp_fu_495_p1;
wire [31:0] grp_fu_495_p2;
wire [2:0] grp_fu_500_p0;
wire [2:0] grp_fu_500_p2;
wire [31:0] grp_fu_509_p2;
wire [31:0] grp_fu_514_p2;
wire [21:0] grp_fu_529_p0;
wire [21:0] grp_fu_529_p1;
wire [21:0] grp_fu_529_p2;
wire [31:0] grp_fu_538_p0;
wire [31:0] grp_fu_538_p2;
wire [33:0] grp_fu_567_p0;
wire [33:0] grp_fu_567_p1;
wire [33:0] grp_fu_567_p2;
wire [31:0] grp_fu_583_p2;
wire [31:0] grp_fu_631_p1;
wire [31:0] grp_fu_631_p2;
wire [16:0] grp_fu_643_p0;
wire [16:0] grp_fu_643_p1;
wire [16:0] grp_fu_643_p2;
wire [31:0] grp_fu_652_p0;
wire [31:0] grp_fu_652_p2;
wire icmp_ln768_fu_284_p2;
wire icmp_ln850_fu_412_p2;
wire lhs_V_4_fu_237_p2;
wire [26:0] lhs_V_fu_368_p3;
wire newsignbit_fu_227_p2;
wire [3:0] op_0;
wire [7:0] op_1;
wire op_10_V_fu_322_p3;
wire [1:0] op_11;
wire [1:0] op_12;
wire [31:0] op_14;
wire [15:0] op_15;
wire [15:0] op_19;
wire [15:0] op_2;
wire [31:0] op_29;
wire op_29_ap_vld;
wire op_3_V_fu_197_p1;
wire [7:0] op_4;
wire [7:0] op_5;
wire op_6_V_fu_261_p2;
wire [7:0] op_7;
wire [19:0] op_8_V_fu_361_p3;
wire [1:0] op_9;
wire or_ln340_fu_317_p2;
wire or_ln785_fu_302_p2;
wire overflow_fu_311_p2;
wire p_Result_1_fu_456_p3;
wire p_Result_2_fu_601_p3;
wire p_Result_s_12_fu_438_p3;
wire [1:0] r_fu_596_p3;
wire ret_V_10_fu_450_p2;
wire [31:0] ret_V_13_fu_472_p3;
wire [31:0] ret_V_15_fu_621_p3;
wire [32:0] rhs_4_fu_556_p3;
wire [4:0] select_ln1192_fu_328_p3;
wire [2:0] select_ln69_fu_479_p3;
wire [31:0] select_ln850_1_fu_615_p3;
wire [31:0] select_ln850_fu_466_p3;
wire [1:0] sext_ln1192_fu_340_p0;
wire [7:0] sext_ln215_fu_205_p0;
wire [31:0] sext_ln781_fu_505_p1;
wire [31:0] sext_ln831_fu_403_p1;
wire \shl_32s_32ns_32_7_1_U11.ce ;
wire \shl_32s_32ns_32_7_1_U11.clk ;
wire [31:0] \shl_32s_32ns_32_7_1_U11.din0 ;
wire [31:0] \shl_32s_32ns_32_7_1_U11.din1 ;
wire [31:0] \shl_32s_32ns_32_7_1_U11.din1_cast ;
wire [31:0] \shl_32s_32ns_32_7_1_U11.din1_mask ;
wire [31:0] \shl_32s_32ns_32_7_1_U11.dout ;
wire \shl_32s_32ns_32_7_1_U11.reset ;
wire signbit_1_fu_247_p2;
wire \sub_22ns_22ns_22_2_1_U12.ce ;
wire \sub_22ns_22ns_22_2_1_U12.clk ;
wire [21:0] \sub_22ns_22ns_22_2_1_U12.din0 ;
wire [21:0] \sub_22ns_22ns_22_2_1_U12.din1 ;
wire [21:0] \sub_22ns_22ns_22_2_1_U12.dout ;
wire \sub_22ns_22ns_22_2_1_U12.reset ;
wire [21:0] \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.a ;
wire [21:0] \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.ain_s0 ;
wire [21:0] \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.b ;
wire [21:0] \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.bin_s0 ;
wire \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.ce ;
wire \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.clk ;
wire \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.facout_s1 ;
wire \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.facout_s2 ;
wire [10:0] \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.fas_s1 ;
wire [10:0] \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.fas_s2 ;
wire \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.reset ;
wire [21:0] \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.s ;
wire [10:0] \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.u1.a ;
wire [10:0] \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.u1.b ;
wire \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.u1.cin ;
wire \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.u1.cout ;
wire [10:0] \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.u1.s ;
wire [10:0] \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.u2.a ;
wire [10:0] \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.u2.b ;
wire \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.u2.cin ;
wire \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.u2.cout ;
wire [10:0] \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.u2.s ;
wire \sub_28s_28ns_28_2_1_U5.ce ;
wire \sub_28s_28ns_28_2_1_U5.clk ;
wire [27:0] \sub_28s_28ns_28_2_1_U5.din0 ;
wire [27:0] \sub_28s_28ns_28_2_1_U5.din1 ;
wire [27:0] \sub_28s_28ns_28_2_1_U5.dout ;
wire \sub_28s_28ns_28_2_1_U5.reset ;
wire [27:0] \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.a ;
wire [27:0] \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.ain_s0 ;
wire [27:0] \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.b ;
wire [27:0] \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.bin_s0 ;
wire \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.ce ;
wire \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.clk ;
wire \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.facout_s1 ;
wire \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.facout_s2 ;
wire [13:0] \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.fas_s1 ;
wire [13:0] \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.fas_s2 ;
wire \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.reset ;
wire [27:0] \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.s ;
wire [13:0] \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.u1.a ;
wire [13:0] \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.u1.b ;
wire \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.u1.cin ;
wire \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.u1.cout ;
wire [13:0] \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.u1.s ;
wire [13:0] \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.u2.a ;
wire [13:0] \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.u2.b ;
wire \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.u2.cin ;
wire \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.u2.cout ;
wire [13:0] \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.u2.s ;
wire \sub_32ns_32ns_32_2_1_U7.ce ;
wire \sub_32ns_32ns_32_2_1_U7.clk ;
wire [31:0] \sub_32ns_32ns_32_2_1_U7.din0 ;
wire [31:0] \sub_32ns_32ns_32_2_1_U7.din1 ;
wire [31:0] \sub_32ns_32ns_32_2_1_U7.dout ;
wire \sub_32ns_32ns_32_2_1_U7.reset ;
wire [31:0] \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.a ;
wire [31:0] \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.ain_s0 ;
wire [31:0] \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.b ;
wire [31:0] \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.bin_s0 ;
wire \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.ce ;
wire \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.clk ;
wire \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.facout_s1 ;
wire \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.facout_s2 ;
wire [15:0] \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.fas_s1 ;
wire [15:0] \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.fas_s2 ;
wire \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.reset ;
wire [31:0] \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.s ;
wire [15:0] \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.u1.a ;
wire [15:0] \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.u1.b ;
wire \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.u1.cin ;
wire \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.u1.cout ;
wire [15:0] \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.u1.s ;
wire [15:0] \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.u2.a ;
wire [15:0] \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.u2.b ;
wire \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.u2.cin ;
wire \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.u2.cout ;
wire [15:0] \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.u2.s ;
wire [5:0] tmp_4_fu_344_p3;
wire tmp_6_fu_608_p3;
wire tmp_fu_431_p3;
wire trunc_ln1346_1_fu_217_p1;
wire [7:0] trunc_ln1346_fu_213_p0;
wire trunc_ln1346_fu_213_p1;
wire trunc_ln213_1_fu_257_p1;
wire trunc_ln213_fu_201_p1;
wire [2:0] trunc_ln728_fu_253_p1;
wire [1:0] trunc_ln798_1_fu_592_p1;
wire [1:0] trunc_ln798_fu_588_p1;
wire [1:0] trunc_ln851_1_fu_463_p0;
wire trunc_ln851_1_fu_463_p1;
wire [18:0] trunc_ln851_fu_399_p1;
wire xor_ln785_fu_306_p2;
wire [15:0] zext_ln878_1_fu_243_p1;
wire [15:0] zext_ln878_fu_233_p1;


assign _040_ = ap_CS_fsm[18] & _044_;
assign _041_ = ap_CS_fsm[18] & p_Result_4_reg_820;
assign _042_ = _045_ & ap_CS_fsm[0];
assign _043_ = ap_start & ap_CS_fsm[0];
assign and_ln353_fu_445_p2 = ret_V_9_reg_786[27] & icmp_ln850_reg_804;
assign overflow_fu_311_p2 = xor_ln785_fu_306_p2 & or_ln785_fu_302_p2;
assign xor_ln785_fu_306_p2 = ~ p_Result_3_reg_704;
assign _044_ = ~ p_Result_4_reg_820;
assign _045_ = ~ ap_start;
always @(posedge \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.clk )
\add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.bin_s1  <= _047_;
always @(posedge \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.clk )
\add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.ain_s1  <= _046_;
always @(posedge \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.clk )
\add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.sum_s1  <= _049_;
always @(posedge \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.clk )
\add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.carry_s1  <= _048_;
assign _047_ = \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.ce  ? \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.b [9:5] : \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.bin_s1 ;
assign _046_ = \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.ce  ? \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.a [9:5] : \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.ain_s1 ;
assign _048_ = \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.ce  ? \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.facout_s1  : \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.carry_s1 ;
assign _049_ = \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.ce  ? \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.fas_s1  : \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.sum_s1 ;
assign _050_ = \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.u1.a  + \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.u1.b ;
assign { \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.u1.cout , \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.u1.s  } = _050_ + \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.u1.cin ;
assign _051_ = \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.u2.a  + \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.u2.b ;
assign { \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.u2.cout , \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.u2.s  } = _051_ + \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.u2.cin ;
always @(posedge \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.clk )
\add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.bin_s1  <= _053_;
always @(posedge \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.clk )
\add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.ain_s1  <= _052_;
always @(posedge \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.clk )
\add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.sum_s1  <= _055_;
always @(posedge \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.clk )
\add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.carry_s1  <= _054_;
assign _053_ = \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.ce  ? \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.b [16:8] : \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.bin_s1 ;
assign _052_ = \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.ce  ? \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.a [16:8] : \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.ain_s1 ;
assign _054_ = \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.ce  ? \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.facout_s1  : \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.carry_s1 ;
assign _055_ = \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.ce  ? \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.fas_s1  : \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.sum_s1 ;
assign _056_ = \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.u1.a  + \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.u1.b ;
assign { \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.u1.cout , \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.u1.s  } = _056_ + \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.u1.cin ;
assign _057_ = \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.u2.a  + \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.u2.b ;
assign { \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.u2.cout , \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.u2.s  } = _057_ + \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.u2.cin ;
always @(posedge \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.clk )
\add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.bin_s1  <= _059_;
always @(posedge \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.clk )
\add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.ain_s1  <= _058_;
always @(posedge \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.clk )
\add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.sum_s1  <= _061_;
always @(posedge \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.clk )
\add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.carry_s1  <= _060_;
assign _059_ = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.ce  ? \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.b [31:16] : \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.bin_s1 ;
assign _058_ = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.ce  ? \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.a [31:16] : \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.ain_s1 ;
assign _060_ = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.ce  ? \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.facout_s1  : \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.carry_s1 ;
assign _061_ = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.ce  ? \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.fas_s1  : \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.sum_s1 ;
assign _062_ = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.a  + \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.b ;
assign { \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.cout , \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.s  } = _062_ + \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.cin ;
assign _063_ = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.a  + \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.b ;
assign { \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.cout , \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.s  } = _063_ + \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.cin ;
always @(posedge \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.clk )
\add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.bin_s1  <= _065_;
always @(posedge \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.clk )
\add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.ain_s1  <= _064_;
always @(posedge \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.clk )
\add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.sum_s1  <= _067_;
always @(posedge \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.clk )
\add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.carry_s1  <= _066_;
assign _065_ = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.ce  ? \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.b [31:16] : \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.bin_s1 ;
assign _064_ = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.ce  ? \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.a [31:16] : \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.ain_s1 ;
assign _066_ = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.ce  ? \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.facout_s1  : \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.carry_s1 ;
assign _067_ = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.ce  ? \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.fas_s1  : \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.sum_s1 ;
assign _068_ = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.a  + \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.b ;
assign { \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.cout , \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.s  } = _068_ + \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.cin ;
assign _069_ = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.a  + \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.b ;
assign { \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.cout , \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.s  } = _069_ + \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.cin ;
always @(posedge \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.clk )
\add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.bin_s1  <= _071_;
always @(posedge \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.clk )
\add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.ain_s1  <= _070_;
always @(posedge \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.clk )
\add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.sum_s1  <= _073_;
always @(posedge \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.clk )
\add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.carry_s1  <= _072_;
assign _071_ = \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.ce  ? \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.b [31:16] : \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.bin_s1 ;
assign _070_ = \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.ce  ? \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.a [31:16] : \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.ain_s1 ;
assign _072_ = \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.ce  ? \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.facout_s1  : \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.carry_s1 ;
assign _073_ = \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.ce  ? \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.fas_s1  : \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.sum_s1 ;
assign _074_ = \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.u1.a  + \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.u1.b ;
assign { \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.u1.cout , \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.u1.s  } = _074_ + \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.u1.cin ;
assign _075_ = \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.u2.a  + \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.u2.b ;
assign { \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.u2.cout , \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.u2.s  } = _075_ + \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.u2.cin ;
always @(posedge \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.clk )
\add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.bin_s1  <= _077_;
always @(posedge \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.clk )
\add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.ain_s1  <= _076_;
always @(posedge \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.clk )
\add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.sum_s1  <= _079_;
always @(posedge \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.clk )
\add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.carry_s1  <= _078_;
assign _077_ = \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.ce  ? \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.b [31:16] : \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.bin_s1 ;
assign _076_ = \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.ce  ? \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.a [31:16] : \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.ain_s1 ;
assign _078_ = \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.ce  ? \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.facout_s1  : \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.carry_s1 ;
assign _079_ = \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.ce  ? \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.fas_s1  : \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.sum_s1 ;
assign _080_ = \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.u1.a  + \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.u1.b ;
assign { \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.u1.cout , \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.u1.s  } = _080_ + \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.u1.cin ;
assign _081_ = \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.u2.a  + \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.u2.b ;
assign { \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.u2.cout , \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.u2.s  } = _081_ + \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.u2.cin ;
always @(posedge \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.clk )
\add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.bin_s1  <= _083_;
always @(posedge \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.clk )
\add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.ain_s1  <= _082_;
always @(posedge \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.clk )
\add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.sum_s1  <= _085_;
always @(posedge \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.clk )
\add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.carry_s1  <= _084_;
assign _083_ = \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.ce  ? \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.b [31:16] : \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.bin_s1 ;
assign _082_ = \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.ce  ? \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.a [31:16] : \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.ain_s1 ;
assign _084_ = \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.ce  ? \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.facout_s1  : \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.carry_s1 ;
assign _085_ = \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.ce  ? \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.fas_s1  : \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.sum_s1 ;
assign _086_ = \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.u1.a  + \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.u1.b ;
assign { \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.u1.cout , \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.u1.s  } = _086_ + \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.u1.cin ;
assign _087_ = \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.u2.a  + \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.u2.b ;
assign { \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.u2.cout , \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.u2.s  } = _087_ + \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.u2.cin ;
always @(posedge \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.clk )
\add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.bin_s1  <= _089_;
always @(posedge \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.clk )
\add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.ain_s1  <= _088_;
always @(posedge \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.clk )
\add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.sum_s1  <= _091_;
always @(posedge \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.clk )
\add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.carry_s1  <= _090_;
assign _089_ = \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.ce  ? \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.b [31:16] : \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.bin_s1 ;
assign _088_ = \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.ce  ? \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.a [31:16] : \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.ain_s1 ;
assign _090_ = \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.ce  ? \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.facout_s1  : \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.carry_s1 ;
assign _091_ = \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.ce  ? \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.fas_s1  : \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.sum_s1 ;
assign _092_ = \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.u1.a  + \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.u1.b ;
assign { \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.u1.cout , \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.u1.s  } = _092_ + \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.u1.cin ;
assign _093_ = \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.u2.a  + \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.u2.b ;
assign { \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.u2.cout , \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.u2.s  } = _093_ + \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.u2.cin ;
always @(posedge \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.clk )
\add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.bin_s1  <= _095_;
always @(posedge \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.clk )
\add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.ain_s1  <= _094_;
always @(posedge \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.clk )
\add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.sum_s1  <= _097_;
always @(posedge \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.clk )
\add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.carry_s1  <= _096_;
assign _095_ = \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.ce  ? \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.b [33:17] : \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.bin_s1 ;
assign _094_ = \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.ce  ? \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.a [33:17] : \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.ain_s1 ;
assign _096_ = \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.ce  ? \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.facout_s1  : \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.carry_s1 ;
assign _097_ = \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.ce  ? \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.fas_s1  : \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.sum_s1 ;
assign _098_ = \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.u1.a  + \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.u1.b ;
assign { \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.u1.cout , \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.u1.s  } = _098_ + \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.u1.cin ;
assign _099_ = \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.u2.a  + \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.u2.b ;
assign { \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.u2.cout , \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.u2.s  } = _099_ + \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.u2.cin ;
always @(posedge \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.clk )
\add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.bin_s1  <= _101_;
always @(posedge \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.clk )
\add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.ain_s1  <= _100_;
always @(posedge \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.clk )
\add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.sum_s1  <= _103_;
always @(posedge \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.clk )
\add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.carry_s1  <= _102_;
assign _101_ = \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.ce  ? \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.b [2:1] : \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.bin_s1 ;
assign _100_ = \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.ce  ? \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.a [2:1] : \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.ain_s1 ;
assign _102_ = \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.ce  ? \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.facout_s1  : \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.carry_s1 ;
assign _103_ = \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.ce  ? \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.fas_s1  : \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.sum_s1 ;
assign _104_ = \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.u1.a  + \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.u1.b ;
assign { \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.u1.cout , \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.u1.s  } = _104_ + \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.u1.cin ;
assign _105_ = \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.u2.a  + \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.u2.b ;
assign { \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.u2.cout , \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.u2.s  } = _105_ + \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.u2.cin ;
always @(posedge \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.clk )
\add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.bin_s1  <= _107_;
always @(posedge \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.clk )
\add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.ain_s1  <= _106_;
always @(posedge \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.clk )
\add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.sum_s1  <= _109_;
always @(posedge \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.clk )
\add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.carry_s1  <= _108_;
assign _107_ = \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.ce  ? \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.b [4:2] : \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.bin_s1 ;
assign _106_ = \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.ce  ? \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.a [4:2] : \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.ain_s1 ;
assign _108_ = \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.ce  ? \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.facout_s1  : \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.carry_s1 ;
assign _109_ = \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.ce  ? \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.fas_s1  : \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.sum_s1 ;
assign _110_ = \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.u1.a  + \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.u1.b ;
assign { \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.u1.cout , \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.u1.s  } = _110_ + \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.u1.cin ;
assign _111_ = \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.u2.a  + \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.u2.b ;
assign { \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.u2.cout , \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.u2.s  } = _111_ + \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.u2.cin ;
always @(posedge \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.clk )
\add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.bin_s1  <= _113_;
always @(posedge \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.clk )
\add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.ain_s1  <= _112_;
always @(posedge \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.clk )
\add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.sum_s1  <= _115_;
always @(posedge \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.clk )
\add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.carry_s1  <= _114_;
assign _113_ = \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.ce  ? \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.b [4:2] : \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.bin_s1 ;
assign _112_ = \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.ce  ? \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.a [4:2] : \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.ain_s1 ;
assign _114_ = \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.ce  ? \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.facout_s1  : \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.carry_s1 ;
assign _115_ = \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.ce  ? \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.fas_s1  : \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.sum_s1 ;
assign _116_ = \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.u1.a  + \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.u1.b ;
assign { \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.u1.cout , \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.u1.s  } = _116_ + \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.u1.cin ;
assign _117_ = \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.u2.a  + \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.u2.b ;
assign { \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.u2.cout , \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.u2.s  } = _117_ + \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.u2.cin ;
always @(posedge \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.clk )
\add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.bin_s1  <= _119_;
always @(posedge \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.clk )
\add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.ain_s1  <= _118_;
always @(posedge \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.clk )
\add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.sum_s1  <= _121_;
always @(posedge \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.clk )
\add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.carry_s1  <= _120_;
assign _119_ = \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.ce  ? \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.b [6:3] : \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.bin_s1 ;
assign _118_ = \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.ce  ? \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.a [6:3] : \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.ain_s1 ;
assign _120_ = \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.ce  ? \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.facout_s1  : \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.carry_s1 ;
assign _121_ = \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.ce  ? \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.fas_s1  : \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.sum_s1 ;
assign _122_ = \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.u1.a  + \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.u1.b ;
assign { \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.u1.cout , \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.u1.s  } = _122_ + \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.u1.cin ;
assign _123_ = \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.u2.a  + \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.u2.b ;
assign { \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.u2.cout , \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.u2.s  } = _123_ + \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.u2.cin ;
always @(posedge \ashr_32s_32ns_32_7_1_U10.clk )
\ashr_32s_32ns_32_7_1_U10.dout_array[5]  <= _135_;
always @(posedge \ashr_32s_32ns_32_7_1_U10.clk )
\ashr_32s_32ns_32_7_1_U10.din1_cast_array[5]  <= _129_;
always @(posedge \ashr_32s_32ns_32_7_1_U10.clk )
\ashr_32s_32ns_32_7_1_U10.dout_array[4]  <= _134_;
always @(posedge \ashr_32s_32ns_32_7_1_U10.clk )
\ashr_32s_32ns_32_7_1_U10.din1_cast_array[4]  <= _128_;
always @(posedge \ashr_32s_32ns_32_7_1_U10.clk )
\ashr_32s_32ns_32_7_1_U10.dout_array[3]  <= _133_;
always @(posedge \ashr_32s_32ns_32_7_1_U10.clk )
\ashr_32s_32ns_32_7_1_U10.din1_cast_array[3]  <= _127_;
always @(posedge \ashr_32s_32ns_32_7_1_U10.clk )
\ashr_32s_32ns_32_7_1_U10.dout_array[2]  <= _132_;
always @(posedge \ashr_32s_32ns_32_7_1_U10.clk )
\ashr_32s_32ns_32_7_1_U10.din1_cast_array[2]  <= _126_;
always @(posedge \ashr_32s_32ns_32_7_1_U10.clk )
\ashr_32s_32ns_32_7_1_U10.dout_array[1]  <= _131_;
always @(posedge \ashr_32s_32ns_32_7_1_U10.clk )
\ashr_32s_32ns_32_7_1_U10.din1_cast_array[1]  <= _125_;
always @(posedge \ashr_32s_32ns_32_7_1_U10.clk )
\ashr_32s_32ns_32_7_1_U10.dout_array[0]  <= _130_;
always @(posedge \ashr_32s_32ns_32_7_1_U10.clk )
\ashr_32s_32ns_32_7_1_U10.din1_cast_array[0]  <= _124_;
assign _136_ = \ashr_32s_32ns_32_7_1_U10.ce  ? \ashr_32s_32ns_32_7_1_U10.din1_cast_array[4]  : \ashr_32s_32ns_32_7_1_U10.din1_cast_array[5] ;
assign _129_ = \ashr_32s_32ns_32_7_1_U10.reset  ? 32'd0 : _136_;
assign _137_ = \ashr_32s_32ns_32_7_1_U10.ce  ? _153_ : \ashr_32s_32ns_32_7_1_U10.dout_array[5] ;
assign _135_ = \ashr_32s_32ns_32_7_1_U10.reset  ? 32'd0 : _137_;
assign _138_ = \ashr_32s_32ns_32_7_1_U10.ce  ? \ashr_32s_32ns_32_7_1_U10.din1_cast_array[3]  : \ashr_32s_32ns_32_7_1_U10.din1_cast_array[4] ;
assign _128_ = \ashr_32s_32ns_32_7_1_U10.reset  ? 32'd0 : _138_;
assign _139_ = \ashr_32s_32ns_32_7_1_U10.ce  ? _152_ : \ashr_32s_32ns_32_7_1_U10.dout_array[4] ;
assign _134_ = \ashr_32s_32ns_32_7_1_U10.reset  ? 32'd0 : _139_;
assign _140_ = \ashr_32s_32ns_32_7_1_U10.ce  ? \ashr_32s_32ns_32_7_1_U10.din1_cast_array[2]  : \ashr_32s_32ns_32_7_1_U10.din1_cast_array[3] ;
assign _127_ = \ashr_32s_32ns_32_7_1_U10.reset  ? 32'd0 : _140_;
assign _141_ = \ashr_32s_32ns_32_7_1_U10.ce  ? _151_ : \ashr_32s_32ns_32_7_1_U10.dout_array[3] ;
assign _133_ = \ashr_32s_32ns_32_7_1_U10.reset  ? 32'd0 : _141_;
assign _142_ = \ashr_32s_32ns_32_7_1_U10.ce  ? \ashr_32s_32ns_32_7_1_U10.din1_cast_array[1]  : \ashr_32s_32ns_32_7_1_U10.din1_cast_array[2] ;
assign _126_ = \ashr_32s_32ns_32_7_1_U10.reset  ? 32'd0 : _142_;
assign _143_ = \ashr_32s_32ns_32_7_1_U10.ce  ? _150_ : \ashr_32s_32ns_32_7_1_U10.dout_array[2] ;
assign _132_ = \ashr_32s_32ns_32_7_1_U10.reset  ? 32'd0 : _143_;
assign _144_ = \ashr_32s_32ns_32_7_1_U10.ce  ? \ashr_32s_32ns_32_7_1_U10.din1_cast_array[0]  : \ashr_32s_32ns_32_7_1_U10.din1_cast_array[1] ;
assign _125_ = \ashr_32s_32ns_32_7_1_U10.reset  ? 32'd0 : _144_;
assign _145_ = \ashr_32s_32ns_32_7_1_U10.ce  ? _149_ : \ashr_32s_32ns_32_7_1_U10.dout_array[1] ;
assign _131_ = \ashr_32s_32ns_32_7_1_U10.reset  ? 32'd0 : _145_;
assign _146_ = \ashr_32s_32ns_32_7_1_U10.ce  ? \ashr_32s_32ns_32_7_1_U10.din1  : \ashr_32s_32ns_32_7_1_U10.din1_cast_array[0] ;
assign _124_ = \ashr_32s_32ns_32_7_1_U10.reset  ? 32'd0 : _146_;
assign _147_ = \ashr_32s_32ns_32_7_1_U10.ce  ? _148_ : \ashr_32s_32ns_32_7_1_U10.dout_array[0] ;
assign _130_ = \ashr_32s_32ns_32_7_1_U10.reset  ? 32'd0 : _147_;
assign _148_ = $signed(\ashr_32s_32ns_32_7_1_U10.din0 ) >>> { \ashr_32s_32ns_32_7_1_U10.din1 [31:30], 30'h00000000 };
assign _149_ = $signed(\ashr_32s_32ns_32_7_1_U10.dout_array[0] ) >>> { \ashr_32s_32ns_32_7_1_U10.din1_cast_array[0] [29:25], 25'h0000000 };
assign _150_ = $signed(\ashr_32s_32ns_32_7_1_U10.dout_array[1] ) >>> { \ashr_32s_32ns_32_7_1_U10.din1_cast_array[1] [24:20], 20'h00000 };
assign _151_ = $signed(\ashr_32s_32ns_32_7_1_U10.dout_array[2] ) >>> { \ashr_32s_32ns_32_7_1_U10.din1_cast_array[2] [19:15], 15'h0000 };
assign _152_ = $signed(\ashr_32s_32ns_32_7_1_U10.dout_array[3] ) >>> { \ashr_32s_32ns_32_7_1_U10.din1_cast_array[3] [14:10], 10'h000 };
assign _153_ = $signed(\ashr_32s_32ns_32_7_1_U10.dout_array[4] ) >>> { \ashr_32s_32ns_32_7_1_U10.din1_cast_array[4] [9:5], 5'h00 };
assign \ashr_32s_32ns_32_7_1_U10.dout  = $signed(\ashr_32s_32ns_32_7_1_U10.dout_array[5] ) >>> \ashr_32s_32ns_32_7_1_U10.din1_cast_array[5] [4:0];
always @(posedge \shl_32s_32ns_32_7_1_U11.clk )
\shl_32s_32ns_32_7_1_U11.dout_array[5]  <= _165_;
always @(posedge \shl_32s_32ns_32_7_1_U11.clk )
\shl_32s_32ns_32_7_1_U11.din1_cast_array[5]  <= _159_;
always @(posedge \shl_32s_32ns_32_7_1_U11.clk )
\shl_32s_32ns_32_7_1_U11.dout_array[4]  <= _164_;
always @(posedge \shl_32s_32ns_32_7_1_U11.clk )
\shl_32s_32ns_32_7_1_U11.din1_cast_array[4]  <= _158_;
always @(posedge \shl_32s_32ns_32_7_1_U11.clk )
\shl_32s_32ns_32_7_1_U11.dout_array[3]  <= _163_;
always @(posedge \shl_32s_32ns_32_7_1_U11.clk )
\shl_32s_32ns_32_7_1_U11.din1_cast_array[3]  <= _157_;
always @(posedge \shl_32s_32ns_32_7_1_U11.clk )
\shl_32s_32ns_32_7_1_U11.dout_array[2]  <= _162_;
always @(posedge \shl_32s_32ns_32_7_1_U11.clk )
\shl_32s_32ns_32_7_1_U11.din1_cast_array[2]  <= _156_;
always @(posedge \shl_32s_32ns_32_7_1_U11.clk )
\shl_32s_32ns_32_7_1_U11.dout_array[1]  <= _161_;
always @(posedge \shl_32s_32ns_32_7_1_U11.clk )
\shl_32s_32ns_32_7_1_U11.din1_cast_array[1]  <= _155_;
always @(posedge \shl_32s_32ns_32_7_1_U11.clk )
\shl_32s_32ns_32_7_1_U11.dout_array[0]  <= _160_;
always @(posedge \shl_32s_32ns_32_7_1_U11.clk )
\shl_32s_32ns_32_7_1_U11.din1_cast_array[0]  <= _154_;
assign _166_ = \shl_32s_32ns_32_7_1_U11.ce  ? \shl_32s_32ns_32_7_1_U11.din1_cast_array[4]  : \shl_32s_32ns_32_7_1_U11.din1_cast_array[5] ;
assign _159_ = \shl_32s_32ns_32_7_1_U11.reset  ? 32'd0 : _166_;
assign _167_ = \shl_32s_32ns_32_7_1_U11.ce  ? _183_ : \shl_32s_32ns_32_7_1_U11.dout_array[5] ;
assign _165_ = \shl_32s_32ns_32_7_1_U11.reset  ? 32'd0 : _167_;
assign _168_ = \shl_32s_32ns_32_7_1_U11.ce  ? \shl_32s_32ns_32_7_1_U11.din1_cast_array[3]  : \shl_32s_32ns_32_7_1_U11.din1_cast_array[4] ;
assign _158_ = \shl_32s_32ns_32_7_1_U11.reset  ? 32'd0 : _168_;
assign _169_ = \shl_32s_32ns_32_7_1_U11.ce  ? _182_ : \shl_32s_32ns_32_7_1_U11.dout_array[4] ;
assign _164_ = \shl_32s_32ns_32_7_1_U11.reset  ? 32'd0 : _169_;
assign _170_ = \shl_32s_32ns_32_7_1_U11.ce  ? \shl_32s_32ns_32_7_1_U11.din1_cast_array[2]  : \shl_32s_32ns_32_7_1_U11.din1_cast_array[3] ;
assign _157_ = \shl_32s_32ns_32_7_1_U11.reset  ? 32'd0 : _170_;
assign _171_ = \shl_32s_32ns_32_7_1_U11.ce  ? _181_ : \shl_32s_32ns_32_7_1_U11.dout_array[3] ;
assign _163_ = \shl_32s_32ns_32_7_1_U11.reset  ? 32'd0 : _171_;
assign _172_ = \shl_32s_32ns_32_7_1_U11.ce  ? \shl_32s_32ns_32_7_1_U11.din1_cast_array[1]  : \shl_32s_32ns_32_7_1_U11.din1_cast_array[2] ;
assign _156_ = \shl_32s_32ns_32_7_1_U11.reset  ? 32'd0 : _172_;
assign _173_ = \shl_32s_32ns_32_7_1_U11.ce  ? _180_ : \shl_32s_32ns_32_7_1_U11.dout_array[2] ;
assign _162_ = \shl_32s_32ns_32_7_1_U11.reset  ? 32'd0 : _173_;
assign _174_ = \shl_32s_32ns_32_7_1_U11.ce  ? \shl_32s_32ns_32_7_1_U11.din1_cast_array[0]  : \shl_32s_32ns_32_7_1_U11.din1_cast_array[1] ;
assign _155_ = \shl_32s_32ns_32_7_1_U11.reset  ? 32'd0 : _174_;
assign _175_ = \shl_32s_32ns_32_7_1_U11.ce  ? _179_ : \shl_32s_32ns_32_7_1_U11.dout_array[1] ;
assign _161_ = \shl_32s_32ns_32_7_1_U11.reset  ? 32'd0 : _175_;
assign _176_ = \shl_32s_32ns_32_7_1_U11.ce  ? \shl_32s_32ns_32_7_1_U11.din1  : \shl_32s_32ns_32_7_1_U11.din1_cast_array[0] ;
assign _154_ = \shl_32s_32ns_32_7_1_U11.reset  ? 32'd0 : _176_;
assign _177_ = \shl_32s_32ns_32_7_1_U11.ce  ? _178_ : \shl_32s_32ns_32_7_1_U11.dout_array[0] ;
assign _160_ = \shl_32s_32ns_32_7_1_U11.reset  ? 32'd0 : _177_;
assign _178_ = \shl_32s_32ns_32_7_1_U11.din0  << { \shl_32s_32ns_32_7_1_U11.din1 [31:30], 30'h00000000 };
assign _179_ = \shl_32s_32ns_32_7_1_U11.dout_array[0]  << { \shl_32s_32ns_32_7_1_U11.din1_cast_array[0] [29:25], 25'h0000000 };
assign _180_ = \shl_32s_32ns_32_7_1_U11.dout_array[1]  << { \shl_32s_32ns_32_7_1_U11.din1_cast_array[1] [24:20], 20'h00000 };
assign _181_ = \shl_32s_32ns_32_7_1_U11.dout_array[2]  << { \shl_32s_32ns_32_7_1_U11.din1_cast_array[2] [19:15], 15'h0000 };
assign _182_ = \shl_32s_32ns_32_7_1_U11.dout_array[3]  << { \shl_32s_32ns_32_7_1_U11.din1_cast_array[3] [14:10], 10'h000 };
assign _183_ = \shl_32s_32ns_32_7_1_U11.dout_array[4]  << { \shl_32s_32ns_32_7_1_U11.din1_cast_array[4] [9:5], 5'h00 };
assign \shl_32s_32ns_32_7_1_U11.dout  = \shl_32s_32ns_32_7_1_U11.dout_array[5]  << \shl_32s_32ns_32_7_1_U11.din1_cast_array[5] [4:0];
assign \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.bin_s0  = ~ \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.b ;
always @(posedge \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.clk )
\sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.bin_s1  <= _185_;
always @(posedge \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.clk )
\sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.ain_s1  <= _184_;
always @(posedge \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.clk )
\sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.sum_s1  <= _187_;
always @(posedge \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.clk )
\sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.carry_s1  <= _186_;
assign _185_ = \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.ce  ? \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.bin_s0 [21:11] : \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.bin_s1 ;
assign _184_ = \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.ce  ? \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.a [21:11] : \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.ain_s1 ;
assign _186_ = \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.ce  ? \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.facout_s1  : \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.carry_s1 ;
assign _187_ = \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.ce  ? \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.fas_s1  : \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.sum_s1 ;
assign _188_ = \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.u1.a  + \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.u1.b ;
assign { \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.u1.cout , \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.u1.s  } = _188_ + \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.u1.cin ;
assign _189_ = \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.u2.a  + \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.u2.b ;
assign { \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.u2.cout , \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.u2.s  } = _189_ + \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.u2.cin ;
assign \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.bin_s0  = ~ \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.b ;
always @(posedge \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.clk )
\sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.bin_s1  <= _191_;
always @(posedge \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.clk )
\sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.ain_s1  <= _190_;
always @(posedge \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.clk )
\sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.sum_s1  <= _193_;
always @(posedge \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.clk )
\sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.carry_s1  <= _192_;
assign _191_ = \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.ce  ? \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.bin_s0 [27:14] : \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.bin_s1 ;
assign _190_ = \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.ce  ? \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.a [27:14] : \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.ain_s1 ;
assign _192_ = \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.ce  ? \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.facout_s1  : \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.carry_s1 ;
assign _193_ = \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.ce  ? \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.fas_s1  : \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.sum_s1 ;
assign _194_ = \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.u1.a  + \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.u1.b ;
assign { \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.u1.cout , \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.u1.s  } = _194_ + \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.u1.cin ;
assign _195_ = \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.u2.a  + \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.u2.b ;
assign { \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.u2.cout , \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.u2.s  } = _195_ + \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.u2.cin ;
assign \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.bin_s0  = ~ \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.b ;
always @(posedge \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.clk )
\sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.bin_s1  <= _197_;
always @(posedge \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.clk )
\sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.ain_s1  <= _196_;
always @(posedge \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.clk )
\sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.sum_s1  <= _199_;
always @(posedge \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.clk )
\sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.carry_s1  <= _198_;
assign _197_ = \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.ce  ? \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.bin_s0 [31:16] : \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.bin_s1 ;
assign _196_ = \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.ce  ? \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.a [31:16] : \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.ain_s1 ;
assign _198_ = \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.ce  ? \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.facout_s1  : \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.carry_s1 ;
assign _199_ = \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.ce  ? \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.fas_s1  : \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.sum_s1 ;
assign _200_ = \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.u1.a  + \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.u1.b ;
assign { \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.u1.cout , \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.u1.s  } = _200_ + \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.u1.cin ;
assign _201_ = \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.u2.a  + \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.u2.b ;
assign { \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.u2.cout , \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.u2.s  } = _201_ + \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.u2.cin ;
assign _202_ = op_7 > op_2;
assign _203_ = op_1[0] > op_2;
assign _204_ = | p_Result_s_reg_711;
assign _205_ = | trunc_ln851_reg_792;
assign op_6_V_fu_261_p2 = trunc_ln213_reg_658 | op_4[0];
assign or_ln340_fu_317_p2 = p_Result_3_reg_704 | overflow_fu_311_p2;
assign or_ln785_fu_302_p2 = newsignbit_reg_673 | icmp_ln768_reg_716;
always @(posedge ap_clk)
op_8_V_reg_761[18:0] <= 19'h00000;
always @(posedge ap_clk)
trunc_ln798_reg_918 <= _037_;
always @(posedge ap_clk)
trunc_ln798_1_reg_923 <= _036_;
always @(posedge ap_clk)
sh_reg_835 <= _031_;
always @(posedge ap_clk)
ret_V_9_reg_786 <= _026_;
always @(posedge ap_clk)
trunc_ln851_reg_792 <= _038_;
always @(posedge ap_clk)
sext_ln831_reg_797 <= _030_;
always @(posedge ap_clk)
ret_V_14_reg_906 <= _022_;
always @(posedge ap_clk)
ret_V_9_cast_reg_911 <= _025_;
always @(posedge ap_clk)
ret_V_11_reg_741 <= _019_;
always @(posedge ap_clk)
ret_1_reg_731 <= _018_;
always @(posedge ap_clk)
select_ln1192_reg_736 <= _028_;
always @(posedge ap_clk)
r_reg_933 <= _017_;
always @(posedge ap_clk)
ret_V_15_reg_938 <= _023_;
always @(posedge ap_clk)
p_Result_4_reg_820 <= _015_;
always @(posedge ap_clk)
ret_V_13_reg_825 <= _021_;
always @(posedge ap_clk)
select_ln69_reg_830 <= _029_;
always @(posedge ap_clk)
op_8_V_reg_761[19] <= _013_;
always @(posedge ap_clk)
ret_V_12_reg_776 <= _020_;
always @(posedge ap_clk)
tmp_2_reg_781 <= _033_;
always @(posedge ap_clk)
op_6_V_reg_699 <= _012_;
always @(posedge ap_clk)
p_Result_3_reg_704 <= _014_;
always @(posedge ap_clk)
p_Result_s_reg_711 <= _016_;
always @(posedge ap_clk)
ret_V_reg_881 <= _027_;
always @(posedge ap_clk)
op_16_V_reg_886 <= _010_;
always @(posedge ap_clk)
op_25_V_reg_891 <= _011_;
always @(posedge ap_clk)
trunc_ln213_reg_658 <= _034_;
always @(posedge ap_clk)
newsignbit_reg_673 <= _009_;
always @(posedge ap_clk)
lhs_V_4_reg_679 <= _008_;
always @(posedge ap_clk)
signbit_1_reg_684 <= _032_;
always @(posedge ap_clk)
trunc_ln728_reg_689 <= _035_;
always @(posedge ap_clk)
icmp_ln768_reg_716 <= _006_;
always @(posedge ap_clk)
ret_V_16_reg_958 <= _024_;
always @(posedge ap_clk)
add_ln69_3_reg_963 <= _003_;
always @(posedge ap_clk)
add_ln69_reg_856 <= _004_;
always @(posedge ap_clk)
add_ln69_1_reg_861 <= _002_;
always @(posedge ap_clk)
icmp_ln850_reg_804 <= _007_;
always @(posedge ap_clk)
add_ln691_reg_809 <= _001_;
always @(posedge ap_clk)
add_ln691_1_reg_928 <= _000_;
always @(posedge ap_clk)
ap_CS_fsm <= _005_;
assign _039_ = _043_ ? 2'h2 : 2'h1;
assign _206_ = ap_CS_fsm == 1'h1;
function [23:0] _569_;
input [23:0] a;
input [575:0] b;
input [23:0] s;
case (s)
24'b000000000000000000000001:
_569_ = b[23:0];
24'b000000000000000000000010:
_569_ = b[47:24];
24'b000000000000000000000100:
_569_ = b[71:48];
24'b000000000000000000001000:
_569_ = b[95:72];
24'b000000000000000000010000:
_569_ = b[119:96];
24'b000000000000000000100000:
_569_ = b[143:120];
24'b000000000000000001000000:
_569_ = b[167:144];
24'b000000000000000010000000:
_569_ = b[191:168];
24'b000000000000000100000000:
_569_ = b[215:192];
24'b000000000000001000000000:
_569_ = b[239:216];
24'b000000000000010000000000:
_569_ = b[263:240];
24'b000000000000100000000000:
_569_ = b[287:264];
24'b000000000001000000000000:
_569_ = b[311:288];
24'b000000000010000000000000:
_569_ = b[335:312];
24'b000000000100000000000000:
_569_ = b[359:336];
24'b000000001000000000000000:
_569_ = b[383:360];
24'b000000010000000000000000:
_569_ = b[407:384];
24'b000000100000000000000000:
_569_ = b[431:408];
24'b000001000000000000000000:
_569_ = b[455:432];
24'b000010000000000000000000:
_569_ = b[479:456];
24'b000100000000000000000000:
_569_ = b[503:480];
24'b001000000000000000000000:
_569_ = b[527:504];
24'b010000000000000000000000:
_569_ = b[551:528];
24'b100000000000000000000000:
_569_ = b[575:552];
24'b000000000000000000000000:
_569_ = a;
default:
_569_ = 24'bx;
endcase
endfunction
assign ap_NS_fsm = _569_(24'hxxxxxx, { 22'h000000, _039_, 552'h000004000008000010000020000040000080000100000200000400000800001000002000004000008000010000020000040000080000100000200000400000800000000001 }, { _206_, _229_, _228_, _227_, _226_, _225_, _224_, _223_, _222_, _221_, _220_, _219_, _218_, _217_, _216_, _215_, _214_, _213_, _212_, _211_, _210_, _209_, _208_, _207_ });
assign _207_ = ap_CS_fsm == 24'h800000;
assign _208_ = ap_CS_fsm == 23'h400000;
assign _209_ = ap_CS_fsm == 22'h200000;
assign _210_ = ap_CS_fsm == 21'h100000;
assign _211_ = ap_CS_fsm == 20'h80000;
assign _212_ = ap_CS_fsm == 19'h40000;
assign _213_ = ap_CS_fsm == 18'h20000;
assign _214_ = ap_CS_fsm == 17'h10000;
assign _215_ = ap_CS_fsm == 16'h8000;
assign _216_ = ap_CS_fsm == 15'h4000;
assign _217_ = ap_CS_fsm == 14'h2000;
assign _218_ = ap_CS_fsm == 13'h1000;
assign _219_ = ap_CS_fsm == 12'h800;
assign _220_ = ap_CS_fsm == 11'h400;
assign _221_ = ap_CS_fsm == 10'h200;
assign _222_ = ap_CS_fsm == 9'h100;
assign _223_ = ap_CS_fsm == 8'h80;
assign _224_ = ap_CS_fsm == 7'h40;
assign _225_ = ap_CS_fsm == 6'h20;
assign _226_ = ap_CS_fsm == 5'h10;
assign _227_ = ap_CS_fsm == 4'h8;
assign _228_ = ap_CS_fsm == 3'h4;
assign _229_ = ap_CS_fsm == 2'h2;
assign op_29_ap_vld = ap_CS_fsm[23] ? 1'h1 : 1'h0;
assign ap_idle = _042_ ? 1'h1 : 1'h0;
assign _037_ = _041_ ? grp_fu_509_p2[1:0] : trunc_ln798_reg_918;
assign _036_ = _040_ ? grp_fu_514_p2[1:0] : trunc_ln798_1_reg_923;
assign _031_ = ap_CS_fsm[11] ? grp_fu_425_p2 : sh_reg_835;
assign _030_ = ap_CS_fsm[8] ? { tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781 } : sext_ln831_reg_797;
assign _038_ = ap_CS_fsm[8] ? grp_fu_383_p2[18:0] : trunc_ln851_reg_792;
assign _026_ = ap_CS_fsm[8] ? grp_fu_383_p2 : ret_V_9_reg_786;
assign _025_ = ap_CS_fsm[16] ? grp_fu_567_p2[32:1] : ret_V_9_cast_reg_911;
assign _022_ = ap_CS_fsm[16] ? grp_fu_567_p2 : ret_V_14_reg_906;
assign _019_ = ap_CS_fsm[5] ? grp_fu_336_p2 : ret_V_11_reg_741;
assign _028_ = ap_CS_fsm[3] ? select_ln1192_fu_328_p3 : select_ln1192_reg_736;
assign _018_ = ap_CS_fsm[3] ? grp_fu_296_p2 : ret_1_reg_731;
assign _023_ = ap_CS_fsm[19] ? ret_V_15_fu_621_p3 : ret_V_15_reg_938;
assign _017_ = ap_CS_fsm[19] ? r_fu_596_p3 : r_reg_933;
assign _029_ = ap_CS_fsm[10] ? select_ln69_fu_479_p3 : select_ln69_reg_830;
assign _021_ = ap_CS_fsm[10] ? ret_V_13_fu_472_p3 : ret_V_13_reg_825;
assign _015_ = ap_CS_fsm[10] ? op_14[31] : p_Result_4_reg_820;
assign _033_ = ap_CS_fsm[7] ? grp_fu_355_p2[6:1] : tmp_2_reg_781;
assign _020_ = ap_CS_fsm[7] ? grp_fu_355_p2 : ret_V_12_reg_776;
assign _013_ = ap_CS_fsm[7] ? signbit_1_reg_684 : op_8_V_reg_761[19];
assign _016_ = ap_CS_fsm[1] ? grp_fu_221_p2[9:1] : p_Result_s_reg_711;
assign _014_ = ap_CS_fsm[1] ? grp_fu_221_p2[9] : p_Result_3_reg_704;
assign _012_ = ap_CS_fsm[1] ? op_6_V_fu_261_p2 : op_6_V_reg_699;
assign _011_ = ap_CS_fsm[14] ? grp_fu_538_p2 : op_25_V_reg_891;
assign _010_ = ap_CS_fsm[14] ? grp_fu_529_p2[21:18] : op_16_V_reg_886;
assign _027_ = ap_CS_fsm[14] ? grp_fu_529_p2 : ret_V_reg_881;
assign _035_ = ap_CS_fsm[0] ? op_7[2:0] : trunc_ln728_reg_689;
assign _032_ = ap_CS_fsm[0] ? signbit_1_fu_247_p2 : signbit_1_reg_684;
assign _008_ = ap_CS_fsm[0] ? lhs_V_4_fu_237_p2 : lhs_V_4_reg_679;
assign _009_ = ap_CS_fsm[0] ? newsignbit_fu_227_p2 : newsignbit_reg_673;
assign _034_ = ap_CS_fsm[0] ? op_2[0] : trunc_ln213_reg_658;
assign _006_ = ap_CS_fsm[2] ? icmp_ln768_fu_284_p2 : icmp_ln768_reg_716;
assign _003_ = ap_CS_fsm[21] ? grp_fu_643_p2 : add_ln69_3_reg_963;
assign _024_ = ap_CS_fsm[21] ? grp_fu_631_p2 : ret_V_16_reg_958;
assign _002_ = ap_CS_fsm[12] ? grp_fu_500_p2 : add_ln69_1_reg_861;
assign _004_ = ap_CS_fsm[12] ? grp_fu_495_p2 : add_ln69_reg_856;
assign _001_ = ap_CS_fsm[9] ? grp_fu_406_p2 : add_ln691_reg_809;
assign _007_ = ap_CS_fsm[9] ? icmp_ln850_fu_412_p2 : icmp_ln850_reg_804;
assign _000_ = ap_CS_fsm[18] ? grp_fu_583_p2 : add_ln691_1_reg_928;
assign _005_ = ap_rst ? 24'h000001 : ap_NS_fsm;
assign icmp_ln768_fu_284_p2 = _204_ ? 1'h1 : 1'h0;
assign icmp_ln850_fu_412_p2 = _205_ ? 1'h1 : 1'h0;
assign lhs_V_4_fu_237_p2 = _202_ ? 1'h1 : 1'h0;
assign op_10_V_fu_322_p3 = or_ln340_fu_317_p2 ? p_Result_3_reg_704 : newsignbit_reg_673;
assign r_fu_596_p3 = p_Result_4_reg_820 ? trunc_ln798_reg_918 : trunc_ln798_1_reg_923;
assign ret_V_13_fu_472_p3 = ret_V_12_reg_776[6] ? select_ln850_fu_466_p3 : sext_ln831_reg_797;
assign ret_V_15_fu_621_p3 = ret_V_14_reg_906[33] ? select_ln850_1_fu_615_p3 : ret_V_9_cast_reg_911;
assign select_ln1192_fu_328_p3 = op_10_V_fu_322_p3 ? 5'h1f : 5'h00;
assign select_ln69_fu_479_p3 = ret_V_10_fu_450_p2 ? 3'h7 : 3'h0;
assign select_ln850_1_fu_615_p3 = ret_V_reg_881[18] ? add_ln691_1_reg_928 : ret_V_9_cast_reg_911;
assign select_ln850_fu_466_p3 = op_11[0] ? add_ln691_reg_809 : sext_ln831_reg_797;
assign signbit_1_fu_247_p2 = _203_ ? 1'h1 : 1'h0;
assign newsignbit_fu_227_p2 = op_5[0] ^ op_7[0];
assign ret_V_10_fu_450_p2 = ret_V_9_reg_786[19] ^ and_ln353_fu_445_p2;
assign ap_CS_fsm_state1 = ap_CS_fsm[0];
assign ap_CS_fsm_state10 = ap_CS_fsm[9];
assign ap_CS_fsm_state11 = ap_CS_fsm[10];
assign ap_CS_fsm_state12 = ap_CS_fsm[11];
assign ap_CS_fsm_state13 = ap_CS_fsm[12];
assign ap_CS_fsm_state14 = ap_CS_fsm[13];
assign ap_CS_fsm_state15 = ap_CS_fsm[14];
assign ap_CS_fsm_state16 = ap_CS_fsm[15];
assign ap_CS_fsm_state17 = ap_CS_fsm[16];
assign ap_CS_fsm_state18 = ap_CS_fsm[17];
assign ap_CS_fsm_state19 = ap_CS_fsm[18];
assign ap_CS_fsm_state2 = ap_CS_fsm[1];
assign ap_CS_fsm_state20 = ap_CS_fsm[19];
assign ap_CS_fsm_state21 = ap_CS_fsm[20];
assign ap_CS_fsm_state22 = ap_CS_fsm[21];
assign ap_CS_fsm_state23 = ap_CS_fsm[22];
assign ap_CS_fsm_state24 = ap_CS_fsm[23];
assign ap_CS_fsm_state3 = ap_CS_fsm[2];
assign ap_CS_fsm_state4 = ap_CS_fsm[3];
assign ap_CS_fsm_state5 = ap_CS_fsm[4];
assign ap_CS_fsm_state6 = ap_CS_fsm[5];
assign ap_CS_fsm_state7 = ap_CS_fsm[6];
assign ap_CS_fsm_state8 = ap_CS_fsm[7];
assign ap_CS_fsm_state9 = ap_CS_fsm[8];
assign ap_done = op_29_ap_vld;
assign ap_ready = op_29_ap_vld;
assign grp_fu_221_p0 = { 2'h0, op_7 };
assign grp_fu_221_p1 = { op_5[7], op_5[7], op_5 };
assign grp_fu_296_p0 = { op_0[3], op_0 };
assign grp_fu_296_p1 = { 4'h0, op_6_V_reg_699 };
assign grp_fu_355_p0 = { ret_V_11_reg_741[4], ret_V_11_reg_741, 1'h0 };
assign grp_fu_355_p1 = { op_11[1], op_11[1], op_11[1], op_11[1], op_11[1], op_11 };
assign grp_fu_383_p0 = { op_4[7], op_4, 19'h00000 };
assign grp_fu_383_p1 = { 8'h00, signbit_1_reg_684, 19'h00000 };
assign grp_fu_406_p0 = { tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781 };
assign grp_fu_495_p1 = { op_15[15], op_15[15], op_15[15], op_15[15], op_15[15], op_15[15], op_15[15], op_15[15], op_15[15], op_15[15], op_15[15], op_15[15], op_15[15], op_15[15], op_15[15], op_15[15], op_15 };
assign grp_fu_500_p0 = { op_12[1], op_12 };
assign grp_fu_529_p0 = { trunc_ln728_reg_689, 19'h00000 };
assign grp_fu_529_p1 = { 2'h0, op_8_V_reg_761 };
assign grp_fu_538_p0 = { add_ln69_1_reg_861[2], add_ln69_1_reg_861[2], add_ln69_1_reg_861[2], add_ln69_1_reg_861[2], add_ln69_1_reg_861[2], add_ln69_1_reg_861[2], add_ln69_1_reg_861[2], add_ln69_1_reg_861[2], add_ln69_1_reg_861[2], add_ln69_1_reg_861[2], add_ln69_1_reg_861[2], add_ln69_1_reg_861[2], add_ln69_1_reg_861[2], add_ln69_1_reg_861[2], add_ln69_1_reg_861[2], add_ln69_1_reg_861[2], add_ln69_1_reg_861[2], add_ln69_1_reg_861[2], add_ln69_1_reg_861[2], add_ln69_1_reg_861[2], add_ln69_1_reg_861[2], add_ln69_1_reg_861[2], add_ln69_1_reg_861[2], add_ln69_1_reg_861[2], add_ln69_1_reg_861[2], add_ln69_1_reg_861[2], add_ln69_1_reg_861[2], add_ln69_1_reg_861[2], add_ln69_1_reg_861[2], add_ln69_1_reg_861 };
assign grp_fu_567_p0 = { op_25_V_reg_891[31], op_25_V_reg_891, 1'h0 };
assign grp_fu_567_p1 = { op_16_V_reg_886[3], op_16_V_reg_886[3], op_16_V_reg_886[3], op_16_V_reg_886[3], op_16_V_reg_886[3], op_16_V_reg_886[3], op_16_V_reg_886[3], op_16_V_reg_886[3], op_16_V_reg_886[3], op_16_V_reg_886[3], op_16_V_reg_886[3], op_16_V_reg_886[3], op_16_V_reg_886[3], op_16_V_reg_886[3], op_16_V_reg_886[3], op_16_V_reg_886[3], op_16_V_reg_886[3], op_16_V_reg_886[3], op_16_V_reg_886[3], op_16_V_reg_886[3], op_16_V_reg_886[3], op_16_V_reg_886[3], op_16_V_reg_886[3], op_16_V_reg_886[3], op_16_V_reg_886[3], op_16_V_reg_886[3], op_16_V_reg_886[3], op_16_V_reg_886[3], op_16_V_reg_886[3], op_16_V_reg_886[3], op_16_V_reg_886 };
assign grp_fu_631_p1 = { 31'h00000000, lhs_V_4_reg_679 };
assign grp_fu_643_p0 = { op_19[15], op_19 };
assign grp_fu_643_p1 = { r_reg_933[1], r_reg_933[1], r_reg_933[1], r_reg_933[1], r_reg_933[1], r_reg_933[1], r_reg_933[1], r_reg_933[1], r_reg_933[1], r_reg_933[1], r_reg_933[1], r_reg_933[1], r_reg_933[1], r_reg_933[1], r_reg_933[1], r_reg_933 };
assign grp_fu_652_p0 = { add_ln69_3_reg_963[16], add_ln69_3_reg_963[16], add_ln69_3_reg_963[16], add_ln69_3_reg_963[16], add_ln69_3_reg_963[16], add_ln69_3_reg_963[16], add_ln69_3_reg_963[16], add_ln69_3_reg_963[16], add_ln69_3_reg_963[16], add_ln69_3_reg_963[16], add_ln69_3_reg_963[16], add_ln69_3_reg_963[16], add_ln69_3_reg_963[16], add_ln69_3_reg_963[16], add_ln69_3_reg_963[16], add_ln69_3_reg_963 };
assign lhs_V_fu_368_p3 = { op_4, 19'h00000 };
assign op_29 = grp_fu_652_p2;
assign op_3_V_fu_197_p1 = op_1[0];
assign op_8_V_fu_361_p3 = { signbit_1_reg_684, 19'h00000 };
assign p_Result_1_fu_456_p3 = ret_V_12_reg_776[6];
assign p_Result_2_fu_601_p3 = ret_V_14_reg_906[33];
assign p_Result_s_12_fu_438_p3 = ret_V_9_reg_786[27];
assign rhs_4_fu_556_p3 = { op_25_V_reg_891, 1'h0 };
assign sext_ln1192_fu_340_p0 = op_11;
assign sext_ln215_fu_205_p0 = op_5;
assign sext_ln781_fu_505_p1 = { op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9 };
assign sext_ln831_fu_403_p1 = { tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781 };
assign tmp_4_fu_344_p3 = { ret_V_11_reg_741, 1'h0 };
assign tmp_6_fu_608_p3 = ret_V_reg_881[18];
assign tmp_fu_431_p3 = ret_V_9_reg_786[19];
assign trunc_ln1346_1_fu_217_p1 = op_7[0];
assign trunc_ln1346_fu_213_p0 = op_5;
assign trunc_ln1346_fu_213_p1 = op_5[0];
assign trunc_ln213_1_fu_257_p1 = op_4[0];
assign trunc_ln213_fu_201_p1 = op_2[0];
assign trunc_ln728_fu_253_p1 = op_7[2:0];
assign trunc_ln798_1_fu_592_p1 = grp_fu_514_p2[1:0];
assign trunc_ln798_fu_588_p1 = grp_fu_509_p2[1:0];
assign trunc_ln851_1_fu_463_p0 = op_11;
assign trunc_ln851_1_fu_463_p1 = op_11[0];
assign trunc_ln851_fu_399_p1 = grp_fu_383_p2[18:0];
assign zext_ln878_1_fu_243_p1 = { 15'h0000, op_1[0] };
assign zext_ln878_fu_233_p1 = { 8'h00, op_7 };
assign \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.ain_s0  = \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.a ;
assign \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.s  = { \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.fas_s2 , \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.sum_s1  };
assign \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.u2.a  = \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.ain_s1 ;
assign \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.u2.b  = \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.bin_s1 ;
assign \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.u2.cin  = \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.carry_s1 ;
assign \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.facout_s2  = \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.u2.cout ;
assign \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.fas_s2  = \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.u2.s ;
assign \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.u1.a  = \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.a [15:0];
assign \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.u1.b  = \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.bin_s0 [15:0];
assign \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.u1.cin  = 1'h1;
assign \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.facout_s1  = \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.u1.cout ;
assign \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.fas_s1  = \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.u1.s ;
assign \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.a  = \sub_32ns_32ns_32_2_1_U7.din0 ;
assign \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.b  = \sub_32ns_32ns_32_2_1_U7.din1 ;
assign \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.ce  = \sub_32ns_32ns_32_2_1_U7.ce ;
assign \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.clk  = \sub_32ns_32ns_32_2_1_U7.clk ;
assign \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.reset  = \sub_32ns_32ns_32_2_1_U7.reset ;
assign \sub_32ns_32ns_32_2_1_U7.dout  = \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.s ;
assign \sub_32ns_32ns_32_2_1_U7.ce  = 1'h1;
assign \sub_32ns_32ns_32_2_1_U7.clk  = ap_clk;
assign \sub_32ns_32ns_32_2_1_U7.din0  = 32'd0;
assign \sub_32ns_32ns_32_2_1_U7.din1  = op_14;
assign grp_fu_425_p2 = \sub_32ns_32ns_32_2_1_U7.dout ;
assign \sub_32ns_32ns_32_2_1_U7.reset  = ap_rst;
assign \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.ain_s0  = \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.a ;
assign \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.s  = { \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.fas_s2 , \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.sum_s1  };
assign \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.u2.a  = \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.ain_s1 ;
assign \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.u2.b  = \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.bin_s1 ;
assign \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.u2.cin  = \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.carry_s1 ;
assign \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.facout_s2  = \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.u2.cout ;
assign \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.fas_s2  = \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.u2.s ;
assign \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.u1.a  = \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.a [13:0];
assign \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.u1.b  = \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.bin_s0 [13:0];
assign \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.u1.cin  = 1'h1;
assign \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.facout_s1  = \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.u1.cout ;
assign \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.fas_s1  = \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.u1.s ;
assign \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.a  = \sub_28s_28ns_28_2_1_U5.din0 ;
assign \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.b  = \sub_28s_28ns_28_2_1_U5.din1 ;
assign \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.ce  = \sub_28s_28ns_28_2_1_U5.ce ;
assign \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.clk  = \sub_28s_28ns_28_2_1_U5.clk ;
assign \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.reset  = \sub_28s_28ns_28_2_1_U5.reset ;
assign \sub_28s_28ns_28_2_1_U5.dout  = \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.s ;
assign \sub_28s_28ns_28_2_1_U5.ce  = 1'h1;
assign \sub_28s_28ns_28_2_1_U5.clk  = ap_clk;
assign \sub_28s_28ns_28_2_1_U5.din0  = { op_4[7], op_4, 19'h00000 };
assign \sub_28s_28ns_28_2_1_U5.din1  = { 8'h00, signbit_1_reg_684, 19'h00000 };
assign grp_fu_383_p2 = \sub_28s_28ns_28_2_1_U5.dout ;
assign \sub_28s_28ns_28_2_1_U5.reset  = ap_rst;
assign \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.ain_s0  = \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.a ;
assign \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.s  = { \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.fas_s2 , \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.sum_s1  };
assign \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.u2.a  = \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.ain_s1 ;
assign \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.u2.b  = \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.bin_s1 ;
assign \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.u2.cin  = \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.carry_s1 ;
assign \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.facout_s2  = \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.u2.cout ;
assign \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.fas_s2  = \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.u2.s ;
assign \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.u1.a  = \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.a [10:0];
assign \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.u1.b  = \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.bin_s0 [10:0];
assign \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.u1.cin  = 1'h1;
assign \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.facout_s1  = \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.u1.cout ;
assign \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.fas_s1  = \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.u1.s ;
assign \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.a  = \sub_22ns_22ns_22_2_1_U12.din0 ;
assign \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.b  = \sub_22ns_22ns_22_2_1_U12.din1 ;
assign \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.ce  = \sub_22ns_22ns_22_2_1_U12.ce ;
assign \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.clk  = \sub_22ns_22ns_22_2_1_U12.clk ;
assign \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.reset  = \sub_22ns_22ns_22_2_1_U12.reset ;
assign \sub_22ns_22ns_22_2_1_U12.dout  = \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.s ;
assign \sub_22ns_22ns_22_2_1_U12.ce  = 1'h1;
assign \sub_22ns_22ns_22_2_1_U12.clk  = ap_clk;
assign \sub_22ns_22ns_22_2_1_U12.din0  = { trunc_ln728_reg_689, 19'h00000 };
assign \sub_22ns_22ns_22_2_1_U12.din1  = { 2'h0, op_8_V_reg_761 };
assign grp_fu_529_p2 = \sub_22ns_22ns_22_2_1_U12.dout ;
assign \sub_22ns_22ns_22_2_1_U12.reset  = ap_rst;
assign \shl_32s_32ns_32_7_1_U11.din1_cast  = \shl_32s_32ns_32_7_1_U11.din1 ;
assign \shl_32s_32ns_32_7_1_U11.din1_mask  = 32'd31;
assign \shl_32s_32ns_32_7_1_U11.ce  = 1'h1;
assign \shl_32s_32ns_32_7_1_U11.clk  = ap_clk;
assign \shl_32s_32ns_32_7_1_U11.din0  = { op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9 };
assign \shl_32s_32ns_32_7_1_U11.din1  = op_14;
assign grp_fu_514_p2 = \shl_32s_32ns_32_7_1_U11.dout ;
assign \shl_32s_32ns_32_7_1_U11.reset  = ap_rst;
assign \ashr_32s_32ns_32_7_1_U10.din1_cast  = \ashr_32s_32ns_32_7_1_U10.din1 ;
assign \ashr_32s_32ns_32_7_1_U10.din1_mask  = 32'd31;
assign \ashr_32s_32ns_32_7_1_U10.ce  = 1'h1;
assign \ashr_32s_32ns_32_7_1_U10.clk  = ap_clk;
assign \ashr_32s_32ns_32_7_1_U10.din0  = { op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9 };
assign \ashr_32s_32ns_32_7_1_U10.din1  = sh_reg_835;
assign grp_fu_509_p2 = \ashr_32s_32ns_32_7_1_U10.dout ;
assign \ashr_32s_32ns_32_7_1_U10.reset  = ap_rst;
assign \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.ain_s0  = \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.a ;
assign \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.bin_s0  = \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.b ;
assign \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.s  = { \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.fas_s2 , \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.sum_s1  };
assign \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.u2.a  = \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.ain_s1 ;
assign \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.u2.b  = \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.bin_s1 ;
assign \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.u2.cin  = \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.carry_s1 ;
assign \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.facout_s2  = \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.u2.cout ;
assign \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.fas_s2  = \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.u2.s ;
assign \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.u1.a  = \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.a [2:0];
assign \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.u1.b  = \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.b [2:0];
assign \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.u1.cin  = 1'h0;
assign \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.facout_s1  = \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.u1.cout ;
assign \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.fas_s1  = \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.u1.s ;
assign \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.a  = \add_7s_7s_7_2_1_U4.din0 ;
assign \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.b  = \add_7s_7s_7_2_1_U4.din1 ;
assign \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.ce  = \add_7s_7s_7_2_1_U4.ce ;
assign \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.clk  = \add_7s_7s_7_2_1_U4.clk ;
assign \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.reset  = \add_7s_7s_7_2_1_U4.reset ;
assign \add_7s_7s_7_2_1_U4.dout  = \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.s ;
assign \add_7s_7s_7_2_1_U4.ce  = 1'h1;
assign \add_7s_7s_7_2_1_U4.clk  = ap_clk;
assign \add_7s_7s_7_2_1_U4.din0  = { ret_V_11_reg_741[4], ret_V_11_reg_741, 1'h0 };
assign \add_7s_7s_7_2_1_U4.din1  = { op_11[1], op_11[1], op_11[1], op_11[1], op_11[1], op_11 };
assign grp_fu_355_p2 = \add_7s_7s_7_2_1_U4.dout ;
assign \add_7s_7s_7_2_1_U4.reset  = ap_rst;
assign \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.ain_s0  = \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.a ;
assign \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.bin_s0  = \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.b ;
assign \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.s  = { \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.fas_s2 , \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.sum_s1  };
assign \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.u2.a  = \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.ain_s1 ;
assign \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.u2.b  = \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.bin_s1 ;
assign \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.u2.cin  = \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.carry_s1 ;
assign \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.facout_s2  = \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.u2.cout ;
assign \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.fas_s2  = \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.u2.s ;
assign \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.u1.a  = \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.a [1:0];
assign \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.u1.b  = \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.b [1:0];
assign \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.u1.cin  = 1'h0;
assign \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.facout_s1  = \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.u1.cout ;
assign \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.fas_s1  = \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.u1.s ;
assign \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.a  = \add_5s_5ns_5_2_1_U2.din0 ;
assign \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.b  = \add_5s_5ns_5_2_1_U2.din1 ;
assign \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.ce  = \add_5s_5ns_5_2_1_U2.ce ;
assign \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.clk  = \add_5s_5ns_5_2_1_U2.clk ;
assign \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.reset  = \add_5s_5ns_5_2_1_U2.reset ;
assign \add_5s_5ns_5_2_1_U2.dout  = \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.s ;
assign \add_5s_5ns_5_2_1_U2.ce  = 1'h1;
assign \add_5s_5ns_5_2_1_U2.clk  = ap_clk;
assign \add_5s_5ns_5_2_1_U2.din0  = { op_0[3], op_0 };
assign \add_5s_5ns_5_2_1_U2.din1  = { 4'h0, op_6_V_reg_699 };
assign grp_fu_296_p2 = \add_5s_5ns_5_2_1_U2.dout ;
assign \add_5s_5ns_5_2_1_U2.reset  = ap_rst;
assign \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.ain_s0  = \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.a ;
assign \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.bin_s0  = \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.b ;
assign \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.s  = { \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.fas_s2 , \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.sum_s1  };
assign \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.u2.a  = \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.ain_s1 ;
assign \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.u2.b  = \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.bin_s1 ;
assign \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.u2.cin  = \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.carry_s1 ;
assign \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.facout_s2  = \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.u2.cout ;
assign \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.fas_s2  = \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.u2.s ;
assign \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.u1.a  = \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.a [1:0];
assign \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.u1.b  = \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.b [1:0];
assign \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.u1.cin  = 1'h0;
assign \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.facout_s1  = \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.u1.cout ;
assign \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.fas_s1  = \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.u1.s ;
assign \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.a  = \add_5ns_5ns_5_2_1_U3.din0 ;
assign \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.b  = \add_5ns_5ns_5_2_1_U3.din1 ;
assign \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.ce  = \add_5ns_5ns_5_2_1_U3.ce ;
assign \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.clk  = \add_5ns_5ns_5_2_1_U3.clk ;
assign \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.reset  = \add_5ns_5ns_5_2_1_U3.reset ;
assign \add_5ns_5ns_5_2_1_U3.dout  = \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.s ;
assign \add_5ns_5ns_5_2_1_U3.ce  = 1'h1;
assign \add_5ns_5ns_5_2_1_U3.clk  = ap_clk;
assign \add_5ns_5ns_5_2_1_U3.din0  = ret_1_reg_731;
assign \add_5ns_5ns_5_2_1_U3.din1  = select_ln1192_reg_736;
assign grp_fu_336_p2 = \add_5ns_5ns_5_2_1_U3.dout ;
assign \add_5ns_5ns_5_2_1_U3.reset  = ap_rst;
assign \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.ain_s0  = \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.a ;
assign \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.bin_s0  = \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.b ;
assign \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.s  = { \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.fas_s2 , \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.sum_s1  };
assign \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.u2.a  = \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.ain_s1 ;
assign \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.u2.b  = \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.bin_s1 ;
assign \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.u2.cin  = \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.carry_s1 ;
assign \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.facout_s2  = \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.u2.cout ;
assign \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.fas_s2  = \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.u2.s ;
assign \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.u1.a  = \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.a [0];
assign \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.u1.b  = \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.b [0];
assign \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.u1.cin  = 1'h0;
assign \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.facout_s1  = \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.u1.cout ;
assign \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.fas_s1  = \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.u1.s ;
assign \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.a  = \add_3s_3ns_3_2_1_U9.din0 ;
assign \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.b  = \add_3s_3ns_3_2_1_U9.din1 ;
assign \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.ce  = \add_3s_3ns_3_2_1_U9.ce ;
assign \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.clk  = \add_3s_3ns_3_2_1_U9.clk ;
assign \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.reset  = \add_3s_3ns_3_2_1_U9.reset ;
assign \add_3s_3ns_3_2_1_U9.dout  = \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.s ;
assign \add_3s_3ns_3_2_1_U9.ce  = 1'h1;
assign \add_3s_3ns_3_2_1_U9.clk  = ap_clk;
assign \add_3s_3ns_3_2_1_U9.din0  = { op_12[1], op_12 };
assign \add_3s_3ns_3_2_1_U9.din1  = select_ln69_reg_830;
assign grp_fu_500_p2 = \add_3s_3ns_3_2_1_U9.dout ;
assign \add_3s_3ns_3_2_1_U9.reset  = ap_rst;
assign \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.ain_s0  = \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.a ;
assign \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.bin_s0  = \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.b ;
assign \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.s  = { \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.fas_s2 , \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.sum_s1  };
assign \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.u2.a  = \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.ain_s1 ;
assign \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.u2.b  = \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.bin_s1 ;
assign \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.u2.cin  = \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.carry_s1 ;
assign \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.facout_s2  = \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.u2.cout ;
assign \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.fas_s2  = \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.u2.s ;
assign \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.u1.a  = \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.a [16:0];
assign \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.u1.b  = \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.b [16:0];
assign \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.u1.cin  = 1'h0;
assign \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.facout_s1  = \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.u1.cout ;
assign \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.fas_s1  = \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.u1.s ;
assign \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.a  = \add_34s_34s_34_2_1_U14.din0 ;
assign \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.b  = \add_34s_34s_34_2_1_U14.din1 ;
assign \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.ce  = \add_34s_34s_34_2_1_U14.ce ;
assign \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.clk  = \add_34s_34s_34_2_1_U14.clk ;
assign \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.reset  = \add_34s_34s_34_2_1_U14.reset ;
assign \add_34s_34s_34_2_1_U14.dout  = \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.s ;
assign \add_34s_34s_34_2_1_U14.ce  = 1'h1;
assign \add_34s_34s_34_2_1_U14.clk  = ap_clk;
assign \add_34s_34s_34_2_1_U14.din0  = { op_25_V_reg_891[31], op_25_V_reg_891, 1'h0 };
assign \add_34s_34s_34_2_1_U14.din1  = { op_16_V_reg_886[3], op_16_V_reg_886[3], op_16_V_reg_886[3], op_16_V_reg_886[3], op_16_V_reg_886[3], op_16_V_reg_886[3], op_16_V_reg_886[3], op_16_V_reg_886[3], op_16_V_reg_886[3], op_16_V_reg_886[3], op_16_V_reg_886[3], op_16_V_reg_886[3], op_16_V_reg_886[3], op_16_V_reg_886[3], op_16_V_reg_886[3], op_16_V_reg_886[3], op_16_V_reg_886[3], op_16_V_reg_886[3], op_16_V_reg_886[3], op_16_V_reg_886[3], op_16_V_reg_886[3], op_16_V_reg_886[3], op_16_V_reg_886[3], op_16_V_reg_886[3], op_16_V_reg_886[3], op_16_V_reg_886[3], op_16_V_reg_886[3], op_16_V_reg_886[3], op_16_V_reg_886[3], op_16_V_reg_886[3], op_16_V_reg_886 };
assign grp_fu_567_p2 = \add_34s_34s_34_2_1_U14.dout ;
assign \add_34s_34s_34_2_1_U14.reset  = ap_rst;
assign \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.ain_s0  = \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.a ;
assign \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.bin_s0  = \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.b ;
assign \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.s  = { \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.fas_s2 , \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.sum_s1  };
assign \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.u2.a  = \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.ain_s1 ;
assign \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.u2.b  = \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.bin_s1 ;
assign \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.u2.cin  = \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.carry_s1 ;
assign \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.facout_s2  = \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.u2.cout ;
assign \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.fas_s2  = \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.u2.s ;
assign \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.u1.a  = \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.a [15:0];
assign \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.u1.b  = \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.b [15:0];
assign \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.u1.cin  = 1'h0;
assign \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.facout_s1  = \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.u1.cout ;
assign \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.fas_s1  = \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.u1.s ;
assign \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.a  = \add_32s_32ns_32_2_1_U6.din0 ;
assign \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.b  = \add_32s_32ns_32_2_1_U6.din1 ;
assign \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.ce  = \add_32s_32ns_32_2_1_U6.ce ;
assign \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.clk  = \add_32s_32ns_32_2_1_U6.clk ;
assign \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.reset  = \add_32s_32ns_32_2_1_U6.reset ;
assign \add_32s_32ns_32_2_1_U6.dout  = \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.s ;
assign \add_32s_32ns_32_2_1_U6.ce  = 1'h1;
assign \add_32s_32ns_32_2_1_U6.clk  = ap_clk;
assign \add_32s_32ns_32_2_1_U6.din0  = { tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781 };
assign \add_32s_32ns_32_2_1_U6.din1  = 32'd1;
assign grp_fu_406_p2 = \add_32s_32ns_32_2_1_U6.dout ;
assign \add_32s_32ns_32_2_1_U6.reset  = ap_rst;
assign \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.ain_s0  = \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.a ;
assign \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.bin_s0  = \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.b ;
assign \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.s  = { \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.fas_s2 , \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.sum_s1  };
assign \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.u2.a  = \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.ain_s1 ;
assign \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.u2.b  = \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.bin_s1 ;
assign \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.u2.cin  = \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.carry_s1 ;
assign \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.facout_s2  = \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.u2.cout ;
assign \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.fas_s2  = \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.u2.s ;
assign \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.u1.a  = \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.a [15:0];
assign \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.u1.b  = \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.b [15:0];
assign \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.u1.cin  = 1'h0;
assign \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.facout_s1  = \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.u1.cout ;
assign \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.fas_s1  = \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.u1.s ;
assign \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.a  = \add_32s_32ns_32_2_1_U18.din0 ;
assign \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.b  = \add_32s_32ns_32_2_1_U18.din1 ;
assign \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.ce  = \add_32s_32ns_32_2_1_U18.ce ;
assign \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.clk  = \add_32s_32ns_32_2_1_U18.clk ;
assign \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.reset  = \add_32s_32ns_32_2_1_U18.reset ;
assign \add_32s_32ns_32_2_1_U18.dout  = \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.s ;
assign \add_32s_32ns_32_2_1_U18.ce  = 1'h1;
assign \add_32s_32ns_32_2_1_U18.clk  = ap_clk;
assign \add_32s_32ns_32_2_1_U18.din0  = { add_ln69_3_reg_963[16], add_ln69_3_reg_963[16], add_ln69_3_reg_963[16], add_ln69_3_reg_963[16], add_ln69_3_reg_963[16], add_ln69_3_reg_963[16], add_ln69_3_reg_963[16], add_ln69_3_reg_963[16], add_ln69_3_reg_963[16], add_ln69_3_reg_963[16], add_ln69_3_reg_963[16], add_ln69_3_reg_963[16], add_ln69_3_reg_963[16], add_ln69_3_reg_963[16], add_ln69_3_reg_963[16], add_ln69_3_reg_963 };
assign \add_32s_32ns_32_2_1_U18.din1  = ret_V_16_reg_958;
assign grp_fu_652_p2 = \add_32s_32ns_32_2_1_U18.dout ;
assign \add_32s_32ns_32_2_1_U18.reset  = ap_rst;
assign \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.ain_s0  = \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.a ;
assign \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.bin_s0  = \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.b ;
assign \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.s  = { \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.fas_s2 , \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.sum_s1  };
assign \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.u2.a  = \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.ain_s1 ;
assign \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.u2.b  = \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.bin_s1 ;
assign \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.u2.cin  = \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.carry_s1 ;
assign \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.facout_s2  = \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.u2.cout ;
assign \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.fas_s2  = \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.u2.s ;
assign \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.u1.a  = \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.a [15:0];
assign \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.u1.b  = \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.b [15:0];
assign \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.u1.cin  = 1'h0;
assign \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.facout_s1  = \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.u1.cout ;
assign \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.fas_s1  = \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.u1.s ;
assign \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.a  = \add_32s_32ns_32_2_1_U13.din0 ;
assign \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.b  = \add_32s_32ns_32_2_1_U13.din1 ;
assign \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.ce  = \add_32s_32ns_32_2_1_U13.ce ;
assign \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.clk  = \add_32s_32ns_32_2_1_U13.clk ;
assign \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.reset  = \add_32s_32ns_32_2_1_U13.reset ;
assign \add_32s_32ns_32_2_1_U13.dout  = \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.s ;
assign \add_32s_32ns_32_2_1_U13.ce  = 1'h1;
assign \add_32s_32ns_32_2_1_U13.clk  = ap_clk;
assign \add_32s_32ns_32_2_1_U13.din0  = { add_ln69_1_reg_861[2], add_ln69_1_reg_861[2], add_ln69_1_reg_861[2], add_ln69_1_reg_861[2], add_ln69_1_reg_861[2], add_ln69_1_reg_861[2], add_ln69_1_reg_861[2], add_ln69_1_reg_861[2], add_ln69_1_reg_861[2], add_ln69_1_reg_861[2], add_ln69_1_reg_861[2], add_ln69_1_reg_861[2], add_ln69_1_reg_861[2], add_ln69_1_reg_861[2], add_ln69_1_reg_861[2], add_ln69_1_reg_861[2], add_ln69_1_reg_861[2], add_ln69_1_reg_861[2], add_ln69_1_reg_861[2], add_ln69_1_reg_861[2], add_ln69_1_reg_861[2], add_ln69_1_reg_861[2], add_ln69_1_reg_861[2], add_ln69_1_reg_861[2], add_ln69_1_reg_861[2], add_ln69_1_reg_861[2], add_ln69_1_reg_861[2], add_ln69_1_reg_861[2], add_ln69_1_reg_861[2], add_ln69_1_reg_861 };
assign \add_32s_32ns_32_2_1_U13.din1  = add_ln69_reg_856;
assign grp_fu_538_p2 = \add_32s_32ns_32_2_1_U13.dout ;
assign \add_32s_32ns_32_2_1_U13.reset  = ap_rst;
assign \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.ain_s0  = \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.a ;
assign \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.bin_s0  = \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.b ;
assign \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.s  = { \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.fas_s2 , \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.sum_s1  };
assign \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.u2.a  = \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.ain_s1 ;
assign \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.u2.b  = \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.bin_s1 ;
assign \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.u2.cin  = \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.carry_s1 ;
assign \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.facout_s2  = \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.u2.cout ;
assign \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.fas_s2  = \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.u2.s ;
assign \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.u1.a  = \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.a [15:0];
assign \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.u1.b  = \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.b [15:0];
assign \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.u1.cin  = 1'h0;
assign \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.facout_s1  = \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.u1.cout ;
assign \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.fas_s1  = \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.u1.s ;
assign \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.a  = \add_32ns_32s_32_2_1_U8.din0 ;
assign \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.b  = \add_32ns_32s_32_2_1_U8.din1 ;
assign \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.ce  = \add_32ns_32s_32_2_1_U8.ce ;
assign \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.clk  = \add_32ns_32s_32_2_1_U8.clk ;
assign \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.reset  = \add_32ns_32s_32_2_1_U8.reset ;
assign \add_32ns_32s_32_2_1_U8.dout  = \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.s ;
assign \add_32ns_32s_32_2_1_U8.ce  = 1'h1;
assign \add_32ns_32s_32_2_1_U8.clk  = ap_clk;
assign \add_32ns_32s_32_2_1_U8.din0  = ret_V_13_reg_825;
assign \add_32ns_32s_32_2_1_U8.din1  = { op_15[15], op_15[15], op_15[15], op_15[15], op_15[15], op_15[15], op_15[15], op_15[15], op_15[15], op_15[15], op_15[15], op_15[15], op_15[15], op_15[15], op_15[15], op_15[15], op_15 };
assign grp_fu_495_p2 = \add_32ns_32s_32_2_1_U8.dout ;
assign \add_32ns_32s_32_2_1_U8.reset  = ap_rst;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.ain_s0  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.a ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.bin_s0  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.b ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.s  = { \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.fas_s2 , \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.sum_s1  };
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.a  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.ain_s1 ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.b  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.bin_s1 ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.cin  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.carry_s1 ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.facout_s2  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.cout ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.fas_s2  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.s ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.a  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.a [15:0];
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.b  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.b [15:0];
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.cin  = 1'h0;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.facout_s1  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.cout ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.fas_s1  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.s ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.a  = \add_32ns_32ns_32_2_1_U16.din0 ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.b  = \add_32ns_32ns_32_2_1_U16.din1 ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.ce  = \add_32ns_32ns_32_2_1_U16.ce ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.clk  = \add_32ns_32ns_32_2_1_U16.clk ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.reset  = \add_32ns_32ns_32_2_1_U16.reset ;
assign \add_32ns_32ns_32_2_1_U16.dout  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.s ;
assign \add_32ns_32ns_32_2_1_U16.ce  = 1'h1;
assign \add_32ns_32ns_32_2_1_U16.clk  = ap_clk;
assign \add_32ns_32ns_32_2_1_U16.din0  = ret_V_15_reg_938;
assign \add_32ns_32ns_32_2_1_U16.din1  = { 31'h00000000, lhs_V_4_reg_679 };
assign grp_fu_631_p2 = \add_32ns_32ns_32_2_1_U16.dout ;
assign \add_32ns_32ns_32_2_1_U16.reset  = ap_rst;
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.ain_s0  = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.a ;
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.bin_s0  = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.b ;
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.s  = { \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.fas_s2 , \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.sum_s1  };
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.a  = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.ain_s1 ;
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.b  = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.bin_s1 ;
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.cin  = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.carry_s1 ;
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.facout_s2  = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.cout ;
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.fas_s2  = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.s ;
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.a  = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.a [15:0];
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.b  = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.b [15:0];
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.cin  = 1'h0;
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.facout_s1  = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.cout ;
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.fas_s1  = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.s ;
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.a  = \add_32ns_32ns_32_2_1_U15.din0 ;
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.b  = \add_32ns_32ns_32_2_1_U15.din1 ;
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.ce  = \add_32ns_32ns_32_2_1_U15.ce ;
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.clk  = \add_32ns_32ns_32_2_1_U15.clk ;
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.reset  = \add_32ns_32ns_32_2_1_U15.reset ;
assign \add_32ns_32ns_32_2_1_U15.dout  = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.s ;
assign \add_32ns_32ns_32_2_1_U15.ce  = 1'h1;
assign \add_32ns_32ns_32_2_1_U15.clk  = ap_clk;
assign \add_32ns_32ns_32_2_1_U15.din0  = ret_V_9_cast_reg_911;
assign \add_32ns_32ns_32_2_1_U15.din1  = 32'd1;
assign grp_fu_583_p2 = \add_32ns_32ns_32_2_1_U15.dout ;
assign \add_32ns_32ns_32_2_1_U15.reset  = ap_rst;
assign \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.ain_s0  = \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.a ;
assign \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.bin_s0  = \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.b ;
assign \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.s  = { \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.fas_s2 , \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.sum_s1  };
assign \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.u2.a  = \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.ain_s1 ;
assign \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.u2.b  = \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.bin_s1 ;
assign \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.u2.cin  = \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.carry_s1 ;
assign \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.facout_s2  = \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.u2.cout ;
assign \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.fas_s2  = \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.u2.s ;
assign \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.u1.a  = \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.a [7:0];
assign \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.u1.b  = \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.b [7:0];
assign \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.u1.cin  = 1'h0;
assign \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.facout_s1  = \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.u1.cout ;
assign \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.fas_s1  = \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.u1.s ;
assign \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.a  = \add_17s_17s_17_2_1_U17.din0 ;
assign \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.b  = \add_17s_17s_17_2_1_U17.din1 ;
assign \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.ce  = \add_17s_17s_17_2_1_U17.ce ;
assign \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.clk  = \add_17s_17s_17_2_1_U17.clk ;
assign \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.reset  = \add_17s_17s_17_2_1_U17.reset ;
assign \add_17s_17s_17_2_1_U17.dout  = \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.s ;
assign \add_17s_17s_17_2_1_U17.ce  = 1'h1;
assign \add_17s_17s_17_2_1_U17.clk  = ap_clk;
assign \add_17s_17s_17_2_1_U17.din0  = { op_19[15], op_19 };
assign \add_17s_17s_17_2_1_U17.din1  = { r_reg_933[1], r_reg_933[1], r_reg_933[1], r_reg_933[1], r_reg_933[1], r_reg_933[1], r_reg_933[1], r_reg_933[1], r_reg_933[1], r_reg_933[1], r_reg_933[1], r_reg_933[1], r_reg_933[1], r_reg_933[1], r_reg_933[1], r_reg_933 };
assign grp_fu_643_p2 = \add_17s_17s_17_2_1_U17.dout ;
assign \add_17s_17s_17_2_1_U17.reset  = ap_rst;
assign \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.ain_s0  = \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.a ;
assign \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.bin_s0  = \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.b ;
assign \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.s  = { \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.fas_s2 , \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.sum_s1  };
assign \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.u2.a  = \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.ain_s1 ;
assign \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.u2.b  = \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.bin_s1 ;
assign \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.u2.cin  = \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.carry_s1 ;
assign \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.facout_s2  = \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.u2.cout ;
assign \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.fas_s2  = \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.u2.s ;
assign \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.u1.a  = \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.a [4:0];
assign \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.u1.b  = \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.b [4:0];
assign \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.u1.cin  = 1'h0;
assign \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.facout_s1  = \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.u1.cout ;
assign \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.fas_s1  = \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.u1.s ;
assign \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.a  = \add_10ns_10s_10_2_1_U1.din0 ;
assign \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.b  = \add_10ns_10s_10_2_1_U1.din1 ;
assign \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.ce  = \add_10ns_10s_10_2_1_U1.ce ;
assign \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.clk  = \add_10ns_10s_10_2_1_U1.clk ;
assign \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.reset  = \add_10ns_10s_10_2_1_U1.reset ;
assign \add_10ns_10s_10_2_1_U1.dout  = \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.s ;
assign \add_10ns_10s_10_2_1_U1.ce  = 1'h1;
assign \add_10ns_10s_10_2_1_U1.clk  = ap_clk;
assign \add_10ns_10s_10_2_1_U1.din0  = { 2'h0, op_7 };
assign \add_10ns_10s_10_2_1_U1.din1  = { op_5[7], op_5[7], op_5 };
assign grp_fu_221_p2 = \add_10ns_10s_10_2_1_U1.dout ;
assign \add_10ns_10s_10_2_1_U1.reset  = ap_rst;
endmodule


// Machine B:
// Processed by function `add_clk_enable_signal` in `verilog_tricks.py`.
// Processed by function `remove_reset_signal` in `verilog_tricks.py`.
module top_B (
  ap_clk,
  ap_start,
  ap_done,
  ap_idle,
  ap_ready,
  op_0,
  op_1,
  op_2,
  op_4,
  op_5,
  op_7,
  op_9,
  op_11,
  op_12,
  op_14,
  op_15,
  op_19,
  op_29,
  op_29_ap_vld,
clk_enable
);
input clk_enable;


input ap_clk;
wire ap_rst;
assign ap_rst = op_29_ap_vld;
input ap_start;
input [3:0] op_0;
input [7:0] op_1;
input [1:0] op_11;
input [1:0] op_12;
input [31:0] op_14;
input [15:0] op_15;
input [15:0] op_19;
input [15:0] op_2;
input [7:0] op_4;
input [7:0] op_5;
input [7:0] op_7;
input [1:0] op_9;
output ap_done;
output ap_idle;
output ap_ready;
output [31:0] op_29;
output op_29_ap_vld;


reg [4:0] \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.ain_s1 ;
reg [4:0] \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.bin_s1 ;
reg \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.carry_s1 ;
reg [4:0] \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.sum_s1 ;
reg [8:0] \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.ain_s1 ;
reg [8:0] \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.bin_s1 ;
reg \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.carry_s1 ;
reg [7:0] \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.sum_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.ain_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.bin_s1 ;
reg \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.carry_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.sum_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.ain_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.bin_s1 ;
reg \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.carry_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.sum_s1 ;
reg [15:0] \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.ain_s1 ;
reg [15:0] \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.bin_s1 ;
reg \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.carry_s1 ;
reg [15:0] \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.sum_s1 ;
reg [15:0] \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.ain_s1 ;
reg [15:0] \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.bin_s1 ;
reg \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.carry_s1 ;
reg [15:0] \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.sum_s1 ;
reg [15:0] \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.ain_s1 ;
reg [15:0] \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.bin_s1 ;
reg \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.carry_s1 ;
reg [15:0] \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.sum_s1 ;
reg [15:0] \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.ain_s1 ;
reg [15:0] \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.bin_s1 ;
reg \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.carry_s1 ;
reg [15:0] \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.sum_s1 ;
reg [16:0] \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.ain_s1 ;
reg [16:0] \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.bin_s1 ;
reg \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.carry_s1 ;
reg [16:0] \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.sum_s1 ;
reg [1:0] \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.ain_s1 ;
reg [1:0] \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.bin_s1 ;
reg \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.carry_s1 ;
reg \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.sum_s1 ;
reg [2:0] \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.ain_s1 ;
reg [2:0] \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.bin_s1 ;
reg \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.carry_s1 ;
reg [1:0] \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.sum_s1 ;
reg [2:0] \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.ain_s1 ;
reg [2:0] \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.bin_s1 ;
reg \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.carry_s1 ;
reg [1:0] \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.sum_s1 ;
reg [3:0] \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.ain_s1 ;
reg [3:0] \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.bin_s1 ;
reg \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.carry_s1 ;
reg [2:0] \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.sum_s1 ;
reg [31:0] add_ln691_1_reg_928;
reg [31:0] add_ln691_reg_809;
reg [2:0] add_ln69_1_reg_861;
reg [16:0] add_ln69_3_reg_963;
reg [31:0] add_ln69_reg_856;
reg [23:0] ap_CS_fsm = 24'h000001;
reg [31:0] \ashr_32s_32ns_32_7_1_U10.din1_cast_array[0] ;
reg [31:0] \ashr_32s_32ns_32_7_1_U10.din1_cast_array[1] ;
reg [31:0] \ashr_32s_32ns_32_7_1_U10.din1_cast_array[2] ;
reg [31:0] \ashr_32s_32ns_32_7_1_U10.din1_cast_array[3] ;
reg [31:0] \ashr_32s_32ns_32_7_1_U10.din1_cast_array[4] ;
reg [31:0] \ashr_32s_32ns_32_7_1_U10.din1_cast_array[5] ;
reg [31:0] \ashr_32s_32ns_32_7_1_U10.dout_array[0] ;
reg [31:0] \ashr_32s_32ns_32_7_1_U10.dout_array[1] ;
reg [31:0] \ashr_32s_32ns_32_7_1_U10.dout_array[2] ;
reg [31:0] \ashr_32s_32ns_32_7_1_U10.dout_array[3] ;
reg [31:0] \ashr_32s_32ns_32_7_1_U10.dout_array[4] ;
reg [31:0] \ashr_32s_32ns_32_7_1_U10.dout_array[5] ;
reg icmp_ln768_reg_716;
reg icmp_ln850_reg_804;
reg lhs_V_4_reg_679;
reg newsignbit_reg_673;
reg [3:0] op_16_V_reg_886;
reg [31:0] op_25_V_reg_891;
reg op_6_V_reg_699;
reg [19:0] op_8_V_reg_761;
reg p_Result_3_reg_704;
reg p_Result_4_reg_820;
reg [8:0] p_Result_s_reg_711;
reg [1:0] r_reg_933;
reg [4:0] ret_1_reg_731;
reg [4:0] ret_V_11_reg_741;
reg [6:0] ret_V_12_reg_776;
reg [31:0] ret_V_13_reg_825;
reg [33:0] ret_V_14_reg_906;
reg [31:0] ret_V_15_reg_938;
reg [31:0] ret_V_16_reg_958;
reg [31:0] ret_V_9_cast_reg_911;
reg [27:0] ret_V_9_reg_786;
reg [21:0] ret_V_reg_881;
reg [4:0] select_ln1192_reg_736;
reg [2:0] select_ln69_reg_830;
reg [31:0] sext_ln831_reg_797;
reg [31:0] sh_reg_835;
reg [31:0] \shl_32s_32ns_32_7_1_U11.din1_cast_array[0] ;
reg [31:0] \shl_32s_32ns_32_7_1_U11.din1_cast_array[1] ;
reg [31:0] \shl_32s_32ns_32_7_1_U11.din1_cast_array[2] ;
reg [31:0] \shl_32s_32ns_32_7_1_U11.din1_cast_array[3] ;
reg [31:0] \shl_32s_32ns_32_7_1_U11.din1_cast_array[4] ;
reg [31:0] \shl_32s_32ns_32_7_1_U11.din1_cast_array[5] ;
reg [31:0] \shl_32s_32ns_32_7_1_U11.dout_array[0] ;
reg [31:0] \shl_32s_32ns_32_7_1_U11.dout_array[1] ;
reg [31:0] \shl_32s_32ns_32_7_1_U11.dout_array[2] ;
reg [31:0] \shl_32s_32ns_32_7_1_U11.dout_array[3] ;
reg [31:0] \shl_32s_32ns_32_7_1_U11.dout_array[4] ;
reg [31:0] \shl_32s_32ns_32_7_1_U11.dout_array[5] ;
reg signbit_1_reg_684;
reg [10:0] \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.ain_s1 ;
reg [10:0] \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.bin_s1 ;
reg \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.carry_s1 ;
reg [10:0] \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.sum_s1 ;
reg [13:0] \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.ain_s1 ;
reg [13:0] \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.bin_s1 ;
reg \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.carry_s1 ;
reg [13:0] \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.sum_s1 ;
reg [15:0] \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.ain_s1 ;
reg [15:0] \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.bin_s1 ;
reg \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.carry_s1 ;
reg [15:0] \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.sum_s1 ;
reg [5:0] tmp_2_reg_781;
reg trunc_ln213_reg_658;
reg [2:0] trunc_ln728_reg_689;
reg [1:0] trunc_ln798_1_reg_923;
reg [1:0] trunc_ln798_reg_918;
reg [18:0] trunc_ln851_reg_792;
wire [31:0] _000_;
wire [31:0] _001_;
wire [2:0] _002_;
wire [16:0] _003_;
wire [31:0] _004_;
wire [23:0] _005_;
wire _006_;
wire _007_;
wire _008_;
wire _009_;
wire [3:0] _010_;
wire [31:0] _011_;
wire _012_;
wire _013_;
wire _014_;
wire _015_;
wire [8:0] _016_;
wire [1:0] _017_;
wire [4:0] _018_;
wire [4:0] _019_;
wire [6:0] _020_;
wire [31:0] _021_;
wire [33:0] _022_;
wire [31:0] _023_;
wire [31:0] _024_;
wire [31:0] _025_;
wire [27:0] _026_;
wire [21:0] _027_;
wire [4:0] _028_;
wire [2:0] _029_;
wire [31:0] _030_;
wire [31:0] _031_;
wire _032_;
wire [5:0] _033_;
wire _034_;
wire [2:0] _035_;
wire [1:0] _036_;
wire [1:0] _037_;
wire [18:0] _038_;
wire [1:0] _039_;
wire _040_;
wire _041_;
wire _042_;
wire _043_;
wire _044_;
wire _045_;
wire [4:0] _046_;
wire [4:0] _047_;
wire _048_;
wire [4:0] _049_;
wire [5:0] _050_;
wire [5:0] _051_;
wire [8:0] _052_;
wire [8:0] _053_;
wire _054_;
wire [7:0] _055_;
wire [8:0] _056_;
wire [9:0] _057_;
wire [15:0] _058_;
wire [15:0] _059_;
wire _060_;
wire [15:0] _061_;
wire [16:0] _062_;
wire [16:0] _063_;
wire [15:0] _064_;
wire [15:0] _065_;
wire _066_;
wire [15:0] _067_;
wire [16:0] _068_;
wire [16:0] _069_;
wire [15:0] _070_;
wire [15:0] _071_;
wire _072_;
wire [15:0] _073_;
wire [16:0] _074_;
wire [16:0] _075_;
wire [15:0] _076_;
wire [15:0] _077_;
wire _078_;
wire [15:0] _079_;
wire [16:0] _080_;
wire [16:0] _081_;
wire [15:0] _082_;
wire [15:0] _083_;
wire _084_;
wire [15:0] _085_;
wire [16:0] _086_;
wire [16:0] _087_;
wire [15:0] _088_;
wire [15:0] _089_;
wire _090_;
wire [15:0] _091_;
wire [16:0] _092_;
wire [16:0] _093_;
wire [16:0] _094_;
wire [16:0] _095_;
wire _096_;
wire [16:0] _097_;
wire [17:0] _098_;
wire [17:0] _099_;
wire [1:0] _100_;
wire [1:0] _101_;
wire _102_;
wire _103_;
wire [1:0] _104_;
wire [2:0] _105_;
wire [2:0] _106_;
wire [2:0] _107_;
wire _108_;
wire [1:0] _109_;
wire [2:0] _110_;
wire [3:0] _111_;
wire [2:0] _112_;
wire [2:0] _113_;
wire _114_;
wire [1:0] _115_;
wire [2:0] _116_;
wire [3:0] _117_;
wire [3:0] _118_;
wire [3:0] _119_;
wire _120_;
wire [2:0] _121_;
wire [3:0] _122_;
wire [4:0] _123_;
wire [31:0] _124_;
wire [31:0] _125_;
wire [31:0] _126_;
wire [31:0] _127_;
wire [31:0] _128_;
wire [31:0] _129_;
wire [31:0] _130_;
wire [31:0] _131_;
wire [31:0] _132_;
wire [31:0] _133_;
wire [31:0] _134_;
wire [31:0] _135_;
wire [31:0] _136_;
wire [31:0] _137_;
wire [31:0] _138_;
wire [31:0] _139_;
wire [31:0] _140_;
wire [31:0] _141_;
wire [31:0] _142_;
wire [31:0] _143_;
wire [31:0] _144_;
wire [31:0] _145_;
wire [31:0] _146_;
wire [31:0] _147_;
wire [31:0] _148_;
wire [31:0] _149_;
wire [31:0] _150_;
wire [31:0] _151_;
wire [31:0] _152_;
wire [31:0] _153_;
wire [31:0] _154_;
wire [31:0] _155_;
wire [31:0] _156_;
wire [31:0] _157_;
wire [31:0] _158_;
wire [31:0] _159_;
wire [31:0] _160_;
wire [31:0] _161_;
wire [31:0] _162_;
wire [31:0] _163_;
wire [31:0] _164_;
wire [31:0] _165_;
wire [31:0] _166_;
wire [31:0] _167_;
wire [31:0] _168_;
wire [31:0] _169_;
wire [31:0] _170_;
wire [31:0] _171_;
wire [31:0] _172_;
wire [31:0] _173_;
wire [31:0] _174_;
wire [31:0] _175_;
wire [31:0] _176_;
wire [31:0] _177_;
wire [31:0] _178_;
wire [31:0] _179_;
wire [31:0] _180_;
wire [31:0] _181_;
wire [31:0] _182_;
wire [31:0] _183_;
wire [10:0] _184_;
wire [10:0] _185_;
wire _186_;
wire [10:0] _187_;
wire [11:0] _188_;
wire [11:0] _189_;
wire [13:0] _190_;
wire [13:0] _191_;
wire _192_;
wire [13:0] _193_;
wire [14:0] _194_;
wire [14:0] _195_;
wire [15:0] _196_;
wire [15:0] _197_;
wire _198_;
wire [15:0] _199_;
wire [16:0] _200_;
wire [16:0] _201_;
wire _202_;
wire _203_;
wire _204_;
wire _205_;
wire _206_;
wire _207_;
wire _208_;
wire _209_;
wire _210_;
wire _211_;
wire _212_;
wire _213_;
wire _214_;
wire _215_;
wire _216_;
wire _217_;
wire _218_;
wire _219_;
wire _220_;
wire _221_;
wire _222_;
wire _223_;
wire _224_;
wire _225_;
wire _226_;
wire _227_;
wire _228_;
wire _229_;
wire \add_10ns_10s_10_2_1_U1.ce ;
wire \add_10ns_10s_10_2_1_U1.clk ;
wire [9:0] \add_10ns_10s_10_2_1_U1.din0 ;
wire [9:0] \add_10ns_10s_10_2_1_U1.din1 ;
wire [9:0] \add_10ns_10s_10_2_1_U1.dout ;
wire \add_10ns_10s_10_2_1_U1.reset ;
wire [9:0] \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.a ;
wire [9:0] \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.ain_s0 ;
wire [9:0] \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.b ;
wire [9:0] \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.bin_s0 ;
wire \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.ce ;
wire \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.clk ;
wire \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.facout_s1 ;
wire \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.facout_s2 ;
wire [4:0] \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.fas_s1 ;
wire [4:0] \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.fas_s2 ;
wire \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.reset ;
wire [9:0] \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.s ;
wire [4:0] \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.u1.a ;
wire [4:0] \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.u1.b ;
wire \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.u1.cin ;
wire \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.u1.cout ;
wire [4:0] \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.u1.s ;
wire [4:0] \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.u2.a ;
wire [4:0] \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.u2.b ;
wire \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.u2.cin ;
wire \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.u2.cout ;
wire [4:0] \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.u2.s ;
wire \add_17s_17s_17_2_1_U17.ce ;
wire \add_17s_17s_17_2_1_U17.clk ;
wire [16:0] \add_17s_17s_17_2_1_U17.din0 ;
wire [16:0] \add_17s_17s_17_2_1_U17.din1 ;
wire [16:0] \add_17s_17s_17_2_1_U17.dout ;
wire \add_17s_17s_17_2_1_U17.reset ;
wire [16:0] \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.a ;
wire [16:0] \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.ain_s0 ;
wire [16:0] \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.b ;
wire [16:0] \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.bin_s0 ;
wire \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.ce ;
wire \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.clk ;
wire \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.facout_s1 ;
wire \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.facout_s2 ;
wire [7:0] \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.fas_s1 ;
wire [8:0] \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.fas_s2 ;
wire \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.reset ;
wire [16:0] \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.s ;
wire [7:0] \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.u1.a ;
wire [7:0] \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.u1.b ;
wire \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.u1.cin ;
wire \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.u1.cout ;
wire [7:0] \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.u1.s ;
wire [8:0] \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.u2.a ;
wire [8:0] \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.u2.b ;
wire \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.u2.cin ;
wire \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.u2.cout ;
wire [8:0] \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.u2.s ;
wire \add_32ns_32ns_32_2_1_U15.ce ;
wire \add_32ns_32ns_32_2_1_U15.clk ;
wire [31:0] \add_32ns_32ns_32_2_1_U15.din0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U15.din1 ;
wire [31:0] \add_32ns_32ns_32_2_1_U15.dout ;
wire \add_32ns_32ns_32_2_1_U15.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.a ;
wire [31:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.ain_s0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.b ;
wire [31:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.bin_s0 ;
wire \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.ce ;
wire \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.clk ;
wire \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.facout_s1 ;
wire \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.facout_s2 ;
wire [15:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.fas_s1 ;
wire [15:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.fas_s2 ;
wire \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.b ;
wire \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.cin ;
wire \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.b ;
wire \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.cin ;
wire \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.s ;
wire \add_32ns_32ns_32_2_1_U16.ce ;
wire \add_32ns_32ns_32_2_1_U16.clk ;
wire [31:0] \add_32ns_32ns_32_2_1_U16.din0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U16.din1 ;
wire [31:0] \add_32ns_32ns_32_2_1_U16.dout ;
wire \add_32ns_32ns_32_2_1_U16.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.a ;
wire [31:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.ain_s0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.b ;
wire [31:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.bin_s0 ;
wire \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.ce ;
wire \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.clk ;
wire \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.facout_s1 ;
wire \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.facout_s2 ;
wire [15:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.fas_s1 ;
wire [15:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.fas_s2 ;
wire \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.b ;
wire \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.cin ;
wire \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.b ;
wire \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.cin ;
wire \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.s ;
wire \add_32ns_32s_32_2_1_U8.ce ;
wire \add_32ns_32s_32_2_1_U8.clk ;
wire [31:0] \add_32ns_32s_32_2_1_U8.din0 ;
wire [31:0] \add_32ns_32s_32_2_1_U8.din1 ;
wire [31:0] \add_32ns_32s_32_2_1_U8.dout ;
wire \add_32ns_32s_32_2_1_U8.reset ;
wire [31:0] \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.a ;
wire [31:0] \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.ain_s0 ;
wire [31:0] \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.b ;
wire [31:0] \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.bin_s0 ;
wire \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.ce ;
wire \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.clk ;
wire \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.facout_s1 ;
wire \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.facout_s2 ;
wire [15:0] \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.fas_s1 ;
wire [15:0] \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.fas_s2 ;
wire \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.reset ;
wire [31:0] \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.s ;
wire [15:0] \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.u1.a ;
wire [15:0] \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.u1.b ;
wire \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.u1.cin ;
wire \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.u1.cout ;
wire [15:0] \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.u1.s ;
wire [15:0] \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.u2.a ;
wire [15:0] \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.u2.b ;
wire \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.u2.cin ;
wire \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.u2.cout ;
wire [15:0] \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.u2.s ;
wire \add_32s_32ns_32_2_1_U13.ce ;
wire \add_32s_32ns_32_2_1_U13.clk ;
wire [31:0] \add_32s_32ns_32_2_1_U13.din0 ;
wire [31:0] \add_32s_32ns_32_2_1_U13.din1 ;
wire [31:0] \add_32s_32ns_32_2_1_U13.dout ;
wire \add_32s_32ns_32_2_1_U13.reset ;
wire [31:0] \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.a ;
wire [31:0] \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.ain_s0 ;
wire [31:0] \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.b ;
wire [31:0] \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.bin_s0 ;
wire \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.ce ;
wire \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.clk ;
wire \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.facout_s1 ;
wire \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.facout_s2 ;
wire [15:0] \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.fas_s1 ;
wire [15:0] \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.fas_s2 ;
wire \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.reset ;
wire [31:0] \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.s ;
wire [15:0] \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.u1.a ;
wire [15:0] \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.u1.b ;
wire \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.u1.cin ;
wire \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.u1.cout ;
wire [15:0] \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.u1.s ;
wire [15:0] \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.u2.a ;
wire [15:0] \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.u2.b ;
wire \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.u2.cin ;
wire \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.u2.cout ;
wire [15:0] \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.u2.s ;
wire \add_32s_32ns_32_2_1_U18.ce ;
wire \add_32s_32ns_32_2_1_U18.clk ;
wire [31:0] \add_32s_32ns_32_2_1_U18.din0 ;
wire [31:0] \add_32s_32ns_32_2_1_U18.din1 ;
wire [31:0] \add_32s_32ns_32_2_1_U18.dout ;
wire \add_32s_32ns_32_2_1_U18.reset ;
wire [31:0] \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.a ;
wire [31:0] \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.ain_s0 ;
wire [31:0] \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.b ;
wire [31:0] \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.bin_s0 ;
wire \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.ce ;
wire \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.clk ;
wire \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.facout_s1 ;
wire \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.facout_s2 ;
wire [15:0] \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.fas_s1 ;
wire [15:0] \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.fas_s2 ;
wire \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.reset ;
wire [31:0] \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.s ;
wire [15:0] \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.u1.a ;
wire [15:0] \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.u1.b ;
wire \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.u1.cin ;
wire \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.u1.cout ;
wire [15:0] \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.u1.s ;
wire [15:0] \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.u2.a ;
wire [15:0] \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.u2.b ;
wire \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.u2.cin ;
wire \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.u2.cout ;
wire [15:0] \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.u2.s ;
wire \add_32s_32ns_32_2_1_U6.ce ;
wire \add_32s_32ns_32_2_1_U6.clk ;
wire [31:0] \add_32s_32ns_32_2_1_U6.din0 ;
wire [31:0] \add_32s_32ns_32_2_1_U6.din1 ;
wire [31:0] \add_32s_32ns_32_2_1_U6.dout ;
wire \add_32s_32ns_32_2_1_U6.reset ;
wire [31:0] \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.a ;
wire [31:0] \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.ain_s0 ;
wire [31:0] \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.b ;
wire [31:0] \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.bin_s0 ;
wire \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.ce ;
wire \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.clk ;
wire \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.facout_s1 ;
wire \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.facout_s2 ;
wire [15:0] \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.fas_s1 ;
wire [15:0] \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.fas_s2 ;
wire \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.reset ;
wire [31:0] \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.s ;
wire [15:0] \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.u1.a ;
wire [15:0] \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.u1.b ;
wire \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.u1.cin ;
wire \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.u1.cout ;
wire [15:0] \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.u1.s ;
wire [15:0] \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.u2.a ;
wire [15:0] \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.u2.b ;
wire \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.u2.cin ;
wire \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.u2.cout ;
wire [15:0] \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.u2.s ;
wire \add_34s_34s_34_2_1_U14.ce ;
wire \add_34s_34s_34_2_1_U14.clk ;
wire [33:0] \add_34s_34s_34_2_1_U14.din0 ;
wire [33:0] \add_34s_34s_34_2_1_U14.din1 ;
wire [33:0] \add_34s_34s_34_2_1_U14.dout ;
wire \add_34s_34s_34_2_1_U14.reset ;
wire [33:0] \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.a ;
wire [33:0] \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.ain_s0 ;
wire [33:0] \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.b ;
wire [33:0] \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.bin_s0 ;
wire \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.ce ;
wire \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.clk ;
wire \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.facout_s1 ;
wire \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.facout_s2 ;
wire [16:0] \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.fas_s1 ;
wire [16:0] \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.fas_s2 ;
wire \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.reset ;
wire [33:0] \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.s ;
wire [16:0] \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.u1.a ;
wire [16:0] \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.u1.b ;
wire \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.u1.cin ;
wire \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.u1.cout ;
wire [16:0] \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.u1.s ;
wire [16:0] \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.u2.a ;
wire [16:0] \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.u2.b ;
wire \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.u2.cin ;
wire \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.u2.cout ;
wire [16:0] \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.u2.s ;
wire \add_3s_3ns_3_2_1_U9.ce ;
wire \add_3s_3ns_3_2_1_U9.clk ;
wire [2:0] \add_3s_3ns_3_2_1_U9.din0 ;
wire [2:0] \add_3s_3ns_3_2_1_U9.din1 ;
wire [2:0] \add_3s_3ns_3_2_1_U9.dout ;
wire \add_3s_3ns_3_2_1_U9.reset ;
wire [2:0] \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.a ;
wire [2:0] \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.ain_s0 ;
wire [2:0] \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.b ;
wire [2:0] \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.bin_s0 ;
wire \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.ce ;
wire \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.clk ;
wire \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.facout_s1 ;
wire \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.facout_s2 ;
wire \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.fas_s1 ;
wire [1:0] \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.fas_s2 ;
wire \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.reset ;
wire [2:0] \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.s ;
wire \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.u1.a ;
wire \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.u1.b ;
wire \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.u1.cin ;
wire \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.u1.cout ;
wire \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.u1.s ;
wire [1:0] \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.u2.a ;
wire [1:0] \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.u2.b ;
wire \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.u2.cin ;
wire \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.u2.cout ;
wire [1:0] \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.u2.s ;
wire \add_5ns_5ns_5_2_1_U3.ce ;
wire \add_5ns_5ns_5_2_1_U3.clk ;
wire [4:0] \add_5ns_5ns_5_2_1_U3.din0 ;
wire [4:0] \add_5ns_5ns_5_2_1_U3.din1 ;
wire [4:0] \add_5ns_5ns_5_2_1_U3.dout ;
wire \add_5ns_5ns_5_2_1_U3.reset ;
wire [4:0] \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.a ;
wire [4:0] \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.ain_s0 ;
wire [4:0] \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.b ;
wire [4:0] \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.bin_s0 ;
wire \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.ce ;
wire \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.clk ;
wire \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.facout_s1 ;
wire \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.facout_s2 ;
wire [1:0] \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.fas_s1 ;
wire [2:0] \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.fas_s2 ;
wire \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.reset ;
wire [4:0] \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.s ;
wire [1:0] \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.u1.a ;
wire [1:0] \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.u1.b ;
wire \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.u1.cin ;
wire \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.u1.cout ;
wire [1:0] \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.u1.s ;
wire [2:0] \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.u2.a ;
wire [2:0] \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.u2.b ;
wire \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.u2.cin ;
wire \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.u2.cout ;
wire [2:0] \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.u2.s ;
wire \add_5s_5ns_5_2_1_U2.ce ;
wire \add_5s_5ns_5_2_1_U2.clk ;
wire [4:0] \add_5s_5ns_5_2_1_U2.din0 ;
wire [4:0] \add_5s_5ns_5_2_1_U2.din1 ;
wire [4:0] \add_5s_5ns_5_2_1_U2.dout ;
wire \add_5s_5ns_5_2_1_U2.reset ;
wire [4:0] \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.a ;
wire [4:0] \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.ain_s0 ;
wire [4:0] \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.b ;
wire [4:0] \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.bin_s0 ;
wire \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.ce ;
wire \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.clk ;
wire \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.facout_s1 ;
wire \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.facout_s2 ;
wire [1:0] \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.fas_s1 ;
wire [2:0] \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.fas_s2 ;
wire \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.reset ;
wire [4:0] \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.s ;
wire [1:0] \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.u1.a ;
wire [1:0] \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.u1.b ;
wire \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.u1.cin ;
wire \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.u1.cout ;
wire [1:0] \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.u1.s ;
wire [2:0] \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.u2.a ;
wire [2:0] \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.u2.b ;
wire \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.u2.cin ;
wire \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.u2.cout ;
wire [2:0] \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.u2.s ;
wire \add_7s_7s_7_2_1_U4.ce ;
wire \add_7s_7s_7_2_1_U4.clk ;
wire [6:0] \add_7s_7s_7_2_1_U4.din0 ;
wire [6:0] \add_7s_7s_7_2_1_U4.din1 ;
wire [6:0] \add_7s_7s_7_2_1_U4.dout ;
wire \add_7s_7s_7_2_1_U4.reset ;
wire [6:0] \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.a ;
wire [6:0] \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.ain_s0 ;
wire [6:0] \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.b ;
wire [6:0] \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.bin_s0 ;
wire \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.ce ;
wire \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.clk ;
wire \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.facout_s1 ;
wire \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.facout_s2 ;
wire [2:0] \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.fas_s1 ;
wire [3:0] \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.fas_s2 ;
wire \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.reset ;
wire [6:0] \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.s ;
wire [2:0] \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.u1.a ;
wire [2:0] \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.u1.b ;
wire \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.u1.cin ;
wire \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.u1.cout ;
wire [2:0] \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.u1.s ;
wire [3:0] \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.u2.a ;
wire [3:0] \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.u2.b ;
wire \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.u2.cin ;
wire \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.u2.cout ;
wire [3:0] \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.u2.s ;
wire and_ln353_fu_445_p2;
wire ap_CS_fsm_state1;
wire ap_CS_fsm_state10;
wire ap_CS_fsm_state11;
wire ap_CS_fsm_state12;
wire ap_CS_fsm_state13;
wire ap_CS_fsm_state14;
wire ap_CS_fsm_state15;
wire ap_CS_fsm_state16;
wire ap_CS_fsm_state17;
wire ap_CS_fsm_state18;
wire ap_CS_fsm_state19;
wire ap_CS_fsm_state2;
wire ap_CS_fsm_state20;
wire ap_CS_fsm_state21;
wire ap_CS_fsm_state22;
wire ap_CS_fsm_state23;
wire ap_CS_fsm_state24;
wire ap_CS_fsm_state3;
wire ap_CS_fsm_state4;
wire ap_CS_fsm_state5;
wire ap_CS_fsm_state6;
wire ap_CS_fsm_state7;
wire ap_CS_fsm_state8;
wire ap_CS_fsm_state9;
wire [23:0] ap_NS_fsm;
wire ap_clk;
wire ap_done;
wire ap_idle;
wire ap_ready;
wire ap_rst;
wire ap_start;
wire \ashr_32s_32ns_32_7_1_U10.ce ;
wire \ashr_32s_32ns_32_7_1_U10.clk ;
wire [31:0] \ashr_32s_32ns_32_7_1_U10.din0 ;
wire [31:0] \ashr_32s_32ns_32_7_1_U10.din1 ;
wire [31:0] \ashr_32s_32ns_32_7_1_U10.din1_cast ;
wire [31:0] \ashr_32s_32ns_32_7_1_U10.din1_mask ;
wire [31:0] \ashr_32s_32ns_32_7_1_U10.dout ;
wire \ashr_32s_32ns_32_7_1_U10.reset ;
wire [9:0] grp_fu_221_p0;
wire [9:0] grp_fu_221_p1;
wire [9:0] grp_fu_221_p2;
wire [4:0] grp_fu_296_p0;
wire [4:0] grp_fu_296_p1;
wire [4:0] grp_fu_296_p2;
wire [4:0] grp_fu_336_p2;
wire [6:0] grp_fu_355_p0;
wire [6:0] grp_fu_355_p1;
wire [6:0] grp_fu_355_p2;
wire [27:0] grp_fu_383_p0;
wire [27:0] grp_fu_383_p1;
wire [27:0] grp_fu_383_p2;
wire [31:0] grp_fu_406_p0;
wire [31:0] grp_fu_406_p2;
wire [31:0] grp_fu_425_p2;
wire [31:0] grp_fu_495_p1;
wire [31:0] grp_fu_495_p2;
wire [2:0] grp_fu_500_p0;
wire [2:0] grp_fu_500_p2;
wire [31:0] grp_fu_509_p2;
wire [31:0] grp_fu_514_p2;
wire [21:0] grp_fu_529_p0;
wire [21:0] grp_fu_529_p1;
wire [21:0] grp_fu_529_p2;
wire [31:0] grp_fu_538_p0;
wire [31:0] grp_fu_538_p2;
wire [33:0] grp_fu_567_p0;
wire [33:0] grp_fu_567_p1;
wire [33:0] grp_fu_567_p2;
wire [31:0] grp_fu_583_p2;
wire [31:0] grp_fu_631_p1;
wire [31:0] grp_fu_631_p2;
wire [16:0] grp_fu_643_p0;
wire [16:0] grp_fu_643_p1;
wire [16:0] grp_fu_643_p2;
wire [31:0] grp_fu_652_p0;
wire [31:0] grp_fu_652_p2;
wire icmp_ln768_fu_284_p2;
wire icmp_ln850_fu_412_p2;
wire lhs_V_4_fu_237_p2;
wire [26:0] lhs_V_fu_368_p3;
wire newsignbit_fu_227_p2;
wire [3:0] op_0;
wire [7:0] op_1;
wire op_10_V_fu_322_p3;
wire [1:0] op_11;
wire [1:0] op_12;
wire [31:0] op_14;
wire [15:0] op_15;
wire [15:0] op_19;
wire [15:0] op_2;
wire [31:0] op_29;
wire op_29_ap_vld;
wire op_3_V_fu_197_p1;
wire [7:0] op_4;
wire [7:0] op_5;
wire op_6_V_fu_261_p2;
wire [7:0] op_7;
wire [19:0] op_8_V_fu_361_p3;
wire [1:0] op_9;
wire or_ln340_fu_317_p2;
wire or_ln785_fu_302_p2;
wire overflow_fu_311_p2;
wire p_Result_1_fu_456_p3;
wire p_Result_2_fu_601_p3;
wire p_Result_s_12_fu_438_p3;
wire [1:0] r_fu_596_p3;
wire ret_V_10_fu_450_p2;
wire [31:0] ret_V_13_fu_472_p3;
wire [31:0] ret_V_15_fu_621_p3;
wire [32:0] rhs_4_fu_556_p3;
wire [4:0] select_ln1192_fu_328_p3;
wire [2:0] select_ln69_fu_479_p3;
wire [31:0] select_ln850_1_fu_615_p3;
wire [31:0] select_ln850_fu_466_p3;
wire [1:0] sext_ln1192_fu_340_p0;
wire [7:0] sext_ln215_fu_205_p0;
wire [31:0] sext_ln781_fu_505_p1;
wire [31:0] sext_ln831_fu_403_p1;
wire \shl_32s_32ns_32_7_1_U11.ce ;
wire \shl_32s_32ns_32_7_1_U11.clk ;
wire [31:0] \shl_32s_32ns_32_7_1_U11.din0 ;
wire [31:0] \shl_32s_32ns_32_7_1_U11.din1 ;
wire [31:0] \shl_32s_32ns_32_7_1_U11.din1_cast ;
wire [31:0] \shl_32s_32ns_32_7_1_U11.din1_mask ;
wire [31:0] \shl_32s_32ns_32_7_1_U11.dout ;
wire \shl_32s_32ns_32_7_1_U11.reset ;
wire signbit_1_fu_247_p2;
wire \sub_22ns_22ns_22_2_1_U12.ce ;
wire \sub_22ns_22ns_22_2_1_U12.clk ;
wire [21:0] \sub_22ns_22ns_22_2_1_U12.din0 ;
wire [21:0] \sub_22ns_22ns_22_2_1_U12.din1 ;
wire [21:0] \sub_22ns_22ns_22_2_1_U12.dout ;
wire \sub_22ns_22ns_22_2_1_U12.reset ;
wire [21:0] \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.a ;
wire [21:0] \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.ain_s0 ;
wire [21:0] \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.b ;
wire [21:0] \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.bin_s0 ;
wire \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.ce ;
wire \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.clk ;
wire \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.facout_s1 ;
wire \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.facout_s2 ;
wire [10:0] \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.fas_s1 ;
wire [10:0] \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.fas_s2 ;
wire \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.reset ;
wire [21:0] \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.s ;
wire [10:0] \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.u1.a ;
wire [10:0] \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.u1.b ;
wire \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.u1.cin ;
wire \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.u1.cout ;
wire [10:0] \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.u1.s ;
wire [10:0] \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.u2.a ;
wire [10:0] \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.u2.b ;
wire \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.u2.cin ;
wire \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.u2.cout ;
wire [10:0] \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.u2.s ;
wire \sub_28s_28ns_28_2_1_U5.ce ;
wire \sub_28s_28ns_28_2_1_U5.clk ;
wire [27:0] \sub_28s_28ns_28_2_1_U5.din0 ;
wire [27:0] \sub_28s_28ns_28_2_1_U5.din1 ;
wire [27:0] \sub_28s_28ns_28_2_1_U5.dout ;
wire \sub_28s_28ns_28_2_1_U5.reset ;
wire [27:0] \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.a ;
wire [27:0] \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.ain_s0 ;
wire [27:0] \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.b ;
wire [27:0] \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.bin_s0 ;
wire \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.ce ;
wire \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.clk ;
wire \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.facout_s1 ;
wire \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.facout_s2 ;
wire [13:0] \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.fas_s1 ;
wire [13:0] \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.fas_s2 ;
wire \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.reset ;
wire [27:0] \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.s ;
wire [13:0] \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.u1.a ;
wire [13:0] \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.u1.b ;
wire \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.u1.cin ;
wire \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.u1.cout ;
wire [13:0] \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.u1.s ;
wire [13:0] \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.u2.a ;
wire [13:0] \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.u2.b ;
wire \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.u2.cin ;
wire \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.u2.cout ;
wire [13:0] \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.u2.s ;
wire \sub_32ns_32ns_32_2_1_U7.ce ;
wire \sub_32ns_32ns_32_2_1_U7.clk ;
wire [31:0] \sub_32ns_32ns_32_2_1_U7.din0 ;
wire [31:0] \sub_32ns_32ns_32_2_1_U7.din1 ;
wire [31:0] \sub_32ns_32ns_32_2_1_U7.dout ;
wire \sub_32ns_32ns_32_2_1_U7.reset ;
wire [31:0] \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.a ;
wire [31:0] \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.ain_s0 ;
wire [31:0] \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.b ;
wire [31:0] \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.bin_s0 ;
wire \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.ce ;
wire \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.clk ;
wire \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.facout_s1 ;
wire \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.facout_s2 ;
wire [15:0] \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.fas_s1 ;
wire [15:0] \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.fas_s2 ;
wire \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.reset ;
wire [31:0] \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.s ;
wire [15:0] \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.u1.a ;
wire [15:0] \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.u1.b ;
wire \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.u1.cin ;
wire \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.u1.cout ;
wire [15:0] \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.u1.s ;
wire [15:0] \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.u2.a ;
wire [15:0] \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.u2.b ;
wire \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.u2.cin ;
wire \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.u2.cout ;
wire [15:0] \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.u2.s ;
wire [5:0] tmp_4_fu_344_p3;
wire tmp_6_fu_608_p3;
wire tmp_fu_431_p3;
wire trunc_ln1346_1_fu_217_p1;
wire [7:0] trunc_ln1346_fu_213_p0;
wire trunc_ln1346_fu_213_p1;
wire trunc_ln213_1_fu_257_p1;
wire trunc_ln213_fu_201_p1;
wire [2:0] trunc_ln728_fu_253_p1;
wire [1:0] trunc_ln798_1_fu_592_p1;
wire [1:0] trunc_ln798_fu_588_p1;
wire [1:0] trunc_ln851_1_fu_463_p0;
wire trunc_ln851_1_fu_463_p1;
wire [18:0] trunc_ln851_fu_399_p1;
wire xor_ln785_fu_306_p2;
wire [15:0] zext_ln878_1_fu_243_p1;
wire [15:0] zext_ln878_fu_233_p1;


assign _040_ = ap_CS_fsm[18] & _044_;
assign _041_ = ap_CS_fsm[18] & p_Result_4_reg_820;
assign _042_ = _045_ & ap_CS_fsm[0];
assign _043_ = ap_start & ap_CS_fsm[0];
assign and_ln353_fu_445_p2 = ret_V_9_reg_786[27] & icmp_ln850_reg_804;
assign overflow_fu_311_p2 = xor_ln785_fu_306_p2 & or_ln785_fu_302_p2;
assign xor_ln785_fu_306_p2 = ~ p_Result_3_reg_704;
assign _044_ = ~ p_Result_4_reg_820;
assign _045_ = ~ ap_start;
always @(posedge \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.clk )
\add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.bin_s1  <= _047_;
always @(posedge \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.clk )
\add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.ain_s1  <= _046_;
always @(posedge \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.clk )
\add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.sum_s1  <= _049_;
always @(posedge \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.clk )
\add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.carry_s1  <= _048_;
assign _047_ = \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.ce  ? \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.b [9:5] : \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.bin_s1 ;
assign _046_ = \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.ce  ? \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.a [9:5] : \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.ain_s1 ;
assign _048_ = \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.ce  ? \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.facout_s1  : \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.carry_s1 ;
assign _049_ = \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.ce  ? \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.fas_s1  : \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.sum_s1 ;
assign _050_ = \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.u1.a  + \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.u1.b ;
assign { \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.u1.cout , \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.u1.s  } = _050_ + \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.u1.cin ;
assign _051_ = \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.u2.a  + \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.u2.b ;
assign { \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.u2.cout , \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.u2.s  } = _051_ + \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.u2.cin ;
always @(posedge \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.clk )
\add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.bin_s1  <= _053_;
always @(posedge \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.clk )
\add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.ain_s1  <= _052_;
always @(posedge \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.clk )
\add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.sum_s1  <= _055_;
always @(posedge \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.clk )
\add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.carry_s1  <= _054_;
assign _053_ = \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.ce  ? \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.b [16:8] : \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.bin_s1 ;
assign _052_ = \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.ce  ? \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.a [16:8] : \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.ain_s1 ;
assign _054_ = \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.ce  ? \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.facout_s1  : \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.carry_s1 ;
assign _055_ = \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.ce  ? \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.fas_s1  : \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.sum_s1 ;
assign _056_ = \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.u1.a  + \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.u1.b ;
assign { \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.u1.cout , \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.u1.s  } = _056_ + \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.u1.cin ;
assign _057_ = \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.u2.a  + \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.u2.b ;
assign { \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.u2.cout , \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.u2.s  } = _057_ + \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.u2.cin ;
always @(posedge \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.clk )
\add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.bin_s1  <= _059_;
always @(posedge \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.clk )
\add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.ain_s1  <= _058_;
always @(posedge \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.clk )
\add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.sum_s1  <= _061_;
always @(posedge \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.clk )
\add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.carry_s1  <= _060_;
assign _059_ = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.ce  ? \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.b [31:16] : \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.bin_s1 ;
assign _058_ = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.ce  ? \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.a [31:16] : \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.ain_s1 ;
assign _060_ = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.ce  ? \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.facout_s1  : \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.carry_s1 ;
assign _061_ = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.ce  ? \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.fas_s1  : \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.sum_s1 ;
assign _062_ = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.a  + \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.b ;
assign { \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.cout , \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.s  } = _062_ + \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.cin ;
assign _063_ = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.a  + \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.b ;
assign { \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.cout , \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.s  } = _063_ + \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.cin ;
always @(posedge \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.clk )
\add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.bin_s1  <= _065_;
always @(posedge \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.clk )
\add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.ain_s1  <= _064_;
always @(posedge \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.clk )
\add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.sum_s1  <= _067_;
always @(posedge \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.clk )
\add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.carry_s1  <= _066_;
assign _065_ = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.ce  ? \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.b [31:16] : \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.bin_s1 ;
assign _064_ = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.ce  ? \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.a [31:16] : \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.ain_s1 ;
assign _066_ = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.ce  ? \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.facout_s1  : \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.carry_s1 ;
assign _067_ = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.ce  ? \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.fas_s1  : \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.sum_s1 ;
assign _068_ = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.a  + \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.b ;
assign { \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.cout , \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.s  } = _068_ + \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.cin ;
assign _069_ = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.a  + \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.b ;
assign { \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.cout , \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.s  } = _069_ + \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.cin ;
always @(posedge \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.clk )
\add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.bin_s1  <= _071_;
always @(posedge \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.clk )
\add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.ain_s1  <= _070_;
always @(posedge \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.clk )
\add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.sum_s1  <= _073_;
always @(posedge \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.clk )
\add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.carry_s1  <= _072_;
assign _071_ = \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.ce  ? \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.b [31:16] : \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.bin_s1 ;
assign _070_ = \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.ce  ? \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.a [31:16] : \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.ain_s1 ;
assign _072_ = \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.ce  ? \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.facout_s1  : \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.carry_s1 ;
assign _073_ = \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.ce  ? \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.fas_s1  : \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.sum_s1 ;
assign _074_ = \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.u1.a  + \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.u1.b ;
assign { \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.u1.cout , \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.u1.s  } = _074_ + \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.u1.cin ;
assign _075_ = \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.u2.a  + \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.u2.b ;
assign { \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.u2.cout , \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.u2.s  } = _075_ + \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.u2.cin ;
always @(posedge \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.clk )
\add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.bin_s1  <= _077_;
always @(posedge \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.clk )
\add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.ain_s1  <= _076_;
always @(posedge \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.clk )
\add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.sum_s1  <= _079_;
always @(posedge \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.clk )
\add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.carry_s1  <= _078_;
assign _077_ = \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.ce  ? \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.b [31:16] : \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.bin_s1 ;
assign _076_ = \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.ce  ? \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.a [31:16] : \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.ain_s1 ;
assign _078_ = \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.ce  ? \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.facout_s1  : \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.carry_s1 ;
assign _079_ = \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.ce  ? \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.fas_s1  : \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.sum_s1 ;
assign _080_ = \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.u1.a  + \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.u1.b ;
assign { \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.u1.cout , \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.u1.s  } = _080_ + \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.u1.cin ;
assign _081_ = \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.u2.a  + \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.u2.b ;
assign { \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.u2.cout , \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.u2.s  } = _081_ + \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.u2.cin ;
always @(posedge \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.clk )
\add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.bin_s1  <= _083_;
always @(posedge \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.clk )
\add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.ain_s1  <= _082_;
always @(posedge \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.clk )
\add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.sum_s1  <= _085_;
always @(posedge \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.clk )
\add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.carry_s1  <= _084_;
assign _083_ = \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.ce  ? \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.b [31:16] : \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.bin_s1 ;
assign _082_ = \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.ce  ? \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.a [31:16] : \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.ain_s1 ;
assign _084_ = \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.ce  ? \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.facout_s1  : \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.carry_s1 ;
assign _085_ = \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.ce  ? \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.fas_s1  : \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.sum_s1 ;
assign _086_ = \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.u1.a  + \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.u1.b ;
assign { \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.u1.cout , \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.u1.s  } = _086_ + \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.u1.cin ;
assign _087_ = \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.u2.a  + \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.u2.b ;
assign { \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.u2.cout , \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.u2.s  } = _087_ + \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.u2.cin ;
always @(posedge \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.clk )
\add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.bin_s1  <= _089_;
always @(posedge \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.clk )
\add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.ain_s1  <= _088_;
always @(posedge \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.clk )
\add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.sum_s1  <= _091_;
always @(posedge \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.clk )
\add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.carry_s1  <= _090_;
assign _089_ = \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.ce  ? \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.b [31:16] : \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.bin_s1 ;
assign _088_ = \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.ce  ? \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.a [31:16] : \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.ain_s1 ;
assign _090_ = \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.ce  ? \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.facout_s1  : \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.carry_s1 ;
assign _091_ = \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.ce  ? \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.fas_s1  : \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.sum_s1 ;
assign _092_ = \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.u1.a  + \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.u1.b ;
assign { \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.u1.cout , \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.u1.s  } = _092_ + \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.u1.cin ;
assign _093_ = \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.u2.a  + \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.u2.b ;
assign { \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.u2.cout , \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.u2.s  } = _093_ + \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.u2.cin ;
always @(posedge \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.clk )
\add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.bin_s1  <= _095_;
always @(posedge \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.clk )
\add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.ain_s1  <= _094_;
always @(posedge \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.clk )
\add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.sum_s1  <= _097_;
always @(posedge \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.clk )
\add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.carry_s1  <= _096_;
assign _095_ = \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.ce  ? \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.b [33:17] : \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.bin_s1 ;
assign _094_ = \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.ce  ? \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.a [33:17] : \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.ain_s1 ;
assign _096_ = \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.ce  ? \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.facout_s1  : \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.carry_s1 ;
assign _097_ = \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.ce  ? \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.fas_s1  : \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.sum_s1 ;
assign _098_ = \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.u1.a  + \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.u1.b ;
assign { \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.u1.cout , \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.u1.s  } = _098_ + \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.u1.cin ;
assign _099_ = \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.u2.a  + \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.u2.b ;
assign { \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.u2.cout , \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.u2.s  } = _099_ + \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.u2.cin ;
always @(posedge \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.clk )
\add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.bin_s1  <= _101_;
always @(posedge \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.clk )
\add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.ain_s1  <= _100_;
always @(posedge \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.clk )
\add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.sum_s1  <= _103_;
always @(posedge \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.clk )
\add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.carry_s1  <= _102_;
assign _101_ = \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.ce  ? \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.b [2:1] : \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.bin_s1 ;
assign _100_ = \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.ce  ? \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.a [2:1] : \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.ain_s1 ;
assign _102_ = \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.ce  ? \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.facout_s1  : \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.carry_s1 ;
assign _103_ = \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.ce  ? \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.fas_s1  : \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.sum_s1 ;
assign _104_ = \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.u1.a  + \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.u1.b ;
assign { \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.u1.cout , \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.u1.s  } = _104_ + \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.u1.cin ;
assign _105_ = \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.u2.a  + \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.u2.b ;
assign { \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.u2.cout , \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.u2.s  } = _105_ + \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.u2.cin ;
always @(posedge \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.clk )
\add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.bin_s1  <= _107_;
always @(posedge \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.clk )
\add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.ain_s1  <= _106_;
always @(posedge \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.clk )
\add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.sum_s1  <= _109_;
always @(posedge \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.clk )
\add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.carry_s1  <= _108_;
assign _107_ = \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.ce  ? \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.b [4:2] : \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.bin_s1 ;
assign _106_ = \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.ce  ? \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.a [4:2] : \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.ain_s1 ;
assign _108_ = \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.ce  ? \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.facout_s1  : \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.carry_s1 ;
assign _109_ = \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.ce  ? \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.fas_s1  : \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.sum_s1 ;
assign _110_ = \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.u1.a  + \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.u1.b ;
assign { \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.u1.cout , \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.u1.s  } = _110_ + \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.u1.cin ;
assign _111_ = \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.u2.a  + \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.u2.b ;
assign { \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.u2.cout , \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.u2.s  } = _111_ + \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.u2.cin ;
always @(posedge \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.clk )
\add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.bin_s1  <= _113_;
always @(posedge \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.clk )
\add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.ain_s1  <= _112_;
always @(posedge \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.clk )
\add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.sum_s1  <= _115_;
always @(posedge \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.clk )
\add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.carry_s1  <= _114_;
assign _113_ = \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.ce  ? \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.b [4:2] : \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.bin_s1 ;
assign _112_ = \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.ce  ? \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.a [4:2] : \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.ain_s1 ;
assign _114_ = \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.ce  ? \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.facout_s1  : \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.carry_s1 ;
assign _115_ = \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.ce  ? \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.fas_s1  : \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.sum_s1 ;
assign _116_ = \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.u1.a  + \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.u1.b ;
assign { \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.u1.cout , \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.u1.s  } = _116_ + \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.u1.cin ;
assign _117_ = \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.u2.a  + \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.u2.b ;
assign { \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.u2.cout , \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.u2.s  } = _117_ + \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.u2.cin ;
always @(posedge \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.clk )
\add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.bin_s1  <= _119_;
always @(posedge \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.clk )
\add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.ain_s1  <= _118_;
always @(posedge \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.clk )
\add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.sum_s1  <= _121_;
always @(posedge \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.clk )
\add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.carry_s1  <= _120_;
assign _119_ = \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.ce  ? \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.b [6:3] : \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.bin_s1 ;
assign _118_ = \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.ce  ? \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.a [6:3] : \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.ain_s1 ;
assign _120_ = \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.ce  ? \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.facout_s1  : \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.carry_s1 ;
assign _121_ = \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.ce  ? \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.fas_s1  : \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.sum_s1 ;
assign _122_ = \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.u1.a  + \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.u1.b ;
assign { \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.u1.cout , \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.u1.s  } = _122_ + \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.u1.cin ;
assign _123_ = \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.u2.a  + \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.u2.b ;
assign { \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.u2.cout , \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.u2.s  } = _123_ + \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.u2.cin ;
always @(posedge \ashr_32s_32ns_32_7_1_U10.clk )
\ashr_32s_32ns_32_7_1_U10.dout_array[5]  <= _135_;
always @(posedge \ashr_32s_32ns_32_7_1_U10.clk )
\ashr_32s_32ns_32_7_1_U10.din1_cast_array[5]  <= _129_;
always @(posedge \ashr_32s_32ns_32_7_1_U10.clk )
\ashr_32s_32ns_32_7_1_U10.dout_array[4]  <= _134_;
always @(posedge \ashr_32s_32ns_32_7_1_U10.clk )
\ashr_32s_32ns_32_7_1_U10.din1_cast_array[4]  <= _128_;
always @(posedge \ashr_32s_32ns_32_7_1_U10.clk )
\ashr_32s_32ns_32_7_1_U10.dout_array[3]  <= _133_;
always @(posedge \ashr_32s_32ns_32_7_1_U10.clk )
\ashr_32s_32ns_32_7_1_U10.din1_cast_array[3]  <= _127_;
always @(posedge \ashr_32s_32ns_32_7_1_U10.clk )
\ashr_32s_32ns_32_7_1_U10.dout_array[2]  <= _132_;
always @(posedge \ashr_32s_32ns_32_7_1_U10.clk )
\ashr_32s_32ns_32_7_1_U10.din1_cast_array[2]  <= _126_;
always @(posedge \ashr_32s_32ns_32_7_1_U10.clk )
\ashr_32s_32ns_32_7_1_U10.dout_array[1]  <= _131_;
always @(posedge \ashr_32s_32ns_32_7_1_U10.clk )
\ashr_32s_32ns_32_7_1_U10.din1_cast_array[1]  <= _125_;
always @(posedge \ashr_32s_32ns_32_7_1_U10.clk )
\ashr_32s_32ns_32_7_1_U10.dout_array[0]  <= _130_;
always @(posedge \ashr_32s_32ns_32_7_1_U10.clk )
\ashr_32s_32ns_32_7_1_U10.din1_cast_array[0]  <= _124_;
assign _136_ = \ashr_32s_32ns_32_7_1_U10.ce  ? \ashr_32s_32ns_32_7_1_U10.din1_cast_array[4]  : \ashr_32s_32ns_32_7_1_U10.din1_cast_array[5] ;
assign _129_ = \ashr_32s_32ns_32_7_1_U10.reset  ? 32'd0 : _136_;
assign _137_ = \ashr_32s_32ns_32_7_1_U10.ce  ? _153_ : \ashr_32s_32ns_32_7_1_U10.dout_array[5] ;
assign _135_ = \ashr_32s_32ns_32_7_1_U10.reset  ? 32'd0 : _137_;
assign _138_ = \ashr_32s_32ns_32_7_1_U10.ce  ? \ashr_32s_32ns_32_7_1_U10.din1_cast_array[3]  : \ashr_32s_32ns_32_7_1_U10.din1_cast_array[4] ;
assign _128_ = \ashr_32s_32ns_32_7_1_U10.reset  ? 32'd0 : _138_;
assign _139_ = \ashr_32s_32ns_32_7_1_U10.ce  ? _152_ : \ashr_32s_32ns_32_7_1_U10.dout_array[4] ;
assign _134_ = \ashr_32s_32ns_32_7_1_U10.reset  ? 32'd0 : _139_;
assign _140_ = \ashr_32s_32ns_32_7_1_U10.ce  ? \ashr_32s_32ns_32_7_1_U10.din1_cast_array[2]  : \ashr_32s_32ns_32_7_1_U10.din1_cast_array[3] ;
assign _127_ = \ashr_32s_32ns_32_7_1_U10.reset  ? 32'd0 : _140_;
assign _141_ = \ashr_32s_32ns_32_7_1_U10.ce  ? _151_ : \ashr_32s_32ns_32_7_1_U10.dout_array[3] ;
assign _133_ = \ashr_32s_32ns_32_7_1_U10.reset  ? 32'd0 : _141_;
assign _142_ = \ashr_32s_32ns_32_7_1_U10.ce  ? \ashr_32s_32ns_32_7_1_U10.din1_cast_array[1]  : \ashr_32s_32ns_32_7_1_U10.din1_cast_array[2] ;
assign _126_ = \ashr_32s_32ns_32_7_1_U10.reset  ? 32'd0 : _142_;
assign _143_ = \ashr_32s_32ns_32_7_1_U10.ce  ? _150_ : \ashr_32s_32ns_32_7_1_U10.dout_array[2] ;
assign _132_ = \ashr_32s_32ns_32_7_1_U10.reset  ? 32'd0 : _143_;
assign _144_ = \ashr_32s_32ns_32_7_1_U10.ce  ? \ashr_32s_32ns_32_7_1_U10.din1_cast_array[0]  : \ashr_32s_32ns_32_7_1_U10.din1_cast_array[1] ;
assign _125_ = \ashr_32s_32ns_32_7_1_U10.reset  ? 32'd0 : _144_;
assign _145_ = \ashr_32s_32ns_32_7_1_U10.ce  ? _149_ : \ashr_32s_32ns_32_7_1_U10.dout_array[1] ;
assign _131_ = \ashr_32s_32ns_32_7_1_U10.reset  ? 32'd0 : _145_;
assign _146_ = \ashr_32s_32ns_32_7_1_U10.ce  ? \ashr_32s_32ns_32_7_1_U10.din1  : \ashr_32s_32ns_32_7_1_U10.din1_cast_array[0] ;
assign _124_ = \ashr_32s_32ns_32_7_1_U10.reset  ? 32'd0 : _146_;
assign _147_ = \ashr_32s_32ns_32_7_1_U10.ce  ? _148_ : \ashr_32s_32ns_32_7_1_U10.dout_array[0] ;
assign _130_ = \ashr_32s_32ns_32_7_1_U10.reset  ? 32'd0 : _147_;
assign _148_ = $signed(\ashr_32s_32ns_32_7_1_U10.din0 ) >>> { \ashr_32s_32ns_32_7_1_U10.din1 [31:30], 30'h00000000 };
assign _149_ = $signed(\ashr_32s_32ns_32_7_1_U10.dout_array[0] ) >>> { \ashr_32s_32ns_32_7_1_U10.din1_cast_array[0] [29:25], 25'h0000000 };
assign _150_ = $signed(\ashr_32s_32ns_32_7_1_U10.dout_array[1] ) >>> { \ashr_32s_32ns_32_7_1_U10.din1_cast_array[1] [24:20], 20'h00000 };
assign _151_ = $signed(\ashr_32s_32ns_32_7_1_U10.dout_array[2] ) >>> { \ashr_32s_32ns_32_7_1_U10.din1_cast_array[2] [19:15], 15'h0000 };
assign _152_ = $signed(\ashr_32s_32ns_32_7_1_U10.dout_array[3] ) >>> { \ashr_32s_32ns_32_7_1_U10.din1_cast_array[3] [14:10], 10'h000 };
assign _153_ = $signed(\ashr_32s_32ns_32_7_1_U10.dout_array[4] ) >>> { \ashr_32s_32ns_32_7_1_U10.din1_cast_array[4] [9:5], 5'h00 };
assign \ashr_32s_32ns_32_7_1_U10.dout  = $signed(\ashr_32s_32ns_32_7_1_U10.dout_array[5] ) >>> \ashr_32s_32ns_32_7_1_U10.din1_cast_array[5] [4:0];
always @(posedge \shl_32s_32ns_32_7_1_U11.clk )
\shl_32s_32ns_32_7_1_U11.dout_array[5]  <= _165_;
always @(posedge \shl_32s_32ns_32_7_1_U11.clk )
\shl_32s_32ns_32_7_1_U11.din1_cast_array[5]  <= _159_;
always @(posedge \shl_32s_32ns_32_7_1_U11.clk )
\shl_32s_32ns_32_7_1_U11.dout_array[4]  <= _164_;
always @(posedge \shl_32s_32ns_32_7_1_U11.clk )
\shl_32s_32ns_32_7_1_U11.din1_cast_array[4]  <= _158_;
always @(posedge \shl_32s_32ns_32_7_1_U11.clk )
\shl_32s_32ns_32_7_1_U11.dout_array[3]  <= _163_;
always @(posedge \shl_32s_32ns_32_7_1_U11.clk )
\shl_32s_32ns_32_7_1_U11.din1_cast_array[3]  <= _157_;
always @(posedge \shl_32s_32ns_32_7_1_U11.clk )
\shl_32s_32ns_32_7_1_U11.dout_array[2]  <= _162_;
always @(posedge \shl_32s_32ns_32_7_1_U11.clk )
\shl_32s_32ns_32_7_1_U11.din1_cast_array[2]  <= _156_;
always @(posedge \shl_32s_32ns_32_7_1_U11.clk )
\shl_32s_32ns_32_7_1_U11.dout_array[1]  <= _161_;
always @(posedge \shl_32s_32ns_32_7_1_U11.clk )
\shl_32s_32ns_32_7_1_U11.din1_cast_array[1]  <= _155_;
always @(posedge \shl_32s_32ns_32_7_1_U11.clk )
\shl_32s_32ns_32_7_1_U11.dout_array[0]  <= _160_;
always @(posedge \shl_32s_32ns_32_7_1_U11.clk )
\shl_32s_32ns_32_7_1_U11.din1_cast_array[0]  <= _154_;
assign _166_ = \shl_32s_32ns_32_7_1_U11.ce  ? \shl_32s_32ns_32_7_1_U11.din1_cast_array[4]  : \shl_32s_32ns_32_7_1_U11.din1_cast_array[5] ;
assign _159_ = \shl_32s_32ns_32_7_1_U11.reset  ? 32'd0 : _166_;
assign _167_ = \shl_32s_32ns_32_7_1_U11.ce  ? _183_ : \shl_32s_32ns_32_7_1_U11.dout_array[5] ;
assign _165_ = \shl_32s_32ns_32_7_1_U11.reset  ? 32'd0 : _167_;
assign _168_ = \shl_32s_32ns_32_7_1_U11.ce  ? \shl_32s_32ns_32_7_1_U11.din1_cast_array[3]  : \shl_32s_32ns_32_7_1_U11.din1_cast_array[4] ;
assign _158_ = \shl_32s_32ns_32_7_1_U11.reset  ? 32'd0 : _168_;
assign _169_ = \shl_32s_32ns_32_7_1_U11.ce  ? _182_ : \shl_32s_32ns_32_7_1_U11.dout_array[4] ;
assign _164_ = \shl_32s_32ns_32_7_1_U11.reset  ? 32'd0 : _169_;
assign _170_ = \shl_32s_32ns_32_7_1_U11.ce  ? \shl_32s_32ns_32_7_1_U11.din1_cast_array[2]  : \shl_32s_32ns_32_7_1_U11.din1_cast_array[3] ;
assign _157_ = \shl_32s_32ns_32_7_1_U11.reset  ? 32'd0 : _170_;
assign _171_ = \shl_32s_32ns_32_7_1_U11.ce  ? _181_ : \shl_32s_32ns_32_7_1_U11.dout_array[3] ;
assign _163_ = \shl_32s_32ns_32_7_1_U11.reset  ? 32'd0 : _171_;
assign _172_ = \shl_32s_32ns_32_7_1_U11.ce  ? \shl_32s_32ns_32_7_1_U11.din1_cast_array[1]  : \shl_32s_32ns_32_7_1_U11.din1_cast_array[2] ;
assign _156_ = \shl_32s_32ns_32_7_1_U11.reset  ? 32'd0 : _172_;
assign _173_ = \shl_32s_32ns_32_7_1_U11.ce  ? _180_ : \shl_32s_32ns_32_7_1_U11.dout_array[2] ;
assign _162_ = \shl_32s_32ns_32_7_1_U11.reset  ? 32'd0 : _173_;
assign _174_ = \shl_32s_32ns_32_7_1_U11.ce  ? \shl_32s_32ns_32_7_1_U11.din1_cast_array[0]  : \shl_32s_32ns_32_7_1_U11.din1_cast_array[1] ;
assign _155_ = \shl_32s_32ns_32_7_1_U11.reset  ? 32'd0 : _174_;
assign _175_ = \shl_32s_32ns_32_7_1_U11.ce  ? _179_ : \shl_32s_32ns_32_7_1_U11.dout_array[1] ;
assign _161_ = \shl_32s_32ns_32_7_1_U11.reset  ? 32'd0 : _175_;
assign _176_ = \shl_32s_32ns_32_7_1_U11.ce  ? \shl_32s_32ns_32_7_1_U11.din1  : \shl_32s_32ns_32_7_1_U11.din1_cast_array[0] ;
assign _154_ = \shl_32s_32ns_32_7_1_U11.reset  ? 32'd0 : _176_;
assign _177_ = \shl_32s_32ns_32_7_1_U11.ce  ? _178_ : \shl_32s_32ns_32_7_1_U11.dout_array[0] ;
assign _160_ = \shl_32s_32ns_32_7_1_U11.reset  ? 32'd0 : _177_;
assign _178_ = \shl_32s_32ns_32_7_1_U11.din0  << { \shl_32s_32ns_32_7_1_U11.din1 [31:30], 30'h00000000 };
assign _179_ = \shl_32s_32ns_32_7_1_U11.dout_array[0]  << { \shl_32s_32ns_32_7_1_U11.din1_cast_array[0] [29:25], 25'h0000000 };
assign _180_ = \shl_32s_32ns_32_7_1_U11.dout_array[1]  << { \shl_32s_32ns_32_7_1_U11.din1_cast_array[1] [24:20], 20'h00000 };
assign _181_ = \shl_32s_32ns_32_7_1_U11.dout_array[2]  << { \shl_32s_32ns_32_7_1_U11.din1_cast_array[2] [19:15], 15'h0000 };
assign _182_ = \shl_32s_32ns_32_7_1_U11.dout_array[3]  << { \shl_32s_32ns_32_7_1_U11.din1_cast_array[3] [14:10], 10'h000 };
assign _183_ = \shl_32s_32ns_32_7_1_U11.dout_array[4]  << { \shl_32s_32ns_32_7_1_U11.din1_cast_array[4] [9:5], 5'h00 };
assign \shl_32s_32ns_32_7_1_U11.dout  = \shl_32s_32ns_32_7_1_U11.dout_array[5]  << \shl_32s_32ns_32_7_1_U11.din1_cast_array[5] [4:0];
assign \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.bin_s0  = ~ \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.b ;
always @(posedge \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.clk )
\sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.bin_s1  <= _185_;
always @(posedge \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.clk )
\sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.ain_s1  <= _184_;
always @(posedge \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.clk )
\sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.sum_s1  <= _187_;
always @(posedge \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.clk )
\sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.carry_s1  <= _186_;
assign _185_ = \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.ce  ? \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.bin_s0 [21:11] : \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.bin_s1 ;
assign _184_ = \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.ce  ? \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.a [21:11] : \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.ain_s1 ;
assign _186_ = \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.ce  ? \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.facout_s1  : \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.carry_s1 ;
assign _187_ = \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.ce  ? \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.fas_s1  : \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.sum_s1 ;
assign _188_ = \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.u1.a  + \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.u1.b ;
assign { \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.u1.cout , \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.u1.s  } = _188_ + \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.u1.cin ;
assign _189_ = \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.u2.a  + \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.u2.b ;
assign { \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.u2.cout , \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.u2.s  } = _189_ + \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.u2.cin ;
assign \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.bin_s0  = ~ \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.b ;
always @(posedge \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.clk )
\sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.bin_s1  <= _191_;
always @(posedge \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.clk )
\sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.ain_s1  <= _190_;
always @(posedge \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.clk )
\sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.sum_s1  <= _193_;
always @(posedge \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.clk )
\sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.carry_s1  <= _192_;
assign _191_ = \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.ce  ? \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.bin_s0 [27:14] : \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.bin_s1 ;
assign _190_ = \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.ce  ? \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.a [27:14] : \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.ain_s1 ;
assign _192_ = \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.ce  ? \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.facout_s1  : \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.carry_s1 ;
assign _193_ = \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.ce  ? \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.fas_s1  : \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.sum_s1 ;
assign _194_ = \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.u1.a  + \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.u1.b ;
assign { \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.u1.cout , \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.u1.s  } = _194_ + \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.u1.cin ;
assign _195_ = \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.u2.a  + \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.u2.b ;
assign { \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.u2.cout , \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.u2.s  } = _195_ + \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.u2.cin ;
assign \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.bin_s0  = ~ \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.b ;
always @(posedge \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.clk )
\sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.bin_s1  <= _197_;
always @(posedge \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.clk )
\sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.ain_s1  <= _196_;
always @(posedge \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.clk )
\sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.sum_s1  <= _199_;
always @(posedge \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.clk )
\sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.carry_s1  <= _198_;
assign _197_ = \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.ce  ? \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.bin_s0 [31:16] : \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.bin_s1 ;
assign _196_ = \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.ce  ? \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.a [31:16] : \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.ain_s1 ;
assign _198_ = \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.ce  ? \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.facout_s1  : \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.carry_s1 ;
assign _199_ = \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.ce  ? \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.fas_s1  : \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.sum_s1 ;
assign _200_ = \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.u1.a  + \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.u1.b ;
assign { \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.u1.cout , \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.u1.s  } = _200_ + \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.u1.cin ;
assign _201_ = \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.u2.a  + \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.u2.b ;
assign { \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.u2.cout , \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.u2.s  } = _201_ + \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.u2.cin ;
assign _202_ = op_7 > op_2;
assign _203_ = op_1[0] > op_2;
assign _204_ = | p_Result_s_reg_711;
assign _205_ = | trunc_ln851_reg_792;
assign op_6_V_fu_261_p2 = trunc_ln213_reg_658 | op_4[0];
assign or_ln340_fu_317_p2 = p_Result_3_reg_704 | overflow_fu_311_p2;
assign or_ln785_fu_302_p2 = newsignbit_reg_673 | icmp_ln768_reg_716;
always @(posedge ap_clk)
op_8_V_reg_761[18:0] <= 19'h00000;
always @(posedge ap_clk)
trunc_ln798_reg_918 <= _037_;
always @(posedge ap_clk)
trunc_ln798_1_reg_923 <= _036_;
always @(posedge ap_clk)
sh_reg_835 <= _031_;
always @(posedge ap_clk)
ret_V_9_reg_786 <= _026_;
always @(posedge ap_clk)
trunc_ln851_reg_792 <= _038_;
always @(posedge ap_clk)
sext_ln831_reg_797 <= _030_;
always @(posedge ap_clk)
ret_V_14_reg_906 <= _022_;
always @(posedge ap_clk)
ret_V_9_cast_reg_911 <= _025_;
always @(posedge ap_clk)
ret_V_11_reg_741 <= _019_;
always @(posedge ap_clk)
ret_1_reg_731 <= _018_;
always @(posedge ap_clk)
select_ln1192_reg_736 <= _028_;
always @(posedge ap_clk)
r_reg_933 <= _017_;
always @(posedge ap_clk)
ret_V_15_reg_938 <= _023_;
always @(posedge ap_clk)
p_Result_4_reg_820 <= _015_;
always @(posedge ap_clk)
ret_V_13_reg_825 <= _021_;
always @(posedge ap_clk)
select_ln69_reg_830 <= _029_;
always @(posedge ap_clk)
op_8_V_reg_761[19] <= _013_;
always @(posedge ap_clk)
ret_V_12_reg_776 <= _020_;
always @(posedge ap_clk)
tmp_2_reg_781 <= _033_;
always @(posedge ap_clk)
op_6_V_reg_699 <= _012_;
always @(posedge ap_clk)
p_Result_3_reg_704 <= _014_;
always @(posedge ap_clk)
p_Result_s_reg_711 <= _016_;
always @(posedge ap_clk)
ret_V_reg_881 <= _027_;
always @(posedge ap_clk)
op_16_V_reg_886 <= _010_;
always @(posedge ap_clk)
op_25_V_reg_891 <= _011_;
always @(posedge ap_clk)
trunc_ln213_reg_658 <= _034_;
always @(posedge ap_clk)
newsignbit_reg_673 <= _009_;
always @(posedge ap_clk)
lhs_V_4_reg_679 <= _008_;
always @(posedge ap_clk)
signbit_1_reg_684 <= _032_;
always @(posedge ap_clk)
trunc_ln728_reg_689 <= _035_;
always @(posedge ap_clk)
icmp_ln768_reg_716 <= _006_;
always @(posedge ap_clk)
ret_V_16_reg_958 <= _024_;
always @(posedge ap_clk)
add_ln69_3_reg_963 <= _003_;
always @(posedge ap_clk)
add_ln69_reg_856 <= _004_;
always @(posedge ap_clk)
add_ln69_1_reg_861 <= _002_;
always @(posedge ap_clk)
icmp_ln850_reg_804 <= _007_;
always @(posedge ap_clk)
add_ln691_reg_809 <= _001_;
always @(posedge ap_clk)
add_ln691_1_reg_928 <= _000_;
always @(posedge ap_clk)
ap_CS_fsm <= _005_;
assign _039_ = _043_ ? 2'h2 : 2'h1;
assign _206_ = ap_CS_fsm == 1'h1;
function [23:0] _569_;
input [23:0] a;
input [575:0] b;
input [23:0] s;
case (s)
24'b000000000000000000000001:
_569_ = b[23:0];
24'b000000000000000000000010:
_569_ = b[47:24];
24'b000000000000000000000100:
_569_ = b[71:48];
24'b000000000000000000001000:
_569_ = b[95:72];
24'b000000000000000000010000:
_569_ = b[119:96];
24'b000000000000000000100000:
_569_ = b[143:120];
24'b000000000000000001000000:
_569_ = b[167:144];
24'b000000000000000010000000:
_569_ = b[191:168];
24'b000000000000000100000000:
_569_ = b[215:192];
24'b000000000000001000000000:
_569_ = b[239:216];
24'b000000000000010000000000:
_569_ = b[263:240];
24'b000000000000100000000000:
_569_ = b[287:264];
24'b000000000001000000000000:
_569_ = b[311:288];
24'b000000000010000000000000:
_569_ = b[335:312];
24'b000000000100000000000000:
_569_ = b[359:336];
24'b000000001000000000000000:
_569_ = b[383:360];
24'b000000010000000000000000:
_569_ = b[407:384];
24'b000000100000000000000000:
_569_ = b[431:408];
24'b000001000000000000000000:
_569_ = b[455:432];
24'b000010000000000000000000:
_569_ = b[479:456];
24'b000100000000000000000000:
_569_ = b[503:480];
24'b001000000000000000000000:
_569_ = b[527:504];
24'b010000000000000000000000:
_569_ = b[551:528];
24'b100000000000000000000000:
_569_ = b[575:552];
24'b000000000000000000000000:
_569_ = a;
default:
_569_ = 24'bx;
endcase
endfunction
assign ap_NS_fsm = _569_(24'hxxxxxx, { 22'h000000, _039_, 552'h000004000008000010000020000040000080000100000200000400000800001000002000004000008000010000020000040000080000100000200000400000800000000001 }, { _206_, _229_, _228_, _227_, _226_, _225_, _224_, _223_, _222_, _221_, _220_, _219_, _218_, _217_, _216_, _215_, _214_, _213_, _212_, _211_, _210_, _209_, _208_, _207_ });
assign _207_ = ap_CS_fsm == 24'h800000;
assign _208_ = ap_CS_fsm == 23'h400000;
assign _209_ = ap_CS_fsm == 22'h200000;
assign _210_ = ap_CS_fsm == 21'h100000;
assign _211_ = ap_CS_fsm == 20'h80000;
assign _212_ = ap_CS_fsm == 19'h40000;
assign _213_ = ap_CS_fsm == 18'h20000;
assign _214_ = ap_CS_fsm == 17'h10000;
assign _215_ = ap_CS_fsm == 16'h8000;
assign _216_ = ap_CS_fsm == 15'h4000;
assign _217_ = ap_CS_fsm == 14'h2000;
assign _218_ = ap_CS_fsm == 13'h1000;
assign _219_ = ap_CS_fsm == 12'h800;
assign _220_ = ap_CS_fsm == 11'h400;
assign _221_ = ap_CS_fsm == 10'h200;
assign _222_ = ap_CS_fsm == 9'h100;
assign _223_ = ap_CS_fsm == 8'h80;
assign _224_ = ap_CS_fsm == 7'h40;
assign _225_ = ap_CS_fsm == 6'h20;
assign _226_ = ap_CS_fsm == 5'h10;
assign _227_ = ap_CS_fsm == 4'h8;
assign _228_ = ap_CS_fsm == 3'h4;
assign _229_ = ap_CS_fsm == 2'h2;
assign op_29_ap_vld = ap_CS_fsm[23] ? 1'h1 : 1'h0;
assign ap_idle = _042_ ? 1'h1 : 1'h0;
assign _037_ = _041_ ? grp_fu_509_p2[1:0] : trunc_ln798_reg_918;
assign _036_ = _040_ ? grp_fu_514_p2[1:0] : trunc_ln798_1_reg_923;
assign _031_ = ap_CS_fsm[11] ? grp_fu_425_p2 : sh_reg_835;
assign _030_ = ap_CS_fsm[8] ? { tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781 } : sext_ln831_reg_797;
assign _038_ = ap_CS_fsm[8] ? grp_fu_383_p2[18:0] : trunc_ln851_reg_792;
assign _026_ = ap_CS_fsm[8] ? grp_fu_383_p2 : ret_V_9_reg_786;
assign _025_ = ap_CS_fsm[16] ? grp_fu_567_p2[32:1] : ret_V_9_cast_reg_911;
assign _022_ = ap_CS_fsm[16] ? grp_fu_567_p2 : ret_V_14_reg_906;
assign _019_ = ap_CS_fsm[5] ? grp_fu_336_p2 : ret_V_11_reg_741;
assign _028_ = ap_CS_fsm[3] ? select_ln1192_fu_328_p3 : select_ln1192_reg_736;
assign _018_ = ap_CS_fsm[3] ? grp_fu_296_p2 : ret_1_reg_731;
assign _023_ = ap_CS_fsm[19] ? ret_V_15_fu_621_p3 : ret_V_15_reg_938;
assign _017_ = ap_CS_fsm[19] ? r_fu_596_p3 : r_reg_933;
assign _029_ = ap_CS_fsm[10] ? select_ln69_fu_479_p3 : select_ln69_reg_830;
assign _021_ = ap_CS_fsm[10] ? ret_V_13_fu_472_p3 : ret_V_13_reg_825;
assign _015_ = ap_CS_fsm[10] ? op_14[31] : p_Result_4_reg_820;
assign _033_ = ap_CS_fsm[7] ? grp_fu_355_p2[6:1] : tmp_2_reg_781;
assign _020_ = ap_CS_fsm[7] ? grp_fu_355_p2 : ret_V_12_reg_776;
assign _013_ = ap_CS_fsm[7] ? signbit_1_reg_684 : op_8_V_reg_761[19];
assign _016_ = ap_CS_fsm[1] ? grp_fu_221_p2[9:1] : p_Result_s_reg_711;
assign _014_ = ap_CS_fsm[1] ? grp_fu_221_p2[9] : p_Result_3_reg_704;
assign _012_ = ap_CS_fsm[1] ? op_6_V_fu_261_p2 : op_6_V_reg_699;
assign _011_ = ap_CS_fsm[14] ? grp_fu_538_p2 : op_25_V_reg_891;
assign _010_ = ap_CS_fsm[14] ? grp_fu_529_p2[21:18] : op_16_V_reg_886;
assign _027_ = ap_CS_fsm[14] ? grp_fu_529_p2 : ret_V_reg_881;
assign _035_ = ap_CS_fsm[0] ? op_7[2:0] : trunc_ln728_reg_689;
assign _032_ = ap_CS_fsm[0] ? signbit_1_fu_247_p2 : signbit_1_reg_684;
assign _008_ = ap_CS_fsm[0] ? lhs_V_4_fu_237_p2 : lhs_V_4_reg_679;
assign _009_ = ap_CS_fsm[0] ? newsignbit_fu_227_p2 : newsignbit_reg_673;
assign _034_ = ap_CS_fsm[0] ? op_2[0] : trunc_ln213_reg_658;
assign _006_ = ap_CS_fsm[2] ? icmp_ln768_fu_284_p2 : icmp_ln768_reg_716;
assign _003_ = ap_CS_fsm[21] ? grp_fu_643_p2 : add_ln69_3_reg_963;
assign _024_ = ap_CS_fsm[21] ? grp_fu_631_p2 : ret_V_16_reg_958;
assign _002_ = ap_CS_fsm[12] ? grp_fu_500_p2 : add_ln69_1_reg_861;
assign _004_ = ap_CS_fsm[12] ? grp_fu_495_p2 : add_ln69_reg_856;
assign _001_ = ap_CS_fsm[9] ? grp_fu_406_p2 : add_ln691_reg_809;
assign _007_ = ap_CS_fsm[9] ? icmp_ln850_fu_412_p2 : icmp_ln850_reg_804;
assign _000_ = ap_CS_fsm[18] ? grp_fu_583_p2 : add_ln691_1_reg_928;
assign _005_ = ap_rst ? 24'h000001 : ap_NS_fsm;
assign icmp_ln768_fu_284_p2 = _204_ ? 1'h1 : 1'h0;
assign icmp_ln850_fu_412_p2 = _205_ ? 1'h1 : 1'h0;
assign lhs_V_4_fu_237_p2 = _202_ ? 1'h1 : 1'h0;
assign op_10_V_fu_322_p3 = or_ln340_fu_317_p2 ? p_Result_3_reg_704 : newsignbit_reg_673;
assign r_fu_596_p3 = p_Result_4_reg_820 ? trunc_ln798_reg_918 : trunc_ln798_1_reg_923;
assign ret_V_13_fu_472_p3 = ret_V_12_reg_776[6] ? select_ln850_fu_466_p3 : sext_ln831_reg_797;
assign ret_V_15_fu_621_p3 = ret_V_14_reg_906[33] ? select_ln850_1_fu_615_p3 : ret_V_9_cast_reg_911;
assign select_ln1192_fu_328_p3 = op_10_V_fu_322_p3 ? 5'h1f : 5'h00;
assign select_ln69_fu_479_p3 = ret_V_10_fu_450_p2 ? 3'h7 : 3'h0;
assign select_ln850_1_fu_615_p3 = ret_V_reg_881[18] ? add_ln691_1_reg_928 : ret_V_9_cast_reg_911;
assign select_ln850_fu_466_p3 = op_11[0] ? add_ln691_reg_809 : sext_ln831_reg_797;
assign signbit_1_fu_247_p2 = _203_ ? 1'h1 : 1'h0;
assign newsignbit_fu_227_p2 = op_5[0] ^ op_7[0];
assign ret_V_10_fu_450_p2 = ret_V_9_reg_786[19] ^ and_ln353_fu_445_p2;
assign ap_CS_fsm_state1 = ap_CS_fsm[0];
assign ap_CS_fsm_state10 = ap_CS_fsm[9];
assign ap_CS_fsm_state11 = ap_CS_fsm[10];
assign ap_CS_fsm_state12 = ap_CS_fsm[11];
assign ap_CS_fsm_state13 = ap_CS_fsm[12];
assign ap_CS_fsm_state14 = ap_CS_fsm[13];
assign ap_CS_fsm_state15 = ap_CS_fsm[14];
assign ap_CS_fsm_state16 = ap_CS_fsm[15];
assign ap_CS_fsm_state17 = ap_CS_fsm[16];
assign ap_CS_fsm_state18 = ap_CS_fsm[17];
assign ap_CS_fsm_state19 = ap_CS_fsm[18];
assign ap_CS_fsm_state2 = ap_CS_fsm[1];
assign ap_CS_fsm_state20 = ap_CS_fsm[19];
assign ap_CS_fsm_state21 = ap_CS_fsm[20];
assign ap_CS_fsm_state22 = ap_CS_fsm[21];
assign ap_CS_fsm_state23 = ap_CS_fsm[22];
assign ap_CS_fsm_state24 = ap_CS_fsm[23];
assign ap_CS_fsm_state3 = ap_CS_fsm[2];
assign ap_CS_fsm_state4 = ap_CS_fsm[3];
assign ap_CS_fsm_state5 = ap_CS_fsm[4];
assign ap_CS_fsm_state6 = ap_CS_fsm[5];
assign ap_CS_fsm_state7 = ap_CS_fsm[6];
assign ap_CS_fsm_state8 = ap_CS_fsm[7];
assign ap_CS_fsm_state9 = ap_CS_fsm[8];
assign ap_done = op_29_ap_vld;
assign ap_ready = op_29_ap_vld;
assign grp_fu_221_p0 = { 2'h0, op_7 };
assign grp_fu_221_p1 = { op_5[7], op_5[7], op_5 };
assign grp_fu_296_p0 = { op_0[3], op_0 };
assign grp_fu_296_p1 = { 4'h0, op_6_V_reg_699 };
assign grp_fu_355_p0 = { ret_V_11_reg_741[4], ret_V_11_reg_741, 1'h0 };
assign grp_fu_355_p1 = { op_11[1], op_11[1], op_11[1], op_11[1], op_11[1], op_11 };
assign grp_fu_383_p0 = { op_4[7], op_4, 19'h00000 };
assign grp_fu_383_p1 = { 8'h00, signbit_1_reg_684, 19'h00000 };
assign grp_fu_406_p0 = { tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781 };
assign grp_fu_495_p1 = { op_15[15], op_15[15], op_15[15], op_15[15], op_15[15], op_15[15], op_15[15], op_15[15], op_15[15], op_15[15], op_15[15], op_15[15], op_15[15], op_15[15], op_15[15], op_15[15], op_15 };
assign grp_fu_500_p0 = { op_12[1], op_12 };
assign grp_fu_529_p0 = { trunc_ln728_reg_689, 19'h00000 };
assign grp_fu_529_p1 = { 2'h0, op_8_V_reg_761 };
assign grp_fu_538_p0 = { add_ln69_1_reg_861[2], add_ln69_1_reg_861[2], add_ln69_1_reg_861[2], add_ln69_1_reg_861[2], add_ln69_1_reg_861[2], add_ln69_1_reg_861[2], add_ln69_1_reg_861[2], add_ln69_1_reg_861[2], add_ln69_1_reg_861[2], add_ln69_1_reg_861[2], add_ln69_1_reg_861[2], add_ln69_1_reg_861[2], add_ln69_1_reg_861[2], add_ln69_1_reg_861[2], add_ln69_1_reg_861[2], add_ln69_1_reg_861[2], add_ln69_1_reg_861[2], add_ln69_1_reg_861[2], add_ln69_1_reg_861[2], add_ln69_1_reg_861[2], add_ln69_1_reg_861[2], add_ln69_1_reg_861[2], add_ln69_1_reg_861[2], add_ln69_1_reg_861[2], add_ln69_1_reg_861[2], add_ln69_1_reg_861[2], add_ln69_1_reg_861[2], add_ln69_1_reg_861[2], add_ln69_1_reg_861[2], add_ln69_1_reg_861 };
assign grp_fu_567_p0 = { op_25_V_reg_891[31], op_25_V_reg_891, 1'h0 };
assign grp_fu_567_p1 = { op_16_V_reg_886[3], op_16_V_reg_886[3], op_16_V_reg_886[3], op_16_V_reg_886[3], op_16_V_reg_886[3], op_16_V_reg_886[3], op_16_V_reg_886[3], op_16_V_reg_886[3], op_16_V_reg_886[3], op_16_V_reg_886[3], op_16_V_reg_886[3], op_16_V_reg_886[3], op_16_V_reg_886[3], op_16_V_reg_886[3], op_16_V_reg_886[3], op_16_V_reg_886[3], op_16_V_reg_886[3], op_16_V_reg_886[3], op_16_V_reg_886[3], op_16_V_reg_886[3], op_16_V_reg_886[3], op_16_V_reg_886[3], op_16_V_reg_886[3], op_16_V_reg_886[3], op_16_V_reg_886[3], op_16_V_reg_886[3], op_16_V_reg_886[3], op_16_V_reg_886[3], op_16_V_reg_886[3], op_16_V_reg_886[3], op_16_V_reg_886 };
assign grp_fu_631_p1 = { 31'h00000000, lhs_V_4_reg_679 };
assign grp_fu_643_p0 = { op_19[15], op_19 };
assign grp_fu_643_p1 = { r_reg_933[1], r_reg_933[1], r_reg_933[1], r_reg_933[1], r_reg_933[1], r_reg_933[1], r_reg_933[1], r_reg_933[1], r_reg_933[1], r_reg_933[1], r_reg_933[1], r_reg_933[1], r_reg_933[1], r_reg_933[1], r_reg_933[1], r_reg_933 };
assign grp_fu_652_p0 = { add_ln69_3_reg_963[16], add_ln69_3_reg_963[16], add_ln69_3_reg_963[16], add_ln69_3_reg_963[16], add_ln69_3_reg_963[16], add_ln69_3_reg_963[16], add_ln69_3_reg_963[16], add_ln69_3_reg_963[16], add_ln69_3_reg_963[16], add_ln69_3_reg_963[16], add_ln69_3_reg_963[16], add_ln69_3_reg_963[16], add_ln69_3_reg_963[16], add_ln69_3_reg_963[16], add_ln69_3_reg_963[16], add_ln69_3_reg_963 };
assign lhs_V_fu_368_p3 = { op_4, 19'h00000 };
assign op_29 = grp_fu_652_p2;
assign op_3_V_fu_197_p1 = op_1[0];
assign op_8_V_fu_361_p3 = { signbit_1_reg_684, 19'h00000 };
assign p_Result_1_fu_456_p3 = ret_V_12_reg_776[6];
assign p_Result_2_fu_601_p3 = ret_V_14_reg_906[33];
assign p_Result_s_12_fu_438_p3 = ret_V_9_reg_786[27];
assign rhs_4_fu_556_p3 = { op_25_V_reg_891, 1'h0 };
assign sext_ln1192_fu_340_p0 = op_11;
assign sext_ln215_fu_205_p0 = op_5;
assign sext_ln781_fu_505_p1 = { op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9 };
assign sext_ln831_fu_403_p1 = { tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781 };
assign tmp_4_fu_344_p3 = { ret_V_11_reg_741, 1'h0 };
assign tmp_6_fu_608_p3 = ret_V_reg_881[18];
assign tmp_fu_431_p3 = ret_V_9_reg_786[19];
assign trunc_ln1346_1_fu_217_p1 = op_7[0];
assign trunc_ln1346_fu_213_p0 = op_5;
assign trunc_ln1346_fu_213_p1 = op_5[0];
assign trunc_ln213_1_fu_257_p1 = op_4[0];
assign trunc_ln213_fu_201_p1 = op_2[0];
assign trunc_ln728_fu_253_p1 = op_7[2:0];
assign trunc_ln798_1_fu_592_p1 = grp_fu_514_p2[1:0];
assign trunc_ln798_fu_588_p1 = grp_fu_509_p2[1:0];
assign trunc_ln851_1_fu_463_p0 = op_11;
assign trunc_ln851_1_fu_463_p1 = op_11[0];
assign trunc_ln851_fu_399_p1 = grp_fu_383_p2[18:0];
assign zext_ln878_1_fu_243_p1 = { 15'h0000, op_1[0] };
assign zext_ln878_fu_233_p1 = { 8'h00, op_7 };
assign \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.ain_s0  = \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.a ;
assign \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.s  = { \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.fas_s2 , \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.sum_s1  };
assign \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.u2.a  = \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.ain_s1 ;
assign \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.u2.b  = \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.bin_s1 ;
assign \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.u2.cin  = \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.carry_s1 ;
assign \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.facout_s2  = \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.u2.cout ;
assign \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.fas_s2  = \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.u2.s ;
assign \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.u1.a  = \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.a [15:0];
assign \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.u1.b  = \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.bin_s0 [15:0];
assign \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.u1.cin  = 1'h1;
assign \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.facout_s1  = \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.u1.cout ;
assign \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.fas_s1  = \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.u1.s ;
assign \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.a  = \sub_32ns_32ns_32_2_1_U7.din0 ;
assign \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.b  = \sub_32ns_32ns_32_2_1_U7.din1 ;
assign \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.ce  = \sub_32ns_32ns_32_2_1_U7.ce ;
assign \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.clk  = \sub_32ns_32ns_32_2_1_U7.clk ;
assign \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.reset  = \sub_32ns_32ns_32_2_1_U7.reset ;
assign \sub_32ns_32ns_32_2_1_U7.dout  = \sub_32ns_32ns_32_2_1_U7.top_sub_32ns_32ns_32_2_1_Adder_6_U.s ;
assign \sub_32ns_32ns_32_2_1_U7.ce  = 1'h1;
assign \sub_32ns_32ns_32_2_1_U7.clk  = ap_clk;
assign \sub_32ns_32ns_32_2_1_U7.din0  = 32'd0;
assign \sub_32ns_32ns_32_2_1_U7.din1  = op_14;
assign grp_fu_425_p2 = \sub_32ns_32ns_32_2_1_U7.dout ;
assign \sub_32ns_32ns_32_2_1_U7.reset  = ap_rst;
assign \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.ain_s0  = \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.a ;
assign \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.s  = { \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.fas_s2 , \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.sum_s1  };
assign \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.u2.a  = \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.ain_s1 ;
assign \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.u2.b  = \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.bin_s1 ;
assign \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.u2.cin  = \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.carry_s1 ;
assign \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.facout_s2  = \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.u2.cout ;
assign \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.fas_s2  = \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.u2.s ;
assign \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.u1.a  = \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.a [13:0];
assign \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.u1.b  = \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.bin_s0 [13:0];
assign \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.u1.cin  = 1'h1;
assign \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.facout_s1  = \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.u1.cout ;
assign \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.fas_s1  = \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.u1.s ;
assign \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.a  = \sub_28s_28ns_28_2_1_U5.din0 ;
assign \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.b  = \sub_28s_28ns_28_2_1_U5.din1 ;
assign \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.ce  = \sub_28s_28ns_28_2_1_U5.ce ;
assign \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.clk  = \sub_28s_28ns_28_2_1_U5.clk ;
assign \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.reset  = \sub_28s_28ns_28_2_1_U5.reset ;
assign \sub_28s_28ns_28_2_1_U5.dout  = \sub_28s_28ns_28_2_1_U5.top_sub_28s_28ns_28_2_1_Adder_4_U.s ;
assign \sub_28s_28ns_28_2_1_U5.ce  = 1'h1;
assign \sub_28s_28ns_28_2_1_U5.clk  = ap_clk;
assign \sub_28s_28ns_28_2_1_U5.din0  = { op_4[7], op_4, 19'h00000 };
assign \sub_28s_28ns_28_2_1_U5.din1  = { 8'h00, signbit_1_reg_684, 19'h00000 };
assign grp_fu_383_p2 = \sub_28s_28ns_28_2_1_U5.dout ;
assign \sub_28s_28ns_28_2_1_U5.reset  = ap_rst;
assign \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.ain_s0  = \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.a ;
assign \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.s  = { \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.fas_s2 , \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.sum_s1  };
assign \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.u2.a  = \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.ain_s1 ;
assign \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.u2.b  = \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.bin_s1 ;
assign \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.u2.cin  = \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.carry_s1 ;
assign \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.facout_s2  = \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.u2.cout ;
assign \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.fas_s2  = \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.u2.s ;
assign \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.u1.a  = \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.a [10:0];
assign \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.u1.b  = \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.bin_s0 [10:0];
assign \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.u1.cin  = 1'h1;
assign \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.facout_s1  = \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.u1.cout ;
assign \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.fas_s1  = \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.u1.s ;
assign \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.a  = \sub_22ns_22ns_22_2_1_U12.din0 ;
assign \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.b  = \sub_22ns_22ns_22_2_1_U12.din1 ;
assign \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.ce  = \sub_22ns_22ns_22_2_1_U12.ce ;
assign \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.clk  = \sub_22ns_22ns_22_2_1_U12.clk ;
assign \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.reset  = \sub_22ns_22ns_22_2_1_U12.reset ;
assign \sub_22ns_22ns_22_2_1_U12.dout  = \sub_22ns_22ns_22_2_1_U12.top_sub_22ns_22ns_22_2_1_Adder_9_U.s ;
assign \sub_22ns_22ns_22_2_1_U12.ce  = 1'h1;
assign \sub_22ns_22ns_22_2_1_U12.clk  = ap_clk;
assign \sub_22ns_22ns_22_2_1_U12.din0  = { trunc_ln728_reg_689, 19'h00000 };
assign \sub_22ns_22ns_22_2_1_U12.din1  = { 2'h0, op_8_V_reg_761 };
assign grp_fu_529_p2 = \sub_22ns_22ns_22_2_1_U12.dout ;
assign \sub_22ns_22ns_22_2_1_U12.reset  = ap_rst;
assign \shl_32s_32ns_32_7_1_U11.din1_cast  = \shl_32s_32ns_32_7_1_U11.din1 ;
assign \shl_32s_32ns_32_7_1_U11.din1_mask  = 32'd31;
assign \shl_32s_32ns_32_7_1_U11.ce  = 1'h1;
assign \shl_32s_32ns_32_7_1_U11.clk  = ap_clk;
assign \shl_32s_32ns_32_7_1_U11.din0  = { op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9 };
assign \shl_32s_32ns_32_7_1_U11.din1  = op_14;
assign grp_fu_514_p2 = \shl_32s_32ns_32_7_1_U11.dout ;
assign \shl_32s_32ns_32_7_1_U11.reset  = ap_rst;
assign \ashr_32s_32ns_32_7_1_U10.din1_cast  = \ashr_32s_32ns_32_7_1_U10.din1 ;
assign \ashr_32s_32ns_32_7_1_U10.din1_mask  = 32'd31;
assign \ashr_32s_32ns_32_7_1_U10.ce  = 1'h1;
assign \ashr_32s_32ns_32_7_1_U10.clk  = ap_clk;
assign \ashr_32s_32ns_32_7_1_U10.din0  = { op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9[1], op_9 };
assign \ashr_32s_32ns_32_7_1_U10.din1  = sh_reg_835;
assign grp_fu_509_p2 = \ashr_32s_32ns_32_7_1_U10.dout ;
assign \ashr_32s_32ns_32_7_1_U10.reset  = ap_rst;
assign \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.ain_s0  = \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.a ;
assign \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.bin_s0  = \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.b ;
assign \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.s  = { \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.fas_s2 , \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.sum_s1  };
assign \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.u2.a  = \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.ain_s1 ;
assign \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.u2.b  = \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.bin_s1 ;
assign \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.u2.cin  = \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.carry_s1 ;
assign \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.facout_s2  = \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.u2.cout ;
assign \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.fas_s2  = \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.u2.s ;
assign \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.u1.a  = \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.a [2:0];
assign \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.u1.b  = \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.b [2:0];
assign \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.u1.cin  = 1'h0;
assign \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.facout_s1  = \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.u1.cout ;
assign \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.fas_s1  = \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.u1.s ;
assign \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.a  = \add_7s_7s_7_2_1_U4.din0 ;
assign \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.b  = \add_7s_7s_7_2_1_U4.din1 ;
assign \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.ce  = \add_7s_7s_7_2_1_U4.ce ;
assign \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.clk  = \add_7s_7s_7_2_1_U4.clk ;
assign \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.reset  = \add_7s_7s_7_2_1_U4.reset ;
assign \add_7s_7s_7_2_1_U4.dout  = \add_7s_7s_7_2_1_U4.top_add_7s_7s_7_2_1_Adder_3_U.s ;
assign \add_7s_7s_7_2_1_U4.ce  = 1'h1;
assign \add_7s_7s_7_2_1_U4.clk  = ap_clk;
assign \add_7s_7s_7_2_1_U4.din0  = { ret_V_11_reg_741[4], ret_V_11_reg_741, 1'h0 };
assign \add_7s_7s_7_2_1_U4.din1  = { op_11[1], op_11[1], op_11[1], op_11[1], op_11[1], op_11 };
assign grp_fu_355_p2 = \add_7s_7s_7_2_1_U4.dout ;
assign \add_7s_7s_7_2_1_U4.reset  = ap_rst;
assign \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.ain_s0  = \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.a ;
assign \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.bin_s0  = \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.b ;
assign \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.s  = { \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.fas_s2 , \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.sum_s1  };
assign \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.u2.a  = \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.ain_s1 ;
assign \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.u2.b  = \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.bin_s1 ;
assign \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.u2.cin  = \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.carry_s1 ;
assign \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.facout_s2  = \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.u2.cout ;
assign \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.fas_s2  = \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.u2.s ;
assign \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.u1.a  = \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.a [1:0];
assign \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.u1.b  = \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.b [1:0];
assign \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.u1.cin  = 1'h0;
assign \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.facout_s1  = \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.u1.cout ;
assign \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.fas_s1  = \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.u1.s ;
assign \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.a  = \add_5s_5ns_5_2_1_U2.din0 ;
assign \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.b  = \add_5s_5ns_5_2_1_U2.din1 ;
assign \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.ce  = \add_5s_5ns_5_2_1_U2.ce ;
assign \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.clk  = \add_5s_5ns_5_2_1_U2.clk ;
assign \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.reset  = \add_5s_5ns_5_2_1_U2.reset ;
assign \add_5s_5ns_5_2_1_U2.dout  = \add_5s_5ns_5_2_1_U2.top_add_5s_5ns_5_2_1_Adder_1_U.s ;
assign \add_5s_5ns_5_2_1_U2.ce  = 1'h1;
assign \add_5s_5ns_5_2_1_U2.clk  = ap_clk;
assign \add_5s_5ns_5_2_1_U2.din0  = { op_0[3], op_0 };
assign \add_5s_5ns_5_2_1_U2.din1  = { 4'h0, op_6_V_reg_699 };
assign grp_fu_296_p2 = \add_5s_5ns_5_2_1_U2.dout ;
assign \add_5s_5ns_5_2_1_U2.reset  = ap_rst;
assign \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.ain_s0  = \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.a ;
assign \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.bin_s0  = \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.b ;
assign \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.s  = { \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.fas_s2 , \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.sum_s1  };
assign \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.u2.a  = \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.ain_s1 ;
assign \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.u2.b  = \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.bin_s1 ;
assign \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.u2.cin  = \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.carry_s1 ;
assign \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.facout_s2  = \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.u2.cout ;
assign \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.fas_s2  = \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.u2.s ;
assign \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.u1.a  = \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.a [1:0];
assign \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.u1.b  = \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.b [1:0];
assign \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.u1.cin  = 1'h0;
assign \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.facout_s1  = \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.u1.cout ;
assign \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.fas_s1  = \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.u1.s ;
assign \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.a  = \add_5ns_5ns_5_2_1_U3.din0 ;
assign \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.b  = \add_5ns_5ns_5_2_1_U3.din1 ;
assign \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.ce  = \add_5ns_5ns_5_2_1_U3.ce ;
assign \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.clk  = \add_5ns_5ns_5_2_1_U3.clk ;
assign \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.reset  = \add_5ns_5ns_5_2_1_U3.reset ;
assign \add_5ns_5ns_5_2_1_U3.dout  = \add_5ns_5ns_5_2_1_U3.top_add_5ns_5ns_5_2_1_Adder_2_U.s ;
assign \add_5ns_5ns_5_2_1_U3.ce  = 1'h1;
assign \add_5ns_5ns_5_2_1_U3.clk  = ap_clk;
assign \add_5ns_5ns_5_2_1_U3.din0  = ret_1_reg_731;
assign \add_5ns_5ns_5_2_1_U3.din1  = select_ln1192_reg_736;
assign grp_fu_336_p2 = \add_5ns_5ns_5_2_1_U3.dout ;
assign \add_5ns_5ns_5_2_1_U3.reset  = ap_rst;
assign \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.ain_s0  = \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.a ;
assign \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.bin_s0  = \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.b ;
assign \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.s  = { \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.fas_s2 , \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.sum_s1  };
assign \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.u2.a  = \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.ain_s1 ;
assign \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.u2.b  = \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.bin_s1 ;
assign \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.u2.cin  = \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.carry_s1 ;
assign \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.facout_s2  = \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.u2.cout ;
assign \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.fas_s2  = \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.u2.s ;
assign \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.u1.a  = \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.a [0];
assign \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.u1.b  = \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.b [0];
assign \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.u1.cin  = 1'h0;
assign \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.facout_s1  = \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.u1.cout ;
assign \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.fas_s1  = \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.u1.s ;
assign \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.a  = \add_3s_3ns_3_2_1_U9.din0 ;
assign \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.b  = \add_3s_3ns_3_2_1_U9.din1 ;
assign \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.ce  = \add_3s_3ns_3_2_1_U9.ce ;
assign \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.clk  = \add_3s_3ns_3_2_1_U9.clk ;
assign \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.reset  = \add_3s_3ns_3_2_1_U9.reset ;
assign \add_3s_3ns_3_2_1_U9.dout  = \add_3s_3ns_3_2_1_U9.top_add_3s_3ns_3_2_1_Adder_8_U.s ;
assign \add_3s_3ns_3_2_1_U9.ce  = 1'h1;
assign \add_3s_3ns_3_2_1_U9.clk  = ap_clk;
assign \add_3s_3ns_3_2_1_U9.din0  = { op_12[1], op_12 };
assign \add_3s_3ns_3_2_1_U9.din1  = select_ln69_reg_830;
assign grp_fu_500_p2 = \add_3s_3ns_3_2_1_U9.dout ;
assign \add_3s_3ns_3_2_1_U9.reset  = ap_rst;
assign \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.ain_s0  = \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.a ;
assign \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.bin_s0  = \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.b ;
assign \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.s  = { \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.fas_s2 , \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.sum_s1  };
assign \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.u2.a  = \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.ain_s1 ;
assign \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.u2.b  = \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.bin_s1 ;
assign \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.u2.cin  = \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.carry_s1 ;
assign \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.facout_s2  = \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.u2.cout ;
assign \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.fas_s2  = \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.u2.s ;
assign \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.u1.a  = \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.a [16:0];
assign \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.u1.b  = \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.b [16:0];
assign \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.u1.cin  = 1'h0;
assign \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.facout_s1  = \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.u1.cout ;
assign \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.fas_s1  = \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.u1.s ;
assign \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.a  = \add_34s_34s_34_2_1_U14.din0 ;
assign \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.b  = \add_34s_34s_34_2_1_U14.din1 ;
assign \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.ce  = \add_34s_34s_34_2_1_U14.ce ;
assign \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.clk  = \add_34s_34s_34_2_1_U14.clk ;
assign \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.reset  = \add_34s_34s_34_2_1_U14.reset ;
assign \add_34s_34s_34_2_1_U14.dout  = \add_34s_34s_34_2_1_U14.top_add_34s_34s_34_2_1_Adder_10_U.s ;
assign \add_34s_34s_34_2_1_U14.ce  = 1'h1;
assign \add_34s_34s_34_2_1_U14.clk  = ap_clk;
assign \add_34s_34s_34_2_1_U14.din0  = { op_25_V_reg_891[31], op_25_V_reg_891, 1'h0 };
assign \add_34s_34s_34_2_1_U14.din1  = { op_16_V_reg_886[3], op_16_V_reg_886[3], op_16_V_reg_886[3], op_16_V_reg_886[3], op_16_V_reg_886[3], op_16_V_reg_886[3], op_16_V_reg_886[3], op_16_V_reg_886[3], op_16_V_reg_886[3], op_16_V_reg_886[3], op_16_V_reg_886[3], op_16_V_reg_886[3], op_16_V_reg_886[3], op_16_V_reg_886[3], op_16_V_reg_886[3], op_16_V_reg_886[3], op_16_V_reg_886[3], op_16_V_reg_886[3], op_16_V_reg_886[3], op_16_V_reg_886[3], op_16_V_reg_886[3], op_16_V_reg_886[3], op_16_V_reg_886[3], op_16_V_reg_886[3], op_16_V_reg_886[3], op_16_V_reg_886[3], op_16_V_reg_886[3], op_16_V_reg_886[3], op_16_V_reg_886[3], op_16_V_reg_886[3], op_16_V_reg_886 };
assign grp_fu_567_p2 = \add_34s_34s_34_2_1_U14.dout ;
assign \add_34s_34s_34_2_1_U14.reset  = ap_rst;
assign \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.ain_s0  = \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.a ;
assign \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.bin_s0  = \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.b ;
assign \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.s  = { \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.fas_s2 , \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.sum_s1  };
assign \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.u2.a  = \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.ain_s1 ;
assign \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.u2.b  = \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.bin_s1 ;
assign \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.u2.cin  = \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.carry_s1 ;
assign \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.facout_s2  = \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.u2.cout ;
assign \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.fas_s2  = \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.u2.s ;
assign \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.u1.a  = \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.a [15:0];
assign \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.u1.b  = \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.b [15:0];
assign \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.u1.cin  = 1'h0;
assign \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.facout_s1  = \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.u1.cout ;
assign \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.fas_s1  = \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.u1.s ;
assign \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.a  = \add_32s_32ns_32_2_1_U6.din0 ;
assign \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.b  = \add_32s_32ns_32_2_1_U6.din1 ;
assign \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.ce  = \add_32s_32ns_32_2_1_U6.ce ;
assign \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.clk  = \add_32s_32ns_32_2_1_U6.clk ;
assign \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.reset  = \add_32s_32ns_32_2_1_U6.reset ;
assign \add_32s_32ns_32_2_1_U6.dout  = \add_32s_32ns_32_2_1_U6.top_add_32s_32ns_32_2_1_Adder_5_U.s ;
assign \add_32s_32ns_32_2_1_U6.ce  = 1'h1;
assign \add_32s_32ns_32_2_1_U6.clk  = ap_clk;
assign \add_32s_32ns_32_2_1_U6.din0  = { tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781[5], tmp_2_reg_781 };
assign \add_32s_32ns_32_2_1_U6.din1  = 32'd1;
assign grp_fu_406_p2 = \add_32s_32ns_32_2_1_U6.dout ;
assign \add_32s_32ns_32_2_1_U6.reset  = ap_rst;
assign \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.ain_s0  = \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.a ;
assign \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.bin_s0  = \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.b ;
assign \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.s  = { \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.fas_s2 , \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.sum_s1  };
assign \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.u2.a  = \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.ain_s1 ;
assign \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.u2.b  = \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.bin_s1 ;
assign \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.u2.cin  = \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.carry_s1 ;
assign \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.facout_s2  = \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.u2.cout ;
assign \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.fas_s2  = \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.u2.s ;
assign \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.u1.a  = \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.a [15:0];
assign \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.u1.b  = \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.b [15:0];
assign \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.u1.cin  = 1'h0;
assign \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.facout_s1  = \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.u1.cout ;
assign \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.fas_s1  = \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.u1.s ;
assign \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.a  = \add_32s_32ns_32_2_1_U18.din0 ;
assign \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.b  = \add_32s_32ns_32_2_1_U18.din1 ;
assign \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.ce  = \add_32s_32ns_32_2_1_U18.ce ;
assign \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.clk  = \add_32s_32ns_32_2_1_U18.clk ;
assign \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.reset  = \add_32s_32ns_32_2_1_U18.reset ;
assign \add_32s_32ns_32_2_1_U18.dout  = \add_32s_32ns_32_2_1_U18.top_add_32s_32ns_32_2_1_Adder_5_U.s ;
assign \add_32s_32ns_32_2_1_U18.ce  = 1'h1;
assign \add_32s_32ns_32_2_1_U18.clk  = ap_clk;
assign \add_32s_32ns_32_2_1_U18.din0  = { add_ln69_3_reg_963[16], add_ln69_3_reg_963[16], add_ln69_3_reg_963[16], add_ln69_3_reg_963[16], add_ln69_3_reg_963[16], add_ln69_3_reg_963[16], add_ln69_3_reg_963[16], add_ln69_3_reg_963[16], add_ln69_3_reg_963[16], add_ln69_3_reg_963[16], add_ln69_3_reg_963[16], add_ln69_3_reg_963[16], add_ln69_3_reg_963[16], add_ln69_3_reg_963[16], add_ln69_3_reg_963[16], add_ln69_3_reg_963 };
assign \add_32s_32ns_32_2_1_U18.din1  = ret_V_16_reg_958;
assign grp_fu_652_p2 = \add_32s_32ns_32_2_1_U18.dout ;
assign \add_32s_32ns_32_2_1_U18.reset  = ap_rst;
assign \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.ain_s0  = \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.a ;
assign \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.bin_s0  = \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.b ;
assign \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.s  = { \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.fas_s2 , \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.sum_s1  };
assign \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.u2.a  = \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.ain_s1 ;
assign \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.u2.b  = \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.bin_s1 ;
assign \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.u2.cin  = \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.carry_s1 ;
assign \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.facout_s2  = \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.u2.cout ;
assign \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.fas_s2  = \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.u2.s ;
assign \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.u1.a  = \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.a [15:0];
assign \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.u1.b  = \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.b [15:0];
assign \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.u1.cin  = 1'h0;
assign \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.facout_s1  = \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.u1.cout ;
assign \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.fas_s1  = \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.u1.s ;
assign \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.a  = \add_32s_32ns_32_2_1_U13.din0 ;
assign \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.b  = \add_32s_32ns_32_2_1_U13.din1 ;
assign \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.ce  = \add_32s_32ns_32_2_1_U13.ce ;
assign \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.clk  = \add_32s_32ns_32_2_1_U13.clk ;
assign \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.reset  = \add_32s_32ns_32_2_1_U13.reset ;
assign \add_32s_32ns_32_2_1_U13.dout  = \add_32s_32ns_32_2_1_U13.top_add_32s_32ns_32_2_1_Adder_5_U.s ;
assign \add_32s_32ns_32_2_1_U13.ce  = 1'h1;
assign \add_32s_32ns_32_2_1_U13.clk  = ap_clk;
assign \add_32s_32ns_32_2_1_U13.din0  = { add_ln69_1_reg_861[2], add_ln69_1_reg_861[2], add_ln69_1_reg_861[2], add_ln69_1_reg_861[2], add_ln69_1_reg_861[2], add_ln69_1_reg_861[2], add_ln69_1_reg_861[2], add_ln69_1_reg_861[2], add_ln69_1_reg_861[2], add_ln69_1_reg_861[2], add_ln69_1_reg_861[2], add_ln69_1_reg_861[2], add_ln69_1_reg_861[2], add_ln69_1_reg_861[2], add_ln69_1_reg_861[2], add_ln69_1_reg_861[2], add_ln69_1_reg_861[2], add_ln69_1_reg_861[2], add_ln69_1_reg_861[2], add_ln69_1_reg_861[2], add_ln69_1_reg_861[2], add_ln69_1_reg_861[2], add_ln69_1_reg_861[2], add_ln69_1_reg_861[2], add_ln69_1_reg_861[2], add_ln69_1_reg_861[2], add_ln69_1_reg_861[2], add_ln69_1_reg_861[2], add_ln69_1_reg_861[2], add_ln69_1_reg_861 };
assign \add_32s_32ns_32_2_1_U13.din1  = add_ln69_reg_856;
assign grp_fu_538_p2 = \add_32s_32ns_32_2_1_U13.dout ;
assign \add_32s_32ns_32_2_1_U13.reset  = ap_rst;
assign \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.ain_s0  = \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.a ;
assign \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.bin_s0  = \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.b ;
assign \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.s  = { \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.fas_s2 , \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.sum_s1  };
assign \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.u2.a  = \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.ain_s1 ;
assign \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.u2.b  = \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.bin_s1 ;
assign \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.u2.cin  = \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.carry_s1 ;
assign \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.facout_s2  = \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.u2.cout ;
assign \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.fas_s2  = \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.u2.s ;
assign \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.u1.a  = \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.a [15:0];
assign \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.u1.b  = \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.b [15:0];
assign \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.u1.cin  = 1'h0;
assign \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.facout_s1  = \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.u1.cout ;
assign \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.fas_s1  = \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.u1.s ;
assign \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.a  = \add_32ns_32s_32_2_1_U8.din0 ;
assign \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.b  = \add_32ns_32s_32_2_1_U8.din1 ;
assign \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.ce  = \add_32ns_32s_32_2_1_U8.ce ;
assign \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.clk  = \add_32ns_32s_32_2_1_U8.clk ;
assign \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.reset  = \add_32ns_32s_32_2_1_U8.reset ;
assign \add_32ns_32s_32_2_1_U8.dout  = \add_32ns_32s_32_2_1_U8.top_add_32ns_32s_32_2_1_Adder_7_U.s ;
assign \add_32ns_32s_32_2_1_U8.ce  = 1'h1;
assign \add_32ns_32s_32_2_1_U8.clk  = ap_clk;
assign \add_32ns_32s_32_2_1_U8.din0  = ret_V_13_reg_825;
assign \add_32ns_32s_32_2_1_U8.din1  = { op_15[15], op_15[15], op_15[15], op_15[15], op_15[15], op_15[15], op_15[15], op_15[15], op_15[15], op_15[15], op_15[15], op_15[15], op_15[15], op_15[15], op_15[15], op_15[15], op_15 };
assign grp_fu_495_p2 = \add_32ns_32s_32_2_1_U8.dout ;
assign \add_32ns_32s_32_2_1_U8.reset  = ap_rst;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.ain_s0  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.a ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.bin_s0  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.b ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.s  = { \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.fas_s2 , \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.sum_s1  };
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.a  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.ain_s1 ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.b  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.bin_s1 ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.cin  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.carry_s1 ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.facout_s2  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.cout ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.fas_s2  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.s ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.a  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.a [15:0];
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.b  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.b [15:0];
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.cin  = 1'h0;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.facout_s1  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.cout ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.fas_s1  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.s ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.a  = \add_32ns_32ns_32_2_1_U16.din0 ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.b  = \add_32ns_32ns_32_2_1_U16.din1 ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.ce  = \add_32ns_32ns_32_2_1_U16.ce ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.clk  = \add_32ns_32ns_32_2_1_U16.clk ;
assign \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.reset  = \add_32ns_32ns_32_2_1_U16.reset ;
assign \add_32ns_32ns_32_2_1_U16.dout  = \add_32ns_32ns_32_2_1_U16.top_add_32ns_32ns_32_2_1_Adder_11_U.s ;
assign \add_32ns_32ns_32_2_1_U16.ce  = 1'h1;
assign \add_32ns_32ns_32_2_1_U16.clk  = ap_clk;
assign \add_32ns_32ns_32_2_1_U16.din0  = ret_V_15_reg_938;
assign \add_32ns_32ns_32_2_1_U16.din1  = { 31'h00000000, lhs_V_4_reg_679 };
assign grp_fu_631_p2 = \add_32ns_32ns_32_2_1_U16.dout ;
assign \add_32ns_32ns_32_2_1_U16.reset  = ap_rst;
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.ain_s0  = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.a ;
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.bin_s0  = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.b ;
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.s  = { \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.fas_s2 , \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.sum_s1  };
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.a  = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.ain_s1 ;
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.b  = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.bin_s1 ;
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.cin  = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.carry_s1 ;
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.facout_s2  = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.cout ;
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.fas_s2  = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.u2.s ;
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.a  = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.a [15:0];
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.b  = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.b [15:0];
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.cin  = 1'h0;
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.facout_s1  = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.cout ;
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.fas_s1  = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.u1.s ;
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.a  = \add_32ns_32ns_32_2_1_U15.din0 ;
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.b  = \add_32ns_32ns_32_2_1_U15.din1 ;
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.ce  = \add_32ns_32ns_32_2_1_U15.ce ;
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.clk  = \add_32ns_32ns_32_2_1_U15.clk ;
assign \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.reset  = \add_32ns_32ns_32_2_1_U15.reset ;
assign \add_32ns_32ns_32_2_1_U15.dout  = \add_32ns_32ns_32_2_1_U15.top_add_32ns_32ns_32_2_1_Adder_11_U.s ;
assign \add_32ns_32ns_32_2_1_U15.ce  = 1'h1;
assign \add_32ns_32ns_32_2_1_U15.clk  = ap_clk;
assign \add_32ns_32ns_32_2_1_U15.din0  = ret_V_9_cast_reg_911;
assign \add_32ns_32ns_32_2_1_U15.din1  = 32'd1;
assign grp_fu_583_p2 = \add_32ns_32ns_32_2_1_U15.dout ;
assign \add_32ns_32ns_32_2_1_U15.reset  = ap_rst;
assign \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.ain_s0  = \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.a ;
assign \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.bin_s0  = \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.b ;
assign \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.s  = { \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.fas_s2 , \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.sum_s1  };
assign \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.u2.a  = \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.ain_s1 ;
assign \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.u2.b  = \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.bin_s1 ;
assign \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.u2.cin  = \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.carry_s1 ;
assign \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.facout_s2  = \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.u2.cout ;
assign \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.fas_s2  = \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.u2.s ;
assign \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.u1.a  = \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.a [7:0];
assign \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.u1.b  = \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.b [7:0];
assign \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.u1.cin  = 1'h0;
assign \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.facout_s1  = \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.u1.cout ;
assign \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.fas_s1  = \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.u1.s ;
assign \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.a  = \add_17s_17s_17_2_1_U17.din0 ;
assign \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.b  = \add_17s_17s_17_2_1_U17.din1 ;
assign \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.ce  = \add_17s_17s_17_2_1_U17.ce ;
assign \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.clk  = \add_17s_17s_17_2_1_U17.clk ;
assign \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.reset  = \add_17s_17s_17_2_1_U17.reset ;
assign \add_17s_17s_17_2_1_U17.dout  = \add_17s_17s_17_2_1_U17.top_add_17s_17s_17_2_1_Adder_12_U.s ;
assign \add_17s_17s_17_2_1_U17.ce  = 1'h1;
assign \add_17s_17s_17_2_1_U17.clk  = ap_clk;
assign \add_17s_17s_17_2_1_U17.din0  = { op_19[15], op_19 };
assign \add_17s_17s_17_2_1_U17.din1  = { r_reg_933[1], r_reg_933[1], r_reg_933[1], r_reg_933[1], r_reg_933[1], r_reg_933[1], r_reg_933[1], r_reg_933[1], r_reg_933[1], r_reg_933[1], r_reg_933[1], r_reg_933[1], r_reg_933[1], r_reg_933[1], r_reg_933[1], r_reg_933 };
assign grp_fu_643_p2 = \add_17s_17s_17_2_1_U17.dout ;
assign \add_17s_17s_17_2_1_U17.reset  = ap_rst;
assign \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.ain_s0  = \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.a ;
assign \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.bin_s0  = \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.b ;
assign \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.s  = { \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.fas_s2 , \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.sum_s1  };
assign \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.u2.a  = \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.ain_s1 ;
assign \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.u2.b  = \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.bin_s1 ;
assign \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.u2.cin  = \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.carry_s1 ;
assign \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.facout_s2  = \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.u2.cout ;
assign \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.fas_s2  = \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.u2.s ;
assign \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.u1.a  = \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.a [4:0];
assign \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.u1.b  = \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.b [4:0];
assign \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.u1.cin  = 1'h0;
assign \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.facout_s1  = \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.u1.cout ;
assign \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.fas_s1  = \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.u1.s ;
assign \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.a  = \add_10ns_10s_10_2_1_U1.din0 ;
assign \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.b  = \add_10ns_10s_10_2_1_U1.din1 ;
assign \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.ce  = \add_10ns_10s_10_2_1_U1.ce ;
assign \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.clk  = \add_10ns_10s_10_2_1_U1.clk ;
assign \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.reset  = \add_10ns_10s_10_2_1_U1.reset ;
assign \add_10ns_10s_10_2_1_U1.dout  = \add_10ns_10s_10_2_1_U1.top_add_10ns_10s_10_2_1_Adder_0_U.s ;
assign \add_10ns_10s_10_2_1_U1.ce  = 1'h1;
assign \add_10ns_10s_10_2_1_U1.clk  = ap_clk;
assign \add_10ns_10s_10_2_1_U1.din0  = { 2'h0, op_7 };
assign \add_10ns_10s_10_2_1_U1.din1  = { op_5[7], op_5[7], op_5 };
assign grp_fu_221_p2 = \add_10ns_10s_10_2_1_U1.dout ;
assign \add_10ns_10s_10_2_1_U1.reset  = ap_rst;
endmodule


// Product machine:
module top_A_times_top_B (ap_start, op_0, op_1, op_11, op_12, op_14, op_15, op_19, op_2, op_4, op_5, op_7, op_9, ap_clk, unsafe_signal);
input ap_start;
input [3:0] op_0;
input [7:0] op_1;
input [1:0] op_11;
input [1:0] op_12;
input [31:0] op_14;
input [15:0] op_15;
input [15:0] op_19;
input [15:0] op_2;
input [7:0] op_4;
input [7:0] op_5;
input [7:0] op_7;
input [1:0] op_9;
input ap_clk;
output unsafe_signal;
reg _setup;
initial _setup = 1'b0;
always @ (posedge ap_clk) _setup <= 1'b1;
reg ap_start_internal;
always @ (posedge ap_clk) if (!_setup) ap_start_internal <= ap_start;
reg [3:0] op_0_internal;
always @ (posedge ap_clk) if (!_setup) op_0_internal <= op_0;
reg [7:0] op_1_internal;
always @ (posedge ap_clk) if (!_setup) op_1_internal <= op_1;
reg [1:0] op_11_internal;
always @ (posedge ap_clk) if (!_setup) op_11_internal <= op_11;
reg [1:0] op_12_internal;
always @ (posedge ap_clk) if (!_setup) op_12_internal <= op_12;
reg [31:0] op_14_internal;
always @ (posedge ap_clk) if (!_setup) op_14_internal <= op_14;
reg [15:0] op_15_internal;
always @ (posedge ap_clk) if (!_setup) op_15_internal <= op_15;
reg [15:0] op_19_internal;
always @ (posedge ap_clk) if (!_setup) op_19_internal <= op_19;
reg [15:0] op_2_internal;
always @ (posedge ap_clk) if (!_setup) op_2_internal <= op_2;
reg [7:0] op_4_internal;
always @ (posedge ap_clk) if (!_setup) op_4_internal <= op_4;
reg [7:0] op_5_internal;
always @ (posedge ap_clk) if (!_setup) op_5_internal <= op_5;
reg [7:0] op_7_internal;
always @ (posedge ap_clk) if (!_setup) op_7_internal <= op_7;
reg [1:0] op_9_internal;
always @ (posedge ap_clk) if (!_setup) op_9_internal <= op_9;
wire ap_done_A;
wire ap_done_B;
wire ap_done_eq;
assign ap_done_eq = ap_done_A == ap_done_B;
wire ap_idle_A;
wire ap_idle_B;
wire ap_idle_eq;
assign ap_idle_eq = ap_idle_A == ap_idle_B;
wire ap_ready_A;
wire ap_ready_B;
wire ap_ready_eq;
assign ap_ready_eq = ap_ready_A == ap_ready_B;
wire [31:0] op_29_A;
wire [31:0] op_29_B;
wire op_29_eq;
assign op_29_eq = op_29_A == op_29_B;
wire op_29_ap_vld_A;
wire op_29_ap_vld_B;
wire clk_enable_A;
wire clk_enable_B;
assign clk_enable_A = _setup & (~op_29_ap_vld_A | op_29_ap_vld_B);
assign clk_enable_B = _setup;
wire divergent;
assign divergent = ~(ap_done_eq & ap_idle_eq & ap_ready_eq & op_29_eq);
assign unsafe_signal = op_29_ap_vld_A & op_29_ap_vld_B & divergent;
top_A instance_A (
    .ap_clk(ap_clk),
    .clk_enable(clk_enable_A),
    .ap_start(ap_start_internal),
    .op_0(op_0_internal),
    .op_1(op_1_internal),
    .op_11(op_11_internal),
    .op_12(op_12_internal),
    .op_14(op_14_internal),
    .op_15(op_15_internal),
    .op_19(op_19_internal),
    .op_2(op_2_internal),
    .op_4(op_4_internal),
    .op_5(op_5_internal),
    .op_7(op_7_internal),
    .op_9(op_9_internal),
    .ap_done(ap_done_A),
    .ap_idle(ap_idle_A),
    .ap_ready(ap_ready_A),
    .op_29(op_29_A),
    .op_29_ap_vld(op_29_ap_vld_A)
);
top_B instance_B (
    .ap_clk(ap_clk),
    .clk_enable(clk_enable_B),
    .ap_start(ap_start_internal),
    .op_0(op_0_internal),
    .op_1(op_1_internal),
    .op_11(op_11_internal),
    .op_12(op_12_internal),
    .op_14(op_14_internal),
    .op_15(op_15_internal),
    .op_19(op_19_internal),
    .op_2(op_2_internal),
    .op_4(op_4_internal),
    .op_5(op_5_internal),
    .op_7(op_7_internal),
    .op_9(op_9_internal),
    .ap_done(ap_done_B),
    .ap_idle(ap_idle_B),
    .ap_ready(ap_ready_B),
    .op_29(op_29_B),
    .op_29_ap_vld(op_29_ap_vld_B)
);
endmodule
