// Processed by function `construct_kairos` in `verilog_tricks.py`.
// Machine A:
// Processed by function `add_clk_enable_signal` in `verilog_tricks.py`.
// Processed by function `remove_reset_signal` in `verilog_tricks.py`.
module top_A (
  ap_clk,
  ap_start,
  ap_done,
  ap_idle,
  ap_ready,
  op_0,
  op_1,
  op_2,
  op_5,
  op_8,
  op_12,
  op_14,
  op_16,
  op_18,
  op_30,
  op_30_ap_vld,
clk_enable
);
input clk_enable;


input ap_clk;
wire ap_rst;
assign ap_rst = op_30_ap_vld;
input ap_start;
input [1:0] op_0;
input [3:0] op_1;
input [1:0] op_12;
input op_14;
input [3:0] op_16;
input [3:0] op_18;
input [7:0] op_2;
input [3:0] op_5;
input [3:0] op_8;
output ap_done;
output ap_idle;
output ap_ready;
output [31:0] op_30;
output op_30_ap_vld;


reg [5:0] add_ln69_2_reg_807;
reg [10:0] add_ln69_reg_802;
reg [11:0] ap_CS_fsm = 12'h001;
reg [15:0] \ashr_32s_16ns_32_2_1_U4.din1_cast_array[0] ;
reg [31:0] \ashr_32s_16ns_32_2_1_U4.dout_array[0] ;
reg icmp_ln1499_reg_756;
reg icmp_ln851_3_reg_913;
reg icmp_ln851_reg_734;
reg isNeg_reg_791;
reg lhs_V_2_reg_817;
reg [3:0] op_7_V_reg_771;
reg p_Result_8_reg_850;
reg [5:0] r_reg_891;
reg [2:0] ret_V_11_reg_828;
reg [11:0] ret_V_19_reg_722;
reg [9:0] ret_V_20_reg_766;
reg [2:0] ret_V_24_reg_843;
reg [10:0] ret_V_25_reg_835;
reg [10:0] ret_V_26_reg_855;
reg [10:0] ret_V_27_reg_896;
reg [34:0] ret_V_28_reg_901;
reg [31:0] ret_V_30_cast_reg_906;
reg [1:0] ret_V_3_reg_744;
reg [9:0] ret_V_8_reg_776;
reg [9:0] ret_V_reg_727;
reg [2:0] ret_reg_786;
reg [10:0] select_ln1192_reg_812;
reg [31:0] select_ln1368_reg_822;
reg [3:0] sh_V_1_reg_860;
reg [15:0] \shl_32s_16ns_32_2_1_U5.din1_cast_array[0] ;
reg [31:0] \shl_32s_16ns_32_2_1_U5.dout_array[0] ;
reg [31:0] shl_ln1299_reg_739;
reg [3:0] trunc_ln1348_1_reg_761;
reg [2:0] trunc_ln546_reg_881;
reg [5:0] trunc_ln769_reg_886;
reg [1:0] trunc_ln851_1_reg_751;
reg [1:0] trunc_ln851_2_reg_781;
reg [4:0] ush_reg_797;
wire [5:0] _000_;
wire [10:0] _001_;
wire [11:0] _002_;
wire _003_;
wire _004_;
wire _005_;
wire _006_;
wire _007_;
wire [3:0] _008_;
wire _009_;
wire [5:0] _010_;
wire [2:0] _011_;
wire [11:0] _012_;
wire [9:0] _013_;
wire [2:0] _014_;
wire [10:0] _015_;
wire [10:0] _016_;
wire [10:0] _017_;
wire [34:0] _018_;
wire [31:0] _019_;
wire [1:0] _020_;
wire [9:0] _021_;
wire [9:0] _022_;
wire [2:0] _023_;
wire [10:0] _024_;
wire [31:0] _025_;
wire [3:0] _026_;
wire [31:0] _027_;
wire [3:0] _028_;
wire [2:0] _029_;
wire [5:0] _030_;
wire [1:0] _031_;
wire [1:0] _032_;
wire [4:0] _033_;
wire [1:0] _034_;
wire _035_;
wire _036_;
wire _037_;
wire _038_;
wire _039_;
wire _040_;
wire _041_;
wire _042_;
wire _043_;
wire _044_;
wire _045_;
wire [15:0] _046_;
wire [31:0] _047_;
wire [15:0] _048_;
wire [31:0] _049_;
wire [31:0] _050_;
wire [15:0] _051_;
wire [31:0] _052_;
wire [15:0] _053_;
wire [31:0] _054_;
wire [31:0] _055_;
wire _056_;
wire _057_;
wire _058_;
wire _059_;
wire _060_;
wire _061_;
wire _062_;
wire _063_;
wire _064_;
wire _065_;
wire _066_;
wire _067_;
wire _068_;
wire _069_;
wire [31:0] add_ln691_1_fu_703_p2;
wire [10:0] add_ln691_fu_564_p2;
wire [2:0] add_ln69_1_fu_441_p2;
wire [5:0] add_ln69_2_fu_451_p2;
wire [10:0] add_ln69_fu_435_p2;
wire ap_CS_fsm_state1;
wire ap_CS_fsm_state10;
wire ap_CS_fsm_state11;
wire ap_CS_fsm_state12;
wire ap_CS_fsm_state2;
wire ap_CS_fsm_state3;
wire ap_CS_fsm_state4;
wire ap_CS_fsm_state5;
wire ap_CS_fsm_state6;
wire ap_CS_fsm_state7;
wire ap_CS_fsm_state8;
wire ap_CS_fsm_state9;
wire [11:0] ap_NS_fsm;
wire ap_clk;
wire ap_done;
wire ap_idle;
wire ap_ready;
wire ap_rst;
wire ap_start;
wire \ashr_32s_16ns_32_2_1_U4.ce ;
wire \ashr_32s_16ns_32_2_1_U4.clk ;
wire [31:0] \ashr_32s_16ns_32_2_1_U4.din0 ;
wire [31:0] \ashr_32s_16ns_32_2_1_U4.din1 ;
wire [15:0] \ashr_32s_16ns_32_2_1_U4.din1_cast ;
wire [15:0] \ashr_32s_16ns_32_2_1_U4.din1_mask ;
wire [31:0] \ashr_32s_16ns_32_2_1_U4.dout ;
wire \ashr_32s_16ns_32_2_1_U4.reset ;
wire [31:0] \ashr_32s_32s_32_1_1_U3.din0 ;
wire [31:0] \ashr_32s_32s_32_1_1_U3.din1 ;
wire [31:0] \ashr_32s_32s_32_1_1_U3.din1_cast ;
wire [31:0] \ashr_32s_32s_32_1_1_U3.dout ;
wire [31:0] ashr_ln1333_fu_484_p2;
wire [3:0] conv_i_i_i329_fu_474_p0;
wire [31:0] conv_i_i_i329_fu_474_p1;
wire [31:0] grp_fu_601_p1;
wire [31:0] grp_fu_601_p2;
wire [31:0] grp_fu_614_p1;
wire [31:0] grp_fu_614_p2;
wire icmp_ln1499_fu_243_p2;
wire icmp_ln851_1_fu_285_p2;
wire icmp_ln851_2_fu_378_p2;
wire icmp_ln851_3_fu_690_p2;
wire icmp_ln851_fu_209_p2;
wire [11:0] lhs_V_1_fu_318_p3;
wire [3:0] lhs_V_2_fu_465_p0;
wire lhs_V_2_fu_465_p2;
wire [1:0] op_0;
wire [3:0] op_1;
wire [1:0] op_12;
wire op_14;
wire [3:0] op_16;
wire [3:0] op_18;
wire [7:0] op_2;
wire [10:0] op_24_V_fu_510_p2;
wire [10:0] op_27_V_fu_641_p2;
wire [31:0] op_30;
wire op_30_ap_vld;
wire [3:0] op_5;
wire [3:0] op_7_V_fu_313_p2;
wire [3:0] op_8;
wire p_Result_1_fu_278_p3;
wire p_Result_3_fu_371_p3;
wire p_Result_4_fu_520_p3;
wire p_Result_6_fu_557_p3;
wire p_Result_7_fu_696_p3;
wire p_Result_s_fu_253_p3;
wire [5:0] r_fu_631_p3;
wire [2:0] ret_V_12_fu_530_p2;
wire [11:0] ret_V_19_fu_189_p2;
wire [9:0] ret_V_20_fu_271_p3;
wire [1:0] ret_V_21_fu_302_p3;
wire [11:0] ret_V_22_fu_326_p2;
wire [10:0] ret_V_23_fu_397_p3;
wire [2:0] ret_V_24_fu_542_p3;
wire [10:0] ret_V_25_fu_515_p2;
wire [10:0] ret_V_26_fu_575_p3;
wire [10:0] ret_V_27_fu_649_p2;
wire [34:0] ret_V_28_fu_670_p2;
wire [9:0] ret_V_2_fu_260_p2;
wire [1:0] ret_V_5_fu_290_p2;
wire [10:0] ret_V_9_fu_383_p2;
wire [2:0] ret_fu_354_p2;
wire [9:0] rhs_fu_177_p3;
wire [10:0] select_ln1192_fu_457_p3;
wire [31:0] select_ln1368_fu_490_p3;
wire [1:0] select_ln850_1_fu_295_p3;
wire [10:0] select_ln850_2_fu_389_p3;
wire [2:0] select_ln850_3_fu_535_p3;
wire [10:0] select_ln850_4_fu_569_p3;
wire [31:0] select_ln850_5_fu_708_p3;
wire [9:0] select_ln850_fu_265_p3;
wire [34:0] sext_ln1192_1_fu_666_p1;
wire [10:0] sext_ln1192_fu_646_p1;
wire [3:0] sext_ln1299_fu_219_p0;
wire [2:0] sext_ln1346_1_fu_350_p1;
wire [2:0] sext_ln1346_fu_346_p1;
wire [31:0] sext_ln1367_fu_471_p1;
wire [4:0] sext_ln1386_fu_408_p1;
wire [3:0] sext_ln14_fu_582_p1;
wire [10:0] sext_ln21_fu_405_p1;
wire [5:0] sext_ln546_1_fu_628_p1;
wire [15:0] sext_ln546_2_fu_607_p1;
wire [15:0] sext_ln546_fu_594_p1;
wire [5:0] sext_ln69_1_fu_447_p1;
wire [10:0] sext_ln69_2_fu_507_p1;
wire [10:0] sext_ln69_3_fu_637_p1;
wire [2:0] sext_ln69_fu_431_p1;
wire [3:0] sext_ln703_1_fu_655_p0;
wire [34:0] sext_ln703_1_fu_655_p1;
wire [3:0] sext_ln703_fu_173_p0;
wire [11:0] sext_ln703_fu_173_p1;
wire [31:0] sext_ln781_fu_591_p1;
wire [10:0] sext_ln831_fu_368_p1;
wire [3:0] sh_V_1_fu_585_p2;
wire \shl_32s_16ns_32_2_1_U5.ce ;
wire \shl_32s_16ns_32_2_1_U5.clk ;
wire [31:0] \shl_32s_16ns_32_2_1_U5.din0 ;
wire [31:0] \shl_32s_16ns_32_2_1_U5.din1 ;
wire [15:0] \shl_32s_16ns_32_2_1_U5.din1_cast ;
wire [15:0] \shl_32s_16ns_32_2_1_U5.din1_mask ;
wire [31:0] \shl_32s_16ns_32_2_1_U5.dout ;
wire \shl_32s_16ns_32_2_1_U5.reset ;
wire [31:0] \shl_32s_32s_32_1_1_U2.din0 ;
wire [31:0] \shl_32s_32s_32_1_1_U2.din1 ;
wire [31:0] \shl_32s_32s_32_1_1_U2.din1_cast ;
wire [31:0] \shl_32s_32s_32_1_1_U2.dout ;
wire [31:0] \shl_32s_8ns_32_1_1_U1.din0 ;
wire [31:0] \shl_32s_8ns_32_1_1_U1.din1 ;
wire [7:0] \shl_32s_8ns_32_1_1_U1.din1_cast ;
wire [31:0] \shl_32s_8ns_32_1_1_U1.dout ;
wire [31:0] shl_ln1299_1_fu_478_p2;
wire [31:0] shl_ln1299_fu_223_p0;
wire [31:0] shl_ln1299_fu_223_p1;
wire [31:0] shl_ln1299_fu_223_p2;
wire [4:0] sub_ln1367_fu_411_p2;
wire [12:0] tmp_fu_659_p3;
wire [3:0] trunc_ln1348_1_fu_249_p1;
wire [3:0] trunc_ln1348_fu_309_p1;
wire [2:0] trunc_ln546_fu_620_p1;
wire [5:0] trunc_ln769_fu_624_p1;
wire [1:0] trunc_ln851_1_fu_239_p1;
wire [1:0] trunc_ln851_2_fu_342_p1;
wire trunc_ln851_3_fu_527_p1;
wire [3:0] trunc_ln851_4_fu_686_p0;
wire [1:0] trunc_ln851_4_fu_686_p1;
wire [3:0] trunc_ln851_fu_205_p0;
wire [1:0] trunc_ln851_fu_205_p1;
wire [4:0] ush_fu_417_p3;
wire [11:0] zext_ln1192_fu_185_p1;
wire [2:0] zext_ln69_fu_428_p1;
wire [5:0] zext_ln769_fu_424_p1;


assign add_ln691_1_fu_703_p2 = ret_V_30_cast_reg_906 + 1'h1;
assign add_ln691_fu_564_p2 = ret_V_25_reg_835 + 1'h1;
assign add_ln69_1_fu_441_p2 = $signed(op_12) + $signed({ 1'h0, icmp_ln1499_reg_756 });
assign add_ln69_2_fu_451_p2 = $signed(add_ln69_1_fu_441_p2) + $signed({ 1'h0, op_8 });
assign add_ln69_fu_435_p2 = $signed(ret_V_23_fu_397_p3) + $signed(ret_reg_786);
assign op_24_V_fu_510_p2 = $signed(add_ln69_2_reg_807) + $signed(add_ln69_reg_802);
assign op_27_V_fu_641_p2 = $signed(ret_V_26_reg_855) + $signed(op_16);
assign ret_V_12_fu_530_p2 = ret_V_11_reg_828 + 1'h1;
assign ret_V_19_fu_189_p2 = $signed({ 1'h0, op_2, 2'h0 }) + $signed(op_1);
assign ret_V_25_fu_515_p2 = op_24_V_fu_510_p2 + select_ln1192_reg_812;
assign ret_V_27_fu_649_p2 = $signed(op_27_V_fu_641_p2) + $signed(r_reg_891);
assign { ret_V_28_fu_670_p2[34], ret_V_28_fu_670_p2[12:0] } = $signed({ ret_V_27_reg_896, 2'h0 }) + $signed(op_18);
assign ret_V_2_fu_260_p2 = ret_V_reg_727 + 1'h1;
assign ret_V_5_fu_290_p2 = ret_V_3_reg_744 + 1'h1;
assign ret_V_9_fu_383_p2 = $signed(ret_V_8_reg_776) + $signed(2'h1);
assign ret_fu_354_p2 = $signed(ret_V_21_fu_302_p3) + $signed(op_0);
assign _035_ = ap_CS_fsm[5] & p_Result_8_reg_850;
assign _036_ = ap_CS_fsm[7] & p_Result_8_reg_850;
assign _037_ = ap_CS_fsm[7] & _040_;
assign _038_ = ap_CS_fsm[0] & _041_;
assign _039_ = ap_CS_fsm[0] & ap_start;
assign op_7_V_fu_313_p2 = ret_V_20_fu_271_p3[3:0] & trunc_ln1348_1_reg_761;
assign ret_V_22_fu_326_p2[2] = ~ ret_V_20_fu_271_p3[0];
assign _040_ = ~ p_Result_8_reg_850;
assign _041_ = ~ ap_start;
assign _042_ = ! trunc_ln851_1_reg_751;
assign _043_ = ! trunc_ln851_2_reg_781;
assign _044_ = ! op_1[1:0];
assign _045_ = op_5 == 2'h2;
always @(posedge \ashr_32s_16ns_32_2_1_U4.clk )
\ashr_32s_16ns_32_2_1_U4.dout_array[0]  <= _047_;
always @(posedge \ashr_32s_16ns_32_2_1_U4.clk )
\ashr_32s_16ns_32_2_1_U4.din1_cast_array[0]  <= _046_;
assign _048_ = \ashr_32s_16ns_32_2_1_U4.ce  ? \ashr_32s_16ns_32_2_1_U4.din1 [15:0] : \ashr_32s_16ns_32_2_1_U4.din1_cast_array[0] ;
assign _046_ = \ashr_32s_16ns_32_2_1_U4.reset  ? 16'h0000 : _048_;
assign _049_ = \ashr_32s_16ns_32_2_1_U4.ce  ? _050_ : \ashr_32s_16ns_32_2_1_U4.dout_array[0] ;
assign _047_ = \ashr_32s_16ns_32_2_1_U4.reset  ? 32'd0 : _049_;
assign _050_ = $signed(\ashr_32s_16ns_32_2_1_U4.din0 ) >>> { \ashr_32s_16ns_32_2_1_U4.din1 [15:8], 8'h00 };
assign \ashr_32s_16ns_32_2_1_U4.dout  = $signed(\ashr_32s_16ns_32_2_1_U4.dout_array[0] ) >>> \ashr_32s_16ns_32_2_1_U4.din1_cast_array[0] [7:0];
assign \ashr_32s_32s_32_1_1_U3.dout  = $signed(\ashr_32s_32s_32_1_1_U3.din0 ) >>> \ashr_32s_32s_32_1_1_U3.din1 ;
always @(posedge \shl_32s_16ns_32_2_1_U5.clk )
\shl_32s_16ns_32_2_1_U5.dout_array[0]  <= _052_;
always @(posedge \shl_32s_16ns_32_2_1_U5.clk )
\shl_32s_16ns_32_2_1_U5.din1_cast_array[0]  <= _051_;
assign _053_ = \shl_32s_16ns_32_2_1_U5.ce  ? \shl_32s_16ns_32_2_1_U5.din1 [15:0] : \shl_32s_16ns_32_2_1_U5.din1_cast_array[0] ;
assign _051_ = \shl_32s_16ns_32_2_1_U5.reset  ? 16'h0000 : _053_;
assign _054_ = \shl_32s_16ns_32_2_1_U5.ce  ? _055_ : \shl_32s_16ns_32_2_1_U5.dout_array[0] ;
assign _052_ = \shl_32s_16ns_32_2_1_U5.reset  ? 32'd0 : _054_;
assign _055_ = \shl_32s_16ns_32_2_1_U5.din0  << { \shl_32s_16ns_32_2_1_U5.din1 [15:8], 8'h00 };
assign \shl_32s_16ns_32_2_1_U5.dout  = \shl_32s_16ns_32_2_1_U5.dout_array[0]  << \shl_32s_16ns_32_2_1_U5.din1_cast_array[0] [7:0];
assign \shl_32s_32s_32_1_1_U2.dout  = \shl_32s_32s_32_1_1_U2.din0  << \shl_32s_32s_32_1_1_U2.din1 ;
assign \shl_32s_8ns_32_1_1_U1.dout  = \shl_32s_8ns_32_1_1_U1.din0  << \shl_32s_8ns_32_1_1_U1.din1 [7:0];
assign _056_ = op_2 != 1'h1;
assign _057_ = | op_18[1:0];
always @(posedge ap_clk)
trunc_ln769_reg_886 <= _030_;
always @(posedge ap_clk)
trunc_ln546_reg_881 <= _029_;
always @(posedge ap_clk)
sh_V_1_reg_860 <= _026_;
always @(posedge ap_clk)
ret_V_27_reg_896 <= _017_;
always @(posedge ap_clk)
r_reg_891 <= _010_;
always @(posedge ap_clk)
ret_V_24_reg_843 <= _014_;
always @(posedge ap_clk)
p_Result_8_reg_850 <= _009_;
always @(posedge ap_clk)
ret_V_26_reg_855 <= _016_;
always @(posedge ap_clk)
lhs_V_2_reg_817 <= _007_;
always @(posedge ap_clk)
select_ln1368_reg_822 <= _025_;
always @(posedge ap_clk)
ret_V_11_reg_828 <= _011_;
always @(posedge ap_clk)
ret_V_25_reg_835 <= _015_;
always @(posedge ap_clk)
ret_V_20_reg_766 <= _013_;
always @(posedge ap_clk)
op_7_V_reg_771 <= _008_;
always @(posedge ap_clk)
ret_V_8_reg_776 <= _021_;
always @(posedge ap_clk)
trunc_ln851_2_reg_781 <= _032_;
always @(posedge ap_clk)
ret_reg_786 <= _023_;
always @(posedge ap_clk)
isNeg_reg_791 <= _006_;
always @(posedge ap_clk)
ret_V_28_reg_901 <= _018_;
always @(posedge ap_clk)
ret_V_30_cast_reg_906 <= _019_;
always @(posedge ap_clk)
icmp_ln851_3_reg_913 <= _004_;
always @(posedge ap_clk)
ret_V_19_reg_722 <= _012_;
always @(posedge ap_clk)
ret_V_reg_727 <= _022_;
always @(posedge ap_clk)
icmp_ln851_reg_734 <= _005_;
always @(posedge ap_clk)
shl_ln1299_reg_739 <= _027_;
always @(posedge ap_clk)
ret_V_3_reg_744 <= _020_;
always @(posedge ap_clk)
trunc_ln851_1_reg_751 <= _031_;
always @(posedge ap_clk)
icmp_ln1499_reg_756 <= _003_;
always @(posedge ap_clk)
trunc_ln1348_1_reg_761 <= _028_;
always @(posedge ap_clk)
ush_reg_797 <= _033_;
always @(posedge ap_clk)
add_ln69_reg_802 <= _001_;
always @(posedge ap_clk)
add_ln69_2_reg_807 <= _000_;
always @(posedge ap_clk)
select_ln1192_reg_812 <= _024_;
always @(posedge ap_clk)
ap_CS_fsm <= _002_;
assign _034_ = _039_ ? 2'h2 : 2'h1;
assign _058_ = ap_CS_fsm == 1'h1;
function [11:0] _156_;
input [11:0] a;
input [143:0] b;
input [11:0] s;
case (s)
12'b000000000001:
_156_ = b[11:0];
12'b000000000010:
_156_ = b[23:12];
12'b000000000100:
_156_ = b[35:24];
12'b000000001000:
_156_ = b[47:36];
12'b000000010000:
_156_ = b[59:48];
12'b000000100000:
_156_ = b[71:60];
12'b000001000000:
_156_ = b[83:72];
12'b000010000000:
_156_ = b[95:84];
12'b000100000000:
_156_ = b[107:96];
12'b001000000000:
_156_ = b[119:108];
12'b010000000000:
_156_ = b[131:120];
12'b100000000000:
_156_ = b[143:132];
12'b000000000000:
_156_ = a;
default:
_156_ = 12'bx;
endcase
endfunction
assign ap_NS_fsm = _156_(12'hxxx, { 10'h000, _034_, 132'h004008010020040080100200400800001 }, { _058_, _069_, _068_, _067_, _066_, _065_, _064_, _063_, _062_, _061_, _060_, _059_ });
assign _059_ = ap_CS_fsm == 12'h800;
assign _060_ = ap_CS_fsm == 11'h400;
assign _061_ = ap_CS_fsm == 10'h200;
assign _062_ = ap_CS_fsm == 9'h100;
assign _063_ = ap_CS_fsm == 8'h80;
assign _064_ = ap_CS_fsm == 7'h40;
assign _065_ = ap_CS_fsm == 6'h20;
assign _066_ = ap_CS_fsm == 5'h10;
assign _067_ = ap_CS_fsm == 4'h8;
assign _068_ = ap_CS_fsm == 3'h4;
assign _069_ = ap_CS_fsm == 2'h2;
assign op_30_ap_vld = ap_CS_fsm[11] ? 1'h1 : 1'h0;
assign ap_idle = _038_ ? 1'h1 : 1'h0;
assign _030_ = _037_ ? grp_fu_614_p2[5:0] : trunc_ln769_reg_886;
assign _029_ = _036_ ? grp_fu_601_p2[2:0] : trunc_ln546_reg_881;
assign _026_ = _035_ ? sh_V_1_fu_585_p2 : sh_V_1_reg_860;
assign _017_ = ap_CS_fsm[9] ? ret_V_27_fu_649_p2 : ret_V_27_reg_896;
assign _010_ = ap_CS_fsm[8] ? r_fu_631_p3 : r_reg_891;
assign _016_ = ap_CS_fsm[4] ? ret_V_26_fu_575_p3 : ret_V_26_reg_855;
assign _009_ = ap_CS_fsm[4] ? ret_V_24_fu_542_p3[2] : p_Result_8_reg_850;
assign _014_ = ap_CS_fsm[4] ? ret_V_24_fu_542_p3 : ret_V_24_reg_843;
assign _015_ = ap_CS_fsm[3] ? ret_V_25_fu_515_p2 : ret_V_25_reg_835;
assign _011_ = ap_CS_fsm[3] ? select_ln1368_fu_490_p3[3:1] : ret_V_11_reg_828;
assign _025_ = ap_CS_fsm[3] ? select_ln1368_fu_490_p3 : select_ln1368_reg_822;
assign _007_ = ap_CS_fsm[3] ? lhs_V_2_fu_465_p2 : lhs_V_2_reg_817;
assign _006_ = ap_CS_fsm[1] ? op_7_V_fu_313_p2[3] : isNeg_reg_791;
assign _023_ = ap_CS_fsm[1] ? ret_fu_354_p2 : ret_reg_786;
assign _032_ = ap_CS_fsm[1] ? 2'h0 : trunc_ln851_2_reg_781;
assign _021_ = ap_CS_fsm[1] ? { ret_V_20_fu_271_p3[9:1], ret_V_22_fu_326_p2[2] } : ret_V_8_reg_776;
assign _008_ = ap_CS_fsm[1] ? op_7_V_fu_313_p2 : op_7_V_reg_771;
assign _013_ = ap_CS_fsm[1] ? ret_V_20_fu_271_p3 : ret_V_20_reg_766;
assign _004_ = ap_CS_fsm[10] ? icmp_ln851_3_fu_690_p2 : icmp_ln851_3_reg_913;
assign _019_ = ap_CS_fsm[10] ? { ret_V_28_fu_670_p2[34], ret_V_28_fu_670_p2[34], ret_V_28_fu_670_p2[34], ret_V_28_fu_670_p2[34], ret_V_28_fu_670_p2[34], ret_V_28_fu_670_p2[34], ret_V_28_fu_670_p2[34], ret_V_28_fu_670_p2[34], ret_V_28_fu_670_p2[34], ret_V_28_fu_670_p2[34], ret_V_28_fu_670_p2[34], ret_V_28_fu_670_p2[34], ret_V_28_fu_670_p2[34], ret_V_28_fu_670_p2[34], ret_V_28_fu_670_p2[34], ret_V_28_fu_670_p2[34], ret_V_28_fu_670_p2[34], ret_V_28_fu_670_p2[34], ret_V_28_fu_670_p2[34], ret_V_28_fu_670_p2[34], ret_V_28_fu_670_p2[34], ret_V_28_fu_670_p2[12:2] } : ret_V_30_cast_reg_906;
assign _018_ = ap_CS_fsm[10] ? { ret_V_28_fu_670_p2[34], ret_V_28_fu_670_p2[34], ret_V_28_fu_670_p2[34], ret_V_28_fu_670_p2[34], ret_V_28_fu_670_p2[34], ret_V_28_fu_670_p2[34], ret_V_28_fu_670_p2[34], ret_V_28_fu_670_p2[34], ret_V_28_fu_670_p2[34], ret_V_28_fu_670_p2[34], ret_V_28_fu_670_p2[34], ret_V_28_fu_670_p2[34], ret_V_28_fu_670_p2[34], ret_V_28_fu_670_p2[34], ret_V_28_fu_670_p2[34], ret_V_28_fu_670_p2[34], ret_V_28_fu_670_p2[34], ret_V_28_fu_670_p2[34], ret_V_28_fu_670_p2[34], ret_V_28_fu_670_p2[34], ret_V_28_fu_670_p2[34], ret_V_28_fu_670_p2[34], ret_V_28_fu_670_p2[12:0] } : ret_V_28_reg_901;
assign _028_ = ap_CS_fsm[0] ? op_2[3:0] : trunc_ln1348_1_reg_761;
assign _003_ = ap_CS_fsm[0] ? icmp_ln1499_fu_243_p2 : icmp_ln1499_reg_756;
assign _031_ = ap_CS_fsm[0] ? shl_ln1299_fu_223_p2[1:0] : trunc_ln851_1_reg_751;
assign _020_ = ap_CS_fsm[0] ? shl_ln1299_fu_223_p2[3:2] : ret_V_3_reg_744;
assign _027_ = ap_CS_fsm[0] ? shl_ln1299_fu_223_p2 : shl_ln1299_reg_739;
assign _005_ = ap_CS_fsm[0] ? icmp_ln851_fu_209_p2 : icmp_ln851_reg_734;
assign _022_ = ap_CS_fsm[0] ? ret_V_19_fu_189_p2[11:2] : ret_V_reg_727;
assign _012_ = ap_CS_fsm[0] ? ret_V_19_fu_189_p2 : ret_V_19_reg_722;
assign _024_ = ap_CS_fsm[2] ? select_ln1192_fu_457_p3 : select_ln1192_reg_812;
assign _000_ = ap_CS_fsm[2] ? add_ln69_2_fu_451_p2 : add_ln69_2_reg_807;
assign _001_ = ap_CS_fsm[2] ? add_ln69_fu_435_p2 : add_ln69_reg_802;
assign _033_ = ap_CS_fsm[2] ? ush_fu_417_p3 : ush_reg_797;
assign _002_ = ap_rst ? 12'h001 : ap_NS_fsm;
assign sh_V_1_fu_585_p2 = $signed(1'h0) - $signed(ret_V_24_reg_843);
assign sub_ln1367_fu_411_p2 = $signed(1'h0) - $signed(op_7_V_reg_771);
assign icmp_ln1499_fu_243_p2 = _056_ ? 1'h1 : 1'h0;
assign icmp_ln851_1_fu_285_p2 = _042_ ? 1'h1 : 1'h0;
assign icmp_ln851_2_fu_378_p2 = _043_ ? 1'h1 : 1'h0;
assign icmp_ln851_3_fu_690_p2 = _057_ ? 1'h1 : 1'h0;
assign icmp_ln851_fu_209_p2 = _044_ ? 1'h1 : 1'h0;
assign lhs_V_2_fu_465_p2 = _045_ ? 1'h1 : 1'h0;
assign op_30 = ret_V_28_reg_901[34] ? select_ln850_5_fu_708_p3 : ret_V_30_cast_reg_906;
assign r_fu_631_p3 = p_Result_8_reg_850 ? { trunc_ln546_reg_881[2], trunc_ln546_reg_881[2], trunc_ln546_reg_881[2], trunc_ln546_reg_881 } : trunc_ln769_reg_886;
assign ret_V_20_fu_271_p3 = ret_V_19_reg_722[11] ? select_ln850_fu_265_p3 : ret_V_reg_727;
assign ret_V_21_fu_302_p3 = shl_ln1299_reg_739[3] ? select_ln850_1_fu_295_p3 : ret_V_3_reg_744;
assign ret_V_23_fu_397_p3 = ret_V_20_reg_766[9] ? select_ln850_2_fu_389_p3 : { ret_V_8_reg_776[9], ret_V_8_reg_776 };
assign ret_V_24_fu_542_p3 = select_ln1368_reg_822[3] ? select_ln850_3_fu_535_p3 : ret_V_11_reg_828;
assign ret_V_26_fu_575_p3 = ret_V_25_reg_835[10] ? select_ln850_4_fu_569_p3 : { 1'h0, ret_V_25_reg_835[9:0] };
assign select_ln1192_fu_457_p3 = op_14 ? 11'h7ff : 11'h000;
assign select_ln1368_fu_490_p3 = isNeg_reg_791 ? shl_ln1299_1_fu_478_p2 : ashr_ln1333_fu_484_p2;
assign select_ln850_1_fu_295_p3 = icmp_ln851_1_fu_285_p2 ? ret_V_3_reg_744 : ret_V_5_fu_290_p2;
assign select_ln850_2_fu_389_p3 = icmp_ln851_2_fu_378_p2 ? { ret_V_8_reg_776[9], ret_V_8_reg_776 } : ret_V_9_fu_383_p2;
assign select_ln850_3_fu_535_p3 = select_ln1368_reg_822[0] ? ret_V_12_fu_530_p2 : ret_V_11_reg_828;
assign select_ln850_4_fu_569_p3 = lhs_V_2_reg_817 ? add_ln691_fu_564_p2 : { 1'h1, ret_V_25_reg_835[9:0] };
assign select_ln850_5_fu_708_p3 = icmp_ln851_3_reg_913 ? add_ln691_1_fu_703_p2 : ret_V_30_cast_reg_906;
assign select_ln850_fu_265_p3 = icmp_ln851_reg_734 ? ret_V_reg_727 : ret_V_2_fu_260_p2;
assign ush_fu_417_p3 = isNeg_reg_791 ? sub_ln1367_fu_411_p2 : { op_7_V_reg_771[3], op_7_V_reg_771 };
assign ap_CS_fsm_state1 = ap_CS_fsm[0];
assign ap_CS_fsm_state10 = ap_CS_fsm[9];
assign ap_CS_fsm_state11 = ap_CS_fsm[10];
assign ap_CS_fsm_state12 = ap_CS_fsm[11];
assign ap_CS_fsm_state2 = ap_CS_fsm[1];
assign ap_CS_fsm_state3 = ap_CS_fsm[2];
assign ap_CS_fsm_state4 = ap_CS_fsm[3];
assign ap_CS_fsm_state5 = ap_CS_fsm[4];
assign ap_CS_fsm_state6 = ap_CS_fsm[5];
assign ap_CS_fsm_state7 = ap_CS_fsm[6];
assign ap_CS_fsm_state8 = ap_CS_fsm[7];
assign ap_CS_fsm_state9 = ap_CS_fsm[8];
assign ap_done = op_30_ap_vld;
assign ap_ready = op_30_ap_vld;
assign conv_i_i_i329_fu_474_p0 = op_5;
assign conv_i_i_i329_fu_474_p1 = { op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5 };
assign grp_fu_601_p1 = { 16'h0000, sh_V_1_reg_860[3], sh_V_1_reg_860[3], sh_V_1_reg_860[3], sh_V_1_reg_860[3], sh_V_1_reg_860[3], sh_V_1_reg_860[3], sh_V_1_reg_860[3], sh_V_1_reg_860[3], sh_V_1_reg_860[3], sh_V_1_reg_860[3], sh_V_1_reg_860[3], sh_V_1_reg_860[3], sh_V_1_reg_860 };
assign grp_fu_614_p1 = { 16'h0000, ret_V_24_reg_843[2], ret_V_24_reg_843[2], ret_V_24_reg_843[2], ret_V_24_reg_843[2], ret_V_24_reg_843[2], ret_V_24_reg_843[2], ret_V_24_reg_843[2], ret_V_24_reg_843[2], ret_V_24_reg_843[2], ret_V_24_reg_843[2], ret_V_24_reg_843[2], ret_V_24_reg_843[2], ret_V_24_reg_843[2], ret_V_24_reg_843 };
assign lhs_V_1_fu_318_p3 = { ret_V_20_fu_271_p3, 2'h0 };
assign lhs_V_2_fu_465_p0 = op_5;
assign p_Result_1_fu_278_p3 = shl_ln1299_reg_739[3];
assign p_Result_3_fu_371_p3 = ret_V_20_reg_766[9];
assign p_Result_4_fu_520_p3 = select_ln1368_reg_822[3];
assign p_Result_6_fu_557_p3 = ret_V_25_reg_835[10];
assign p_Result_7_fu_696_p3 = ret_V_28_reg_901[34];
assign p_Result_s_fu_253_p3 = ret_V_19_reg_722[11];
assign ret_V_22_fu_326_p2[1:0] = 2'h0;
assign ret_V_22_fu_326_p2[11:3] = ret_V_20_fu_271_p3[9:1];
assign ret_V_28_fu_670_p2[33:13] = { ret_V_28_fu_670_p2[34], ret_V_28_fu_670_p2[34], ret_V_28_fu_670_p2[34], ret_V_28_fu_670_p2[34], ret_V_28_fu_670_p2[34], ret_V_28_fu_670_p2[34], ret_V_28_fu_670_p2[34], ret_V_28_fu_670_p2[34], ret_V_28_fu_670_p2[34], ret_V_28_fu_670_p2[34], ret_V_28_fu_670_p2[34], ret_V_28_fu_670_p2[34], ret_V_28_fu_670_p2[34], ret_V_28_fu_670_p2[34], ret_V_28_fu_670_p2[34], ret_V_28_fu_670_p2[34], ret_V_28_fu_670_p2[34], ret_V_28_fu_670_p2[34], ret_V_28_fu_670_p2[34], ret_V_28_fu_670_p2[34], ret_V_28_fu_670_p2[34] };
assign rhs_fu_177_p3 = { op_2, 2'h0 };
assign sext_ln1192_1_fu_666_p1 = { ret_V_27_reg_896[10], ret_V_27_reg_896[10], ret_V_27_reg_896[10], ret_V_27_reg_896[10], ret_V_27_reg_896[10], ret_V_27_reg_896[10], ret_V_27_reg_896[10], ret_V_27_reg_896[10], ret_V_27_reg_896[10], ret_V_27_reg_896[10], ret_V_27_reg_896[10], ret_V_27_reg_896[10], ret_V_27_reg_896[10], ret_V_27_reg_896[10], ret_V_27_reg_896[10], ret_V_27_reg_896[10], ret_V_27_reg_896[10], ret_V_27_reg_896[10], ret_V_27_reg_896[10], ret_V_27_reg_896[10], ret_V_27_reg_896[10], ret_V_27_reg_896[10], ret_V_27_reg_896, 2'h0 };
assign sext_ln1192_fu_646_p1 = { r_reg_891[5], r_reg_891[5], r_reg_891[5], r_reg_891[5], r_reg_891[5], r_reg_891 };
assign sext_ln1299_fu_219_p0 = op_1;
assign sext_ln1346_1_fu_350_p1 = { ret_V_21_fu_302_p3[1], ret_V_21_fu_302_p3 };
assign sext_ln1346_fu_346_p1 = { op_0[1], op_0 };
assign sext_ln1367_fu_471_p1 = { ush_reg_797[4], ush_reg_797[4], ush_reg_797[4], ush_reg_797[4], ush_reg_797[4], ush_reg_797[4], ush_reg_797[4], ush_reg_797[4], ush_reg_797[4], ush_reg_797[4], ush_reg_797[4], ush_reg_797[4], ush_reg_797[4], ush_reg_797[4], ush_reg_797[4], ush_reg_797[4], ush_reg_797[4], ush_reg_797[4], ush_reg_797[4], ush_reg_797[4], ush_reg_797[4], ush_reg_797[4], ush_reg_797[4], ush_reg_797[4], ush_reg_797[4], ush_reg_797[4], ush_reg_797[4], ush_reg_797 };
assign sext_ln1386_fu_408_p1 = { op_7_V_reg_771[3], op_7_V_reg_771 };
assign sext_ln14_fu_582_p1 = { ret_V_24_reg_843[2], ret_V_24_reg_843 };
assign sext_ln21_fu_405_p1 = { ret_reg_786[2], ret_reg_786[2], ret_reg_786[2], ret_reg_786[2], ret_reg_786[2], ret_reg_786[2], ret_reg_786[2], ret_reg_786[2], ret_reg_786 };
assign sext_ln546_1_fu_628_p1 = { trunc_ln546_reg_881[2], trunc_ln546_reg_881[2], trunc_ln546_reg_881[2], trunc_ln546_reg_881 };
assign sext_ln546_2_fu_607_p1 = { ret_V_24_reg_843[2], ret_V_24_reg_843[2], ret_V_24_reg_843[2], ret_V_24_reg_843[2], ret_V_24_reg_843[2], ret_V_24_reg_843[2], ret_V_24_reg_843[2], ret_V_24_reg_843[2], ret_V_24_reg_843[2], ret_V_24_reg_843[2], ret_V_24_reg_843[2], ret_V_24_reg_843[2], ret_V_24_reg_843[2], ret_V_24_reg_843 };
assign sext_ln546_fu_594_p1 = { sh_V_1_reg_860[3], sh_V_1_reg_860[3], sh_V_1_reg_860[3], sh_V_1_reg_860[3], sh_V_1_reg_860[3], sh_V_1_reg_860[3], sh_V_1_reg_860[3], sh_V_1_reg_860[3], sh_V_1_reg_860[3], sh_V_1_reg_860[3], sh_V_1_reg_860[3], sh_V_1_reg_860[3], sh_V_1_reg_860 };
assign sext_ln69_1_fu_447_p1 = { add_ln69_1_fu_441_p2[2], add_ln69_1_fu_441_p2[2], add_ln69_1_fu_441_p2[2], add_ln69_1_fu_441_p2 };
assign sext_ln69_2_fu_507_p1 = { add_ln69_2_reg_807[5], add_ln69_2_reg_807[5], add_ln69_2_reg_807[5], add_ln69_2_reg_807[5], add_ln69_2_reg_807[5], add_ln69_2_reg_807 };
assign sext_ln69_3_fu_637_p1 = { op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16 };
assign sext_ln69_fu_431_p1 = { op_12[1], op_12 };
assign sext_ln703_1_fu_655_p0 = op_18;
assign sext_ln703_1_fu_655_p1 = { op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18 };
assign sext_ln703_fu_173_p0 = op_1;
assign sext_ln703_fu_173_p1 = { op_1[3], op_1[3], op_1[3], op_1[3], op_1[3], op_1[3], op_1[3], op_1[3], op_1 };
assign sext_ln781_fu_591_p1 = { ret_V_24_reg_843[2], ret_V_24_reg_843[2], ret_V_24_reg_843[2], ret_V_24_reg_843[2], ret_V_24_reg_843[2], ret_V_24_reg_843[2], ret_V_24_reg_843[2], ret_V_24_reg_843[2], ret_V_24_reg_843[2], ret_V_24_reg_843[2], ret_V_24_reg_843[2], ret_V_24_reg_843[2], ret_V_24_reg_843[2], ret_V_24_reg_843[2], ret_V_24_reg_843[2], ret_V_24_reg_843[2], ret_V_24_reg_843[2], ret_V_24_reg_843[2], ret_V_24_reg_843[2], ret_V_24_reg_843[2], ret_V_24_reg_843[2], ret_V_24_reg_843[2], ret_V_24_reg_843[2], ret_V_24_reg_843[2], ret_V_24_reg_843[2], ret_V_24_reg_843[2], ret_V_24_reg_843[2], ret_V_24_reg_843[2], ret_V_24_reg_843[2], ret_V_24_reg_843 };
assign sext_ln831_fu_368_p1 = { ret_V_8_reg_776[9], ret_V_8_reg_776 };
assign shl_ln1299_fu_223_p0 = { op_1[3], op_1[3], op_1[3], op_1[3], op_1[3], op_1[3], op_1[3], op_1[3], op_1[3], op_1[3], op_1[3], op_1[3], op_1[3], op_1[3], op_1[3], op_1[3], op_1[3], op_1[3], op_1[3], op_1[3], op_1[3], op_1[3], op_1[3], op_1[3], op_1[3], op_1[3], op_1[3], op_1[3], op_1 };
assign shl_ln1299_fu_223_p1 = { 24'h000000, op_2 };
assign tmp_fu_659_p3 = { ret_V_27_reg_896, 2'h0 };
assign trunc_ln1348_1_fu_249_p1 = op_2[3:0];
assign trunc_ln1348_fu_309_p1 = ret_V_20_fu_271_p3[3:0];
assign trunc_ln546_fu_620_p1 = grp_fu_601_p2[2:0];
assign trunc_ln769_fu_624_p1 = grp_fu_614_p2[5:0];
assign trunc_ln851_1_fu_239_p1 = shl_ln1299_fu_223_p2[1:0];
assign trunc_ln851_2_fu_342_p1 = 2'h0;
assign trunc_ln851_3_fu_527_p1 = select_ln1368_reg_822[0];
assign trunc_ln851_4_fu_686_p0 = op_18;
assign trunc_ln851_4_fu_686_p1 = op_18[1:0];
assign trunc_ln851_fu_205_p0 = op_1;
assign trunc_ln851_fu_205_p1 = op_1[1:0];
assign zext_ln1192_fu_185_p1 = { 2'h0, op_2, 2'h0 };
assign zext_ln69_fu_428_p1 = { 2'h0, icmp_ln1499_reg_756 };
assign zext_ln769_fu_424_p1 = { 2'h0, op_8 };
assign \shl_32s_8ns_32_1_1_U1.din1_cast  = \shl_32s_8ns_32_1_1_U1.din1 [7:0];
assign \shl_32s_8ns_32_1_1_U1.din0  = { op_1[3], op_1[3], op_1[3], op_1[3], op_1[3], op_1[3], op_1[3], op_1[3], op_1[3], op_1[3], op_1[3], op_1[3], op_1[3], op_1[3], op_1[3], op_1[3], op_1[3], op_1[3], op_1[3], op_1[3], op_1[3], op_1[3], op_1[3], op_1[3], op_1[3], op_1[3], op_1[3], op_1[3], op_1 };
assign \shl_32s_8ns_32_1_1_U1.din1  = { 24'h000000, op_2 };
assign shl_ln1299_fu_223_p2 = \shl_32s_8ns_32_1_1_U1.dout ;
assign \shl_32s_32s_32_1_1_U2.din1_cast  = \shl_32s_32s_32_1_1_U2.din1 ;
assign \shl_32s_32s_32_1_1_U2.din0  = { op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5 };
assign \shl_32s_32s_32_1_1_U2.din1  = { ush_reg_797[4], ush_reg_797[4], ush_reg_797[4], ush_reg_797[4], ush_reg_797[4], ush_reg_797[4], ush_reg_797[4], ush_reg_797[4], ush_reg_797[4], ush_reg_797[4], ush_reg_797[4], ush_reg_797[4], ush_reg_797[4], ush_reg_797[4], ush_reg_797[4], ush_reg_797[4], ush_reg_797[4], ush_reg_797[4], ush_reg_797[4], ush_reg_797[4], ush_reg_797[4], ush_reg_797[4], ush_reg_797[4], ush_reg_797[4], ush_reg_797[4], ush_reg_797[4], ush_reg_797[4], ush_reg_797 };
assign shl_ln1299_1_fu_478_p2 = \shl_32s_32s_32_1_1_U2.dout ;
assign \shl_32s_16ns_32_2_1_U5.din1_cast  = \shl_32s_16ns_32_2_1_U5.din1 [15:0];
assign \shl_32s_16ns_32_2_1_U5.din1_mask  = 16'h00ff;
assign \shl_32s_16ns_32_2_1_U5.ce  = 1'h1;
assign \shl_32s_16ns_32_2_1_U5.clk  = ap_clk;
assign \shl_32s_16ns_32_2_1_U5.din0  = { ret_V_24_reg_843[2], ret_V_24_reg_843[2], ret_V_24_reg_843[2], ret_V_24_reg_843[2], ret_V_24_reg_843[2], ret_V_24_reg_843[2], ret_V_24_reg_843[2], ret_V_24_reg_843[2], ret_V_24_reg_843[2], ret_V_24_reg_843[2], ret_V_24_reg_843[2], ret_V_24_reg_843[2], ret_V_24_reg_843[2], ret_V_24_reg_843[2], ret_V_24_reg_843[2], ret_V_24_reg_843[2], ret_V_24_reg_843[2], ret_V_24_reg_843[2], ret_V_24_reg_843[2], ret_V_24_reg_843[2], ret_V_24_reg_843[2], ret_V_24_reg_843[2], ret_V_24_reg_843[2], ret_V_24_reg_843[2], ret_V_24_reg_843[2], ret_V_24_reg_843[2], ret_V_24_reg_843[2], ret_V_24_reg_843[2], ret_V_24_reg_843[2], ret_V_24_reg_843 };
assign \shl_32s_16ns_32_2_1_U5.din1  = { 16'h0000, ret_V_24_reg_843[2], ret_V_24_reg_843[2], ret_V_24_reg_843[2], ret_V_24_reg_843[2], ret_V_24_reg_843[2], ret_V_24_reg_843[2], ret_V_24_reg_843[2], ret_V_24_reg_843[2], ret_V_24_reg_843[2], ret_V_24_reg_843[2], ret_V_24_reg_843[2], ret_V_24_reg_843[2], ret_V_24_reg_843[2], ret_V_24_reg_843 };
assign grp_fu_614_p2 = \shl_32s_16ns_32_2_1_U5.dout ;
assign \shl_32s_16ns_32_2_1_U5.reset  = ap_rst;
assign \ashr_32s_32s_32_1_1_U3.din1_cast  = \ashr_32s_32s_32_1_1_U3.din1 ;
assign \ashr_32s_32s_32_1_1_U3.din0  = { op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5 };
assign \ashr_32s_32s_32_1_1_U3.din1  = { ush_reg_797[4], ush_reg_797[4], ush_reg_797[4], ush_reg_797[4], ush_reg_797[4], ush_reg_797[4], ush_reg_797[4], ush_reg_797[4], ush_reg_797[4], ush_reg_797[4], ush_reg_797[4], ush_reg_797[4], ush_reg_797[4], ush_reg_797[4], ush_reg_797[4], ush_reg_797[4], ush_reg_797[4], ush_reg_797[4], ush_reg_797[4], ush_reg_797[4], ush_reg_797[4], ush_reg_797[4], ush_reg_797[4], ush_reg_797[4], ush_reg_797[4], ush_reg_797[4], ush_reg_797[4], ush_reg_797 };
assign ashr_ln1333_fu_484_p2 = \ashr_32s_32s_32_1_1_U3.dout ;
assign \ashr_32s_16ns_32_2_1_U4.din1_cast  = \ashr_32s_16ns_32_2_1_U4.din1 [15:0];
assign \ashr_32s_16ns_32_2_1_U4.din1_mask  = 16'h00ff;
assign \ashr_32s_16ns_32_2_1_U4.ce  = 1'h1;
assign \ashr_32s_16ns_32_2_1_U4.clk  = ap_clk;
assign \ashr_32s_16ns_32_2_1_U4.din0  = { ret_V_24_reg_843[2], ret_V_24_reg_843[2], ret_V_24_reg_843[2], ret_V_24_reg_843[2], ret_V_24_reg_843[2], ret_V_24_reg_843[2], ret_V_24_reg_843[2], ret_V_24_reg_843[2], ret_V_24_reg_843[2], ret_V_24_reg_843[2], ret_V_24_reg_843[2], ret_V_24_reg_843[2], ret_V_24_reg_843[2], ret_V_24_reg_843[2], ret_V_24_reg_843[2], ret_V_24_reg_843[2], ret_V_24_reg_843[2], ret_V_24_reg_843[2], ret_V_24_reg_843[2], ret_V_24_reg_843[2], ret_V_24_reg_843[2], ret_V_24_reg_843[2], ret_V_24_reg_843[2], ret_V_24_reg_843[2], ret_V_24_reg_843[2], ret_V_24_reg_843[2], ret_V_24_reg_843[2], ret_V_24_reg_843[2], ret_V_24_reg_843[2], ret_V_24_reg_843 };
assign \ashr_32s_16ns_32_2_1_U4.din1  = { 16'h0000, sh_V_1_reg_860[3], sh_V_1_reg_860[3], sh_V_1_reg_860[3], sh_V_1_reg_860[3], sh_V_1_reg_860[3], sh_V_1_reg_860[3], sh_V_1_reg_860[3], sh_V_1_reg_860[3], sh_V_1_reg_860[3], sh_V_1_reg_860[3], sh_V_1_reg_860[3], sh_V_1_reg_860[3], sh_V_1_reg_860 };
assign grp_fu_601_p2 = \ashr_32s_16ns_32_2_1_U4.dout ;
assign \ashr_32s_16ns_32_2_1_U4.reset  = ap_rst;
endmodule


// Machine B:
// Processed by function `add_clk_enable_signal` in `verilog_tricks.py`.
// Processed by function `remove_reset_signal` in `verilog_tricks.py`.
module top_B (
  ap_clk,
  ap_start,
  ap_done,
  ap_idle,
  ap_ready,
  op_0,
  op_1,
  op_2,
  op_5,
  op_8,
  op_12,
  op_14,
  op_16,
  op_18,
  op_30,
  op_30_ap_vld,
clk_enable
);
input clk_enable;


input ap_clk;
wire ap_rst;
assign ap_rst = op_30_ap_vld;
input ap_start;
input [1:0] op_0;
input [3:0] op_1;
input [1:0] op_12;
input op_14;
input [3:0] op_16;
input [3:0] op_18;
input [7:0] op_2;
input [3:0] op_5;
input [3:0] op_8;
output ap_done;
output ap_idle;
output ap_ready;
output [31:0] op_30;
output op_30_ap_vld;


reg [4:0] \add_10ns_10ns_10_2_1_U3.top_add_10ns_10ns_10_2_1_Adder_1_U.ain_s1 ;
reg [4:0] \add_10ns_10ns_10_2_1_U3.top_add_10ns_10ns_10_2_1_Adder_1_U.bin_s1 ;
reg \add_10ns_10ns_10_2_1_U3.top_add_10ns_10ns_10_2_1_Adder_1_U.carry_s1 ;
reg [4:0] \add_10ns_10ns_10_2_1_U3.top_add_10ns_10ns_10_2_1_Adder_1_U.sum_s1 ;
reg [5:0] \add_11ns_11ns_11_2_1_U14.top_add_11ns_11ns_11_2_1_Adder_9_U.ain_s1 ;
reg [5:0] \add_11ns_11ns_11_2_1_U14.top_add_11ns_11ns_11_2_1_Adder_9_U.bin_s1 ;
reg \add_11ns_11ns_11_2_1_U14.top_add_11ns_11ns_11_2_1_Adder_9_U.carry_s1 ;
reg [4:0] \add_11ns_11ns_11_2_1_U14.top_add_11ns_11ns_11_2_1_Adder_9_U.sum_s1 ;
reg [5:0] \add_11ns_11ns_11_2_1_U16.top_add_11ns_11ns_11_2_1_Adder_9_U.ain_s1 ;
reg [5:0] \add_11ns_11ns_11_2_1_U16.top_add_11ns_11ns_11_2_1_Adder_9_U.bin_s1 ;
reg \add_11ns_11ns_11_2_1_U16.top_add_11ns_11ns_11_2_1_Adder_9_U.carry_s1 ;
reg [4:0] \add_11ns_11ns_11_2_1_U16.top_add_11ns_11ns_11_2_1_Adder_9_U.sum_s1 ;
reg [5:0] \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_7_U.ain_s1 ;
reg [5:0] \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_7_U.bin_s1 ;
reg \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_7_U.carry_s1 ;
reg [4:0] \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_7_U.sum_s1 ;
reg [5:0] \add_11ns_11s_11_2_1_U20.top_add_11ns_11s_11_2_1_Adder_7_U.ain_s1 ;
reg [5:0] \add_11ns_11s_11_2_1_U20.top_add_11ns_11s_11_2_1_Adder_7_U.bin_s1 ;
reg \add_11ns_11s_11_2_1_U20.top_add_11ns_11s_11_2_1_Adder_7_U.carry_s1 ;
reg [4:0] \add_11ns_11s_11_2_1_U20.top_add_11ns_11s_11_2_1_Adder_7_U.sum_s1 ;
reg [5:0] \add_11ns_11s_11_2_1_U21.top_add_11ns_11s_11_2_1_Adder_7_U.ain_s1 ;
reg [5:0] \add_11ns_11s_11_2_1_U21.top_add_11ns_11s_11_2_1_Adder_7_U.bin_s1 ;
reg \add_11ns_11s_11_2_1_U21.top_add_11ns_11s_11_2_1_Adder_7_U.carry_s1 ;
reg [4:0] \add_11ns_11s_11_2_1_U21.top_add_11ns_11s_11_2_1_Adder_7_U.sum_s1 ;
reg [5:0] \add_11s_11ns_11_2_1_U13.top_add_11s_11ns_11_2_1_Adder_4_U.ain_s1 ;
reg [5:0] \add_11s_11ns_11_2_1_U13.top_add_11s_11ns_11_2_1_Adder_4_U.bin_s1 ;
reg \add_11s_11ns_11_2_1_U13.top_add_11s_11ns_11_2_1_Adder_4_U.carry_s1 ;
reg [4:0] \add_11s_11ns_11_2_1_U13.top_add_11s_11ns_11_2_1_Adder_4_U.sum_s1 ;
reg [5:0] \add_11s_11ns_11_2_1_U6.top_add_11s_11ns_11_2_1_Adder_4_U.ain_s1 ;
reg [5:0] \add_11s_11ns_11_2_1_U6.top_add_11s_11ns_11_2_1_Adder_4_U.bin_s1 ;
reg \add_11s_11ns_11_2_1_U6.top_add_11s_11ns_11_2_1_Adder_4_U.carry_s1 ;
reg [4:0] \add_11s_11ns_11_2_1_U6.top_add_11s_11ns_11_2_1_Adder_4_U.sum_s1 ;
reg [5:0] \add_12ns_12s_12_2_1_U1.top_add_12ns_12s_12_2_1_Adder_0_U.ain_s1 ;
reg [5:0] \add_12ns_12s_12_2_1_U1.top_add_12ns_12s_12_2_1_Adder_0_U.bin_s1 ;
reg \add_12ns_12s_12_2_1_U1.top_add_12ns_12s_12_2_1_Adder_0_U.carry_s1 ;
reg [5:0] \add_12ns_12s_12_2_1_U1.top_add_12ns_12s_12_2_1_Adder_0_U.sum_s1 ;
reg \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_3_U.ain_s1 ;
reg \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_3_U.bin_s1 ;
reg \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_3_U.carry_s1 ;
reg \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_3_U.sum_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_13_U.ain_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_13_U.bin_s1 ;
reg \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_13_U.carry_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_13_U.sum_s1 ;
reg [17:0] \add_35s_35s_35_2_1_U22.top_add_35s_35s_35_2_1_Adder_12_U.ain_s1 ;
reg [17:0] \add_35s_35s_35_2_1_U22.top_add_35s_35s_35_2_1_Adder_12_U.bin_s1 ;
reg \add_35s_35s_35_2_1_U22.top_add_35s_35s_35_2_1_Adder_12_U.carry_s1 ;
reg [16:0] \add_35s_35s_35_2_1_U22.top_add_35s_35s_35_2_1_Adder_12_U.sum_s1 ;
reg [1:0] \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_10_U.ain_s1 ;
reg [1:0] \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_10_U.bin_s1 ;
reg \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_10_U.carry_s1 ;
reg \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_10_U.sum_s1 ;
reg [1:0] \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.ain_s1 ;
reg [1:0] \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.bin_s1 ;
reg \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.carry_s1 ;
reg \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.sum_s1 ;
reg [1:0] \add_3s_3s_3_2_1_U9.top_add_3s_3s_3_2_1_Adder_5_U.ain_s1 ;
reg [1:0] \add_3s_3s_3_2_1_U9.top_add_3s_3s_3_2_1_Adder_5_U.bin_s1 ;
reg \add_3s_3s_3_2_1_U9.top_add_3s_3s_3_2_1_Adder_5_U.carry_s1 ;
reg \add_3s_3s_3_2_1_U9.top_add_3s_3s_3_2_1_Adder_5_U.sum_s1 ;
reg [2:0] \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_8_U.ain_s1 ;
reg [2:0] \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_8_U.bin_s1 ;
reg \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_8_U.carry_s1 ;
reg [2:0] \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_8_U.sum_s1 ;
reg [31:0] add_ln691_1_reg_1088;
reg [10:0] add_ln691_reg_990;
reg [2:0] add_ln69_1_reg_897;
reg [5:0] add_ln69_2_reg_922;
reg [10:0] add_ln69_reg_917;
reg [36:0] ap_CS_fsm = 37'h0000000001;
reg [15:0] \ashr_32s_16ns_32_7_1_U18.din1_cast_array[0] ;
reg [15:0] \ashr_32s_16ns_32_7_1_U18.din1_cast_array[1] ;
reg [15:0] \ashr_32s_16ns_32_7_1_U18.din1_cast_array[2] ;
reg [15:0] \ashr_32s_16ns_32_7_1_U18.din1_cast_array[3] ;
reg [15:0] \ashr_32s_16ns_32_7_1_U18.din1_cast_array[4] ;
reg [15:0] \ashr_32s_16ns_32_7_1_U18.din1_cast_array[5] ;
reg [31:0] \ashr_32s_16ns_32_7_1_U18.dout_array[0] ;
reg [31:0] \ashr_32s_16ns_32_7_1_U18.dout_array[1] ;
reg [31:0] \ashr_32s_16ns_32_7_1_U18.dout_array[2] ;
reg [31:0] \ashr_32s_16ns_32_7_1_U18.dout_array[3] ;
reg [31:0] \ashr_32s_16ns_32_7_1_U18.dout_array[4] ;
reg [31:0] \ashr_32s_16ns_32_7_1_U18.dout_array[5] ;
reg [31:0] \ashr_32s_32s_32_7_1_U8.din1_cast_array[0] ;
reg [31:0] \ashr_32s_32s_32_7_1_U8.din1_cast_array[1] ;
reg [31:0] \ashr_32s_32s_32_7_1_U8.din1_cast_array[2] ;
reg [31:0] \ashr_32s_32s_32_7_1_U8.din1_cast_array[3] ;
reg [31:0] \ashr_32s_32s_32_7_1_U8.din1_cast_array[4] ;
reg [31:0] \ashr_32s_32s_32_7_1_U8.din1_cast_array[5] ;
reg [31:0] \ashr_32s_32s_32_7_1_U8.dout_array[0] ;
reg [31:0] \ashr_32s_32s_32_7_1_U8.dout_array[1] ;
reg [31:0] \ashr_32s_32s_32_7_1_U8.dout_array[2] ;
reg [31:0] \ashr_32s_32s_32_7_1_U8.dout_array[3] ;
reg [31:0] \ashr_32s_32s_32_7_1_U8.dout_array[4] ;
reg [31:0] \ashr_32s_32s_32_7_1_U8.dout_array[5] ;
reg [31:0] ashr_ln1333_reg_937;
reg icmp_ln1499_reg_726;
reg icmp_ln851_1_reg_798;
reg icmp_ln851_2_reg_845;
reg icmp_ln851_3_reg_1071;
reg icmp_ln851_reg_711;
reg isNeg_reg_769;
reg lhs_V_2_reg_833;
reg [10:0] op_24_V_reg_942;
reg [10:0] op_27_V_reg_1046;
reg [3:0] op_7_V_reg_764;
reg p_Result_8_reg_985;
reg [5:0] r_reg_1041;
reg [2:0] ret_V_11_reg_958;
reg [2:0] ret_V_12_reg_973;
reg [11:0] ret_V_19_reg_736;
reg [9:0] ret_V_20_reg_753;
reg [1:0] ret_V_21_reg_828;
reg [10:0] ret_V_23_reg_887;
reg [2:0] ret_V_24_reg_978;
reg [10:0] ret_V_25_reg_965;
reg [10:0] ret_V_26_reg_1000;
reg [10:0] ret_V_27_reg_1056;
reg [34:0] ret_V_28_reg_1076;
reg [9:0] ret_V_2_reg_748;
reg [31:0] ret_V_30_cast_reg_1081;
reg [1:0] ret_V_3_reg_780;
reg [1:0] ret_V_5_reg_808;
reg [9:0] ret_V_8_reg_813;
reg [10:0] ret_V_9_reg_862;
reg [9:0] ret_V_reg_741;
reg [2:0] ret_reg_892;
reg [10:0] select_ln1192_reg_947;
reg [31:0] select_ln1368_reg_952;
reg [4:0] sext_ln1386_reg_792;
reg [10:0] sext_ln831_reg_838;
reg [3:0] sh_V_1_reg_1005;
reg [15:0] \shl_32s_16ns_32_7_1_U19.din1_cast_array[0] ;
reg [15:0] \shl_32s_16ns_32_7_1_U19.din1_cast_array[1] ;
reg [15:0] \shl_32s_16ns_32_7_1_U19.din1_cast_array[2] ;
reg [15:0] \shl_32s_16ns_32_7_1_U19.din1_cast_array[3] ;
reg [15:0] \shl_32s_16ns_32_7_1_U19.din1_cast_array[4] ;
reg [15:0] \shl_32s_16ns_32_7_1_U19.din1_cast_array[5] ;
reg [31:0] \shl_32s_16ns_32_7_1_U19.dout_array[0] ;
reg [31:0] \shl_32s_16ns_32_7_1_U19.dout_array[1] ;
reg [31:0] \shl_32s_16ns_32_7_1_U19.dout_array[2] ;
reg [31:0] \shl_32s_16ns_32_7_1_U19.dout_array[3] ;
reg [31:0] \shl_32s_16ns_32_7_1_U19.dout_array[4] ;
reg [31:0] \shl_32s_16ns_32_7_1_U19.dout_array[5] ;
reg [31:0] \shl_32s_32s_32_7_1_U7.din1_cast_array[0] ;
reg [31:0] \shl_32s_32s_32_7_1_U7.din1_cast_array[1] ;
reg [31:0] \shl_32s_32s_32_7_1_U7.din1_cast_array[2] ;
reg [31:0] \shl_32s_32s_32_7_1_U7.din1_cast_array[3] ;
reg [31:0] \shl_32s_32s_32_7_1_U7.din1_cast_array[4] ;
reg [31:0] \shl_32s_32s_32_7_1_U7.din1_cast_array[5] ;
reg [31:0] \shl_32s_32s_32_7_1_U7.dout_array[0] ;
reg [31:0] \shl_32s_32s_32_7_1_U7.dout_array[1] ;
reg [31:0] \shl_32s_32s_32_7_1_U7.dout_array[2] ;
reg [31:0] \shl_32s_32s_32_7_1_U7.dout_array[3] ;
reg [31:0] \shl_32s_32s_32_7_1_U7.dout_array[4] ;
reg [31:0] \shl_32s_32s_32_7_1_U7.dout_array[5] ;
reg [7:0] \shl_32s_8ns_32_7_1_U2.din1_cast_array[0] ;
reg [7:0] \shl_32s_8ns_32_7_1_U2.din1_cast_array[1] ;
reg [7:0] \shl_32s_8ns_32_7_1_U2.din1_cast_array[2] ;
reg [7:0] \shl_32s_8ns_32_7_1_U2.din1_cast_array[3] ;
reg [7:0] \shl_32s_8ns_32_7_1_U2.din1_cast_array[4] ;
reg [7:0] \shl_32s_8ns_32_7_1_U2.din1_cast_array[5] ;
reg [31:0] \shl_32s_8ns_32_7_1_U2.dout_array[0] ;
reg [31:0] \shl_32s_8ns_32_7_1_U2.dout_array[1] ;
reg [31:0] \shl_32s_8ns_32_7_1_U2.dout_array[2] ;
reg [31:0] \shl_32s_8ns_32_7_1_U2.dout_array[3] ;
reg [31:0] \shl_32s_8ns_32_7_1_U2.dout_array[4] ;
reg [31:0] \shl_32s_8ns_32_7_1_U2.dout_array[5] ;
reg [31:0] shl_ln1299_1_reg_932;
reg [31:0] shl_ln1299_reg_775;
reg [1:0] \sub_4ns_4s_4_2_1_U17.top_sub_4ns_4s_4_2_1_Adder_11_U.ain_s1 ;
reg [1:0] \sub_4ns_4s_4_2_1_U17.top_sub_4ns_4s_4_2_1_Adder_11_U.bin_s1 ;
reg \sub_4ns_4s_4_2_1_U17.top_sub_4ns_4s_4_2_1_Adder_11_U.carry_s1 ;
reg [1:0] \sub_4ns_4s_4_2_1_U17.top_sub_4ns_4s_4_2_1_Adder_11_U.sum_s1 ;
reg [2:0] \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.ain_s1 ;
reg [2:0] \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.bin_s1 ;
reg \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.carry_s1 ;
reg [1:0] \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.sum_s1 ;
reg [4:0] sub_ln1367_reg_803;
reg [3:0] trunc_ln1348_1_reg_731;
reg [3:0] trunc_ln1348_reg_759;
reg [2:0] trunc_ln546_reg_1026;
reg [5:0] trunc_ln769_reg_1031;
reg [1:0] trunc_ln851_1_reg_787;
reg [1:0] trunc_ln851_2_reg_818;
reg [4:0] ush_reg_823;
wire [31:0] _000_;
wire [10:0] _001_;
wire [2:0] _002_;
wire [5:0] _003_;
wire [10:0] _004_;
wire [36:0] _005_;
wire [31:0] _006_;
wire _007_;
wire _008_;
wire _009_;
wire _010_;
wire _011_;
wire _012_;
wire _013_;
wire [10:0] _014_;
wire [10:0] _015_;
wire [3:0] _016_;
wire _017_;
wire [5:0] _018_;
wire [2:0] _019_;
wire [2:0] _020_;
wire [11:0] _021_;
wire [9:0] _022_;
wire [1:0] _023_;
wire [10:0] _024_;
wire [2:0] _025_;
wire [10:0] _026_;
wire [10:0] _027_;
wire [10:0] _028_;
wire [34:0] _029_;
wire [9:0] _030_;
wire [31:0] _031_;
wire [1:0] _032_;
wire [1:0] _033_;
wire [9:0] _034_;
wire [10:0] _035_;
wire [9:0] _036_;
wire [2:0] _037_;
wire [10:0] _038_;
wire [31:0] _039_;
wire [4:0] _040_;
wire [10:0] _041_;
wire [3:0] _042_;
wire [31:0] _043_;
wire [31:0] _044_;
wire [4:0] _045_;
wire [3:0] _046_;
wire [3:0] _047_;
wire [2:0] _048_;
wire [5:0] _049_;
wire [1:0] _050_;
wire [1:0] _051_;
wire [4:0] _052_;
wire [1:0] _053_;
wire _054_;
wire _055_;
wire _056_;
wire _057_;
wire _058_;
wire _059_;
wire _060_;
wire _061_;
wire _062_;
wire _063_;
wire _064_;
wire _065_;
wire _066_;
wire _067_;
wire _068_;
wire _069_;
wire _070_;
wire _071_;
wire _072_;
wire [4:0] _073_;
wire [4:0] _074_;
wire _075_;
wire [4:0] _076_;
wire [5:0] _077_;
wire [5:0] _078_;
wire [5:0] _079_;
wire [5:0] _080_;
wire _081_;
wire [4:0] _082_;
wire [5:0] _083_;
wire [6:0] _084_;
wire [5:0] _085_;
wire [5:0] _086_;
wire _087_;
wire [4:0] _088_;
wire [5:0] _089_;
wire [6:0] _090_;
wire [5:0] _091_;
wire [5:0] _092_;
wire _093_;
wire [4:0] _094_;
wire [5:0] _095_;
wire [6:0] _096_;
wire [5:0] _097_;
wire [5:0] _098_;
wire _099_;
wire [4:0] _100_;
wire [5:0] _101_;
wire [6:0] _102_;
wire [5:0] _103_;
wire [5:0] _104_;
wire _105_;
wire [4:0] _106_;
wire [5:0] _107_;
wire [6:0] _108_;
wire [5:0] _109_;
wire [5:0] _110_;
wire _111_;
wire [4:0] _112_;
wire [5:0] _113_;
wire [6:0] _114_;
wire [5:0] _115_;
wire [5:0] _116_;
wire _117_;
wire [4:0] _118_;
wire [5:0] _119_;
wire [6:0] _120_;
wire [5:0] _121_;
wire [5:0] _122_;
wire _123_;
wire [5:0] _124_;
wire [6:0] _125_;
wire [6:0] _126_;
wire _127_;
wire _128_;
wire _129_;
wire _130_;
wire [1:0] _131_;
wire [1:0] _132_;
wire [15:0] _133_;
wire [15:0] _134_;
wire _135_;
wire [15:0] _136_;
wire [16:0] _137_;
wire [16:0] _138_;
wire [17:0] _139_;
wire [17:0] _140_;
wire _141_;
wire [16:0] _142_;
wire [17:0] _143_;
wire [18:0] _144_;
wire [1:0] _145_;
wire [1:0] _146_;
wire _147_;
wire _148_;
wire [1:0] _149_;
wire [2:0] _150_;
wire [1:0] _151_;
wire [1:0] _152_;
wire _153_;
wire _154_;
wire [1:0] _155_;
wire [2:0] _156_;
wire [1:0] _157_;
wire [1:0] _158_;
wire _159_;
wire _160_;
wire [1:0] _161_;
wire [2:0] _162_;
wire [2:0] _163_;
wire [2:0] _164_;
wire _165_;
wire [2:0] _166_;
wire [3:0] _167_;
wire [3:0] _168_;
wire [15:0] _169_;
wire [15:0] _170_;
wire [15:0] _171_;
wire [15:0] _172_;
wire [15:0] _173_;
wire [15:0] _174_;
wire [31:0] _175_;
wire [31:0] _176_;
wire [31:0] _177_;
wire [31:0] _178_;
wire [31:0] _179_;
wire [31:0] _180_;
wire [15:0] _181_;
wire [31:0] _182_;
wire [15:0] _183_;
wire [31:0] _184_;
wire [15:0] _185_;
wire [31:0] _186_;
wire [15:0] _187_;
wire [31:0] _188_;
wire [15:0] _189_;
wire [31:0] _190_;
wire [15:0] _191_;
wire [31:0] _192_;
wire [31:0] _193_;
wire [31:0] _194_;
wire [31:0] _195_;
wire [31:0] _196_;
wire [31:0] _197_;
wire [31:0] _198_;
wire [31:0] _199_;
wire [31:0] _200_;
wire [31:0] _201_;
wire [31:0] _202_;
wire [31:0] _203_;
wire [31:0] _204_;
wire [31:0] _205_;
wire [31:0] _206_;
wire [31:0] _207_;
wire [31:0] _208_;
wire [31:0] _209_;
wire [31:0] _210_;
wire [31:0] _211_;
wire [31:0] _212_;
wire [31:0] _213_;
wire [31:0] _214_;
wire [31:0] _215_;
wire [31:0] _216_;
wire [31:0] _217_;
wire [31:0] _218_;
wire [31:0] _219_;
wire [31:0] _220_;
wire [31:0] _221_;
wire [31:0] _222_;
wire [31:0] _223_;
wire [31:0] _224_;
wire [31:0] _225_;
wire [31:0] _226_;
wire [31:0] _227_;
wire [15:0] _228_;
wire [15:0] _229_;
wire [15:0] _230_;
wire [15:0] _231_;
wire [15:0] _232_;
wire [15:0] _233_;
wire [31:0] _234_;
wire [31:0] _235_;
wire [31:0] _236_;
wire [31:0] _237_;
wire [31:0] _238_;
wire [31:0] _239_;
wire [15:0] _240_;
wire [31:0] _241_;
wire [15:0] _242_;
wire [31:0] _243_;
wire [15:0] _244_;
wire [31:0] _245_;
wire [15:0] _246_;
wire [31:0] _247_;
wire [15:0] _248_;
wire [31:0] _249_;
wire [15:0] _250_;
wire [31:0] _251_;
wire [31:0] _252_;
wire [31:0] _253_;
wire [31:0] _254_;
wire [31:0] _255_;
wire [31:0] _256_;
wire [31:0] _257_;
wire [31:0] _258_;
wire [31:0] _259_;
wire [31:0] _260_;
wire [31:0] _261_;
wire [31:0] _262_;
wire [31:0] _263_;
wire [31:0] _264_;
wire [31:0] _265_;
wire [31:0] _266_;
wire [31:0] _267_;
wire [31:0] _268_;
wire [31:0] _269_;
wire [31:0] _270_;
wire [31:0] _271_;
wire [31:0] _272_;
wire [31:0] _273_;
wire [31:0] _274_;
wire [31:0] _275_;
wire [31:0] _276_;
wire [31:0] _277_;
wire [31:0] _278_;
wire [31:0] _279_;
wire [31:0] _280_;
wire [31:0] _281_;
wire [31:0] _282_;
wire [31:0] _283_;
wire [31:0] _284_;
wire [31:0] _285_;
wire [31:0] _286_;
wire [7:0] _287_;
wire [7:0] _288_;
wire [7:0] _289_;
wire [7:0] _290_;
wire [7:0] _291_;
wire [7:0] _292_;
wire [31:0] _293_;
wire [31:0] _294_;
wire [31:0] _295_;
wire [31:0] _296_;
wire [31:0] _297_;
wire [31:0] _298_;
wire [7:0] _299_;
wire [31:0] _300_;
wire [7:0] _301_;
wire [31:0] _302_;
wire [7:0] _303_;
wire [31:0] _304_;
wire [7:0] _305_;
wire [31:0] _306_;
wire [7:0] _307_;
wire [31:0] _308_;
wire [7:0] _309_;
wire [31:0] _310_;
wire [31:0] _311_;
wire [31:0] _312_;
wire [31:0] _313_;
wire [1:0] _314_;
wire [1:0] _315_;
wire _316_;
wire [1:0] _317_;
wire [2:0] _318_;
wire [2:0] _319_;
wire [2:0] _320_;
wire [2:0] _321_;
wire _322_;
wire [1:0] _323_;
wire [2:0] _324_;
wire [3:0] _325_;
wire _326_;
wire _327_;
wire _328_;
wire _329_;
wire _330_;
wire _331_;
wire _332_;
wire _333_;
wire _334_;
wire _335_;
wire _336_;
wire _337_;
wire _338_;
wire _339_;
wire _340_;
wire _341_;
wire _342_;
wire _343_;
wire _344_;
wire _345_;
wire _346_;
wire _347_;
wire _348_;
wire _349_;
wire _350_;
wire _351_;
wire _352_;
wire _353_;
wire _354_;
wire _355_;
wire _356_;
wire _357_;
wire _358_;
wire _359_;
wire _360_;
wire _361_;
wire _362_;
wire _363_;
wire _364_;
wire \add_10ns_10ns_10_2_1_U3.ce ;
wire \add_10ns_10ns_10_2_1_U3.clk ;
wire [9:0] \add_10ns_10ns_10_2_1_U3.din0 ;
wire [9:0] \add_10ns_10ns_10_2_1_U3.din1 ;
wire [9:0] \add_10ns_10ns_10_2_1_U3.dout ;
wire \add_10ns_10ns_10_2_1_U3.reset ;
wire [9:0] \add_10ns_10ns_10_2_1_U3.top_add_10ns_10ns_10_2_1_Adder_1_U.a ;
wire [9:0] \add_10ns_10ns_10_2_1_U3.top_add_10ns_10ns_10_2_1_Adder_1_U.ain_s0 ;
wire [9:0] \add_10ns_10ns_10_2_1_U3.top_add_10ns_10ns_10_2_1_Adder_1_U.b ;
wire [9:0] \add_10ns_10ns_10_2_1_U3.top_add_10ns_10ns_10_2_1_Adder_1_U.bin_s0 ;
wire \add_10ns_10ns_10_2_1_U3.top_add_10ns_10ns_10_2_1_Adder_1_U.ce ;
wire \add_10ns_10ns_10_2_1_U3.top_add_10ns_10ns_10_2_1_Adder_1_U.clk ;
wire \add_10ns_10ns_10_2_1_U3.top_add_10ns_10ns_10_2_1_Adder_1_U.facout_s1 ;
wire \add_10ns_10ns_10_2_1_U3.top_add_10ns_10ns_10_2_1_Adder_1_U.facout_s2 ;
wire [4:0] \add_10ns_10ns_10_2_1_U3.top_add_10ns_10ns_10_2_1_Adder_1_U.fas_s1 ;
wire [4:0] \add_10ns_10ns_10_2_1_U3.top_add_10ns_10ns_10_2_1_Adder_1_U.fas_s2 ;
wire \add_10ns_10ns_10_2_1_U3.top_add_10ns_10ns_10_2_1_Adder_1_U.reset ;
wire [9:0] \add_10ns_10ns_10_2_1_U3.top_add_10ns_10ns_10_2_1_Adder_1_U.s ;
wire [4:0] \add_10ns_10ns_10_2_1_U3.top_add_10ns_10ns_10_2_1_Adder_1_U.u1.a ;
wire [4:0] \add_10ns_10ns_10_2_1_U3.top_add_10ns_10ns_10_2_1_Adder_1_U.u1.b ;
wire \add_10ns_10ns_10_2_1_U3.top_add_10ns_10ns_10_2_1_Adder_1_U.u1.cin ;
wire \add_10ns_10ns_10_2_1_U3.top_add_10ns_10ns_10_2_1_Adder_1_U.u1.cout ;
wire [4:0] \add_10ns_10ns_10_2_1_U3.top_add_10ns_10ns_10_2_1_Adder_1_U.u1.s ;
wire [4:0] \add_10ns_10ns_10_2_1_U3.top_add_10ns_10ns_10_2_1_Adder_1_U.u2.a ;
wire [4:0] \add_10ns_10ns_10_2_1_U3.top_add_10ns_10ns_10_2_1_Adder_1_U.u2.b ;
wire \add_10ns_10ns_10_2_1_U3.top_add_10ns_10ns_10_2_1_Adder_1_U.u2.cin ;
wire \add_10ns_10ns_10_2_1_U3.top_add_10ns_10ns_10_2_1_Adder_1_U.u2.cout ;
wire [4:0] \add_10ns_10ns_10_2_1_U3.top_add_10ns_10ns_10_2_1_Adder_1_U.u2.s ;
wire \add_11ns_11ns_11_2_1_U14.ce ;
wire \add_11ns_11ns_11_2_1_U14.clk ;
wire [10:0] \add_11ns_11ns_11_2_1_U14.din0 ;
wire [10:0] \add_11ns_11ns_11_2_1_U14.din1 ;
wire [10:0] \add_11ns_11ns_11_2_1_U14.dout ;
wire \add_11ns_11ns_11_2_1_U14.reset ;
wire [10:0] \add_11ns_11ns_11_2_1_U14.top_add_11ns_11ns_11_2_1_Adder_9_U.a ;
wire [10:0] \add_11ns_11ns_11_2_1_U14.top_add_11ns_11ns_11_2_1_Adder_9_U.ain_s0 ;
wire [10:0] \add_11ns_11ns_11_2_1_U14.top_add_11ns_11ns_11_2_1_Adder_9_U.b ;
wire [10:0] \add_11ns_11ns_11_2_1_U14.top_add_11ns_11ns_11_2_1_Adder_9_U.bin_s0 ;
wire \add_11ns_11ns_11_2_1_U14.top_add_11ns_11ns_11_2_1_Adder_9_U.ce ;
wire \add_11ns_11ns_11_2_1_U14.top_add_11ns_11ns_11_2_1_Adder_9_U.clk ;
wire \add_11ns_11ns_11_2_1_U14.top_add_11ns_11ns_11_2_1_Adder_9_U.facout_s1 ;
wire \add_11ns_11ns_11_2_1_U14.top_add_11ns_11ns_11_2_1_Adder_9_U.facout_s2 ;
wire [4:0] \add_11ns_11ns_11_2_1_U14.top_add_11ns_11ns_11_2_1_Adder_9_U.fas_s1 ;
wire [5:0] \add_11ns_11ns_11_2_1_U14.top_add_11ns_11ns_11_2_1_Adder_9_U.fas_s2 ;
wire \add_11ns_11ns_11_2_1_U14.top_add_11ns_11ns_11_2_1_Adder_9_U.reset ;
wire [10:0] \add_11ns_11ns_11_2_1_U14.top_add_11ns_11ns_11_2_1_Adder_9_U.s ;
wire [4:0] \add_11ns_11ns_11_2_1_U14.top_add_11ns_11ns_11_2_1_Adder_9_U.u1.a ;
wire [4:0] \add_11ns_11ns_11_2_1_U14.top_add_11ns_11ns_11_2_1_Adder_9_U.u1.b ;
wire \add_11ns_11ns_11_2_1_U14.top_add_11ns_11ns_11_2_1_Adder_9_U.u1.cin ;
wire \add_11ns_11ns_11_2_1_U14.top_add_11ns_11ns_11_2_1_Adder_9_U.u1.cout ;
wire [4:0] \add_11ns_11ns_11_2_1_U14.top_add_11ns_11ns_11_2_1_Adder_9_U.u1.s ;
wire [5:0] \add_11ns_11ns_11_2_1_U14.top_add_11ns_11ns_11_2_1_Adder_9_U.u2.a ;
wire [5:0] \add_11ns_11ns_11_2_1_U14.top_add_11ns_11ns_11_2_1_Adder_9_U.u2.b ;
wire \add_11ns_11ns_11_2_1_U14.top_add_11ns_11ns_11_2_1_Adder_9_U.u2.cin ;
wire \add_11ns_11ns_11_2_1_U14.top_add_11ns_11ns_11_2_1_Adder_9_U.u2.cout ;
wire [5:0] \add_11ns_11ns_11_2_1_U14.top_add_11ns_11ns_11_2_1_Adder_9_U.u2.s ;
wire \add_11ns_11ns_11_2_1_U16.ce ;
wire \add_11ns_11ns_11_2_1_U16.clk ;
wire [10:0] \add_11ns_11ns_11_2_1_U16.din0 ;
wire [10:0] \add_11ns_11ns_11_2_1_U16.din1 ;
wire [10:0] \add_11ns_11ns_11_2_1_U16.dout ;
wire \add_11ns_11ns_11_2_1_U16.reset ;
wire [10:0] \add_11ns_11ns_11_2_1_U16.top_add_11ns_11ns_11_2_1_Adder_9_U.a ;
wire [10:0] \add_11ns_11ns_11_2_1_U16.top_add_11ns_11ns_11_2_1_Adder_9_U.ain_s0 ;
wire [10:0] \add_11ns_11ns_11_2_1_U16.top_add_11ns_11ns_11_2_1_Adder_9_U.b ;
wire [10:0] \add_11ns_11ns_11_2_1_U16.top_add_11ns_11ns_11_2_1_Adder_9_U.bin_s0 ;
wire \add_11ns_11ns_11_2_1_U16.top_add_11ns_11ns_11_2_1_Adder_9_U.ce ;
wire \add_11ns_11ns_11_2_1_U16.top_add_11ns_11ns_11_2_1_Adder_9_U.clk ;
wire \add_11ns_11ns_11_2_1_U16.top_add_11ns_11ns_11_2_1_Adder_9_U.facout_s1 ;
wire \add_11ns_11ns_11_2_1_U16.top_add_11ns_11ns_11_2_1_Adder_9_U.facout_s2 ;
wire [4:0] \add_11ns_11ns_11_2_1_U16.top_add_11ns_11ns_11_2_1_Adder_9_U.fas_s1 ;
wire [5:0] \add_11ns_11ns_11_2_1_U16.top_add_11ns_11ns_11_2_1_Adder_9_U.fas_s2 ;
wire \add_11ns_11ns_11_2_1_U16.top_add_11ns_11ns_11_2_1_Adder_9_U.reset ;
wire [10:0] \add_11ns_11ns_11_2_1_U16.top_add_11ns_11ns_11_2_1_Adder_9_U.s ;
wire [4:0] \add_11ns_11ns_11_2_1_U16.top_add_11ns_11ns_11_2_1_Adder_9_U.u1.a ;
wire [4:0] \add_11ns_11ns_11_2_1_U16.top_add_11ns_11ns_11_2_1_Adder_9_U.u1.b ;
wire \add_11ns_11ns_11_2_1_U16.top_add_11ns_11ns_11_2_1_Adder_9_U.u1.cin ;
wire \add_11ns_11ns_11_2_1_U16.top_add_11ns_11ns_11_2_1_Adder_9_U.u1.cout ;
wire [4:0] \add_11ns_11ns_11_2_1_U16.top_add_11ns_11ns_11_2_1_Adder_9_U.u1.s ;
wire [5:0] \add_11ns_11ns_11_2_1_U16.top_add_11ns_11ns_11_2_1_Adder_9_U.u2.a ;
wire [5:0] \add_11ns_11ns_11_2_1_U16.top_add_11ns_11ns_11_2_1_Adder_9_U.u2.b ;
wire \add_11ns_11ns_11_2_1_U16.top_add_11ns_11ns_11_2_1_Adder_9_U.u2.cin ;
wire \add_11ns_11ns_11_2_1_U16.top_add_11ns_11ns_11_2_1_Adder_9_U.u2.cout ;
wire [5:0] \add_11ns_11ns_11_2_1_U16.top_add_11ns_11ns_11_2_1_Adder_9_U.u2.s ;
wire \add_11ns_11s_11_2_1_U11.ce ;
wire \add_11ns_11s_11_2_1_U11.clk ;
wire [10:0] \add_11ns_11s_11_2_1_U11.din0 ;
wire [10:0] \add_11ns_11s_11_2_1_U11.din1 ;
wire [10:0] \add_11ns_11s_11_2_1_U11.dout ;
wire \add_11ns_11s_11_2_1_U11.reset ;
wire [10:0] \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_7_U.a ;
wire [10:0] \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_7_U.ain_s0 ;
wire [10:0] \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_7_U.b ;
wire [10:0] \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_7_U.bin_s0 ;
wire \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_7_U.ce ;
wire \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_7_U.clk ;
wire \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_7_U.facout_s1 ;
wire \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_7_U.facout_s2 ;
wire [4:0] \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_7_U.fas_s1 ;
wire [5:0] \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_7_U.fas_s2 ;
wire \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_7_U.reset ;
wire [10:0] \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_7_U.s ;
wire [4:0] \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_7_U.u1.a ;
wire [4:0] \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_7_U.u1.b ;
wire \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_7_U.u1.cin ;
wire \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_7_U.u1.cout ;
wire [4:0] \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_7_U.u1.s ;
wire [5:0] \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_7_U.u2.a ;
wire [5:0] \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_7_U.u2.b ;
wire \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_7_U.u2.cin ;
wire \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_7_U.u2.cout ;
wire [5:0] \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_7_U.u2.s ;
wire \add_11ns_11s_11_2_1_U20.ce ;
wire \add_11ns_11s_11_2_1_U20.clk ;
wire [10:0] \add_11ns_11s_11_2_1_U20.din0 ;
wire [10:0] \add_11ns_11s_11_2_1_U20.din1 ;
wire [10:0] \add_11ns_11s_11_2_1_U20.dout ;
wire \add_11ns_11s_11_2_1_U20.reset ;
wire [10:0] \add_11ns_11s_11_2_1_U20.top_add_11ns_11s_11_2_1_Adder_7_U.a ;
wire [10:0] \add_11ns_11s_11_2_1_U20.top_add_11ns_11s_11_2_1_Adder_7_U.ain_s0 ;
wire [10:0] \add_11ns_11s_11_2_1_U20.top_add_11ns_11s_11_2_1_Adder_7_U.b ;
wire [10:0] \add_11ns_11s_11_2_1_U20.top_add_11ns_11s_11_2_1_Adder_7_U.bin_s0 ;
wire \add_11ns_11s_11_2_1_U20.top_add_11ns_11s_11_2_1_Adder_7_U.ce ;
wire \add_11ns_11s_11_2_1_U20.top_add_11ns_11s_11_2_1_Adder_7_U.clk ;
wire \add_11ns_11s_11_2_1_U20.top_add_11ns_11s_11_2_1_Adder_7_U.facout_s1 ;
wire \add_11ns_11s_11_2_1_U20.top_add_11ns_11s_11_2_1_Adder_7_U.facout_s2 ;
wire [4:0] \add_11ns_11s_11_2_1_U20.top_add_11ns_11s_11_2_1_Adder_7_U.fas_s1 ;
wire [5:0] \add_11ns_11s_11_2_1_U20.top_add_11ns_11s_11_2_1_Adder_7_U.fas_s2 ;
wire \add_11ns_11s_11_2_1_U20.top_add_11ns_11s_11_2_1_Adder_7_U.reset ;
wire [10:0] \add_11ns_11s_11_2_1_U20.top_add_11ns_11s_11_2_1_Adder_7_U.s ;
wire [4:0] \add_11ns_11s_11_2_1_U20.top_add_11ns_11s_11_2_1_Adder_7_U.u1.a ;
wire [4:0] \add_11ns_11s_11_2_1_U20.top_add_11ns_11s_11_2_1_Adder_7_U.u1.b ;
wire \add_11ns_11s_11_2_1_U20.top_add_11ns_11s_11_2_1_Adder_7_U.u1.cin ;
wire \add_11ns_11s_11_2_1_U20.top_add_11ns_11s_11_2_1_Adder_7_U.u1.cout ;
wire [4:0] \add_11ns_11s_11_2_1_U20.top_add_11ns_11s_11_2_1_Adder_7_U.u1.s ;
wire [5:0] \add_11ns_11s_11_2_1_U20.top_add_11ns_11s_11_2_1_Adder_7_U.u2.a ;
wire [5:0] \add_11ns_11s_11_2_1_U20.top_add_11ns_11s_11_2_1_Adder_7_U.u2.b ;
wire \add_11ns_11s_11_2_1_U20.top_add_11ns_11s_11_2_1_Adder_7_U.u2.cin ;
wire \add_11ns_11s_11_2_1_U20.top_add_11ns_11s_11_2_1_Adder_7_U.u2.cout ;
wire [5:0] \add_11ns_11s_11_2_1_U20.top_add_11ns_11s_11_2_1_Adder_7_U.u2.s ;
wire \add_11ns_11s_11_2_1_U21.ce ;
wire \add_11ns_11s_11_2_1_U21.clk ;
wire [10:0] \add_11ns_11s_11_2_1_U21.din0 ;
wire [10:0] \add_11ns_11s_11_2_1_U21.din1 ;
wire [10:0] \add_11ns_11s_11_2_1_U21.dout ;
wire \add_11ns_11s_11_2_1_U21.reset ;
wire [10:0] \add_11ns_11s_11_2_1_U21.top_add_11ns_11s_11_2_1_Adder_7_U.a ;
wire [10:0] \add_11ns_11s_11_2_1_U21.top_add_11ns_11s_11_2_1_Adder_7_U.ain_s0 ;
wire [10:0] \add_11ns_11s_11_2_1_U21.top_add_11ns_11s_11_2_1_Adder_7_U.b ;
wire [10:0] \add_11ns_11s_11_2_1_U21.top_add_11ns_11s_11_2_1_Adder_7_U.bin_s0 ;
wire \add_11ns_11s_11_2_1_U21.top_add_11ns_11s_11_2_1_Adder_7_U.ce ;
wire \add_11ns_11s_11_2_1_U21.top_add_11ns_11s_11_2_1_Adder_7_U.clk ;
wire \add_11ns_11s_11_2_1_U21.top_add_11ns_11s_11_2_1_Adder_7_U.facout_s1 ;
wire \add_11ns_11s_11_2_1_U21.top_add_11ns_11s_11_2_1_Adder_7_U.facout_s2 ;
wire [4:0] \add_11ns_11s_11_2_1_U21.top_add_11ns_11s_11_2_1_Adder_7_U.fas_s1 ;
wire [5:0] \add_11ns_11s_11_2_1_U21.top_add_11ns_11s_11_2_1_Adder_7_U.fas_s2 ;
wire \add_11ns_11s_11_2_1_U21.top_add_11ns_11s_11_2_1_Adder_7_U.reset ;
wire [10:0] \add_11ns_11s_11_2_1_U21.top_add_11ns_11s_11_2_1_Adder_7_U.s ;
wire [4:0] \add_11ns_11s_11_2_1_U21.top_add_11ns_11s_11_2_1_Adder_7_U.u1.a ;
wire [4:0] \add_11ns_11s_11_2_1_U21.top_add_11ns_11s_11_2_1_Adder_7_U.u1.b ;
wire \add_11ns_11s_11_2_1_U21.top_add_11ns_11s_11_2_1_Adder_7_U.u1.cin ;
wire \add_11ns_11s_11_2_1_U21.top_add_11ns_11s_11_2_1_Adder_7_U.u1.cout ;
wire [4:0] \add_11ns_11s_11_2_1_U21.top_add_11ns_11s_11_2_1_Adder_7_U.u1.s ;
wire [5:0] \add_11ns_11s_11_2_1_U21.top_add_11ns_11s_11_2_1_Adder_7_U.u2.a ;
wire [5:0] \add_11ns_11s_11_2_1_U21.top_add_11ns_11s_11_2_1_Adder_7_U.u2.b ;
wire \add_11ns_11s_11_2_1_U21.top_add_11ns_11s_11_2_1_Adder_7_U.u2.cin ;
wire \add_11ns_11s_11_2_1_U21.top_add_11ns_11s_11_2_1_Adder_7_U.u2.cout ;
wire [5:0] \add_11ns_11s_11_2_1_U21.top_add_11ns_11s_11_2_1_Adder_7_U.u2.s ;
wire \add_11s_11ns_11_2_1_U13.ce ;
wire \add_11s_11ns_11_2_1_U13.clk ;
wire [10:0] \add_11s_11ns_11_2_1_U13.din0 ;
wire [10:0] \add_11s_11ns_11_2_1_U13.din1 ;
wire [10:0] \add_11s_11ns_11_2_1_U13.dout ;
wire \add_11s_11ns_11_2_1_U13.reset ;
wire [10:0] \add_11s_11ns_11_2_1_U13.top_add_11s_11ns_11_2_1_Adder_4_U.a ;
wire [10:0] \add_11s_11ns_11_2_1_U13.top_add_11s_11ns_11_2_1_Adder_4_U.ain_s0 ;
wire [10:0] \add_11s_11ns_11_2_1_U13.top_add_11s_11ns_11_2_1_Adder_4_U.b ;
wire [10:0] \add_11s_11ns_11_2_1_U13.top_add_11s_11ns_11_2_1_Adder_4_U.bin_s0 ;
wire \add_11s_11ns_11_2_1_U13.top_add_11s_11ns_11_2_1_Adder_4_U.ce ;
wire \add_11s_11ns_11_2_1_U13.top_add_11s_11ns_11_2_1_Adder_4_U.clk ;
wire \add_11s_11ns_11_2_1_U13.top_add_11s_11ns_11_2_1_Adder_4_U.facout_s1 ;
wire \add_11s_11ns_11_2_1_U13.top_add_11s_11ns_11_2_1_Adder_4_U.facout_s2 ;
wire [4:0] \add_11s_11ns_11_2_1_U13.top_add_11s_11ns_11_2_1_Adder_4_U.fas_s1 ;
wire [5:0] \add_11s_11ns_11_2_1_U13.top_add_11s_11ns_11_2_1_Adder_4_U.fas_s2 ;
wire \add_11s_11ns_11_2_1_U13.top_add_11s_11ns_11_2_1_Adder_4_U.reset ;
wire [10:0] \add_11s_11ns_11_2_1_U13.top_add_11s_11ns_11_2_1_Adder_4_U.s ;
wire [4:0] \add_11s_11ns_11_2_1_U13.top_add_11s_11ns_11_2_1_Adder_4_U.u1.a ;
wire [4:0] \add_11s_11ns_11_2_1_U13.top_add_11s_11ns_11_2_1_Adder_4_U.u1.b ;
wire \add_11s_11ns_11_2_1_U13.top_add_11s_11ns_11_2_1_Adder_4_U.u1.cin ;
wire \add_11s_11ns_11_2_1_U13.top_add_11s_11ns_11_2_1_Adder_4_U.u1.cout ;
wire [4:0] \add_11s_11ns_11_2_1_U13.top_add_11s_11ns_11_2_1_Adder_4_U.u1.s ;
wire [5:0] \add_11s_11ns_11_2_1_U13.top_add_11s_11ns_11_2_1_Adder_4_U.u2.a ;
wire [5:0] \add_11s_11ns_11_2_1_U13.top_add_11s_11ns_11_2_1_Adder_4_U.u2.b ;
wire \add_11s_11ns_11_2_1_U13.top_add_11s_11ns_11_2_1_Adder_4_U.u2.cin ;
wire \add_11s_11ns_11_2_1_U13.top_add_11s_11ns_11_2_1_Adder_4_U.u2.cout ;
wire [5:0] \add_11s_11ns_11_2_1_U13.top_add_11s_11ns_11_2_1_Adder_4_U.u2.s ;
wire \add_11s_11ns_11_2_1_U6.ce ;
wire \add_11s_11ns_11_2_1_U6.clk ;
wire [10:0] \add_11s_11ns_11_2_1_U6.din0 ;
wire [10:0] \add_11s_11ns_11_2_1_U6.din1 ;
wire [10:0] \add_11s_11ns_11_2_1_U6.dout ;
wire \add_11s_11ns_11_2_1_U6.reset ;
wire [10:0] \add_11s_11ns_11_2_1_U6.top_add_11s_11ns_11_2_1_Adder_4_U.a ;
wire [10:0] \add_11s_11ns_11_2_1_U6.top_add_11s_11ns_11_2_1_Adder_4_U.ain_s0 ;
wire [10:0] \add_11s_11ns_11_2_1_U6.top_add_11s_11ns_11_2_1_Adder_4_U.b ;
wire [10:0] \add_11s_11ns_11_2_1_U6.top_add_11s_11ns_11_2_1_Adder_4_U.bin_s0 ;
wire \add_11s_11ns_11_2_1_U6.top_add_11s_11ns_11_2_1_Adder_4_U.ce ;
wire \add_11s_11ns_11_2_1_U6.top_add_11s_11ns_11_2_1_Adder_4_U.clk ;
wire \add_11s_11ns_11_2_1_U6.top_add_11s_11ns_11_2_1_Adder_4_U.facout_s1 ;
wire \add_11s_11ns_11_2_1_U6.top_add_11s_11ns_11_2_1_Adder_4_U.facout_s2 ;
wire [4:0] \add_11s_11ns_11_2_1_U6.top_add_11s_11ns_11_2_1_Adder_4_U.fas_s1 ;
wire [5:0] \add_11s_11ns_11_2_1_U6.top_add_11s_11ns_11_2_1_Adder_4_U.fas_s2 ;
wire \add_11s_11ns_11_2_1_U6.top_add_11s_11ns_11_2_1_Adder_4_U.reset ;
wire [10:0] \add_11s_11ns_11_2_1_U6.top_add_11s_11ns_11_2_1_Adder_4_U.s ;
wire [4:0] \add_11s_11ns_11_2_1_U6.top_add_11s_11ns_11_2_1_Adder_4_U.u1.a ;
wire [4:0] \add_11s_11ns_11_2_1_U6.top_add_11s_11ns_11_2_1_Adder_4_U.u1.b ;
wire \add_11s_11ns_11_2_1_U6.top_add_11s_11ns_11_2_1_Adder_4_U.u1.cin ;
wire \add_11s_11ns_11_2_1_U6.top_add_11s_11ns_11_2_1_Adder_4_U.u1.cout ;
wire [4:0] \add_11s_11ns_11_2_1_U6.top_add_11s_11ns_11_2_1_Adder_4_U.u1.s ;
wire [5:0] \add_11s_11ns_11_2_1_U6.top_add_11s_11ns_11_2_1_Adder_4_U.u2.a ;
wire [5:0] \add_11s_11ns_11_2_1_U6.top_add_11s_11ns_11_2_1_Adder_4_U.u2.b ;
wire \add_11s_11ns_11_2_1_U6.top_add_11s_11ns_11_2_1_Adder_4_U.u2.cin ;
wire \add_11s_11ns_11_2_1_U6.top_add_11s_11ns_11_2_1_Adder_4_U.u2.cout ;
wire [5:0] \add_11s_11ns_11_2_1_U6.top_add_11s_11ns_11_2_1_Adder_4_U.u2.s ;
wire \add_12ns_12s_12_2_1_U1.ce ;
wire \add_12ns_12s_12_2_1_U1.clk ;
wire [11:0] \add_12ns_12s_12_2_1_U1.din0 ;
wire [11:0] \add_12ns_12s_12_2_1_U1.din1 ;
wire [11:0] \add_12ns_12s_12_2_1_U1.dout ;
wire \add_12ns_12s_12_2_1_U1.reset ;
wire [11:0] \add_12ns_12s_12_2_1_U1.top_add_12ns_12s_12_2_1_Adder_0_U.a ;
wire [11:0] \add_12ns_12s_12_2_1_U1.top_add_12ns_12s_12_2_1_Adder_0_U.ain_s0 ;
wire [11:0] \add_12ns_12s_12_2_1_U1.top_add_12ns_12s_12_2_1_Adder_0_U.b ;
wire [11:0] \add_12ns_12s_12_2_1_U1.top_add_12ns_12s_12_2_1_Adder_0_U.bin_s0 ;
wire \add_12ns_12s_12_2_1_U1.top_add_12ns_12s_12_2_1_Adder_0_U.ce ;
wire \add_12ns_12s_12_2_1_U1.top_add_12ns_12s_12_2_1_Adder_0_U.clk ;
wire \add_12ns_12s_12_2_1_U1.top_add_12ns_12s_12_2_1_Adder_0_U.facout_s1 ;
wire \add_12ns_12s_12_2_1_U1.top_add_12ns_12s_12_2_1_Adder_0_U.facout_s2 ;
wire [5:0] \add_12ns_12s_12_2_1_U1.top_add_12ns_12s_12_2_1_Adder_0_U.fas_s1 ;
wire [5:0] \add_12ns_12s_12_2_1_U1.top_add_12ns_12s_12_2_1_Adder_0_U.fas_s2 ;
wire \add_12ns_12s_12_2_1_U1.top_add_12ns_12s_12_2_1_Adder_0_U.reset ;
wire [11:0] \add_12ns_12s_12_2_1_U1.top_add_12ns_12s_12_2_1_Adder_0_U.s ;
wire [5:0] \add_12ns_12s_12_2_1_U1.top_add_12ns_12s_12_2_1_Adder_0_U.u1.a ;
wire [5:0] \add_12ns_12s_12_2_1_U1.top_add_12ns_12s_12_2_1_Adder_0_U.u1.b ;
wire \add_12ns_12s_12_2_1_U1.top_add_12ns_12s_12_2_1_Adder_0_U.u1.cin ;
wire \add_12ns_12s_12_2_1_U1.top_add_12ns_12s_12_2_1_Adder_0_U.u1.cout ;
wire [5:0] \add_12ns_12s_12_2_1_U1.top_add_12ns_12s_12_2_1_Adder_0_U.u1.s ;
wire [5:0] \add_12ns_12s_12_2_1_U1.top_add_12ns_12s_12_2_1_Adder_0_U.u2.a ;
wire [5:0] \add_12ns_12s_12_2_1_U1.top_add_12ns_12s_12_2_1_Adder_0_U.u2.b ;
wire \add_12ns_12s_12_2_1_U1.top_add_12ns_12s_12_2_1_Adder_0_U.u2.cin ;
wire \add_12ns_12s_12_2_1_U1.top_add_12ns_12s_12_2_1_Adder_0_U.u2.cout ;
wire [5:0] \add_12ns_12s_12_2_1_U1.top_add_12ns_12s_12_2_1_Adder_0_U.u2.s ;
wire \add_2ns_2ns_2_2_1_U5.ce ;
wire \add_2ns_2ns_2_2_1_U5.clk ;
wire [1:0] \add_2ns_2ns_2_2_1_U5.din0 ;
wire [1:0] \add_2ns_2ns_2_2_1_U5.din1 ;
wire [1:0] \add_2ns_2ns_2_2_1_U5.dout ;
wire \add_2ns_2ns_2_2_1_U5.reset ;
wire [1:0] \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_3_U.a ;
wire [1:0] \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_3_U.ain_s0 ;
wire [1:0] \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_3_U.b ;
wire [1:0] \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_3_U.bin_s0 ;
wire \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_3_U.ce ;
wire \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_3_U.clk ;
wire \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_3_U.facout_s1 ;
wire \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_3_U.facout_s2 ;
wire \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_3_U.fas_s1 ;
wire \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_3_U.fas_s2 ;
wire \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_3_U.reset ;
wire [1:0] \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_3_U.s ;
wire \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_3_U.u1.a ;
wire \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_3_U.u1.b ;
wire \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_3_U.u1.cin ;
wire \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_3_U.u1.cout ;
wire \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_3_U.u1.s ;
wire \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_3_U.u2.a ;
wire \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_3_U.u2.b ;
wire \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_3_U.u2.cin ;
wire \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_3_U.u2.cout ;
wire \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_3_U.u2.s ;
wire \add_32ns_32ns_32_2_1_U23.ce ;
wire \add_32ns_32ns_32_2_1_U23.clk ;
wire [31:0] \add_32ns_32ns_32_2_1_U23.din0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U23.din1 ;
wire [31:0] \add_32ns_32ns_32_2_1_U23.dout ;
wire \add_32ns_32ns_32_2_1_U23.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_13_U.a ;
wire [31:0] \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_13_U.ain_s0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_13_U.b ;
wire [31:0] \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_13_U.bin_s0 ;
wire \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_13_U.ce ;
wire \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_13_U.clk ;
wire \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_13_U.facout_s1 ;
wire \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_13_U.facout_s2 ;
wire [15:0] \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_13_U.fas_s1 ;
wire [15:0] \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_13_U.fas_s2 ;
wire \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_13_U.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_13_U.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_13_U.u1.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_13_U.u1.b ;
wire \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_13_U.u1.cin ;
wire \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_13_U.u1.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_13_U.u1.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_13_U.u2.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_13_U.u2.b ;
wire \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_13_U.u2.cin ;
wire \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_13_U.u2.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_13_U.u2.s ;
wire \add_35s_35s_35_2_1_U22.ce ;
wire \add_35s_35s_35_2_1_U22.clk ;
wire [34:0] \add_35s_35s_35_2_1_U22.din0 ;
wire [34:0] \add_35s_35s_35_2_1_U22.din1 ;
wire [34:0] \add_35s_35s_35_2_1_U22.dout ;
wire \add_35s_35s_35_2_1_U22.reset ;
wire [34:0] \add_35s_35s_35_2_1_U22.top_add_35s_35s_35_2_1_Adder_12_U.a ;
wire [34:0] \add_35s_35s_35_2_1_U22.top_add_35s_35s_35_2_1_Adder_12_U.ain_s0 ;
wire [34:0] \add_35s_35s_35_2_1_U22.top_add_35s_35s_35_2_1_Adder_12_U.b ;
wire [34:0] \add_35s_35s_35_2_1_U22.top_add_35s_35s_35_2_1_Adder_12_U.bin_s0 ;
wire \add_35s_35s_35_2_1_U22.top_add_35s_35s_35_2_1_Adder_12_U.ce ;
wire \add_35s_35s_35_2_1_U22.top_add_35s_35s_35_2_1_Adder_12_U.clk ;
wire \add_35s_35s_35_2_1_U22.top_add_35s_35s_35_2_1_Adder_12_U.facout_s1 ;
wire \add_35s_35s_35_2_1_U22.top_add_35s_35s_35_2_1_Adder_12_U.facout_s2 ;
wire [16:0] \add_35s_35s_35_2_1_U22.top_add_35s_35s_35_2_1_Adder_12_U.fas_s1 ;
wire [17:0] \add_35s_35s_35_2_1_U22.top_add_35s_35s_35_2_1_Adder_12_U.fas_s2 ;
wire \add_35s_35s_35_2_1_U22.top_add_35s_35s_35_2_1_Adder_12_U.reset ;
wire [34:0] \add_35s_35s_35_2_1_U22.top_add_35s_35s_35_2_1_Adder_12_U.s ;
wire [16:0] \add_35s_35s_35_2_1_U22.top_add_35s_35s_35_2_1_Adder_12_U.u1.a ;
wire [16:0] \add_35s_35s_35_2_1_U22.top_add_35s_35s_35_2_1_Adder_12_U.u1.b ;
wire \add_35s_35s_35_2_1_U22.top_add_35s_35s_35_2_1_Adder_12_U.u1.cin ;
wire \add_35s_35s_35_2_1_U22.top_add_35s_35s_35_2_1_Adder_12_U.u1.cout ;
wire [16:0] \add_35s_35s_35_2_1_U22.top_add_35s_35s_35_2_1_Adder_12_U.u1.s ;
wire [17:0] \add_35s_35s_35_2_1_U22.top_add_35s_35s_35_2_1_Adder_12_U.u2.a ;
wire [17:0] \add_35s_35s_35_2_1_U22.top_add_35s_35s_35_2_1_Adder_12_U.u2.b ;
wire \add_35s_35s_35_2_1_U22.top_add_35s_35s_35_2_1_Adder_12_U.u2.cin ;
wire \add_35s_35s_35_2_1_U22.top_add_35s_35s_35_2_1_Adder_12_U.u2.cout ;
wire [17:0] \add_35s_35s_35_2_1_U22.top_add_35s_35s_35_2_1_Adder_12_U.u2.s ;
wire \add_3ns_3ns_3_2_1_U15.ce ;
wire \add_3ns_3ns_3_2_1_U15.clk ;
wire [2:0] \add_3ns_3ns_3_2_1_U15.din0 ;
wire [2:0] \add_3ns_3ns_3_2_1_U15.din1 ;
wire [2:0] \add_3ns_3ns_3_2_1_U15.dout ;
wire \add_3ns_3ns_3_2_1_U15.reset ;
wire [2:0] \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_10_U.a ;
wire [2:0] \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_10_U.ain_s0 ;
wire [2:0] \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_10_U.b ;
wire [2:0] \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_10_U.bin_s0 ;
wire \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_10_U.ce ;
wire \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_10_U.clk ;
wire \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_10_U.facout_s1 ;
wire \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_10_U.facout_s2 ;
wire \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_10_U.fas_s1 ;
wire [1:0] \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_10_U.fas_s2 ;
wire \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_10_U.reset ;
wire [2:0] \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_10_U.s ;
wire \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_10_U.u1.a ;
wire \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_10_U.u1.b ;
wire \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_10_U.u1.cin ;
wire \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_10_U.u1.cout ;
wire \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_10_U.u1.s ;
wire [1:0] \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_10_U.u2.a ;
wire [1:0] \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_10_U.u2.b ;
wire \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_10_U.u2.cin ;
wire \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_10_U.u2.cout ;
wire [1:0] \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_10_U.u2.s ;
wire \add_3s_3ns_3_2_1_U10.ce ;
wire \add_3s_3ns_3_2_1_U10.clk ;
wire [2:0] \add_3s_3ns_3_2_1_U10.din0 ;
wire [2:0] \add_3s_3ns_3_2_1_U10.din1 ;
wire [2:0] \add_3s_3ns_3_2_1_U10.dout ;
wire \add_3s_3ns_3_2_1_U10.reset ;
wire [2:0] \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.a ;
wire [2:0] \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.ain_s0 ;
wire [2:0] \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.b ;
wire [2:0] \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.bin_s0 ;
wire \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.ce ;
wire \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.clk ;
wire \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.facout_s1 ;
wire \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.facout_s2 ;
wire \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.fas_s1 ;
wire [1:0] \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.fas_s2 ;
wire \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.reset ;
wire [2:0] \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.s ;
wire \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.u1.a ;
wire \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.u1.b ;
wire \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.u1.cin ;
wire \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.u1.cout ;
wire \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.u1.s ;
wire [1:0] \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.u2.a ;
wire [1:0] \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.u2.b ;
wire \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.u2.cin ;
wire \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.u2.cout ;
wire [1:0] \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.u2.s ;
wire \add_3s_3s_3_2_1_U9.ce ;
wire \add_3s_3s_3_2_1_U9.clk ;
wire [2:0] \add_3s_3s_3_2_1_U9.din0 ;
wire [2:0] \add_3s_3s_3_2_1_U9.din1 ;
wire [2:0] \add_3s_3s_3_2_1_U9.dout ;
wire \add_3s_3s_3_2_1_U9.reset ;
wire [2:0] \add_3s_3s_3_2_1_U9.top_add_3s_3s_3_2_1_Adder_5_U.a ;
wire [2:0] \add_3s_3s_3_2_1_U9.top_add_3s_3s_3_2_1_Adder_5_U.ain_s0 ;
wire [2:0] \add_3s_3s_3_2_1_U9.top_add_3s_3s_3_2_1_Adder_5_U.b ;
wire [2:0] \add_3s_3s_3_2_1_U9.top_add_3s_3s_3_2_1_Adder_5_U.bin_s0 ;
wire \add_3s_3s_3_2_1_U9.top_add_3s_3s_3_2_1_Adder_5_U.ce ;
wire \add_3s_3s_3_2_1_U9.top_add_3s_3s_3_2_1_Adder_5_U.clk ;
wire \add_3s_3s_3_2_1_U9.top_add_3s_3s_3_2_1_Adder_5_U.facout_s1 ;
wire \add_3s_3s_3_2_1_U9.top_add_3s_3s_3_2_1_Adder_5_U.facout_s2 ;
wire \add_3s_3s_3_2_1_U9.top_add_3s_3s_3_2_1_Adder_5_U.fas_s1 ;
wire [1:0] \add_3s_3s_3_2_1_U9.top_add_3s_3s_3_2_1_Adder_5_U.fas_s2 ;
wire \add_3s_3s_3_2_1_U9.top_add_3s_3s_3_2_1_Adder_5_U.reset ;
wire [2:0] \add_3s_3s_3_2_1_U9.top_add_3s_3s_3_2_1_Adder_5_U.s ;
wire \add_3s_3s_3_2_1_U9.top_add_3s_3s_3_2_1_Adder_5_U.u1.a ;
wire \add_3s_3s_3_2_1_U9.top_add_3s_3s_3_2_1_Adder_5_U.u1.b ;
wire \add_3s_3s_3_2_1_U9.top_add_3s_3s_3_2_1_Adder_5_U.u1.cin ;
wire \add_3s_3s_3_2_1_U9.top_add_3s_3s_3_2_1_Adder_5_U.u1.cout ;
wire \add_3s_3s_3_2_1_U9.top_add_3s_3s_3_2_1_Adder_5_U.u1.s ;
wire [1:0] \add_3s_3s_3_2_1_U9.top_add_3s_3s_3_2_1_Adder_5_U.u2.a ;
wire [1:0] \add_3s_3s_3_2_1_U9.top_add_3s_3s_3_2_1_Adder_5_U.u2.b ;
wire \add_3s_3s_3_2_1_U9.top_add_3s_3s_3_2_1_Adder_5_U.u2.cin ;
wire \add_3s_3s_3_2_1_U9.top_add_3s_3s_3_2_1_Adder_5_U.u2.cout ;
wire [1:0] \add_3s_3s_3_2_1_U9.top_add_3s_3s_3_2_1_Adder_5_U.u2.s ;
wire \add_6s_6ns_6_2_1_U12.ce ;
wire \add_6s_6ns_6_2_1_U12.clk ;
wire [5:0] \add_6s_6ns_6_2_1_U12.din0 ;
wire [5:0] \add_6s_6ns_6_2_1_U12.din1 ;
wire [5:0] \add_6s_6ns_6_2_1_U12.dout ;
wire \add_6s_6ns_6_2_1_U12.reset ;
wire [5:0] \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_8_U.a ;
wire [5:0] \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_8_U.ain_s0 ;
wire [5:0] \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_8_U.b ;
wire [5:0] \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_8_U.bin_s0 ;
wire \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_8_U.ce ;
wire \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_8_U.clk ;
wire \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_8_U.facout_s1 ;
wire \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_8_U.facout_s2 ;
wire [2:0] \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_8_U.fas_s1 ;
wire [2:0] \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_8_U.fas_s2 ;
wire \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_8_U.reset ;
wire [5:0] \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_8_U.s ;
wire [2:0] \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_8_U.u1.a ;
wire [2:0] \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_8_U.u1.b ;
wire \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_8_U.u1.cin ;
wire \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_8_U.u1.cout ;
wire [2:0] \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_8_U.u1.s ;
wire [2:0] \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_8_U.u2.a ;
wire [2:0] \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_8_U.u2.b ;
wire \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_8_U.u2.cin ;
wire \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_8_U.u2.cout ;
wire [2:0] \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_8_U.u2.s ;
wire ap_CS_fsm_state1;
wire ap_CS_fsm_state10;
wire ap_CS_fsm_state11;
wire ap_CS_fsm_state12;
wire ap_CS_fsm_state13;
wire ap_CS_fsm_state14;
wire ap_CS_fsm_state15;
wire ap_CS_fsm_state16;
wire ap_CS_fsm_state17;
wire ap_CS_fsm_state18;
wire ap_CS_fsm_state19;
wire ap_CS_fsm_state2;
wire ap_CS_fsm_state20;
wire ap_CS_fsm_state21;
wire ap_CS_fsm_state22;
wire ap_CS_fsm_state23;
wire ap_CS_fsm_state29;
wire ap_CS_fsm_state3;
wire ap_CS_fsm_state30;
wire ap_CS_fsm_state31;
wire ap_CS_fsm_state32;
wire ap_CS_fsm_state33;
wire ap_CS_fsm_state34;
wire ap_CS_fsm_state35;
wire ap_CS_fsm_state36;
wire ap_CS_fsm_state37;
wire ap_CS_fsm_state4;
wire ap_CS_fsm_state5;
wire ap_CS_fsm_state6;
wire ap_CS_fsm_state7;
wire ap_CS_fsm_state8;
wire ap_CS_fsm_state9;
wire [36:0] ap_NS_fsm;
wire ap_clk;
wire ap_done;
wire ap_idle;
wire ap_ready;
wire ap_rst;
wire ap_start;
wire \ashr_32s_16ns_32_7_1_U18.ce ;
wire \ashr_32s_16ns_32_7_1_U18.clk ;
wire [31:0] \ashr_32s_16ns_32_7_1_U18.din0 ;
wire [31:0] \ashr_32s_16ns_32_7_1_U18.din1 ;
wire [15:0] \ashr_32s_16ns_32_7_1_U18.din1_cast ;
wire [15:0] \ashr_32s_16ns_32_7_1_U18.din1_mask ;
wire [31:0] \ashr_32s_16ns_32_7_1_U18.dout ;
wire \ashr_32s_16ns_32_7_1_U18.reset ;
wire \ashr_32s_32s_32_7_1_U8.ce ;
wire \ashr_32s_32s_32_7_1_U8.clk ;
wire [31:0] \ashr_32s_32s_32_7_1_U8.din0 ;
wire [31:0] \ashr_32s_32s_32_7_1_U8.din1 ;
wire [31:0] \ashr_32s_32s_32_7_1_U8.din1_cast ;
wire [31:0] \ashr_32s_32s_32_7_1_U8.din1_mask ;
wire [31:0] \ashr_32s_32s_32_7_1_U8.dout ;
wire \ashr_32s_32s_32_7_1_U8.reset ;
wire [3:0] conv_i_i_i329_fu_386_p0;
wire [31:0] conv_i_i_i329_fu_386_p1;
wire [11:0] grp_fu_189_p0;
wire [11:0] grp_fu_189_p1;
wire [11:0] grp_fu_189_p2;
wire [31:0] grp_fu_213_p0;
wire [31:0] grp_fu_213_p1;
wire [31:0] grp_fu_213_p2;
wire [9:0] grp_fu_239_p2;
wire [4:0] grp_fu_296_p1;
wire [4:0] grp_fu_296_p2;
wire [1:0] grp_fu_307_p2;
wire [10:0] grp_fu_377_p0;
wire [10:0] grp_fu_377_p2;
wire [31:0] grp_fu_390_p2;
wire [31:0] grp_fu_396_p2;
wire [2:0] grp_fu_409_p0;
wire [2:0] grp_fu_409_p1;
wire [2:0] grp_fu_409_p2;
wire [2:0] grp_fu_422_p0;
wire [2:0] grp_fu_422_p1;
wire [2:0] grp_fu_422_p2;
wire [10:0] grp_fu_454_p1;
wire [10:0] grp_fu_454_p2;
wire [5:0] grp_fu_462_p0;
wire [5:0] grp_fu_462_p1;
wire [5:0] grp_fu_462_p2;
wire [10:0] grp_fu_471_p0;
wire [10:0] grp_fu_471_p2;
wire [10:0] grp_fu_499_p2;
wire [2:0] grp_fu_503_p2;
wire [10:0] grp_fu_508_p2;
wire [3:0] grp_fu_547_p1;
wire [3:0] grp_fu_547_p2;
wire [31:0] grp_fu_582_p1;
wire [31:0] grp_fu_582_p2;
wire [31:0] grp_fu_595_p1;
wire [31:0] grp_fu_595_p2;
wire [10:0] grp_fu_613_p1;
wire [10:0] grp_fu_613_p2;
wire [10:0] grp_fu_630_p1;
wire [10:0] grp_fu_630_p2;
wire [34:0] grp_fu_650_p0;
wire [34:0] grp_fu_650_p1;
wire [34:0] grp_fu_650_p2;
wire [31:0] grp_fu_676_p2;
wire icmp_ln1499_fu_219_p2;
wire icmp_ln851_1_fu_302_p2;
wire icmp_ln851_2_fu_372_p2;
wire icmp_ln851_3_fu_660_p2;
wire icmp_ln851_fu_199_p2;
wire [11:0] lhs_V_1_fu_312_p3;
wire [3:0] lhs_V_2_fu_363_p0;
wire lhs_V_2_fu_363_p2;
wire [1:0] op_0;
wire [3:0] op_1;
wire [1:0] op_12;
wire op_14;
wire [3:0] op_16;
wire [3:0] op_18;
wire [7:0] op_2;
wire [31:0] op_30;
wire op_30_ap_vld;
wire [3:0] op_5;
wire [3:0] op_7_V_fu_267_p2;
wire [3:0] op_8;
wire p_Result_1_fu_344_p3;
wire p_Result_3_fu_428_p3;
wire p_Result_4_fu_513_p3;
wire p_Result_6_fu_553_p3;
wire p_Result_7_fu_681_p3;
wire p_Result_s_fu_244_p3;
wire [5:0] r_fu_621_p3;
wire [9:0] ret_V_20_fu_256_p3;
wire [1:0] ret_V_21_fu_356_p3;
wire [11:0] ret_V_22_fu_319_p2;
wire [10:0] ret_V_23_fu_440_p3;
wire [2:0] ret_V_24_fu_529_p3;
wire [10:0] ret_V_26_fu_565_p3;
wire [9:0] rhs_fu_177_p3;
wire [10:0] select_ln1192_fu_476_p3;
wire [31:0] select_ln1368_fu_484_p3;
wire [1:0] select_ln850_1_fu_351_p3;
wire [10:0] select_ln850_2_fu_435_p3;
wire [2:0] select_ln850_3_fu_523_p3;
wire [10:0] select_ln850_4_fu_560_p3;
wire [31:0] select_ln850_5_fu_688_p3;
wire [9:0] select_ln850_fu_251_p3;
wire [3:0] sext_ln1299_fu_209_p0;
wire [31:0] sext_ln1367_fu_383_p1;
wire [4:0] sext_ln1386_fu_293_p1;
wire [5:0] sext_ln546_1_fu_618_p1;
wire [15:0] sext_ln546_2_fu_588_p1;
wire [15:0] sext_ln546_fu_575_p1;
wire [3:0] sext_ln703_1_fu_635_p0;
wire [3:0] sext_ln703_fu_173_p0;
wire [31:0] sext_ln781_fu_572_p1;
wire [10:0] sext_ln831_fu_369_p1;
wire \shl_32s_16ns_32_7_1_U19.ce ;
wire \shl_32s_16ns_32_7_1_U19.clk ;
wire [31:0] \shl_32s_16ns_32_7_1_U19.din0 ;
wire [31:0] \shl_32s_16ns_32_7_1_U19.din1 ;
wire [15:0] \shl_32s_16ns_32_7_1_U19.din1_cast ;
wire [15:0] \shl_32s_16ns_32_7_1_U19.din1_mask ;
wire [31:0] \shl_32s_16ns_32_7_1_U19.dout ;
wire \shl_32s_16ns_32_7_1_U19.reset ;
wire \shl_32s_32s_32_7_1_U7.ce ;
wire \shl_32s_32s_32_7_1_U7.clk ;
wire [31:0] \shl_32s_32s_32_7_1_U7.din0 ;
wire [31:0] \shl_32s_32s_32_7_1_U7.din1 ;
wire [31:0] \shl_32s_32s_32_7_1_U7.din1_cast ;
wire [31:0] \shl_32s_32s_32_7_1_U7.din1_mask ;
wire [31:0] \shl_32s_32s_32_7_1_U7.dout ;
wire \shl_32s_32s_32_7_1_U7.reset ;
wire \shl_32s_8ns_32_7_1_U2.ce ;
wire \shl_32s_8ns_32_7_1_U2.clk ;
wire [31:0] \shl_32s_8ns_32_7_1_U2.din0 ;
wire [31:0] \shl_32s_8ns_32_7_1_U2.din1 ;
wire [7:0] \shl_32s_8ns_32_7_1_U2.din1_cast ;
wire [7:0] \shl_32s_8ns_32_7_1_U2.din1_mask ;
wire [31:0] \shl_32s_8ns_32_7_1_U2.dout ;
wire \shl_32s_8ns_32_7_1_U2.reset ;
wire \sub_4ns_4s_4_2_1_U17.ce ;
wire \sub_4ns_4s_4_2_1_U17.clk ;
wire [3:0] \sub_4ns_4s_4_2_1_U17.din0 ;
wire [3:0] \sub_4ns_4s_4_2_1_U17.din1 ;
wire [3:0] \sub_4ns_4s_4_2_1_U17.dout ;
wire \sub_4ns_4s_4_2_1_U17.reset ;
wire [3:0] \sub_4ns_4s_4_2_1_U17.top_sub_4ns_4s_4_2_1_Adder_11_U.a ;
wire [3:0] \sub_4ns_4s_4_2_1_U17.top_sub_4ns_4s_4_2_1_Adder_11_U.ain_s0 ;
wire [3:0] \sub_4ns_4s_4_2_1_U17.top_sub_4ns_4s_4_2_1_Adder_11_U.b ;
wire [3:0] \sub_4ns_4s_4_2_1_U17.top_sub_4ns_4s_4_2_1_Adder_11_U.bin_s0 ;
wire \sub_4ns_4s_4_2_1_U17.top_sub_4ns_4s_4_2_1_Adder_11_U.ce ;
wire \sub_4ns_4s_4_2_1_U17.top_sub_4ns_4s_4_2_1_Adder_11_U.clk ;
wire \sub_4ns_4s_4_2_1_U17.top_sub_4ns_4s_4_2_1_Adder_11_U.facout_s1 ;
wire \sub_4ns_4s_4_2_1_U17.top_sub_4ns_4s_4_2_1_Adder_11_U.facout_s2 ;
wire [1:0] \sub_4ns_4s_4_2_1_U17.top_sub_4ns_4s_4_2_1_Adder_11_U.fas_s1 ;
wire [1:0] \sub_4ns_4s_4_2_1_U17.top_sub_4ns_4s_4_2_1_Adder_11_U.fas_s2 ;
wire \sub_4ns_4s_4_2_1_U17.top_sub_4ns_4s_4_2_1_Adder_11_U.reset ;
wire [3:0] \sub_4ns_4s_4_2_1_U17.top_sub_4ns_4s_4_2_1_Adder_11_U.s ;
wire [1:0] \sub_4ns_4s_4_2_1_U17.top_sub_4ns_4s_4_2_1_Adder_11_U.u1.a ;
wire [1:0] \sub_4ns_4s_4_2_1_U17.top_sub_4ns_4s_4_2_1_Adder_11_U.u1.b ;
wire \sub_4ns_4s_4_2_1_U17.top_sub_4ns_4s_4_2_1_Adder_11_U.u1.cin ;
wire \sub_4ns_4s_4_2_1_U17.top_sub_4ns_4s_4_2_1_Adder_11_U.u1.cout ;
wire [1:0] \sub_4ns_4s_4_2_1_U17.top_sub_4ns_4s_4_2_1_Adder_11_U.u1.s ;
wire [1:0] \sub_4ns_4s_4_2_1_U17.top_sub_4ns_4s_4_2_1_Adder_11_U.u2.a ;
wire [1:0] \sub_4ns_4s_4_2_1_U17.top_sub_4ns_4s_4_2_1_Adder_11_U.u2.b ;
wire \sub_4ns_4s_4_2_1_U17.top_sub_4ns_4s_4_2_1_Adder_11_U.u2.cin ;
wire \sub_4ns_4s_4_2_1_U17.top_sub_4ns_4s_4_2_1_Adder_11_U.u2.cout ;
wire [1:0] \sub_4ns_4s_4_2_1_U17.top_sub_4ns_4s_4_2_1_Adder_11_U.u2.s ;
wire \sub_5ns_5s_5_2_1_U4.ce ;
wire \sub_5ns_5s_5_2_1_U4.clk ;
wire [4:0] \sub_5ns_5s_5_2_1_U4.din0 ;
wire [4:0] \sub_5ns_5s_5_2_1_U4.din1 ;
wire [4:0] \sub_5ns_5s_5_2_1_U4.dout ;
wire \sub_5ns_5s_5_2_1_U4.reset ;
wire [4:0] \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.a ;
wire [4:0] \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.ain_s0 ;
wire [4:0] \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.b ;
wire [4:0] \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.bin_s0 ;
wire \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.ce ;
wire \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.clk ;
wire \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.facout_s1 ;
wire \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.facout_s2 ;
wire [1:0] \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.fas_s1 ;
wire [2:0] \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.fas_s2 ;
wire \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.reset ;
wire [4:0] \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.s ;
wire [1:0] \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.u1.a ;
wire [1:0] \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.u1.b ;
wire \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.u1.cin ;
wire \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.u1.cout ;
wire [1:0] \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.u1.s ;
wire [2:0] \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.u2.a ;
wire [2:0] \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.u2.b ;
wire \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.u2.cin ;
wire \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.u2.cout ;
wire [2:0] \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.u2.s ;
wire [12:0] tmp_fu_639_p3;
wire [3:0] trunc_ln1348_1_fu_225_p1;
wire [3:0] trunc_ln1348_fu_263_p1;
wire [2:0] trunc_ln546_fu_601_p1;
wire [5:0] trunc_ln769_fu_605_p1;
wire [1:0] trunc_ln851_1_fu_289_p1;
wire [1:0] trunc_ln851_2_fu_335_p1;
wire trunc_ln851_3_fu_520_p1;
wire [3:0] trunc_ln851_4_fu_656_p0;
wire [1:0] trunc_ln851_4_fu_656_p1;
wire [3:0] trunc_ln851_fu_195_p0;
wire [1:0] trunc_ln851_fu_195_p1;
wire [4:0] ush_fu_339_p3;


assign _054_ = icmp_ln851_3_reg_1071 & ap_CS_fsm[35];
assign _055_ = ap_CS_fsm[19] & lhs_V_2_reg_833;
assign _056_ = ap_CS_fsm[15] & _065_;
assign _057_ = _066_ & ap_CS_fsm[3];
assign _058_ = p_Result_8_reg_985 & ap_CS_fsm[21];
assign _059_ = ap_CS_fsm[15] & isNeg_reg_769;
assign _060_ = ap_CS_fsm[7] & isNeg_reg_769;
assign _061_ = p_Result_8_reg_985 & ap_CS_fsm[28];
assign _062_ = _067_ & ap_CS_fsm[28];
assign _063_ = _068_ & ap_CS_fsm[0];
assign _064_ = ap_start & ap_CS_fsm[0];
assign op_7_V_fu_267_p2 = trunc_ln1348_reg_759 & trunc_ln1348_1_reg_731;
assign ret_V_22_fu_319_p2[2] = ~ ret_V_20_reg_753[0];
assign _065_ = ~ isNeg_reg_769;
assign _066_ = ~ icmp_ln851_reg_711;
assign _067_ = ~ p_Result_8_reg_985;
assign _068_ = ~ ap_start;
assign _069_ = ! trunc_ln851_1_reg_787;
assign _070_ = ! trunc_ln851_2_reg_818;
assign _071_ = ! op_1[1:0];
assign _072_ = op_5 == 2'h2;
always @(posedge \add_10ns_10ns_10_2_1_U3.top_add_10ns_10ns_10_2_1_Adder_1_U.clk )
\add_10ns_10ns_10_2_1_U3.top_add_10ns_10ns_10_2_1_Adder_1_U.bin_s1  <= _074_;
always @(posedge \add_10ns_10ns_10_2_1_U3.top_add_10ns_10ns_10_2_1_Adder_1_U.clk )
\add_10ns_10ns_10_2_1_U3.top_add_10ns_10ns_10_2_1_Adder_1_U.ain_s1  <= _073_;
always @(posedge \add_10ns_10ns_10_2_1_U3.top_add_10ns_10ns_10_2_1_Adder_1_U.clk )
\add_10ns_10ns_10_2_1_U3.top_add_10ns_10ns_10_2_1_Adder_1_U.sum_s1  <= _076_;
always @(posedge \add_10ns_10ns_10_2_1_U3.top_add_10ns_10ns_10_2_1_Adder_1_U.clk )
\add_10ns_10ns_10_2_1_U3.top_add_10ns_10ns_10_2_1_Adder_1_U.carry_s1  <= _075_;
assign _074_ = \add_10ns_10ns_10_2_1_U3.top_add_10ns_10ns_10_2_1_Adder_1_U.ce  ? \add_10ns_10ns_10_2_1_U3.top_add_10ns_10ns_10_2_1_Adder_1_U.b [9:5] : \add_10ns_10ns_10_2_1_U3.top_add_10ns_10ns_10_2_1_Adder_1_U.bin_s1 ;
assign _073_ = \add_10ns_10ns_10_2_1_U3.top_add_10ns_10ns_10_2_1_Adder_1_U.ce  ? \add_10ns_10ns_10_2_1_U3.top_add_10ns_10ns_10_2_1_Adder_1_U.a [9:5] : \add_10ns_10ns_10_2_1_U3.top_add_10ns_10ns_10_2_1_Adder_1_U.ain_s1 ;
assign _075_ = \add_10ns_10ns_10_2_1_U3.top_add_10ns_10ns_10_2_1_Adder_1_U.ce  ? \add_10ns_10ns_10_2_1_U3.top_add_10ns_10ns_10_2_1_Adder_1_U.facout_s1  : \add_10ns_10ns_10_2_1_U3.top_add_10ns_10ns_10_2_1_Adder_1_U.carry_s1 ;
assign _076_ = \add_10ns_10ns_10_2_1_U3.top_add_10ns_10ns_10_2_1_Adder_1_U.ce  ? \add_10ns_10ns_10_2_1_U3.top_add_10ns_10ns_10_2_1_Adder_1_U.fas_s1  : \add_10ns_10ns_10_2_1_U3.top_add_10ns_10ns_10_2_1_Adder_1_U.sum_s1 ;
assign _077_ = \add_10ns_10ns_10_2_1_U3.top_add_10ns_10ns_10_2_1_Adder_1_U.u1.a  + \add_10ns_10ns_10_2_1_U3.top_add_10ns_10ns_10_2_1_Adder_1_U.u1.b ;
assign { \add_10ns_10ns_10_2_1_U3.top_add_10ns_10ns_10_2_1_Adder_1_U.u1.cout , \add_10ns_10ns_10_2_1_U3.top_add_10ns_10ns_10_2_1_Adder_1_U.u1.s  } = _077_ + \add_10ns_10ns_10_2_1_U3.top_add_10ns_10ns_10_2_1_Adder_1_U.u1.cin ;
assign _078_ = \add_10ns_10ns_10_2_1_U3.top_add_10ns_10ns_10_2_1_Adder_1_U.u2.a  + \add_10ns_10ns_10_2_1_U3.top_add_10ns_10ns_10_2_1_Adder_1_U.u2.b ;
assign { \add_10ns_10ns_10_2_1_U3.top_add_10ns_10ns_10_2_1_Adder_1_U.u2.cout , \add_10ns_10ns_10_2_1_U3.top_add_10ns_10ns_10_2_1_Adder_1_U.u2.s  } = _078_ + \add_10ns_10ns_10_2_1_U3.top_add_10ns_10ns_10_2_1_Adder_1_U.u2.cin ;
always @(posedge \add_11ns_11ns_11_2_1_U14.top_add_11ns_11ns_11_2_1_Adder_9_U.clk )
\add_11ns_11ns_11_2_1_U14.top_add_11ns_11ns_11_2_1_Adder_9_U.bin_s1  <= _080_;
always @(posedge \add_11ns_11ns_11_2_1_U14.top_add_11ns_11ns_11_2_1_Adder_9_U.clk )
\add_11ns_11ns_11_2_1_U14.top_add_11ns_11ns_11_2_1_Adder_9_U.ain_s1  <= _079_;
always @(posedge \add_11ns_11ns_11_2_1_U14.top_add_11ns_11ns_11_2_1_Adder_9_U.clk )
\add_11ns_11ns_11_2_1_U14.top_add_11ns_11ns_11_2_1_Adder_9_U.sum_s1  <= _082_;
always @(posedge \add_11ns_11ns_11_2_1_U14.top_add_11ns_11ns_11_2_1_Adder_9_U.clk )
\add_11ns_11ns_11_2_1_U14.top_add_11ns_11ns_11_2_1_Adder_9_U.carry_s1  <= _081_;
assign _080_ = \add_11ns_11ns_11_2_1_U14.top_add_11ns_11ns_11_2_1_Adder_9_U.ce  ? \add_11ns_11ns_11_2_1_U14.top_add_11ns_11ns_11_2_1_Adder_9_U.b [10:5] : \add_11ns_11ns_11_2_1_U14.top_add_11ns_11ns_11_2_1_Adder_9_U.bin_s1 ;
assign _079_ = \add_11ns_11ns_11_2_1_U14.top_add_11ns_11ns_11_2_1_Adder_9_U.ce  ? \add_11ns_11ns_11_2_1_U14.top_add_11ns_11ns_11_2_1_Adder_9_U.a [10:5] : \add_11ns_11ns_11_2_1_U14.top_add_11ns_11ns_11_2_1_Adder_9_U.ain_s1 ;
assign _081_ = \add_11ns_11ns_11_2_1_U14.top_add_11ns_11ns_11_2_1_Adder_9_U.ce  ? \add_11ns_11ns_11_2_1_U14.top_add_11ns_11ns_11_2_1_Adder_9_U.facout_s1  : \add_11ns_11ns_11_2_1_U14.top_add_11ns_11ns_11_2_1_Adder_9_U.carry_s1 ;
assign _082_ = \add_11ns_11ns_11_2_1_U14.top_add_11ns_11ns_11_2_1_Adder_9_U.ce  ? \add_11ns_11ns_11_2_1_U14.top_add_11ns_11ns_11_2_1_Adder_9_U.fas_s1  : \add_11ns_11ns_11_2_1_U14.top_add_11ns_11ns_11_2_1_Adder_9_U.sum_s1 ;
assign _083_ = \add_11ns_11ns_11_2_1_U14.top_add_11ns_11ns_11_2_1_Adder_9_U.u1.a  + \add_11ns_11ns_11_2_1_U14.top_add_11ns_11ns_11_2_1_Adder_9_U.u1.b ;
assign { \add_11ns_11ns_11_2_1_U14.top_add_11ns_11ns_11_2_1_Adder_9_U.u1.cout , \add_11ns_11ns_11_2_1_U14.top_add_11ns_11ns_11_2_1_Adder_9_U.u1.s  } = _083_ + \add_11ns_11ns_11_2_1_U14.top_add_11ns_11ns_11_2_1_Adder_9_U.u1.cin ;
assign _084_ = \add_11ns_11ns_11_2_1_U14.top_add_11ns_11ns_11_2_1_Adder_9_U.u2.a  + \add_11ns_11ns_11_2_1_U14.top_add_11ns_11ns_11_2_1_Adder_9_U.u2.b ;
assign { \add_11ns_11ns_11_2_1_U14.top_add_11ns_11ns_11_2_1_Adder_9_U.u2.cout , \add_11ns_11ns_11_2_1_U14.top_add_11ns_11ns_11_2_1_Adder_9_U.u2.s  } = _084_ + \add_11ns_11ns_11_2_1_U14.top_add_11ns_11ns_11_2_1_Adder_9_U.u2.cin ;
always @(posedge \add_11ns_11ns_11_2_1_U16.top_add_11ns_11ns_11_2_1_Adder_9_U.clk )
\add_11ns_11ns_11_2_1_U16.top_add_11ns_11ns_11_2_1_Adder_9_U.bin_s1  <= _086_;
always @(posedge \add_11ns_11ns_11_2_1_U16.top_add_11ns_11ns_11_2_1_Adder_9_U.clk )
\add_11ns_11ns_11_2_1_U16.top_add_11ns_11ns_11_2_1_Adder_9_U.ain_s1  <= _085_;
always @(posedge \add_11ns_11ns_11_2_1_U16.top_add_11ns_11ns_11_2_1_Adder_9_U.clk )
\add_11ns_11ns_11_2_1_U16.top_add_11ns_11ns_11_2_1_Adder_9_U.sum_s1  <= _088_;
always @(posedge \add_11ns_11ns_11_2_1_U16.top_add_11ns_11ns_11_2_1_Adder_9_U.clk )
\add_11ns_11ns_11_2_1_U16.top_add_11ns_11ns_11_2_1_Adder_9_U.carry_s1  <= _087_;
assign _086_ = \add_11ns_11ns_11_2_1_U16.top_add_11ns_11ns_11_2_1_Adder_9_U.ce  ? \add_11ns_11ns_11_2_1_U16.top_add_11ns_11ns_11_2_1_Adder_9_U.b [10:5] : \add_11ns_11ns_11_2_1_U16.top_add_11ns_11ns_11_2_1_Adder_9_U.bin_s1 ;
assign _085_ = \add_11ns_11ns_11_2_1_U16.top_add_11ns_11ns_11_2_1_Adder_9_U.ce  ? \add_11ns_11ns_11_2_1_U16.top_add_11ns_11ns_11_2_1_Adder_9_U.a [10:5] : \add_11ns_11ns_11_2_1_U16.top_add_11ns_11ns_11_2_1_Adder_9_U.ain_s1 ;
assign _087_ = \add_11ns_11ns_11_2_1_U16.top_add_11ns_11ns_11_2_1_Adder_9_U.ce  ? \add_11ns_11ns_11_2_1_U16.top_add_11ns_11ns_11_2_1_Adder_9_U.facout_s1  : \add_11ns_11ns_11_2_1_U16.top_add_11ns_11ns_11_2_1_Adder_9_U.carry_s1 ;
assign _088_ = \add_11ns_11ns_11_2_1_U16.top_add_11ns_11ns_11_2_1_Adder_9_U.ce  ? \add_11ns_11ns_11_2_1_U16.top_add_11ns_11ns_11_2_1_Adder_9_U.fas_s1  : \add_11ns_11ns_11_2_1_U16.top_add_11ns_11ns_11_2_1_Adder_9_U.sum_s1 ;
assign _089_ = \add_11ns_11ns_11_2_1_U16.top_add_11ns_11ns_11_2_1_Adder_9_U.u1.a  + \add_11ns_11ns_11_2_1_U16.top_add_11ns_11ns_11_2_1_Adder_9_U.u1.b ;
assign { \add_11ns_11ns_11_2_1_U16.top_add_11ns_11ns_11_2_1_Adder_9_U.u1.cout , \add_11ns_11ns_11_2_1_U16.top_add_11ns_11ns_11_2_1_Adder_9_U.u1.s  } = _089_ + \add_11ns_11ns_11_2_1_U16.top_add_11ns_11ns_11_2_1_Adder_9_U.u1.cin ;
assign _090_ = \add_11ns_11ns_11_2_1_U16.top_add_11ns_11ns_11_2_1_Adder_9_U.u2.a  + \add_11ns_11ns_11_2_1_U16.top_add_11ns_11ns_11_2_1_Adder_9_U.u2.b ;
assign { \add_11ns_11ns_11_2_1_U16.top_add_11ns_11ns_11_2_1_Adder_9_U.u2.cout , \add_11ns_11ns_11_2_1_U16.top_add_11ns_11ns_11_2_1_Adder_9_U.u2.s  } = _090_ + \add_11ns_11ns_11_2_1_U16.top_add_11ns_11ns_11_2_1_Adder_9_U.u2.cin ;
always @(posedge \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_7_U.clk )
\add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_7_U.bin_s1  <= _092_;
always @(posedge \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_7_U.clk )
\add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_7_U.ain_s1  <= _091_;
always @(posedge \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_7_U.clk )
\add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_7_U.sum_s1  <= _094_;
always @(posedge \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_7_U.clk )
\add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_7_U.carry_s1  <= _093_;
assign _092_ = \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_7_U.ce  ? \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_7_U.b [10:5] : \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_7_U.bin_s1 ;
assign _091_ = \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_7_U.ce  ? \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_7_U.a [10:5] : \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_7_U.ain_s1 ;
assign _093_ = \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_7_U.ce  ? \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_7_U.facout_s1  : \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_7_U.carry_s1 ;
assign _094_ = \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_7_U.ce  ? \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_7_U.fas_s1  : \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_7_U.sum_s1 ;
assign _095_ = \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_7_U.u1.a  + \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_7_U.u1.b ;
assign { \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_7_U.u1.cout , \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_7_U.u1.s  } = _095_ + \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_7_U.u1.cin ;
assign _096_ = \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_7_U.u2.a  + \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_7_U.u2.b ;
assign { \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_7_U.u2.cout , \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_7_U.u2.s  } = _096_ + \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_7_U.u2.cin ;
always @(posedge \add_11ns_11s_11_2_1_U20.top_add_11ns_11s_11_2_1_Adder_7_U.clk )
\add_11ns_11s_11_2_1_U20.top_add_11ns_11s_11_2_1_Adder_7_U.bin_s1  <= _098_;
always @(posedge \add_11ns_11s_11_2_1_U20.top_add_11ns_11s_11_2_1_Adder_7_U.clk )
\add_11ns_11s_11_2_1_U20.top_add_11ns_11s_11_2_1_Adder_7_U.ain_s1  <= _097_;
always @(posedge \add_11ns_11s_11_2_1_U20.top_add_11ns_11s_11_2_1_Adder_7_U.clk )
\add_11ns_11s_11_2_1_U20.top_add_11ns_11s_11_2_1_Adder_7_U.sum_s1  <= _100_;
always @(posedge \add_11ns_11s_11_2_1_U20.top_add_11ns_11s_11_2_1_Adder_7_U.clk )
\add_11ns_11s_11_2_1_U20.top_add_11ns_11s_11_2_1_Adder_7_U.carry_s1  <= _099_;
assign _098_ = \add_11ns_11s_11_2_1_U20.top_add_11ns_11s_11_2_1_Adder_7_U.ce  ? \add_11ns_11s_11_2_1_U20.top_add_11ns_11s_11_2_1_Adder_7_U.b [10:5] : \add_11ns_11s_11_2_1_U20.top_add_11ns_11s_11_2_1_Adder_7_U.bin_s1 ;
assign _097_ = \add_11ns_11s_11_2_1_U20.top_add_11ns_11s_11_2_1_Adder_7_U.ce  ? \add_11ns_11s_11_2_1_U20.top_add_11ns_11s_11_2_1_Adder_7_U.a [10:5] : \add_11ns_11s_11_2_1_U20.top_add_11ns_11s_11_2_1_Adder_7_U.ain_s1 ;
assign _099_ = \add_11ns_11s_11_2_1_U20.top_add_11ns_11s_11_2_1_Adder_7_U.ce  ? \add_11ns_11s_11_2_1_U20.top_add_11ns_11s_11_2_1_Adder_7_U.facout_s1  : \add_11ns_11s_11_2_1_U20.top_add_11ns_11s_11_2_1_Adder_7_U.carry_s1 ;
assign _100_ = \add_11ns_11s_11_2_1_U20.top_add_11ns_11s_11_2_1_Adder_7_U.ce  ? \add_11ns_11s_11_2_1_U20.top_add_11ns_11s_11_2_1_Adder_7_U.fas_s1  : \add_11ns_11s_11_2_1_U20.top_add_11ns_11s_11_2_1_Adder_7_U.sum_s1 ;
assign _101_ = \add_11ns_11s_11_2_1_U20.top_add_11ns_11s_11_2_1_Adder_7_U.u1.a  + \add_11ns_11s_11_2_1_U20.top_add_11ns_11s_11_2_1_Adder_7_U.u1.b ;
assign { \add_11ns_11s_11_2_1_U20.top_add_11ns_11s_11_2_1_Adder_7_U.u1.cout , \add_11ns_11s_11_2_1_U20.top_add_11ns_11s_11_2_1_Adder_7_U.u1.s  } = _101_ + \add_11ns_11s_11_2_1_U20.top_add_11ns_11s_11_2_1_Adder_7_U.u1.cin ;
assign _102_ = \add_11ns_11s_11_2_1_U20.top_add_11ns_11s_11_2_1_Adder_7_U.u2.a  + \add_11ns_11s_11_2_1_U20.top_add_11ns_11s_11_2_1_Adder_7_U.u2.b ;
assign { \add_11ns_11s_11_2_1_U20.top_add_11ns_11s_11_2_1_Adder_7_U.u2.cout , \add_11ns_11s_11_2_1_U20.top_add_11ns_11s_11_2_1_Adder_7_U.u2.s  } = _102_ + \add_11ns_11s_11_2_1_U20.top_add_11ns_11s_11_2_1_Adder_7_U.u2.cin ;
always @(posedge \add_11ns_11s_11_2_1_U21.top_add_11ns_11s_11_2_1_Adder_7_U.clk )
\add_11ns_11s_11_2_1_U21.top_add_11ns_11s_11_2_1_Adder_7_U.bin_s1  <= _104_;
always @(posedge \add_11ns_11s_11_2_1_U21.top_add_11ns_11s_11_2_1_Adder_7_U.clk )
\add_11ns_11s_11_2_1_U21.top_add_11ns_11s_11_2_1_Adder_7_U.ain_s1  <= _103_;
always @(posedge \add_11ns_11s_11_2_1_U21.top_add_11ns_11s_11_2_1_Adder_7_U.clk )
\add_11ns_11s_11_2_1_U21.top_add_11ns_11s_11_2_1_Adder_7_U.sum_s1  <= _106_;
always @(posedge \add_11ns_11s_11_2_1_U21.top_add_11ns_11s_11_2_1_Adder_7_U.clk )
\add_11ns_11s_11_2_1_U21.top_add_11ns_11s_11_2_1_Adder_7_U.carry_s1  <= _105_;
assign _104_ = \add_11ns_11s_11_2_1_U21.top_add_11ns_11s_11_2_1_Adder_7_U.ce  ? \add_11ns_11s_11_2_1_U21.top_add_11ns_11s_11_2_1_Adder_7_U.b [10:5] : \add_11ns_11s_11_2_1_U21.top_add_11ns_11s_11_2_1_Adder_7_U.bin_s1 ;
assign _103_ = \add_11ns_11s_11_2_1_U21.top_add_11ns_11s_11_2_1_Adder_7_U.ce  ? \add_11ns_11s_11_2_1_U21.top_add_11ns_11s_11_2_1_Adder_7_U.a [10:5] : \add_11ns_11s_11_2_1_U21.top_add_11ns_11s_11_2_1_Adder_7_U.ain_s1 ;
assign _105_ = \add_11ns_11s_11_2_1_U21.top_add_11ns_11s_11_2_1_Adder_7_U.ce  ? \add_11ns_11s_11_2_1_U21.top_add_11ns_11s_11_2_1_Adder_7_U.facout_s1  : \add_11ns_11s_11_2_1_U21.top_add_11ns_11s_11_2_1_Adder_7_U.carry_s1 ;
assign _106_ = \add_11ns_11s_11_2_1_U21.top_add_11ns_11s_11_2_1_Adder_7_U.ce  ? \add_11ns_11s_11_2_1_U21.top_add_11ns_11s_11_2_1_Adder_7_U.fas_s1  : \add_11ns_11s_11_2_1_U21.top_add_11ns_11s_11_2_1_Adder_7_U.sum_s1 ;
assign _107_ = \add_11ns_11s_11_2_1_U21.top_add_11ns_11s_11_2_1_Adder_7_U.u1.a  + \add_11ns_11s_11_2_1_U21.top_add_11ns_11s_11_2_1_Adder_7_U.u1.b ;
assign { \add_11ns_11s_11_2_1_U21.top_add_11ns_11s_11_2_1_Adder_7_U.u1.cout , \add_11ns_11s_11_2_1_U21.top_add_11ns_11s_11_2_1_Adder_7_U.u1.s  } = _107_ + \add_11ns_11s_11_2_1_U21.top_add_11ns_11s_11_2_1_Adder_7_U.u1.cin ;
assign _108_ = \add_11ns_11s_11_2_1_U21.top_add_11ns_11s_11_2_1_Adder_7_U.u2.a  + \add_11ns_11s_11_2_1_U21.top_add_11ns_11s_11_2_1_Adder_7_U.u2.b ;
assign { \add_11ns_11s_11_2_1_U21.top_add_11ns_11s_11_2_1_Adder_7_U.u2.cout , \add_11ns_11s_11_2_1_U21.top_add_11ns_11s_11_2_1_Adder_7_U.u2.s  } = _108_ + \add_11ns_11s_11_2_1_U21.top_add_11ns_11s_11_2_1_Adder_7_U.u2.cin ;
always @(posedge \add_11s_11ns_11_2_1_U13.top_add_11s_11ns_11_2_1_Adder_4_U.clk )
\add_11s_11ns_11_2_1_U13.top_add_11s_11ns_11_2_1_Adder_4_U.bin_s1  <= _110_;
always @(posedge \add_11s_11ns_11_2_1_U13.top_add_11s_11ns_11_2_1_Adder_4_U.clk )
\add_11s_11ns_11_2_1_U13.top_add_11s_11ns_11_2_1_Adder_4_U.ain_s1  <= _109_;
always @(posedge \add_11s_11ns_11_2_1_U13.top_add_11s_11ns_11_2_1_Adder_4_U.clk )
\add_11s_11ns_11_2_1_U13.top_add_11s_11ns_11_2_1_Adder_4_U.sum_s1  <= _112_;
always @(posedge \add_11s_11ns_11_2_1_U13.top_add_11s_11ns_11_2_1_Adder_4_U.clk )
\add_11s_11ns_11_2_1_U13.top_add_11s_11ns_11_2_1_Adder_4_U.carry_s1  <= _111_;
assign _110_ = \add_11s_11ns_11_2_1_U13.top_add_11s_11ns_11_2_1_Adder_4_U.ce  ? \add_11s_11ns_11_2_1_U13.top_add_11s_11ns_11_2_1_Adder_4_U.b [10:5] : \add_11s_11ns_11_2_1_U13.top_add_11s_11ns_11_2_1_Adder_4_U.bin_s1 ;
assign _109_ = \add_11s_11ns_11_2_1_U13.top_add_11s_11ns_11_2_1_Adder_4_U.ce  ? \add_11s_11ns_11_2_1_U13.top_add_11s_11ns_11_2_1_Adder_4_U.a [10:5] : \add_11s_11ns_11_2_1_U13.top_add_11s_11ns_11_2_1_Adder_4_U.ain_s1 ;
assign _111_ = \add_11s_11ns_11_2_1_U13.top_add_11s_11ns_11_2_1_Adder_4_U.ce  ? \add_11s_11ns_11_2_1_U13.top_add_11s_11ns_11_2_1_Adder_4_U.facout_s1  : \add_11s_11ns_11_2_1_U13.top_add_11s_11ns_11_2_1_Adder_4_U.carry_s1 ;
assign _112_ = \add_11s_11ns_11_2_1_U13.top_add_11s_11ns_11_2_1_Adder_4_U.ce  ? \add_11s_11ns_11_2_1_U13.top_add_11s_11ns_11_2_1_Adder_4_U.fas_s1  : \add_11s_11ns_11_2_1_U13.top_add_11s_11ns_11_2_1_Adder_4_U.sum_s1 ;
assign _113_ = \add_11s_11ns_11_2_1_U13.top_add_11s_11ns_11_2_1_Adder_4_U.u1.a  + \add_11s_11ns_11_2_1_U13.top_add_11s_11ns_11_2_1_Adder_4_U.u1.b ;
assign { \add_11s_11ns_11_2_1_U13.top_add_11s_11ns_11_2_1_Adder_4_U.u1.cout , \add_11s_11ns_11_2_1_U13.top_add_11s_11ns_11_2_1_Adder_4_U.u1.s  } = _113_ + \add_11s_11ns_11_2_1_U13.top_add_11s_11ns_11_2_1_Adder_4_U.u1.cin ;
assign _114_ = \add_11s_11ns_11_2_1_U13.top_add_11s_11ns_11_2_1_Adder_4_U.u2.a  + \add_11s_11ns_11_2_1_U13.top_add_11s_11ns_11_2_1_Adder_4_U.u2.b ;
assign { \add_11s_11ns_11_2_1_U13.top_add_11s_11ns_11_2_1_Adder_4_U.u2.cout , \add_11s_11ns_11_2_1_U13.top_add_11s_11ns_11_2_1_Adder_4_U.u2.s  } = _114_ + \add_11s_11ns_11_2_1_U13.top_add_11s_11ns_11_2_1_Adder_4_U.u2.cin ;
always @(posedge \add_11s_11ns_11_2_1_U6.top_add_11s_11ns_11_2_1_Adder_4_U.clk )
\add_11s_11ns_11_2_1_U6.top_add_11s_11ns_11_2_1_Adder_4_U.bin_s1  <= _116_;
always @(posedge \add_11s_11ns_11_2_1_U6.top_add_11s_11ns_11_2_1_Adder_4_U.clk )
\add_11s_11ns_11_2_1_U6.top_add_11s_11ns_11_2_1_Adder_4_U.ain_s1  <= _115_;
always @(posedge \add_11s_11ns_11_2_1_U6.top_add_11s_11ns_11_2_1_Adder_4_U.clk )
\add_11s_11ns_11_2_1_U6.top_add_11s_11ns_11_2_1_Adder_4_U.sum_s1  <= _118_;
always @(posedge \add_11s_11ns_11_2_1_U6.top_add_11s_11ns_11_2_1_Adder_4_U.clk )
\add_11s_11ns_11_2_1_U6.top_add_11s_11ns_11_2_1_Adder_4_U.carry_s1  <= _117_;
assign _116_ = \add_11s_11ns_11_2_1_U6.top_add_11s_11ns_11_2_1_Adder_4_U.ce  ? \add_11s_11ns_11_2_1_U6.top_add_11s_11ns_11_2_1_Adder_4_U.b [10:5] : \add_11s_11ns_11_2_1_U6.top_add_11s_11ns_11_2_1_Adder_4_U.bin_s1 ;
assign _115_ = \add_11s_11ns_11_2_1_U6.top_add_11s_11ns_11_2_1_Adder_4_U.ce  ? \add_11s_11ns_11_2_1_U6.top_add_11s_11ns_11_2_1_Adder_4_U.a [10:5] : \add_11s_11ns_11_2_1_U6.top_add_11s_11ns_11_2_1_Adder_4_U.ain_s1 ;
assign _117_ = \add_11s_11ns_11_2_1_U6.top_add_11s_11ns_11_2_1_Adder_4_U.ce  ? \add_11s_11ns_11_2_1_U6.top_add_11s_11ns_11_2_1_Adder_4_U.facout_s1  : \add_11s_11ns_11_2_1_U6.top_add_11s_11ns_11_2_1_Adder_4_U.carry_s1 ;
assign _118_ = \add_11s_11ns_11_2_1_U6.top_add_11s_11ns_11_2_1_Adder_4_U.ce  ? \add_11s_11ns_11_2_1_U6.top_add_11s_11ns_11_2_1_Adder_4_U.fas_s1  : \add_11s_11ns_11_2_1_U6.top_add_11s_11ns_11_2_1_Adder_4_U.sum_s1 ;
assign _119_ = \add_11s_11ns_11_2_1_U6.top_add_11s_11ns_11_2_1_Adder_4_U.u1.a  + \add_11s_11ns_11_2_1_U6.top_add_11s_11ns_11_2_1_Adder_4_U.u1.b ;
assign { \add_11s_11ns_11_2_1_U6.top_add_11s_11ns_11_2_1_Adder_4_U.u1.cout , \add_11s_11ns_11_2_1_U6.top_add_11s_11ns_11_2_1_Adder_4_U.u1.s  } = _119_ + \add_11s_11ns_11_2_1_U6.top_add_11s_11ns_11_2_1_Adder_4_U.u1.cin ;
assign _120_ = \add_11s_11ns_11_2_1_U6.top_add_11s_11ns_11_2_1_Adder_4_U.u2.a  + \add_11s_11ns_11_2_1_U6.top_add_11s_11ns_11_2_1_Adder_4_U.u2.b ;
assign { \add_11s_11ns_11_2_1_U6.top_add_11s_11ns_11_2_1_Adder_4_U.u2.cout , \add_11s_11ns_11_2_1_U6.top_add_11s_11ns_11_2_1_Adder_4_U.u2.s  } = _120_ + \add_11s_11ns_11_2_1_U6.top_add_11s_11ns_11_2_1_Adder_4_U.u2.cin ;
always @(posedge \add_12ns_12s_12_2_1_U1.top_add_12ns_12s_12_2_1_Adder_0_U.clk )
\add_12ns_12s_12_2_1_U1.top_add_12ns_12s_12_2_1_Adder_0_U.bin_s1  <= _122_;
always @(posedge \add_12ns_12s_12_2_1_U1.top_add_12ns_12s_12_2_1_Adder_0_U.clk )
\add_12ns_12s_12_2_1_U1.top_add_12ns_12s_12_2_1_Adder_0_U.ain_s1  <= _121_;
always @(posedge \add_12ns_12s_12_2_1_U1.top_add_12ns_12s_12_2_1_Adder_0_U.clk )
\add_12ns_12s_12_2_1_U1.top_add_12ns_12s_12_2_1_Adder_0_U.sum_s1  <= _124_;
always @(posedge \add_12ns_12s_12_2_1_U1.top_add_12ns_12s_12_2_1_Adder_0_U.clk )
\add_12ns_12s_12_2_1_U1.top_add_12ns_12s_12_2_1_Adder_0_U.carry_s1  <= _123_;
assign _122_ = \add_12ns_12s_12_2_1_U1.top_add_12ns_12s_12_2_1_Adder_0_U.ce  ? \add_12ns_12s_12_2_1_U1.top_add_12ns_12s_12_2_1_Adder_0_U.b [11:6] : \add_12ns_12s_12_2_1_U1.top_add_12ns_12s_12_2_1_Adder_0_U.bin_s1 ;
assign _121_ = \add_12ns_12s_12_2_1_U1.top_add_12ns_12s_12_2_1_Adder_0_U.ce  ? \add_12ns_12s_12_2_1_U1.top_add_12ns_12s_12_2_1_Adder_0_U.a [11:6] : \add_12ns_12s_12_2_1_U1.top_add_12ns_12s_12_2_1_Adder_0_U.ain_s1 ;
assign _123_ = \add_12ns_12s_12_2_1_U1.top_add_12ns_12s_12_2_1_Adder_0_U.ce  ? \add_12ns_12s_12_2_1_U1.top_add_12ns_12s_12_2_1_Adder_0_U.facout_s1  : \add_12ns_12s_12_2_1_U1.top_add_12ns_12s_12_2_1_Adder_0_U.carry_s1 ;
assign _124_ = \add_12ns_12s_12_2_1_U1.top_add_12ns_12s_12_2_1_Adder_0_U.ce  ? \add_12ns_12s_12_2_1_U1.top_add_12ns_12s_12_2_1_Adder_0_U.fas_s1  : \add_12ns_12s_12_2_1_U1.top_add_12ns_12s_12_2_1_Adder_0_U.sum_s1 ;
assign _125_ = \add_12ns_12s_12_2_1_U1.top_add_12ns_12s_12_2_1_Adder_0_U.u1.a  + \add_12ns_12s_12_2_1_U1.top_add_12ns_12s_12_2_1_Adder_0_U.u1.b ;
assign { \add_12ns_12s_12_2_1_U1.top_add_12ns_12s_12_2_1_Adder_0_U.u1.cout , \add_12ns_12s_12_2_1_U1.top_add_12ns_12s_12_2_1_Adder_0_U.u1.s  } = _125_ + \add_12ns_12s_12_2_1_U1.top_add_12ns_12s_12_2_1_Adder_0_U.u1.cin ;
assign _126_ = \add_12ns_12s_12_2_1_U1.top_add_12ns_12s_12_2_1_Adder_0_U.u2.a  + \add_12ns_12s_12_2_1_U1.top_add_12ns_12s_12_2_1_Adder_0_U.u2.b ;
assign { \add_12ns_12s_12_2_1_U1.top_add_12ns_12s_12_2_1_Adder_0_U.u2.cout , \add_12ns_12s_12_2_1_U1.top_add_12ns_12s_12_2_1_Adder_0_U.u2.s  } = _126_ + \add_12ns_12s_12_2_1_U1.top_add_12ns_12s_12_2_1_Adder_0_U.u2.cin ;
always @(posedge \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_3_U.clk )
\add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_3_U.bin_s1  <= _128_;
always @(posedge \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_3_U.clk )
\add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_3_U.ain_s1  <= _127_;
always @(posedge \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_3_U.clk )
\add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_3_U.sum_s1  <= _130_;
always @(posedge \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_3_U.clk )
\add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_3_U.carry_s1  <= _129_;
assign _128_ = \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_3_U.ce  ? \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_3_U.b [1] : \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_3_U.bin_s1 ;
assign _127_ = \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_3_U.ce  ? \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_3_U.a [1] : \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_3_U.ain_s1 ;
assign _129_ = \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_3_U.ce  ? \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_3_U.facout_s1  : \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_3_U.carry_s1 ;
assign _130_ = \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_3_U.ce  ? \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_3_U.fas_s1  : \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_3_U.sum_s1 ;
assign _131_ = \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_3_U.u1.a  + \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_3_U.u1.b ;
assign { \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_3_U.u1.cout , \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_3_U.u1.s  } = _131_ + \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_3_U.u1.cin ;
assign _132_ = \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_3_U.u2.a  + \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_3_U.u2.b ;
assign { \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_3_U.u2.cout , \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_3_U.u2.s  } = _132_ + \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_3_U.u2.cin ;
always @(posedge \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_13_U.clk )
\add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_13_U.bin_s1  <= _134_;
always @(posedge \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_13_U.clk )
\add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_13_U.ain_s1  <= _133_;
always @(posedge \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_13_U.clk )
\add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_13_U.sum_s1  <= _136_;
always @(posedge \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_13_U.clk )
\add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_13_U.carry_s1  <= _135_;
assign _134_ = \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_13_U.ce  ? \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_13_U.b [31:16] : \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_13_U.bin_s1 ;
assign _133_ = \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_13_U.ce  ? \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_13_U.a [31:16] : \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_13_U.ain_s1 ;
assign _135_ = \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_13_U.ce  ? \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_13_U.facout_s1  : \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_13_U.carry_s1 ;
assign _136_ = \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_13_U.ce  ? \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_13_U.fas_s1  : \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_13_U.sum_s1 ;
assign _137_ = \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_13_U.u1.a  + \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_13_U.u1.b ;
assign { \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_13_U.u1.cout , \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_13_U.u1.s  } = _137_ + \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_13_U.u1.cin ;
assign _138_ = \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_13_U.u2.a  + \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_13_U.u2.b ;
assign { \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_13_U.u2.cout , \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_13_U.u2.s  } = _138_ + \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_13_U.u2.cin ;
always @(posedge \add_35s_35s_35_2_1_U22.top_add_35s_35s_35_2_1_Adder_12_U.clk )
\add_35s_35s_35_2_1_U22.top_add_35s_35s_35_2_1_Adder_12_U.bin_s1  <= _140_;
always @(posedge \add_35s_35s_35_2_1_U22.top_add_35s_35s_35_2_1_Adder_12_U.clk )
\add_35s_35s_35_2_1_U22.top_add_35s_35s_35_2_1_Adder_12_U.ain_s1  <= _139_;
always @(posedge \add_35s_35s_35_2_1_U22.top_add_35s_35s_35_2_1_Adder_12_U.clk )
\add_35s_35s_35_2_1_U22.top_add_35s_35s_35_2_1_Adder_12_U.sum_s1  <= _142_;
always @(posedge \add_35s_35s_35_2_1_U22.top_add_35s_35s_35_2_1_Adder_12_U.clk )
\add_35s_35s_35_2_1_U22.top_add_35s_35s_35_2_1_Adder_12_U.carry_s1  <= _141_;
assign _140_ = \add_35s_35s_35_2_1_U22.top_add_35s_35s_35_2_1_Adder_12_U.ce  ? \add_35s_35s_35_2_1_U22.top_add_35s_35s_35_2_1_Adder_12_U.b [34:17] : \add_35s_35s_35_2_1_U22.top_add_35s_35s_35_2_1_Adder_12_U.bin_s1 ;
assign _139_ = \add_35s_35s_35_2_1_U22.top_add_35s_35s_35_2_1_Adder_12_U.ce  ? \add_35s_35s_35_2_1_U22.top_add_35s_35s_35_2_1_Adder_12_U.a [34:17] : \add_35s_35s_35_2_1_U22.top_add_35s_35s_35_2_1_Adder_12_U.ain_s1 ;
assign _141_ = \add_35s_35s_35_2_1_U22.top_add_35s_35s_35_2_1_Adder_12_U.ce  ? \add_35s_35s_35_2_1_U22.top_add_35s_35s_35_2_1_Adder_12_U.facout_s1  : \add_35s_35s_35_2_1_U22.top_add_35s_35s_35_2_1_Adder_12_U.carry_s1 ;
assign _142_ = \add_35s_35s_35_2_1_U22.top_add_35s_35s_35_2_1_Adder_12_U.ce  ? \add_35s_35s_35_2_1_U22.top_add_35s_35s_35_2_1_Adder_12_U.fas_s1  : \add_35s_35s_35_2_1_U22.top_add_35s_35s_35_2_1_Adder_12_U.sum_s1 ;
assign _143_ = \add_35s_35s_35_2_1_U22.top_add_35s_35s_35_2_1_Adder_12_U.u1.a  + \add_35s_35s_35_2_1_U22.top_add_35s_35s_35_2_1_Adder_12_U.u1.b ;
assign { \add_35s_35s_35_2_1_U22.top_add_35s_35s_35_2_1_Adder_12_U.u1.cout , \add_35s_35s_35_2_1_U22.top_add_35s_35s_35_2_1_Adder_12_U.u1.s  } = _143_ + \add_35s_35s_35_2_1_U22.top_add_35s_35s_35_2_1_Adder_12_U.u1.cin ;
assign _144_ = \add_35s_35s_35_2_1_U22.top_add_35s_35s_35_2_1_Adder_12_U.u2.a  + \add_35s_35s_35_2_1_U22.top_add_35s_35s_35_2_1_Adder_12_U.u2.b ;
assign { \add_35s_35s_35_2_1_U22.top_add_35s_35s_35_2_1_Adder_12_U.u2.cout , \add_35s_35s_35_2_1_U22.top_add_35s_35s_35_2_1_Adder_12_U.u2.s  } = _144_ + \add_35s_35s_35_2_1_U22.top_add_35s_35s_35_2_1_Adder_12_U.u2.cin ;
always @(posedge \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_10_U.clk )
\add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_10_U.bin_s1  <= _146_;
always @(posedge \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_10_U.clk )
\add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_10_U.ain_s1  <= _145_;
always @(posedge \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_10_U.clk )
\add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_10_U.sum_s1  <= _148_;
always @(posedge \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_10_U.clk )
\add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_10_U.carry_s1  <= _147_;
assign _146_ = \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_10_U.ce  ? \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_10_U.b [2:1] : \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_10_U.bin_s1 ;
assign _145_ = \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_10_U.ce  ? \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_10_U.a [2:1] : \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_10_U.ain_s1 ;
assign _147_ = \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_10_U.ce  ? \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_10_U.facout_s1  : \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_10_U.carry_s1 ;
assign _148_ = \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_10_U.ce  ? \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_10_U.fas_s1  : \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_10_U.sum_s1 ;
assign _149_ = \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_10_U.u1.a  + \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_10_U.u1.b ;
assign { \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_10_U.u1.cout , \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_10_U.u1.s  } = _149_ + \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_10_U.u1.cin ;
assign _150_ = \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_10_U.u2.a  + \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_10_U.u2.b ;
assign { \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_10_U.u2.cout , \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_10_U.u2.s  } = _150_ + \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_10_U.u2.cin ;
always @(posedge \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.clk )
\add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.bin_s1  <= _152_;
always @(posedge \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.clk )
\add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.ain_s1  <= _151_;
always @(posedge \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.clk )
\add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.sum_s1  <= _154_;
always @(posedge \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.clk )
\add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.carry_s1  <= _153_;
assign _152_ = \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.ce  ? \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.b [2:1] : \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.bin_s1 ;
assign _151_ = \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.ce  ? \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.a [2:1] : \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.ain_s1 ;
assign _153_ = \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.ce  ? \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.facout_s1  : \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.carry_s1 ;
assign _154_ = \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.ce  ? \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.fas_s1  : \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.sum_s1 ;
assign _155_ = \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.u1.a  + \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.u1.b ;
assign { \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.u1.cout , \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.u1.s  } = _155_ + \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.u1.cin ;
assign _156_ = \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.u2.a  + \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.u2.b ;
assign { \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.u2.cout , \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.u2.s  } = _156_ + \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.u2.cin ;
always @(posedge \add_3s_3s_3_2_1_U9.top_add_3s_3s_3_2_1_Adder_5_U.clk )
\add_3s_3s_3_2_1_U9.top_add_3s_3s_3_2_1_Adder_5_U.bin_s1  <= _158_;
always @(posedge \add_3s_3s_3_2_1_U9.top_add_3s_3s_3_2_1_Adder_5_U.clk )
\add_3s_3s_3_2_1_U9.top_add_3s_3s_3_2_1_Adder_5_U.ain_s1  <= _157_;
always @(posedge \add_3s_3s_3_2_1_U9.top_add_3s_3s_3_2_1_Adder_5_U.clk )
\add_3s_3s_3_2_1_U9.top_add_3s_3s_3_2_1_Adder_5_U.sum_s1  <= _160_;
always @(posedge \add_3s_3s_3_2_1_U9.top_add_3s_3s_3_2_1_Adder_5_U.clk )
\add_3s_3s_3_2_1_U9.top_add_3s_3s_3_2_1_Adder_5_U.carry_s1  <= _159_;
assign _158_ = \add_3s_3s_3_2_1_U9.top_add_3s_3s_3_2_1_Adder_5_U.ce  ? \add_3s_3s_3_2_1_U9.top_add_3s_3s_3_2_1_Adder_5_U.b [2:1] : \add_3s_3s_3_2_1_U9.top_add_3s_3s_3_2_1_Adder_5_U.bin_s1 ;
assign _157_ = \add_3s_3s_3_2_1_U9.top_add_3s_3s_3_2_1_Adder_5_U.ce  ? \add_3s_3s_3_2_1_U9.top_add_3s_3s_3_2_1_Adder_5_U.a [2:1] : \add_3s_3s_3_2_1_U9.top_add_3s_3s_3_2_1_Adder_5_U.ain_s1 ;
assign _159_ = \add_3s_3s_3_2_1_U9.top_add_3s_3s_3_2_1_Adder_5_U.ce  ? \add_3s_3s_3_2_1_U9.top_add_3s_3s_3_2_1_Adder_5_U.facout_s1  : \add_3s_3s_3_2_1_U9.top_add_3s_3s_3_2_1_Adder_5_U.carry_s1 ;
assign _160_ = \add_3s_3s_3_2_1_U9.top_add_3s_3s_3_2_1_Adder_5_U.ce  ? \add_3s_3s_3_2_1_U9.top_add_3s_3s_3_2_1_Adder_5_U.fas_s1  : \add_3s_3s_3_2_1_U9.top_add_3s_3s_3_2_1_Adder_5_U.sum_s1 ;
assign _161_ = \add_3s_3s_3_2_1_U9.top_add_3s_3s_3_2_1_Adder_5_U.u1.a  + \add_3s_3s_3_2_1_U9.top_add_3s_3s_3_2_1_Adder_5_U.u1.b ;
assign { \add_3s_3s_3_2_1_U9.top_add_3s_3s_3_2_1_Adder_5_U.u1.cout , \add_3s_3s_3_2_1_U9.top_add_3s_3s_3_2_1_Adder_5_U.u1.s  } = _161_ + \add_3s_3s_3_2_1_U9.top_add_3s_3s_3_2_1_Adder_5_U.u1.cin ;
assign _162_ = \add_3s_3s_3_2_1_U9.top_add_3s_3s_3_2_1_Adder_5_U.u2.a  + \add_3s_3s_3_2_1_U9.top_add_3s_3s_3_2_1_Adder_5_U.u2.b ;
assign { \add_3s_3s_3_2_1_U9.top_add_3s_3s_3_2_1_Adder_5_U.u2.cout , \add_3s_3s_3_2_1_U9.top_add_3s_3s_3_2_1_Adder_5_U.u2.s  } = _162_ + \add_3s_3s_3_2_1_U9.top_add_3s_3s_3_2_1_Adder_5_U.u2.cin ;
always @(posedge \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_8_U.clk )
\add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_8_U.bin_s1  <= _164_;
always @(posedge \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_8_U.clk )
\add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_8_U.ain_s1  <= _163_;
always @(posedge \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_8_U.clk )
\add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_8_U.sum_s1  <= _166_;
always @(posedge \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_8_U.clk )
\add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_8_U.carry_s1  <= _165_;
assign _164_ = \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_8_U.ce  ? \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_8_U.b [5:3] : \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_8_U.bin_s1 ;
assign _163_ = \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_8_U.ce  ? \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_8_U.a [5:3] : \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_8_U.ain_s1 ;
assign _165_ = \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_8_U.ce  ? \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_8_U.facout_s1  : \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_8_U.carry_s1 ;
assign _166_ = \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_8_U.ce  ? \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_8_U.fas_s1  : \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_8_U.sum_s1 ;
assign _167_ = \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_8_U.u1.a  + \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_8_U.u1.b ;
assign { \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_8_U.u1.cout , \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_8_U.u1.s  } = _167_ + \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_8_U.u1.cin ;
assign _168_ = \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_8_U.u2.a  + \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_8_U.u2.b ;
assign { \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_8_U.u2.cout , \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_8_U.u2.s  } = _168_ + \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_8_U.u2.cin ;
always @(posedge \ashr_32s_16ns_32_7_1_U18.clk )
\ashr_32s_16ns_32_7_1_U18.dout_array[5]  <= _180_;
always @(posedge \ashr_32s_16ns_32_7_1_U18.clk )
\ashr_32s_16ns_32_7_1_U18.din1_cast_array[5]  <= _174_;
always @(posedge \ashr_32s_16ns_32_7_1_U18.clk )
\ashr_32s_16ns_32_7_1_U18.dout_array[4]  <= _179_;
always @(posedge \ashr_32s_16ns_32_7_1_U18.clk )
\ashr_32s_16ns_32_7_1_U18.din1_cast_array[4]  <= _173_;
always @(posedge \ashr_32s_16ns_32_7_1_U18.clk )
\ashr_32s_16ns_32_7_1_U18.dout_array[3]  <= _178_;
always @(posedge \ashr_32s_16ns_32_7_1_U18.clk )
\ashr_32s_16ns_32_7_1_U18.din1_cast_array[3]  <= _172_;
always @(posedge \ashr_32s_16ns_32_7_1_U18.clk )
\ashr_32s_16ns_32_7_1_U18.dout_array[2]  <= _177_;
always @(posedge \ashr_32s_16ns_32_7_1_U18.clk )
\ashr_32s_16ns_32_7_1_U18.din1_cast_array[2]  <= _171_;
always @(posedge \ashr_32s_16ns_32_7_1_U18.clk )
\ashr_32s_16ns_32_7_1_U18.dout_array[1]  <= _176_;
always @(posedge \ashr_32s_16ns_32_7_1_U18.clk )
\ashr_32s_16ns_32_7_1_U18.din1_cast_array[1]  <= _170_;
always @(posedge \ashr_32s_16ns_32_7_1_U18.clk )
\ashr_32s_16ns_32_7_1_U18.dout_array[0]  <= _175_;
always @(posedge \ashr_32s_16ns_32_7_1_U18.clk )
\ashr_32s_16ns_32_7_1_U18.din1_cast_array[0]  <= _169_;
assign _181_ = \ashr_32s_16ns_32_7_1_U18.ce  ? \ashr_32s_16ns_32_7_1_U18.din1_cast_array[4]  : \ashr_32s_16ns_32_7_1_U18.din1_cast_array[5] ;
assign _174_ = \ashr_32s_16ns_32_7_1_U18.reset  ? 16'h0000 : _181_;
assign _182_ = \ashr_32s_16ns_32_7_1_U18.ce  ? _197_ : \ashr_32s_16ns_32_7_1_U18.dout_array[5] ;
assign _180_ = \ashr_32s_16ns_32_7_1_U18.reset  ? 32'd0 : _182_;
assign _183_ = \ashr_32s_16ns_32_7_1_U18.ce  ? \ashr_32s_16ns_32_7_1_U18.din1_cast_array[3]  : \ashr_32s_16ns_32_7_1_U18.din1_cast_array[4] ;
assign _173_ = \ashr_32s_16ns_32_7_1_U18.reset  ? 16'h0000 : _183_;
assign _184_ = \ashr_32s_16ns_32_7_1_U18.ce  ? _196_ : \ashr_32s_16ns_32_7_1_U18.dout_array[4] ;
assign _179_ = \ashr_32s_16ns_32_7_1_U18.reset  ? 32'd0 : _184_;
assign _185_ = \ashr_32s_16ns_32_7_1_U18.ce  ? \ashr_32s_16ns_32_7_1_U18.din1_cast_array[2]  : \ashr_32s_16ns_32_7_1_U18.din1_cast_array[3] ;
assign _172_ = \ashr_32s_16ns_32_7_1_U18.reset  ? 16'h0000 : _185_;
assign _186_ = \ashr_32s_16ns_32_7_1_U18.ce  ? _195_ : \ashr_32s_16ns_32_7_1_U18.dout_array[3] ;
assign _178_ = \ashr_32s_16ns_32_7_1_U18.reset  ? 32'd0 : _186_;
assign _187_ = \ashr_32s_16ns_32_7_1_U18.ce  ? \ashr_32s_16ns_32_7_1_U18.din1_cast_array[1]  : \ashr_32s_16ns_32_7_1_U18.din1_cast_array[2] ;
assign _171_ = \ashr_32s_16ns_32_7_1_U18.reset  ? 16'h0000 : _187_;
assign _188_ = \ashr_32s_16ns_32_7_1_U18.ce  ? _194_ : \ashr_32s_16ns_32_7_1_U18.dout_array[2] ;
assign _177_ = \ashr_32s_16ns_32_7_1_U18.reset  ? 32'd0 : _188_;
assign _189_ = \ashr_32s_16ns_32_7_1_U18.ce  ? \ashr_32s_16ns_32_7_1_U18.din1_cast_array[0]  : \ashr_32s_16ns_32_7_1_U18.din1_cast_array[1] ;
assign _170_ = \ashr_32s_16ns_32_7_1_U18.reset  ? 16'h0000 : _189_;
assign _190_ = \ashr_32s_16ns_32_7_1_U18.ce  ? _193_ : \ashr_32s_16ns_32_7_1_U18.dout_array[1] ;
assign _176_ = \ashr_32s_16ns_32_7_1_U18.reset  ? 32'd0 : _190_;
assign _191_ = \ashr_32s_16ns_32_7_1_U18.ce  ? \ashr_32s_16ns_32_7_1_U18.din1 [15:0] : \ashr_32s_16ns_32_7_1_U18.din1_cast_array[0] ;
assign _169_ = \ashr_32s_16ns_32_7_1_U18.reset  ? 16'h0000 : _191_;
assign _192_ = \ashr_32s_16ns_32_7_1_U18.ce  ? \ashr_32s_16ns_32_7_1_U18.din0  : \ashr_32s_16ns_32_7_1_U18.dout_array[0] ;
assign _175_ = \ashr_32s_16ns_32_7_1_U18.reset  ? 32'd0 : _192_;
assign _193_ = $signed(\ashr_32s_16ns_32_7_1_U18.dout_array[0] ) >>> { \ashr_32s_16ns_32_7_1_U18.din1_cast_array[0] [15], 15'h0000 };
assign _194_ = $signed(\ashr_32s_16ns_32_7_1_U18.dout_array[1] ) >>> { \ashr_32s_16ns_32_7_1_U18.din1_cast_array[1] [14:12], 12'h000 };
assign _195_ = $signed(\ashr_32s_16ns_32_7_1_U18.dout_array[2] ) >>> { \ashr_32s_16ns_32_7_1_U18.din1_cast_array[2] [11:9], 9'h000 };
assign _196_ = $signed(\ashr_32s_16ns_32_7_1_U18.dout_array[3] ) >>> { \ashr_32s_16ns_32_7_1_U18.din1_cast_array[3] [8:6], 6'h00 };
assign _197_ = $signed(\ashr_32s_16ns_32_7_1_U18.dout_array[4] ) >>> { \ashr_32s_16ns_32_7_1_U18.din1_cast_array[4] [5:3], 3'h0 };
assign \ashr_32s_16ns_32_7_1_U18.dout  = $signed(\ashr_32s_16ns_32_7_1_U18.dout_array[5] ) >>> \ashr_32s_16ns_32_7_1_U18.din1_cast_array[5] [2:0];
always @(posedge \ashr_32s_32s_32_7_1_U8.clk )
\ashr_32s_32s_32_7_1_U8.dout_array[5]  <= _209_;
always @(posedge \ashr_32s_32s_32_7_1_U8.clk )
\ashr_32s_32s_32_7_1_U8.din1_cast_array[5]  <= _203_;
always @(posedge \ashr_32s_32s_32_7_1_U8.clk )
\ashr_32s_32s_32_7_1_U8.dout_array[4]  <= _208_;
always @(posedge \ashr_32s_32s_32_7_1_U8.clk )
\ashr_32s_32s_32_7_1_U8.din1_cast_array[4]  <= _202_;
always @(posedge \ashr_32s_32s_32_7_1_U8.clk )
\ashr_32s_32s_32_7_1_U8.dout_array[3]  <= _207_;
always @(posedge \ashr_32s_32s_32_7_1_U8.clk )
\ashr_32s_32s_32_7_1_U8.din1_cast_array[3]  <= _201_;
always @(posedge \ashr_32s_32s_32_7_1_U8.clk )
\ashr_32s_32s_32_7_1_U8.dout_array[2]  <= _206_;
always @(posedge \ashr_32s_32s_32_7_1_U8.clk )
\ashr_32s_32s_32_7_1_U8.din1_cast_array[2]  <= _200_;
always @(posedge \ashr_32s_32s_32_7_1_U8.clk )
\ashr_32s_32s_32_7_1_U8.dout_array[1]  <= _205_;
always @(posedge \ashr_32s_32s_32_7_1_U8.clk )
\ashr_32s_32s_32_7_1_U8.din1_cast_array[1]  <= _199_;
always @(posedge \ashr_32s_32s_32_7_1_U8.clk )
\ashr_32s_32s_32_7_1_U8.dout_array[0]  <= _204_;
always @(posedge \ashr_32s_32s_32_7_1_U8.clk )
\ashr_32s_32s_32_7_1_U8.din1_cast_array[0]  <= _198_;
assign _198_ = \ashr_32s_32s_32_7_1_U8.reset  ? 32'd0 : _221_;
assign _210_ = \ashr_32s_32s_32_7_1_U8.ce  ? _222_ : \ashr_32s_32s_32_7_1_U8.dout_array[0] ;
assign _204_ = \ashr_32s_32s_32_7_1_U8.reset  ? 32'd0 : _210_;
assign _211_ = \ashr_32s_32s_32_7_1_U8.ce  ? \ashr_32s_32s_32_7_1_U8.din1_cast_array[4]  : \ashr_32s_32s_32_7_1_U8.din1_cast_array[5] ;
assign _203_ = \ashr_32s_32s_32_7_1_U8.reset  ? 32'd0 : _211_;
assign _212_ = \ashr_32s_32s_32_7_1_U8.ce  ? _227_ : \ashr_32s_32s_32_7_1_U8.dout_array[5] ;
assign _209_ = \ashr_32s_32s_32_7_1_U8.reset  ? 32'd0 : _212_;
assign _213_ = \ashr_32s_32s_32_7_1_U8.ce  ? \ashr_32s_32s_32_7_1_U8.din1_cast_array[3]  : \ashr_32s_32s_32_7_1_U8.din1_cast_array[4] ;
assign _202_ = \ashr_32s_32s_32_7_1_U8.reset  ? 32'd0 : _213_;
assign _214_ = \ashr_32s_32s_32_7_1_U8.ce  ? _226_ : \ashr_32s_32s_32_7_1_U8.dout_array[4] ;
assign _208_ = \ashr_32s_32s_32_7_1_U8.reset  ? 32'd0 : _214_;
assign _215_ = \ashr_32s_32s_32_7_1_U8.ce  ? \ashr_32s_32s_32_7_1_U8.din1_cast_array[2]  : \ashr_32s_32s_32_7_1_U8.din1_cast_array[3] ;
assign _201_ = \ashr_32s_32s_32_7_1_U8.reset  ? 32'd0 : _215_;
assign _216_ = \ashr_32s_32s_32_7_1_U8.ce  ? _225_ : \ashr_32s_32s_32_7_1_U8.dout_array[3] ;
assign _207_ = \ashr_32s_32s_32_7_1_U8.reset  ? 32'd0 : _216_;
assign _217_ = \ashr_32s_32s_32_7_1_U8.ce  ? \ashr_32s_32s_32_7_1_U8.din1_cast_array[1]  : \ashr_32s_32s_32_7_1_U8.din1_cast_array[2] ;
assign _200_ = \ashr_32s_32s_32_7_1_U8.reset  ? 32'd0 : _217_;
assign _218_ = \ashr_32s_32s_32_7_1_U8.ce  ? _224_ : \ashr_32s_32s_32_7_1_U8.dout_array[2] ;
assign _206_ = \ashr_32s_32s_32_7_1_U8.reset  ? 32'd0 : _218_;
assign _219_ = \ashr_32s_32s_32_7_1_U8.ce  ? \ashr_32s_32s_32_7_1_U8.din1_cast_array[0]  : \ashr_32s_32s_32_7_1_U8.din1_cast_array[1] ;
assign _199_ = \ashr_32s_32s_32_7_1_U8.reset  ? 32'd0 : _219_;
assign _220_ = \ashr_32s_32s_32_7_1_U8.ce  ? _223_ : \ashr_32s_32s_32_7_1_U8.dout_array[1] ;
assign _205_ = \ashr_32s_32s_32_7_1_U8.reset  ? 32'd0 : _220_;
assign _221_ = \ashr_32s_32s_32_7_1_U8.ce  ? \ashr_32s_32s_32_7_1_U8.din1  : \ashr_32s_32s_32_7_1_U8.din1_cast_array[0] ;
assign _222_ = $signed(\ashr_32s_32s_32_7_1_U8.din0 ) >>> { \ashr_32s_32s_32_7_1_U8.din1 [31:30], 30'h00000000 };
assign _223_ = $signed(\ashr_32s_32s_32_7_1_U8.dout_array[0] ) >>> { \ashr_32s_32s_32_7_1_U8.din1_cast_array[0] [29:25], 25'h0000000 };
assign _224_ = $signed(\ashr_32s_32s_32_7_1_U8.dout_array[1] ) >>> { \ashr_32s_32s_32_7_1_U8.din1_cast_array[1] [24:20], 20'h00000 };
assign _225_ = $signed(\ashr_32s_32s_32_7_1_U8.dout_array[2] ) >>> { \ashr_32s_32s_32_7_1_U8.din1_cast_array[2] [19:15], 15'h0000 };
assign _226_ = $signed(\ashr_32s_32s_32_7_1_U8.dout_array[3] ) >>> { \ashr_32s_32s_32_7_1_U8.din1_cast_array[3] [14:10], 10'h000 };
assign _227_ = $signed(\ashr_32s_32s_32_7_1_U8.dout_array[4] ) >>> { \ashr_32s_32s_32_7_1_U8.din1_cast_array[4] [9:5], 5'h00 };
assign \ashr_32s_32s_32_7_1_U8.dout  = $signed(\ashr_32s_32s_32_7_1_U8.dout_array[5] ) >>> \ashr_32s_32s_32_7_1_U8.din1_cast_array[5] [4:0];
always @(posedge \shl_32s_16ns_32_7_1_U19.clk )
\shl_32s_16ns_32_7_1_U19.dout_array[5]  <= _239_;
always @(posedge \shl_32s_16ns_32_7_1_U19.clk )
\shl_32s_16ns_32_7_1_U19.din1_cast_array[5]  <= _233_;
always @(posedge \shl_32s_16ns_32_7_1_U19.clk )
\shl_32s_16ns_32_7_1_U19.dout_array[4]  <= _238_;
always @(posedge \shl_32s_16ns_32_7_1_U19.clk )
\shl_32s_16ns_32_7_1_U19.din1_cast_array[4]  <= _232_;
always @(posedge \shl_32s_16ns_32_7_1_U19.clk )
\shl_32s_16ns_32_7_1_U19.dout_array[3]  <= _237_;
always @(posedge \shl_32s_16ns_32_7_1_U19.clk )
\shl_32s_16ns_32_7_1_U19.din1_cast_array[3]  <= _231_;
always @(posedge \shl_32s_16ns_32_7_1_U19.clk )
\shl_32s_16ns_32_7_1_U19.dout_array[2]  <= _236_;
always @(posedge \shl_32s_16ns_32_7_1_U19.clk )
\shl_32s_16ns_32_7_1_U19.din1_cast_array[2]  <= _230_;
always @(posedge \shl_32s_16ns_32_7_1_U19.clk )
\shl_32s_16ns_32_7_1_U19.dout_array[1]  <= _235_;
always @(posedge \shl_32s_16ns_32_7_1_U19.clk )
\shl_32s_16ns_32_7_1_U19.din1_cast_array[1]  <= _229_;
always @(posedge \shl_32s_16ns_32_7_1_U19.clk )
\shl_32s_16ns_32_7_1_U19.dout_array[0]  <= _234_;
always @(posedge \shl_32s_16ns_32_7_1_U19.clk )
\shl_32s_16ns_32_7_1_U19.din1_cast_array[0]  <= _228_;
assign _240_ = \shl_32s_16ns_32_7_1_U19.ce  ? \shl_32s_16ns_32_7_1_U19.din1_cast_array[4]  : \shl_32s_16ns_32_7_1_U19.din1_cast_array[5] ;
assign _233_ = \shl_32s_16ns_32_7_1_U19.reset  ? 16'h0000 : _240_;
assign _241_ = \shl_32s_16ns_32_7_1_U19.ce  ? _256_ : \shl_32s_16ns_32_7_1_U19.dout_array[5] ;
assign _239_ = \shl_32s_16ns_32_7_1_U19.reset  ? 32'd0 : _241_;
assign _242_ = \shl_32s_16ns_32_7_1_U19.ce  ? \shl_32s_16ns_32_7_1_U19.din1_cast_array[3]  : \shl_32s_16ns_32_7_1_U19.din1_cast_array[4] ;
assign _232_ = \shl_32s_16ns_32_7_1_U19.reset  ? 16'h0000 : _242_;
assign _243_ = \shl_32s_16ns_32_7_1_U19.ce  ? _255_ : \shl_32s_16ns_32_7_1_U19.dout_array[4] ;
assign _238_ = \shl_32s_16ns_32_7_1_U19.reset  ? 32'd0 : _243_;
assign _244_ = \shl_32s_16ns_32_7_1_U19.ce  ? \shl_32s_16ns_32_7_1_U19.din1_cast_array[2]  : \shl_32s_16ns_32_7_1_U19.din1_cast_array[3] ;
assign _231_ = \shl_32s_16ns_32_7_1_U19.reset  ? 16'h0000 : _244_;
assign _245_ = \shl_32s_16ns_32_7_1_U19.ce  ? _254_ : \shl_32s_16ns_32_7_1_U19.dout_array[3] ;
assign _237_ = \shl_32s_16ns_32_7_1_U19.reset  ? 32'd0 : _245_;
assign _246_ = \shl_32s_16ns_32_7_1_U19.ce  ? \shl_32s_16ns_32_7_1_U19.din1_cast_array[1]  : \shl_32s_16ns_32_7_1_U19.din1_cast_array[2] ;
assign _230_ = \shl_32s_16ns_32_7_1_U19.reset  ? 16'h0000 : _246_;
assign _247_ = \shl_32s_16ns_32_7_1_U19.ce  ? _253_ : \shl_32s_16ns_32_7_1_U19.dout_array[2] ;
assign _236_ = \shl_32s_16ns_32_7_1_U19.reset  ? 32'd0 : _247_;
assign _248_ = \shl_32s_16ns_32_7_1_U19.ce  ? \shl_32s_16ns_32_7_1_U19.din1_cast_array[0]  : \shl_32s_16ns_32_7_1_U19.din1_cast_array[1] ;
assign _229_ = \shl_32s_16ns_32_7_1_U19.reset  ? 16'h0000 : _248_;
assign _249_ = \shl_32s_16ns_32_7_1_U19.ce  ? _252_ : \shl_32s_16ns_32_7_1_U19.dout_array[1] ;
assign _235_ = \shl_32s_16ns_32_7_1_U19.reset  ? 32'd0 : _249_;
assign _250_ = \shl_32s_16ns_32_7_1_U19.ce  ? \shl_32s_16ns_32_7_1_U19.din1 [15:0] : \shl_32s_16ns_32_7_1_U19.din1_cast_array[0] ;
assign _228_ = \shl_32s_16ns_32_7_1_U19.reset  ? 16'h0000 : _250_;
assign _251_ = \shl_32s_16ns_32_7_1_U19.ce  ? \shl_32s_16ns_32_7_1_U19.din0  : \shl_32s_16ns_32_7_1_U19.dout_array[0] ;
assign _234_ = \shl_32s_16ns_32_7_1_U19.reset  ? 32'd0 : _251_;
assign _252_ = \shl_32s_16ns_32_7_1_U19.dout_array[0]  << { \shl_32s_16ns_32_7_1_U19.din1_cast_array[0] [15], 15'h0000 };
assign _253_ = \shl_32s_16ns_32_7_1_U19.dout_array[1]  << { \shl_32s_16ns_32_7_1_U19.din1_cast_array[1] [14:12], 12'h000 };
assign _254_ = \shl_32s_16ns_32_7_1_U19.dout_array[2]  << { \shl_32s_16ns_32_7_1_U19.din1_cast_array[2] [11:9], 9'h000 };
assign _255_ = \shl_32s_16ns_32_7_1_U19.dout_array[3]  << { \shl_32s_16ns_32_7_1_U19.din1_cast_array[3] [8:6], 6'h00 };
assign _256_ = \shl_32s_16ns_32_7_1_U19.dout_array[4]  << { \shl_32s_16ns_32_7_1_U19.din1_cast_array[4] [5:3], 3'h0 };
assign \shl_32s_16ns_32_7_1_U19.dout  = \shl_32s_16ns_32_7_1_U19.dout_array[5]  << \shl_32s_16ns_32_7_1_U19.din1_cast_array[5] [2:0];
always @(posedge \shl_32s_32s_32_7_1_U7.clk )
\shl_32s_32s_32_7_1_U7.dout_array[5]  <= _268_;
always @(posedge \shl_32s_32s_32_7_1_U7.clk )
\shl_32s_32s_32_7_1_U7.din1_cast_array[5]  <= _262_;
always @(posedge \shl_32s_32s_32_7_1_U7.clk )
\shl_32s_32s_32_7_1_U7.dout_array[4]  <= _267_;
always @(posedge \shl_32s_32s_32_7_1_U7.clk )
\shl_32s_32s_32_7_1_U7.din1_cast_array[4]  <= _261_;
always @(posedge \shl_32s_32s_32_7_1_U7.clk )
\shl_32s_32s_32_7_1_U7.dout_array[3]  <= _266_;
always @(posedge \shl_32s_32s_32_7_1_U7.clk )
\shl_32s_32s_32_7_1_U7.din1_cast_array[3]  <= _260_;
always @(posedge \shl_32s_32s_32_7_1_U7.clk )
\shl_32s_32s_32_7_1_U7.dout_array[2]  <= _265_;
always @(posedge \shl_32s_32s_32_7_1_U7.clk )
\shl_32s_32s_32_7_1_U7.din1_cast_array[2]  <= _259_;
always @(posedge \shl_32s_32s_32_7_1_U7.clk )
\shl_32s_32s_32_7_1_U7.dout_array[1]  <= _264_;
always @(posedge \shl_32s_32s_32_7_1_U7.clk )
\shl_32s_32s_32_7_1_U7.din1_cast_array[1]  <= _258_;
always @(posedge \shl_32s_32s_32_7_1_U7.clk )
\shl_32s_32s_32_7_1_U7.dout_array[0]  <= _263_;
always @(posedge \shl_32s_32s_32_7_1_U7.clk )
\shl_32s_32s_32_7_1_U7.din1_cast_array[0]  <= _257_;
assign _269_ = \shl_32s_32s_32_7_1_U7.ce  ? \shl_32s_32s_32_7_1_U7.din1_cast_array[4]  : \shl_32s_32s_32_7_1_U7.din1_cast_array[5] ;
assign _262_ = \shl_32s_32s_32_7_1_U7.reset  ? 32'd0 : _269_;
assign _270_ = \shl_32s_32s_32_7_1_U7.ce  ? _286_ : \shl_32s_32s_32_7_1_U7.dout_array[5] ;
assign _268_ = \shl_32s_32s_32_7_1_U7.reset  ? 32'd0 : _270_;
assign _271_ = \shl_32s_32s_32_7_1_U7.ce  ? \shl_32s_32s_32_7_1_U7.din1_cast_array[3]  : \shl_32s_32s_32_7_1_U7.din1_cast_array[4] ;
assign _261_ = \shl_32s_32s_32_7_1_U7.reset  ? 32'd0 : _271_;
assign _272_ = \shl_32s_32s_32_7_1_U7.ce  ? _285_ : \shl_32s_32s_32_7_1_U7.dout_array[4] ;
assign _267_ = \shl_32s_32s_32_7_1_U7.reset  ? 32'd0 : _272_;
assign _273_ = \shl_32s_32s_32_7_1_U7.ce  ? \shl_32s_32s_32_7_1_U7.din1_cast_array[2]  : \shl_32s_32s_32_7_1_U7.din1_cast_array[3] ;
assign _260_ = \shl_32s_32s_32_7_1_U7.reset  ? 32'd0 : _273_;
assign _274_ = \shl_32s_32s_32_7_1_U7.ce  ? _284_ : \shl_32s_32s_32_7_1_U7.dout_array[3] ;
assign _266_ = \shl_32s_32s_32_7_1_U7.reset  ? 32'd0 : _274_;
assign _275_ = \shl_32s_32s_32_7_1_U7.ce  ? \shl_32s_32s_32_7_1_U7.din1_cast_array[1]  : \shl_32s_32s_32_7_1_U7.din1_cast_array[2] ;
assign _259_ = \shl_32s_32s_32_7_1_U7.reset  ? 32'd0 : _275_;
assign _276_ = \shl_32s_32s_32_7_1_U7.ce  ? _283_ : \shl_32s_32s_32_7_1_U7.dout_array[2] ;
assign _265_ = \shl_32s_32s_32_7_1_U7.reset  ? 32'd0 : _276_;
assign _277_ = \shl_32s_32s_32_7_1_U7.ce  ? \shl_32s_32s_32_7_1_U7.din1_cast_array[0]  : \shl_32s_32s_32_7_1_U7.din1_cast_array[1] ;
assign _258_ = \shl_32s_32s_32_7_1_U7.reset  ? 32'd0 : _277_;
assign _278_ = \shl_32s_32s_32_7_1_U7.ce  ? _282_ : \shl_32s_32s_32_7_1_U7.dout_array[1] ;
assign _264_ = \shl_32s_32s_32_7_1_U7.reset  ? 32'd0 : _278_;
assign _279_ = \shl_32s_32s_32_7_1_U7.ce  ? \shl_32s_32s_32_7_1_U7.din1  : \shl_32s_32s_32_7_1_U7.din1_cast_array[0] ;
assign _257_ = \shl_32s_32s_32_7_1_U7.reset  ? 32'd0 : _279_;
assign _280_ = \shl_32s_32s_32_7_1_U7.ce  ? _281_ : \shl_32s_32s_32_7_1_U7.dout_array[0] ;
assign _263_ = \shl_32s_32s_32_7_1_U7.reset  ? 32'd0 : _280_;
assign _281_ = \shl_32s_32s_32_7_1_U7.din0  << { \shl_32s_32s_32_7_1_U7.din1 [31:30], 30'h00000000 };
assign _282_ = \shl_32s_32s_32_7_1_U7.dout_array[0]  << { \shl_32s_32s_32_7_1_U7.din1_cast_array[0] [29:25], 25'h0000000 };
assign _283_ = \shl_32s_32s_32_7_1_U7.dout_array[1]  << { \shl_32s_32s_32_7_1_U7.din1_cast_array[1] [24:20], 20'h00000 };
assign _284_ = \shl_32s_32s_32_7_1_U7.dout_array[2]  << { \shl_32s_32s_32_7_1_U7.din1_cast_array[2] [19:15], 15'h0000 };
assign _285_ = \shl_32s_32s_32_7_1_U7.dout_array[3]  << { \shl_32s_32s_32_7_1_U7.din1_cast_array[3] [14:10], 10'h000 };
assign _286_ = \shl_32s_32s_32_7_1_U7.dout_array[4]  << { \shl_32s_32s_32_7_1_U7.din1_cast_array[4] [9:5], 5'h00 };
assign \shl_32s_32s_32_7_1_U7.dout  = \shl_32s_32s_32_7_1_U7.dout_array[5]  << \shl_32s_32s_32_7_1_U7.din1_cast_array[5] [4:0];
always @(posedge \shl_32s_8ns_32_7_1_U2.clk )
\shl_32s_8ns_32_7_1_U2.dout_array[5]  <= _298_;
always @(posedge \shl_32s_8ns_32_7_1_U2.clk )
\shl_32s_8ns_32_7_1_U2.din1_cast_array[5]  <= _292_;
always @(posedge \shl_32s_8ns_32_7_1_U2.clk )
\shl_32s_8ns_32_7_1_U2.dout_array[4]  <= _297_;
always @(posedge \shl_32s_8ns_32_7_1_U2.clk )
\shl_32s_8ns_32_7_1_U2.din1_cast_array[4]  <= _291_;
always @(posedge \shl_32s_8ns_32_7_1_U2.clk )
\shl_32s_8ns_32_7_1_U2.dout_array[3]  <= _296_;
always @(posedge \shl_32s_8ns_32_7_1_U2.clk )
\shl_32s_8ns_32_7_1_U2.din1_cast_array[3]  <= _290_;
always @(posedge \shl_32s_8ns_32_7_1_U2.clk )
\shl_32s_8ns_32_7_1_U2.dout_array[2]  <= _295_;
always @(posedge \shl_32s_8ns_32_7_1_U2.clk )
\shl_32s_8ns_32_7_1_U2.din1_cast_array[2]  <= _289_;
always @(posedge \shl_32s_8ns_32_7_1_U2.clk )
\shl_32s_8ns_32_7_1_U2.dout_array[1]  <= _294_;
always @(posedge \shl_32s_8ns_32_7_1_U2.clk )
\shl_32s_8ns_32_7_1_U2.din1_cast_array[1]  <= _288_;
always @(posedge \shl_32s_8ns_32_7_1_U2.clk )
\shl_32s_8ns_32_7_1_U2.dout_array[0]  <= _293_;
always @(posedge \shl_32s_8ns_32_7_1_U2.clk )
\shl_32s_8ns_32_7_1_U2.din1_cast_array[0]  <= _287_;
assign _299_ = \shl_32s_8ns_32_7_1_U2.ce  ? \shl_32s_8ns_32_7_1_U2.din1_cast_array[4]  : \shl_32s_8ns_32_7_1_U2.din1_cast_array[5] ;
assign _292_ = \shl_32s_8ns_32_7_1_U2.reset  ? 8'h00 : _299_;
assign _300_ = \shl_32s_8ns_32_7_1_U2.ce  ? _313_ : \shl_32s_8ns_32_7_1_U2.dout_array[5] ;
assign _298_ = \shl_32s_8ns_32_7_1_U2.reset  ? 32'd0 : _300_;
assign _301_ = \shl_32s_8ns_32_7_1_U2.ce  ? \shl_32s_8ns_32_7_1_U2.din1_cast_array[3]  : \shl_32s_8ns_32_7_1_U2.din1_cast_array[4] ;
assign _291_ = \shl_32s_8ns_32_7_1_U2.reset  ? 8'h00 : _301_;
assign _302_ = \shl_32s_8ns_32_7_1_U2.ce  ? _312_ : \shl_32s_8ns_32_7_1_U2.dout_array[4] ;
assign _297_ = \shl_32s_8ns_32_7_1_U2.reset  ? 32'd0 : _302_;
assign _303_ = \shl_32s_8ns_32_7_1_U2.ce  ? \shl_32s_8ns_32_7_1_U2.din1_cast_array[2]  : \shl_32s_8ns_32_7_1_U2.din1_cast_array[3] ;
assign _290_ = \shl_32s_8ns_32_7_1_U2.reset  ? 8'h00 : _303_;
assign _304_ = \shl_32s_8ns_32_7_1_U2.ce  ? _311_ : \shl_32s_8ns_32_7_1_U2.dout_array[3] ;
assign _296_ = \shl_32s_8ns_32_7_1_U2.reset  ? 32'd0 : _304_;
assign _305_ = \shl_32s_8ns_32_7_1_U2.ce  ? \shl_32s_8ns_32_7_1_U2.din1_cast_array[1]  : \shl_32s_8ns_32_7_1_U2.din1_cast_array[2] ;
assign _289_ = \shl_32s_8ns_32_7_1_U2.reset  ? 8'h00 : _305_;
assign _306_ = \shl_32s_8ns_32_7_1_U2.ce  ? \shl_32s_8ns_32_7_1_U2.dout_array[1]  : \shl_32s_8ns_32_7_1_U2.dout_array[2] ;
assign _295_ = \shl_32s_8ns_32_7_1_U2.reset  ? 32'd0 : _306_;
assign _307_ = \shl_32s_8ns_32_7_1_U2.ce  ? \shl_32s_8ns_32_7_1_U2.din1_cast_array[0]  : \shl_32s_8ns_32_7_1_U2.din1_cast_array[1] ;
assign _288_ = \shl_32s_8ns_32_7_1_U2.reset  ? 8'h00 : _307_;
assign _308_ = \shl_32s_8ns_32_7_1_U2.ce  ? \shl_32s_8ns_32_7_1_U2.dout_array[0]  : \shl_32s_8ns_32_7_1_U2.dout_array[1] ;
assign _294_ = \shl_32s_8ns_32_7_1_U2.reset  ? 32'd0 : _308_;
assign _309_ = \shl_32s_8ns_32_7_1_U2.ce  ? \shl_32s_8ns_32_7_1_U2.din1 [7:0] : \shl_32s_8ns_32_7_1_U2.din1_cast_array[0] ;
assign _287_ = \shl_32s_8ns_32_7_1_U2.reset  ? 8'h00 : _309_;
assign _310_ = \shl_32s_8ns_32_7_1_U2.ce  ? \shl_32s_8ns_32_7_1_U2.din0  : \shl_32s_8ns_32_7_1_U2.dout_array[0] ;
assign _293_ = \shl_32s_8ns_32_7_1_U2.reset  ? 32'd0 : _310_;
assign _311_ = \shl_32s_8ns_32_7_1_U2.dout_array[2]  << { \shl_32s_8ns_32_7_1_U2.din1_cast_array[2] [7:6], 6'h00 };
assign _312_ = \shl_32s_8ns_32_7_1_U2.dout_array[3]  << { \shl_32s_8ns_32_7_1_U2.din1_cast_array[3] [5:4], 4'h0 };
assign _313_ = \shl_32s_8ns_32_7_1_U2.dout_array[4]  << { \shl_32s_8ns_32_7_1_U2.din1_cast_array[4] [3:2], 2'h0 };
assign \shl_32s_8ns_32_7_1_U2.dout  = \shl_32s_8ns_32_7_1_U2.dout_array[5]  << \shl_32s_8ns_32_7_1_U2.din1_cast_array[5] [1:0];
assign \sub_4ns_4s_4_2_1_U17.top_sub_4ns_4s_4_2_1_Adder_11_U.bin_s0  = ~ \sub_4ns_4s_4_2_1_U17.top_sub_4ns_4s_4_2_1_Adder_11_U.b ;
always @(posedge \sub_4ns_4s_4_2_1_U17.top_sub_4ns_4s_4_2_1_Adder_11_U.clk )
\sub_4ns_4s_4_2_1_U17.top_sub_4ns_4s_4_2_1_Adder_11_U.bin_s1  <= _315_;
always @(posedge \sub_4ns_4s_4_2_1_U17.top_sub_4ns_4s_4_2_1_Adder_11_U.clk )
\sub_4ns_4s_4_2_1_U17.top_sub_4ns_4s_4_2_1_Adder_11_U.ain_s1  <= _314_;
always @(posedge \sub_4ns_4s_4_2_1_U17.top_sub_4ns_4s_4_2_1_Adder_11_U.clk )
\sub_4ns_4s_4_2_1_U17.top_sub_4ns_4s_4_2_1_Adder_11_U.sum_s1  <= _317_;
always @(posedge \sub_4ns_4s_4_2_1_U17.top_sub_4ns_4s_4_2_1_Adder_11_U.clk )
\sub_4ns_4s_4_2_1_U17.top_sub_4ns_4s_4_2_1_Adder_11_U.carry_s1  <= _316_;
assign _315_ = \sub_4ns_4s_4_2_1_U17.top_sub_4ns_4s_4_2_1_Adder_11_U.ce  ? \sub_4ns_4s_4_2_1_U17.top_sub_4ns_4s_4_2_1_Adder_11_U.bin_s0 [3:2] : \sub_4ns_4s_4_2_1_U17.top_sub_4ns_4s_4_2_1_Adder_11_U.bin_s1 ;
assign _314_ = \sub_4ns_4s_4_2_1_U17.top_sub_4ns_4s_4_2_1_Adder_11_U.ce  ? \sub_4ns_4s_4_2_1_U17.top_sub_4ns_4s_4_2_1_Adder_11_U.a [3:2] : \sub_4ns_4s_4_2_1_U17.top_sub_4ns_4s_4_2_1_Adder_11_U.ain_s1 ;
assign _316_ = \sub_4ns_4s_4_2_1_U17.top_sub_4ns_4s_4_2_1_Adder_11_U.ce  ? \sub_4ns_4s_4_2_1_U17.top_sub_4ns_4s_4_2_1_Adder_11_U.facout_s1  : \sub_4ns_4s_4_2_1_U17.top_sub_4ns_4s_4_2_1_Adder_11_U.carry_s1 ;
assign _317_ = \sub_4ns_4s_4_2_1_U17.top_sub_4ns_4s_4_2_1_Adder_11_U.ce  ? \sub_4ns_4s_4_2_1_U17.top_sub_4ns_4s_4_2_1_Adder_11_U.fas_s1  : \sub_4ns_4s_4_2_1_U17.top_sub_4ns_4s_4_2_1_Adder_11_U.sum_s1 ;
assign _318_ = \sub_4ns_4s_4_2_1_U17.top_sub_4ns_4s_4_2_1_Adder_11_U.u1.a  + \sub_4ns_4s_4_2_1_U17.top_sub_4ns_4s_4_2_1_Adder_11_U.u1.b ;
assign { \sub_4ns_4s_4_2_1_U17.top_sub_4ns_4s_4_2_1_Adder_11_U.u1.cout , \sub_4ns_4s_4_2_1_U17.top_sub_4ns_4s_4_2_1_Adder_11_U.u1.s  } = _318_ + \sub_4ns_4s_4_2_1_U17.top_sub_4ns_4s_4_2_1_Adder_11_U.u1.cin ;
assign _319_ = \sub_4ns_4s_4_2_1_U17.top_sub_4ns_4s_4_2_1_Adder_11_U.u2.a  + \sub_4ns_4s_4_2_1_U17.top_sub_4ns_4s_4_2_1_Adder_11_U.u2.b ;
assign { \sub_4ns_4s_4_2_1_U17.top_sub_4ns_4s_4_2_1_Adder_11_U.u2.cout , \sub_4ns_4s_4_2_1_U17.top_sub_4ns_4s_4_2_1_Adder_11_U.u2.s  } = _319_ + \sub_4ns_4s_4_2_1_U17.top_sub_4ns_4s_4_2_1_Adder_11_U.u2.cin ;
assign \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.bin_s0  = ~ \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.b ;
always @(posedge \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.clk )
\sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.bin_s1  <= _321_;
always @(posedge \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.clk )
\sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.ain_s1  <= _320_;
always @(posedge \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.clk )
\sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.sum_s1  <= _323_;
always @(posedge \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.clk )
\sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.carry_s1  <= _322_;
assign _321_ = \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.ce  ? \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.bin_s0 [4:2] : \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.bin_s1 ;
assign _320_ = \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.ce  ? \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.a [4:2] : \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.ain_s1 ;
assign _322_ = \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.ce  ? \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.facout_s1  : \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.carry_s1 ;
assign _323_ = \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.ce  ? \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.fas_s1  : \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.sum_s1 ;
assign _324_ = \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.u1.a  + \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.u1.b ;
assign { \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.u1.cout , \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.u1.s  } = _324_ + \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.u1.cin ;
assign _325_ = \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.u2.a  + \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.u2.b ;
assign { \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.u2.cout , \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.u2.s  } = _325_ + \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.u2.cin ;
assign _326_ = op_2 != 1'h1;
assign _327_ = | op_18[1:0];
always @(posedge ap_clk)
trunc_ln769_reg_1031 <= _049_;
always @(posedge ap_clk)
trunc_ln546_reg_1026 <= _048_;
always @(posedge ap_clk)
sub_ln1367_reg_803 <= _045_;
always @(posedge ap_clk)
shl_ln1299_1_reg_932 <= _043_;
always @(posedge ap_clk)
sh_V_1_reg_1005 <= _042_;
always @(posedge ap_clk)
ret_V_9_reg_862 <= _035_;
always @(posedge ap_clk)
ret_V_5_reg_808 <= _033_;
always @(posedge ap_clk)
ret_V_8_reg_813 <= _034_;
always @(posedge ap_clk)
trunc_ln851_2_reg_818 <= _051_;
always @(posedge ap_clk)
ush_reg_823 <= _052_;
always @(posedge ap_clk)
shl_ln1299_reg_775 <= _044_;
always @(posedge ap_clk)
ret_V_3_reg_780 <= _032_;
always @(posedge ap_clk)
trunc_ln851_1_reg_787 <= _050_;
always @(posedge ap_clk)
sext_ln1386_reg_792 <= _040_;
always @(posedge ap_clk)
ret_V_2_reg_748 <= _030_;
always @(posedge ap_clk)
ret_V_28_reg_1076 <= _029_;
always @(posedge ap_clk)
ret_V_30_cast_reg_1081 <= _031_;
always @(posedge ap_clk)
ret_V_27_reg_1056 <= _028_;
always @(posedge ap_clk)
ret_V_26_reg_1000 <= _027_;
always @(posedge ap_clk)
ret_V_25_reg_965 <= _026_;
always @(posedge ap_clk)
ret_V_20_reg_753 <= _022_;
always @(posedge ap_clk)
trunc_ln1348_reg_759 <= _047_;
always @(posedge ap_clk)
ret_V_19_reg_736 <= _021_;
always @(posedge ap_clk)
ret_V_reg_741 <= _036_;
always @(posedge ap_clk)
ret_V_12_reg_973 <= _020_;
always @(posedge ap_clk)
select_ln1368_reg_952 <= _039_;
always @(posedge ap_clk)
ret_V_11_reg_958 <= _019_;
always @(posedge ap_clk)
ret_V_24_reg_978 <= _025_;
always @(posedge ap_clk)
p_Result_8_reg_985 <= _017_;
always @(posedge ap_clk)
r_reg_1041 <= _018_;
always @(posedge ap_clk)
op_27_V_reg_1046 <= _015_;
always @(posedge ap_clk)
op_24_V_reg_942 <= _014_;
always @(posedge ap_clk)
select_ln1192_reg_947 <= _038_;
always @(posedge ap_clk)
op_7_V_reg_764 <= _016_;
always @(posedge ap_clk)
isNeg_reg_769 <= _012_;
always @(posedge ap_clk)
icmp_ln851_3_reg_1071 <= _010_;
always @(posedge ap_clk)
ret_V_21_reg_828 <= _023_;
always @(posedge ap_clk)
lhs_V_2_reg_833 <= _013_;
always @(posedge ap_clk)
sext_ln831_reg_838 <= _041_;
always @(posedge ap_clk)
icmp_ln851_2_reg_845 <= _009_;
always @(posedge ap_clk)
icmp_ln851_1_reg_798 <= _008_;
always @(posedge ap_clk)
icmp_ln851_reg_711 <= _011_;
always @(posedge ap_clk)
icmp_ln1499_reg_726 <= _007_;
always @(posedge ap_clk)
trunc_ln1348_1_reg_731 <= _046_;
always @(posedge ap_clk)
ashr_ln1333_reg_937 <= _006_;
always @(posedge ap_clk)
add_ln69_reg_917 <= _004_;
always @(posedge ap_clk)
add_ln69_2_reg_922 <= _003_;
always @(posedge ap_clk)
ret_V_23_reg_887 <= _024_;
always @(posedge ap_clk)
ret_reg_892 <= _037_;
always @(posedge ap_clk)
add_ln69_1_reg_897 <= _002_;
always @(posedge ap_clk)
add_ln691_reg_990 <= _001_;
always @(posedge ap_clk)
add_ln691_1_reg_1088 <= _000_;
always @(posedge ap_clk)
ap_CS_fsm <= _005_;
assign _053_ = _064_ ? 2'h2 : 2'h1;
assign _328_ = ap_CS_fsm == 1'h1;
function [36:0] _871_;
input [36:0] a;
input [1368:0] b;
input [36:0] s;
case (s)
37'b0000000000000000000000000000000000001:
_871_ = b[36:0];
37'b0000000000000000000000000000000000010:
_871_ = b[73:37];
37'b0000000000000000000000000000000000100:
_871_ = b[110:74];
37'b0000000000000000000000000000000001000:
_871_ = b[147:111];
37'b0000000000000000000000000000000010000:
_871_ = b[184:148];
37'b0000000000000000000000000000000100000:
_871_ = b[221:185];
37'b0000000000000000000000000000001000000:
_871_ = b[258:222];
37'b0000000000000000000000000000010000000:
_871_ = b[295:259];
37'b0000000000000000000000000000100000000:
_871_ = b[332:296];
37'b0000000000000000000000000001000000000:
_871_ = b[369:333];
37'b0000000000000000000000000010000000000:
_871_ = b[406:370];
37'b0000000000000000000000000100000000000:
_871_ = b[443:407];
37'b0000000000000000000000001000000000000:
_871_ = b[480:444];
37'b0000000000000000000000010000000000000:
_871_ = b[517:481];
37'b0000000000000000000000100000000000000:
_871_ = b[554:518];
37'b0000000000000000000001000000000000000:
_871_ = b[591:555];
37'b0000000000000000000010000000000000000:
_871_ = b[628:592];
37'b0000000000000000000100000000000000000:
_871_ = b[665:629];
37'b0000000000000000001000000000000000000:
_871_ = b[702:666];
37'b0000000000000000010000000000000000000:
_871_ = b[739:703];
37'b0000000000000000100000000000000000000:
_871_ = b[776:740];
37'b0000000000000001000000000000000000000:
_871_ = b[813:777];
37'b0000000000000010000000000000000000000:
_871_ = b[850:814];
37'b0000000000000100000000000000000000000:
_871_ = b[887:851];
37'b0000000000001000000000000000000000000:
_871_ = b[924:888];
37'b0000000000010000000000000000000000000:
_871_ = b[961:925];
37'b0000000000100000000000000000000000000:
_871_ = b[998:962];
37'b0000000001000000000000000000000000000:
_871_ = b[1035:999];
37'b0000000010000000000000000000000000000:
_871_ = b[1072:1036];
37'b0000000100000000000000000000000000000:
_871_ = b[1109:1073];
37'b0000001000000000000000000000000000000:
_871_ = b[1146:1110];
37'b0000010000000000000000000000000000000:
_871_ = b[1183:1147];
37'b0000100000000000000000000000000000000:
_871_ = b[1220:1184];
37'b0001000000000000000000000000000000000:
_871_ = b[1257:1221];
37'b0010000000000000000000000000000000000:
_871_ = b[1294:1258];
37'b0100000000000000000000000000000000000:
_871_ = b[1331:1295];
37'b1000000000000000000000000000000000000:
_871_ = b[1368:1332];
37'b0000000000000000000000000000000000000:
_871_ = a;
default:
_871_ = 37'bx;
endcase
endfunction
assign ap_NS_fsm = _871_(37'hxxxxxxxxxx, { 35'h000000000, _053_, 1332'h000000002000000002000000002000000002000000002000000002000000002000000002000000002000000002000000002000000002000000002000000002000000002000000002000000002000000002000000002000000002000000002000000002000000002000000002000000002000000002000000002000000002000000002000000002000000002000000002000000002000000002000000002000000000000000001 }, { _328_, _364_, _363_, _362_, _361_, _360_, _359_, _358_, _357_, _356_, _355_, _354_, _353_, _352_, _351_, _350_, _349_, _348_, _347_, _346_, _345_, _344_, _343_, _342_, _341_, _340_, _339_, _338_, _337_, _336_, _335_, _334_, _333_, _332_, _331_, _330_, _329_ });
assign _329_ = ap_CS_fsm == 37'h1000000000;
assign _330_ = ap_CS_fsm == 36'h800000000;
assign _331_ = ap_CS_fsm == 35'h400000000;
assign _332_ = ap_CS_fsm == 34'h200000000;
assign _333_ = ap_CS_fsm == 33'h100000000;
assign _334_ = ap_CS_fsm == 32'd2147483648;
assign _335_ = ap_CS_fsm == 31'h40000000;
assign _336_ = ap_CS_fsm == 30'h20000000;
assign _337_ = ap_CS_fsm == 29'h10000000;
assign _338_ = ap_CS_fsm == 28'h8000000;
assign _339_ = ap_CS_fsm == 27'h4000000;
assign _340_ = ap_CS_fsm == 26'h2000000;
assign _341_ = ap_CS_fsm == 25'h1000000;
assign _342_ = ap_CS_fsm == 24'h800000;
assign _343_ = ap_CS_fsm == 23'h400000;
assign _344_ = ap_CS_fsm == 22'h200000;
assign _345_ = ap_CS_fsm == 21'h100000;
assign _346_ = ap_CS_fsm == 20'h80000;
assign _347_ = ap_CS_fsm == 19'h40000;
assign _348_ = ap_CS_fsm == 18'h20000;
assign _349_ = ap_CS_fsm == 17'h10000;
assign _350_ = ap_CS_fsm == 16'h8000;
assign _351_ = ap_CS_fsm == 15'h4000;
assign _352_ = ap_CS_fsm == 14'h2000;
assign _353_ = ap_CS_fsm == 13'h1000;
assign _354_ = ap_CS_fsm == 12'h800;
assign _355_ = ap_CS_fsm == 11'h400;
assign _356_ = ap_CS_fsm == 10'h200;
assign _357_ = ap_CS_fsm == 9'h100;
assign _358_ = ap_CS_fsm == 8'h80;
assign _359_ = ap_CS_fsm == 7'h40;
assign _360_ = ap_CS_fsm == 6'h20;
assign _361_ = ap_CS_fsm == 5'h10;
assign _362_ = ap_CS_fsm == 4'h8;
assign _363_ = ap_CS_fsm == 3'h4;
assign _364_ = ap_CS_fsm == 2'h2;
assign op_30_ap_vld = ap_CS_fsm[36] ? 1'h1 : 1'h0;
assign ap_idle = _063_ ? 1'h1 : 1'h0;
assign _049_ = _062_ ? grp_fu_595_p2[5:0] : trunc_ln769_reg_1031;
assign _048_ = _061_ ? grp_fu_582_p2[2:0] : trunc_ln546_reg_1026;
assign _045_ = _060_ ? grp_fu_296_p2 : sub_ln1367_reg_803;
assign _043_ = _059_ ? grp_fu_390_p2 : shl_ln1299_1_reg_932;
assign _042_ = _058_ ? grp_fu_547_p2 : sh_V_1_reg_1005;
assign _035_ = ap_CS_fsm[10] ? grp_fu_377_p2 : ret_V_9_reg_862;
assign _052_ = ap_CS_fsm[8] ? ush_fu_339_p3 : ush_reg_823;
assign _051_ = ap_CS_fsm[8] ? 2'h0 : trunc_ln851_2_reg_818;
assign _034_ = ap_CS_fsm[8] ? { ret_V_20_reg_753[9:1], ret_V_22_fu_319_p2[2] } : ret_V_8_reg_813;
assign _033_ = ap_CS_fsm[8] ? grp_fu_307_p2 : ret_V_5_reg_808;
assign _040_ = ap_CS_fsm[6] ? { op_7_V_reg_764[3], op_7_V_reg_764 } : sext_ln1386_reg_792;
assign _050_ = ap_CS_fsm[6] ? grp_fu_213_p2[1:0] : trunc_ln851_1_reg_787;
assign _032_ = ap_CS_fsm[6] ? grp_fu_213_p2[3:2] : ret_V_3_reg_780;
assign _044_ = ap_CS_fsm[6] ? grp_fu_213_p2 : shl_ln1299_reg_775;
assign _030_ = _057_ ? grp_fu_239_p2 : ret_V_2_reg_748;
assign _031_ = ap_CS_fsm[33] ? grp_fu_650_p2[33:2] : ret_V_30_cast_reg_1081;
assign _029_ = ap_CS_fsm[33] ? grp_fu_650_p2 : ret_V_28_reg_1076;
assign _028_ = ap_CS_fsm[31] ? grp_fu_630_p2 : ret_V_27_reg_1056;
assign _027_ = ap_CS_fsm[20] ? ret_V_26_fu_565_p3 : ret_V_26_reg_1000;
assign _026_ = ap_CS_fsm[17] ? grp_fu_499_p2 : ret_V_25_reg_965;
assign _047_ = ap_CS_fsm[4] ? ret_V_20_fu_256_p3[3:0] : trunc_ln1348_reg_759;
assign _022_ = ap_CS_fsm[4] ? ret_V_20_fu_256_p3 : ret_V_20_reg_753;
assign _036_ = ap_CS_fsm[1] ? grp_fu_189_p2[11:2] : ret_V_reg_741;
assign _021_ = ap_CS_fsm[1] ? grp_fu_189_p2 : ret_V_19_reg_736;
assign _020_ = ap_CS_fsm[18] ? grp_fu_503_p2 : ret_V_12_reg_973;
assign _019_ = ap_CS_fsm[16] ? select_ln1368_fu_484_p3[3:1] : ret_V_11_reg_958;
assign _039_ = ap_CS_fsm[16] ? select_ln1368_fu_484_p3 : select_ln1368_reg_952;
assign _017_ = ap_CS_fsm[19] ? ret_V_24_fu_529_p3[2] : p_Result_8_reg_985;
assign _025_ = ap_CS_fsm[19] ? ret_V_24_fu_529_p3 : ret_V_24_reg_978;
assign _015_ = ap_CS_fsm[29] ? grp_fu_613_p2 : op_27_V_reg_1046;
assign _018_ = ap_CS_fsm[29] ? r_fu_621_p3 : r_reg_1041;
assign _038_ = ap_CS_fsm[15] ? select_ln1192_fu_476_p3 : select_ln1192_reg_947;
assign _014_ = ap_CS_fsm[15] ? grp_fu_471_p2 : op_24_V_reg_942;
assign _012_ = ap_CS_fsm[5] ? op_7_V_fu_267_p2[3] : isNeg_reg_769;
assign _016_ = ap_CS_fsm[5] ? op_7_V_fu_267_p2 : op_7_V_reg_764;
assign _010_ = ap_CS_fsm[32] ? icmp_ln851_3_fu_660_p2 : icmp_ln851_3_reg_1071;
assign _009_ = ap_CS_fsm[9] ? icmp_ln851_2_fu_372_p2 : icmp_ln851_2_reg_845;
assign _041_ = ap_CS_fsm[9] ? { ret_V_8_reg_813[9], ret_V_8_reg_813 } : sext_ln831_reg_838;
assign _013_ = ap_CS_fsm[9] ? lhs_V_2_fu_363_p2 : lhs_V_2_reg_833;
assign _023_ = ap_CS_fsm[9] ? ret_V_21_fu_356_p3 : ret_V_21_reg_828;
assign _008_ = ap_CS_fsm[7] ? icmp_ln851_1_fu_302_p2 : icmp_ln851_1_reg_798;
assign _046_ = ap_CS_fsm[0] ? op_2[3:0] : trunc_ln1348_1_reg_731;
assign _007_ = ap_CS_fsm[0] ? icmp_ln1499_fu_219_p2 : icmp_ln1499_reg_726;
assign _011_ = ap_CS_fsm[0] ? icmp_ln851_fu_199_p2 : icmp_ln851_reg_711;
assign _006_ = _056_ ? grp_fu_396_p2 : ashr_ln1333_reg_937;
assign _003_ = ap_CS_fsm[13] ? grp_fu_462_p2 : add_ln69_2_reg_922;
assign _004_ = ap_CS_fsm[13] ? grp_fu_454_p2 : add_ln69_reg_917;
assign _002_ = ap_CS_fsm[11] ? grp_fu_422_p2 : add_ln69_1_reg_897;
assign _037_ = ap_CS_fsm[11] ? grp_fu_409_p2 : ret_reg_892;
assign _024_ = ap_CS_fsm[11] ? ret_V_23_fu_440_p3 : ret_V_23_reg_887;
assign _001_ = _055_ ? grp_fu_508_p2 : add_ln691_reg_990;
assign _000_ = _054_ ? grp_fu_676_p2 : add_ln691_1_reg_1088;
assign _005_ = ap_rst ? 37'h0000000001 : ap_NS_fsm;
assign icmp_ln1499_fu_219_p2 = _326_ ? 1'h1 : 1'h0;
assign icmp_ln851_1_fu_302_p2 = _069_ ? 1'h1 : 1'h0;
assign icmp_ln851_2_fu_372_p2 = _070_ ? 1'h1 : 1'h0;
assign icmp_ln851_3_fu_660_p2 = _327_ ? 1'h1 : 1'h0;
assign icmp_ln851_fu_199_p2 = _071_ ? 1'h1 : 1'h0;
assign lhs_V_2_fu_363_p2 = _072_ ? 1'h1 : 1'h0;
assign op_30 = ret_V_28_reg_1076[34] ? select_ln850_5_fu_688_p3 : ret_V_30_cast_reg_1081;
assign r_fu_621_p3 = p_Result_8_reg_985 ? { trunc_ln546_reg_1026[2], trunc_ln546_reg_1026[2], trunc_ln546_reg_1026[2], trunc_ln546_reg_1026 } : trunc_ln769_reg_1031;
assign ret_V_20_fu_256_p3 = ret_V_19_reg_736[11] ? select_ln850_fu_251_p3 : ret_V_reg_741;
assign ret_V_21_fu_356_p3 = shl_ln1299_reg_775[3] ? select_ln850_1_fu_351_p3 : ret_V_3_reg_780;
assign ret_V_23_fu_440_p3 = ret_V_20_reg_753[9] ? select_ln850_2_fu_435_p3 : sext_ln831_reg_838;
assign ret_V_24_fu_529_p3 = select_ln1368_reg_952[3] ? select_ln850_3_fu_523_p3 : ret_V_11_reg_958;
assign ret_V_26_fu_565_p3 = ret_V_25_reg_965[10] ? select_ln850_4_fu_560_p3 : { 1'h0, ret_V_25_reg_965[9:0] };
assign select_ln1192_fu_476_p3 = op_14 ? 11'h7ff : 11'h000;
assign select_ln1368_fu_484_p3 = isNeg_reg_769 ? shl_ln1299_1_reg_932 : ashr_ln1333_reg_937;
assign select_ln850_1_fu_351_p3 = icmp_ln851_1_reg_798 ? ret_V_3_reg_780 : ret_V_5_reg_808;
assign select_ln850_2_fu_435_p3 = icmp_ln851_2_reg_845 ? sext_ln831_reg_838 : ret_V_9_reg_862;
assign select_ln850_3_fu_523_p3 = select_ln1368_reg_952[0] ? ret_V_12_reg_973 : ret_V_11_reg_958;
assign select_ln850_4_fu_560_p3 = lhs_V_2_reg_833 ? add_ln691_reg_990 : { 1'h1, ret_V_25_reg_965[9:0] };
assign select_ln850_5_fu_688_p3 = icmp_ln851_3_reg_1071 ? add_ln691_1_reg_1088 : ret_V_30_cast_reg_1081;
assign select_ln850_fu_251_p3 = icmp_ln851_reg_711 ? ret_V_reg_741 : ret_V_2_reg_748;
assign ush_fu_339_p3 = isNeg_reg_769 ? sub_ln1367_reg_803 : sext_ln1386_reg_792;
assign ap_CS_fsm_state1 = ap_CS_fsm[0];
assign ap_CS_fsm_state10 = ap_CS_fsm[9];
assign ap_CS_fsm_state11 = ap_CS_fsm[10];
assign ap_CS_fsm_state12 = ap_CS_fsm[11];
assign ap_CS_fsm_state13 = ap_CS_fsm[12];
assign ap_CS_fsm_state14 = ap_CS_fsm[13];
assign ap_CS_fsm_state15 = ap_CS_fsm[14];
assign ap_CS_fsm_state16 = ap_CS_fsm[15];
assign ap_CS_fsm_state17 = ap_CS_fsm[16];
assign ap_CS_fsm_state18 = ap_CS_fsm[17];
assign ap_CS_fsm_state19 = ap_CS_fsm[18];
assign ap_CS_fsm_state2 = ap_CS_fsm[1];
assign ap_CS_fsm_state20 = ap_CS_fsm[19];
assign ap_CS_fsm_state21 = ap_CS_fsm[20];
assign ap_CS_fsm_state22 = ap_CS_fsm[21];
assign ap_CS_fsm_state23 = ap_CS_fsm[22];
assign ap_CS_fsm_state29 = ap_CS_fsm[28];
assign ap_CS_fsm_state3 = ap_CS_fsm[2];
assign ap_CS_fsm_state30 = ap_CS_fsm[29];
assign ap_CS_fsm_state31 = ap_CS_fsm[30];
assign ap_CS_fsm_state32 = ap_CS_fsm[31];
assign ap_CS_fsm_state33 = ap_CS_fsm[32];
assign ap_CS_fsm_state34 = ap_CS_fsm[33];
assign ap_CS_fsm_state35 = ap_CS_fsm[34];
assign ap_CS_fsm_state36 = ap_CS_fsm[35];
assign ap_CS_fsm_state37 = ap_CS_fsm[36];
assign ap_CS_fsm_state4 = ap_CS_fsm[3];
assign ap_CS_fsm_state5 = ap_CS_fsm[4];
assign ap_CS_fsm_state6 = ap_CS_fsm[5];
assign ap_CS_fsm_state7 = ap_CS_fsm[6];
assign ap_CS_fsm_state8 = ap_CS_fsm[7];
assign ap_CS_fsm_state9 = ap_CS_fsm[8];
assign ap_done = op_30_ap_vld;
assign ap_ready = op_30_ap_vld;
assign conv_i_i_i329_fu_386_p0 = op_5;
assign conv_i_i_i329_fu_386_p1 = { op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5 };
assign grp_fu_189_p0 = { 2'h0, op_2, 2'h0 };
assign grp_fu_189_p1 = { op_1[3], op_1[3], op_1[3], op_1[3], op_1[3], op_1[3], op_1[3], op_1[3], op_1 };
assign grp_fu_213_p0 = { op_1[3], op_1[3], op_1[3], op_1[3], op_1[3], op_1[3], op_1[3], op_1[3], op_1[3], op_1[3], op_1[3], op_1[3], op_1[3], op_1[3], op_1[3], op_1[3], op_1[3], op_1[3], op_1[3], op_1[3], op_1[3], op_1[3], op_1[3], op_1[3], op_1[3], op_1[3], op_1[3], op_1[3], op_1 };
assign grp_fu_213_p1 = { 24'h000000, op_2 };
assign grp_fu_296_p1 = { op_7_V_reg_764[3], op_7_V_reg_764 };
assign grp_fu_377_p0 = { ret_V_8_reg_813[9], ret_V_8_reg_813 };
assign grp_fu_409_p0 = { ret_V_21_reg_828[1], ret_V_21_reg_828 };
assign grp_fu_409_p1 = { op_0[1], op_0 };
assign grp_fu_422_p0 = { op_12[1], op_12 };
assign grp_fu_422_p1 = { 2'h0, icmp_ln1499_reg_726 };
assign grp_fu_454_p1 = { ret_reg_892[2], ret_reg_892[2], ret_reg_892[2], ret_reg_892[2], ret_reg_892[2], ret_reg_892[2], ret_reg_892[2], ret_reg_892[2], ret_reg_892 };
assign grp_fu_462_p0 = { add_ln69_1_reg_897[2], add_ln69_1_reg_897[2], add_ln69_1_reg_897[2], add_ln69_1_reg_897 };
assign grp_fu_462_p1 = { 2'h0, op_8 };
assign grp_fu_471_p0 = { add_ln69_2_reg_922[5], add_ln69_2_reg_922[5], add_ln69_2_reg_922[5], add_ln69_2_reg_922[5], add_ln69_2_reg_922[5], add_ln69_2_reg_922 };
assign grp_fu_547_p1 = { ret_V_24_reg_978[2], ret_V_24_reg_978 };
assign grp_fu_582_p1 = { 16'h0000, sh_V_1_reg_1005[3], sh_V_1_reg_1005[3], sh_V_1_reg_1005[3], sh_V_1_reg_1005[3], sh_V_1_reg_1005[3], sh_V_1_reg_1005[3], sh_V_1_reg_1005[3], sh_V_1_reg_1005[3], sh_V_1_reg_1005[3], sh_V_1_reg_1005[3], sh_V_1_reg_1005[3], sh_V_1_reg_1005[3], sh_V_1_reg_1005 };
assign grp_fu_595_p1 = { 16'h0000, ret_V_24_reg_978[2], ret_V_24_reg_978[2], ret_V_24_reg_978[2], ret_V_24_reg_978[2], ret_V_24_reg_978[2], ret_V_24_reg_978[2], ret_V_24_reg_978[2], ret_V_24_reg_978[2], ret_V_24_reg_978[2], ret_V_24_reg_978[2], ret_V_24_reg_978[2], ret_V_24_reg_978[2], ret_V_24_reg_978[2], ret_V_24_reg_978 };
assign grp_fu_613_p1 = { op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16 };
assign grp_fu_630_p1 = { r_reg_1041[5], r_reg_1041[5], r_reg_1041[5], r_reg_1041[5], r_reg_1041[5], r_reg_1041 };
assign grp_fu_650_p0 = { ret_V_27_reg_1056[10], ret_V_27_reg_1056[10], ret_V_27_reg_1056[10], ret_V_27_reg_1056[10], ret_V_27_reg_1056[10], ret_V_27_reg_1056[10], ret_V_27_reg_1056[10], ret_V_27_reg_1056[10], ret_V_27_reg_1056[10], ret_V_27_reg_1056[10], ret_V_27_reg_1056[10], ret_V_27_reg_1056[10], ret_V_27_reg_1056[10], ret_V_27_reg_1056[10], ret_V_27_reg_1056[10], ret_V_27_reg_1056[10], ret_V_27_reg_1056[10], ret_V_27_reg_1056[10], ret_V_27_reg_1056[10], ret_V_27_reg_1056[10], ret_V_27_reg_1056[10], ret_V_27_reg_1056[10], ret_V_27_reg_1056, 2'h0 };
assign grp_fu_650_p1 = { op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18 };
assign lhs_V_1_fu_312_p3 = { ret_V_20_reg_753, 2'h0 };
assign lhs_V_2_fu_363_p0 = op_5;
assign p_Result_1_fu_344_p3 = shl_ln1299_reg_775[3];
assign p_Result_3_fu_428_p3 = ret_V_20_reg_753[9];
assign p_Result_4_fu_513_p3 = select_ln1368_reg_952[3];
assign p_Result_6_fu_553_p3 = ret_V_25_reg_965[10];
assign p_Result_7_fu_681_p3 = ret_V_28_reg_1076[34];
assign p_Result_s_fu_244_p3 = ret_V_19_reg_736[11];
assign ret_V_22_fu_319_p2[1:0] = 2'h0;
assign ret_V_22_fu_319_p2[11:3] = ret_V_20_reg_753[9:1];
assign rhs_fu_177_p3 = { op_2, 2'h0 };
assign sext_ln1299_fu_209_p0 = op_1;
assign sext_ln1367_fu_383_p1 = { ush_reg_823[4], ush_reg_823[4], ush_reg_823[4], ush_reg_823[4], ush_reg_823[4], ush_reg_823[4], ush_reg_823[4], ush_reg_823[4], ush_reg_823[4], ush_reg_823[4], ush_reg_823[4], ush_reg_823[4], ush_reg_823[4], ush_reg_823[4], ush_reg_823[4], ush_reg_823[4], ush_reg_823[4], ush_reg_823[4], ush_reg_823[4], ush_reg_823[4], ush_reg_823[4], ush_reg_823[4], ush_reg_823[4], ush_reg_823[4], ush_reg_823[4], ush_reg_823[4], ush_reg_823[4], ush_reg_823 };
assign sext_ln1386_fu_293_p1 = { op_7_V_reg_764[3], op_7_V_reg_764 };
assign sext_ln546_1_fu_618_p1 = { trunc_ln546_reg_1026[2], trunc_ln546_reg_1026[2], trunc_ln546_reg_1026[2], trunc_ln546_reg_1026 };
assign sext_ln546_2_fu_588_p1 = { ret_V_24_reg_978[2], ret_V_24_reg_978[2], ret_V_24_reg_978[2], ret_V_24_reg_978[2], ret_V_24_reg_978[2], ret_V_24_reg_978[2], ret_V_24_reg_978[2], ret_V_24_reg_978[2], ret_V_24_reg_978[2], ret_V_24_reg_978[2], ret_V_24_reg_978[2], ret_V_24_reg_978[2], ret_V_24_reg_978[2], ret_V_24_reg_978 };
assign sext_ln546_fu_575_p1 = { sh_V_1_reg_1005[3], sh_V_1_reg_1005[3], sh_V_1_reg_1005[3], sh_V_1_reg_1005[3], sh_V_1_reg_1005[3], sh_V_1_reg_1005[3], sh_V_1_reg_1005[3], sh_V_1_reg_1005[3], sh_V_1_reg_1005[3], sh_V_1_reg_1005[3], sh_V_1_reg_1005[3], sh_V_1_reg_1005[3], sh_V_1_reg_1005 };
assign sext_ln703_1_fu_635_p0 = op_18;
assign sext_ln703_fu_173_p0 = op_1;
assign sext_ln781_fu_572_p1 = { ret_V_24_reg_978[2], ret_V_24_reg_978[2], ret_V_24_reg_978[2], ret_V_24_reg_978[2], ret_V_24_reg_978[2], ret_V_24_reg_978[2], ret_V_24_reg_978[2], ret_V_24_reg_978[2], ret_V_24_reg_978[2], ret_V_24_reg_978[2], ret_V_24_reg_978[2], ret_V_24_reg_978[2], ret_V_24_reg_978[2], ret_V_24_reg_978[2], ret_V_24_reg_978[2], ret_V_24_reg_978[2], ret_V_24_reg_978[2], ret_V_24_reg_978[2], ret_V_24_reg_978[2], ret_V_24_reg_978[2], ret_V_24_reg_978[2], ret_V_24_reg_978[2], ret_V_24_reg_978[2], ret_V_24_reg_978[2], ret_V_24_reg_978[2], ret_V_24_reg_978[2], ret_V_24_reg_978[2], ret_V_24_reg_978[2], ret_V_24_reg_978[2], ret_V_24_reg_978 };
assign sext_ln831_fu_369_p1 = { ret_V_8_reg_813[9], ret_V_8_reg_813 };
assign tmp_fu_639_p3 = { ret_V_27_reg_1056, 2'h0 };
assign trunc_ln1348_1_fu_225_p1 = op_2[3:0];
assign trunc_ln1348_fu_263_p1 = ret_V_20_fu_256_p3[3:0];
assign trunc_ln546_fu_601_p1 = grp_fu_582_p2[2:0];
assign trunc_ln769_fu_605_p1 = grp_fu_595_p2[5:0];
assign trunc_ln851_1_fu_289_p1 = grp_fu_213_p2[1:0];
assign trunc_ln851_2_fu_335_p1 = 2'h0;
assign trunc_ln851_3_fu_520_p1 = select_ln1368_reg_952[0];
assign trunc_ln851_4_fu_656_p0 = op_18;
assign trunc_ln851_4_fu_656_p1 = op_18[1:0];
assign trunc_ln851_fu_195_p0 = op_1;
assign trunc_ln851_fu_195_p1 = op_1[1:0];
assign \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.ain_s0  = \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.a ;
assign \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.s  = { \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.fas_s2 , \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.sum_s1  };
assign \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.u2.a  = \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.ain_s1 ;
assign \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.u2.b  = \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.bin_s1 ;
assign \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.u2.cin  = \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.carry_s1 ;
assign \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.facout_s2  = \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.u2.cout ;
assign \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.fas_s2  = \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.u2.s ;
assign \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.u1.a  = \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.a [1:0];
assign \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.u1.b  = \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.bin_s0 [1:0];
assign \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.u1.cin  = 1'h1;
assign \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.facout_s1  = \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.u1.cout ;
assign \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.fas_s1  = \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.u1.s ;
assign \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.a  = \sub_5ns_5s_5_2_1_U4.din0 ;
assign \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.b  = \sub_5ns_5s_5_2_1_U4.din1 ;
assign \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.ce  = \sub_5ns_5s_5_2_1_U4.ce ;
assign \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.clk  = \sub_5ns_5s_5_2_1_U4.clk ;
assign \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.reset  = \sub_5ns_5s_5_2_1_U4.reset ;
assign \sub_5ns_5s_5_2_1_U4.dout  = \sub_5ns_5s_5_2_1_U4.top_sub_5ns_5s_5_2_1_Adder_2_U.s ;
assign \sub_5ns_5s_5_2_1_U4.ce  = 1'h1;
assign \sub_5ns_5s_5_2_1_U4.clk  = ap_clk;
assign \sub_5ns_5s_5_2_1_U4.din0  = 5'h00;
assign \sub_5ns_5s_5_2_1_U4.din1  = { op_7_V_reg_764[3], op_7_V_reg_764 };
assign grp_fu_296_p2 = \sub_5ns_5s_5_2_1_U4.dout ;
assign \sub_5ns_5s_5_2_1_U4.reset  = ap_rst;
assign \sub_4ns_4s_4_2_1_U17.top_sub_4ns_4s_4_2_1_Adder_11_U.ain_s0  = \sub_4ns_4s_4_2_1_U17.top_sub_4ns_4s_4_2_1_Adder_11_U.a ;
assign \sub_4ns_4s_4_2_1_U17.top_sub_4ns_4s_4_2_1_Adder_11_U.s  = { \sub_4ns_4s_4_2_1_U17.top_sub_4ns_4s_4_2_1_Adder_11_U.fas_s2 , \sub_4ns_4s_4_2_1_U17.top_sub_4ns_4s_4_2_1_Adder_11_U.sum_s1  };
assign \sub_4ns_4s_4_2_1_U17.top_sub_4ns_4s_4_2_1_Adder_11_U.u2.a  = \sub_4ns_4s_4_2_1_U17.top_sub_4ns_4s_4_2_1_Adder_11_U.ain_s1 ;
assign \sub_4ns_4s_4_2_1_U17.top_sub_4ns_4s_4_2_1_Adder_11_U.u2.b  = \sub_4ns_4s_4_2_1_U17.top_sub_4ns_4s_4_2_1_Adder_11_U.bin_s1 ;
assign \sub_4ns_4s_4_2_1_U17.top_sub_4ns_4s_4_2_1_Adder_11_U.u2.cin  = \sub_4ns_4s_4_2_1_U17.top_sub_4ns_4s_4_2_1_Adder_11_U.carry_s1 ;
assign \sub_4ns_4s_4_2_1_U17.top_sub_4ns_4s_4_2_1_Adder_11_U.facout_s2  = \sub_4ns_4s_4_2_1_U17.top_sub_4ns_4s_4_2_1_Adder_11_U.u2.cout ;
assign \sub_4ns_4s_4_2_1_U17.top_sub_4ns_4s_4_2_1_Adder_11_U.fas_s2  = \sub_4ns_4s_4_2_1_U17.top_sub_4ns_4s_4_2_1_Adder_11_U.u2.s ;
assign \sub_4ns_4s_4_2_1_U17.top_sub_4ns_4s_4_2_1_Adder_11_U.u1.a  = \sub_4ns_4s_4_2_1_U17.top_sub_4ns_4s_4_2_1_Adder_11_U.a [1:0];
assign \sub_4ns_4s_4_2_1_U17.top_sub_4ns_4s_4_2_1_Adder_11_U.u1.b  = \sub_4ns_4s_4_2_1_U17.top_sub_4ns_4s_4_2_1_Adder_11_U.bin_s0 [1:0];
assign \sub_4ns_4s_4_2_1_U17.top_sub_4ns_4s_4_2_1_Adder_11_U.u1.cin  = 1'h1;
assign \sub_4ns_4s_4_2_1_U17.top_sub_4ns_4s_4_2_1_Adder_11_U.facout_s1  = \sub_4ns_4s_4_2_1_U17.top_sub_4ns_4s_4_2_1_Adder_11_U.u1.cout ;
assign \sub_4ns_4s_4_2_1_U17.top_sub_4ns_4s_4_2_1_Adder_11_U.fas_s1  = \sub_4ns_4s_4_2_1_U17.top_sub_4ns_4s_4_2_1_Adder_11_U.u1.s ;
assign \sub_4ns_4s_4_2_1_U17.top_sub_4ns_4s_4_2_1_Adder_11_U.a  = \sub_4ns_4s_4_2_1_U17.din0 ;
assign \sub_4ns_4s_4_2_1_U17.top_sub_4ns_4s_4_2_1_Adder_11_U.b  = \sub_4ns_4s_4_2_1_U17.din1 ;
assign \sub_4ns_4s_4_2_1_U17.top_sub_4ns_4s_4_2_1_Adder_11_U.ce  = \sub_4ns_4s_4_2_1_U17.ce ;
assign \sub_4ns_4s_4_2_1_U17.top_sub_4ns_4s_4_2_1_Adder_11_U.clk  = \sub_4ns_4s_4_2_1_U17.clk ;
assign \sub_4ns_4s_4_2_1_U17.top_sub_4ns_4s_4_2_1_Adder_11_U.reset  = \sub_4ns_4s_4_2_1_U17.reset ;
assign \sub_4ns_4s_4_2_1_U17.dout  = \sub_4ns_4s_4_2_1_U17.top_sub_4ns_4s_4_2_1_Adder_11_U.s ;
assign \sub_4ns_4s_4_2_1_U17.ce  = 1'h1;
assign \sub_4ns_4s_4_2_1_U17.clk  = ap_clk;
assign \sub_4ns_4s_4_2_1_U17.din0  = 4'h0;
assign \sub_4ns_4s_4_2_1_U17.din1  = { ret_V_24_reg_978[2], ret_V_24_reg_978 };
assign grp_fu_547_p2 = \sub_4ns_4s_4_2_1_U17.dout ;
assign \sub_4ns_4s_4_2_1_U17.reset  = ap_rst;
assign \shl_32s_8ns_32_7_1_U2.din1_cast  = \shl_32s_8ns_32_7_1_U2.din1 [7:0];
assign \shl_32s_8ns_32_7_1_U2.din1_mask  = 8'h03;
assign \shl_32s_8ns_32_7_1_U2.ce  = 1'h1;
assign \shl_32s_8ns_32_7_1_U2.clk  = ap_clk;
assign \shl_32s_8ns_32_7_1_U2.din0  = { op_1[3], op_1[3], op_1[3], op_1[3], op_1[3], op_1[3], op_1[3], op_1[3], op_1[3], op_1[3], op_1[3], op_1[3], op_1[3], op_1[3], op_1[3], op_1[3], op_1[3], op_1[3], op_1[3], op_1[3], op_1[3], op_1[3], op_1[3], op_1[3], op_1[3], op_1[3], op_1[3], op_1[3], op_1 };
assign \shl_32s_8ns_32_7_1_U2.din1  = { 24'h000000, op_2 };
assign grp_fu_213_p2 = \shl_32s_8ns_32_7_1_U2.dout ;
assign \shl_32s_8ns_32_7_1_U2.reset  = ap_rst;
assign \shl_32s_32s_32_7_1_U7.din1_cast  = \shl_32s_32s_32_7_1_U7.din1 ;
assign \shl_32s_32s_32_7_1_U7.din1_mask  = 32'd31;
assign \shl_32s_32s_32_7_1_U7.ce  = 1'h1;
assign \shl_32s_32s_32_7_1_U7.clk  = ap_clk;
assign \shl_32s_32s_32_7_1_U7.din0  = { op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5 };
assign \shl_32s_32s_32_7_1_U7.din1  = { ush_reg_823[4], ush_reg_823[4], ush_reg_823[4], ush_reg_823[4], ush_reg_823[4], ush_reg_823[4], ush_reg_823[4], ush_reg_823[4], ush_reg_823[4], ush_reg_823[4], ush_reg_823[4], ush_reg_823[4], ush_reg_823[4], ush_reg_823[4], ush_reg_823[4], ush_reg_823[4], ush_reg_823[4], ush_reg_823[4], ush_reg_823[4], ush_reg_823[4], ush_reg_823[4], ush_reg_823[4], ush_reg_823[4], ush_reg_823[4], ush_reg_823[4], ush_reg_823[4], ush_reg_823[4], ush_reg_823 };
assign grp_fu_390_p2 = \shl_32s_32s_32_7_1_U7.dout ;
assign \shl_32s_32s_32_7_1_U7.reset  = ap_rst;
assign \shl_32s_16ns_32_7_1_U19.din1_cast  = \shl_32s_16ns_32_7_1_U19.din1 [15:0];
assign \shl_32s_16ns_32_7_1_U19.din1_mask  = 16'h0007;
assign \shl_32s_16ns_32_7_1_U19.ce  = 1'h1;
assign \shl_32s_16ns_32_7_1_U19.clk  = ap_clk;
assign \shl_32s_16ns_32_7_1_U19.din0  = { ret_V_24_reg_978[2], ret_V_24_reg_978[2], ret_V_24_reg_978[2], ret_V_24_reg_978[2], ret_V_24_reg_978[2], ret_V_24_reg_978[2], ret_V_24_reg_978[2], ret_V_24_reg_978[2], ret_V_24_reg_978[2], ret_V_24_reg_978[2], ret_V_24_reg_978[2], ret_V_24_reg_978[2], ret_V_24_reg_978[2], ret_V_24_reg_978[2], ret_V_24_reg_978[2], ret_V_24_reg_978[2], ret_V_24_reg_978[2], ret_V_24_reg_978[2], ret_V_24_reg_978[2], ret_V_24_reg_978[2], ret_V_24_reg_978[2], ret_V_24_reg_978[2], ret_V_24_reg_978[2], ret_V_24_reg_978[2], ret_V_24_reg_978[2], ret_V_24_reg_978[2], ret_V_24_reg_978[2], ret_V_24_reg_978[2], ret_V_24_reg_978[2], ret_V_24_reg_978 };
assign \shl_32s_16ns_32_7_1_U19.din1  = { 16'h0000, ret_V_24_reg_978[2], ret_V_24_reg_978[2], ret_V_24_reg_978[2], ret_V_24_reg_978[2], ret_V_24_reg_978[2], ret_V_24_reg_978[2], ret_V_24_reg_978[2], ret_V_24_reg_978[2], ret_V_24_reg_978[2], ret_V_24_reg_978[2], ret_V_24_reg_978[2], ret_V_24_reg_978[2], ret_V_24_reg_978[2], ret_V_24_reg_978 };
assign grp_fu_595_p2 = \shl_32s_16ns_32_7_1_U19.dout ;
assign \shl_32s_16ns_32_7_1_U19.reset  = ap_rst;
assign \ashr_32s_32s_32_7_1_U8.din1_cast  = \ashr_32s_32s_32_7_1_U8.din1 ;
assign \ashr_32s_32s_32_7_1_U8.din1_mask  = 32'd31;
assign \ashr_32s_32s_32_7_1_U8.ce  = 1'h1;
assign \ashr_32s_32s_32_7_1_U8.clk  = ap_clk;
assign \ashr_32s_32s_32_7_1_U8.din0  = { op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5[3], op_5 };
assign \ashr_32s_32s_32_7_1_U8.din1  = { ush_reg_823[4], ush_reg_823[4], ush_reg_823[4], ush_reg_823[4], ush_reg_823[4], ush_reg_823[4], ush_reg_823[4], ush_reg_823[4], ush_reg_823[4], ush_reg_823[4], ush_reg_823[4], ush_reg_823[4], ush_reg_823[4], ush_reg_823[4], ush_reg_823[4], ush_reg_823[4], ush_reg_823[4], ush_reg_823[4], ush_reg_823[4], ush_reg_823[4], ush_reg_823[4], ush_reg_823[4], ush_reg_823[4], ush_reg_823[4], ush_reg_823[4], ush_reg_823[4], ush_reg_823[4], ush_reg_823 };
assign grp_fu_396_p2 = \ashr_32s_32s_32_7_1_U8.dout ;
assign \ashr_32s_32s_32_7_1_U8.reset  = ap_rst;
assign \ashr_32s_16ns_32_7_1_U18.din1_cast  = \ashr_32s_16ns_32_7_1_U18.din1 [15:0];
assign \ashr_32s_16ns_32_7_1_U18.din1_mask  = 16'h0007;
assign \ashr_32s_16ns_32_7_1_U18.ce  = 1'h1;
assign \ashr_32s_16ns_32_7_1_U18.clk  = ap_clk;
assign \ashr_32s_16ns_32_7_1_U18.din0  = { ret_V_24_reg_978[2], ret_V_24_reg_978[2], ret_V_24_reg_978[2], ret_V_24_reg_978[2], ret_V_24_reg_978[2], ret_V_24_reg_978[2], ret_V_24_reg_978[2], ret_V_24_reg_978[2], ret_V_24_reg_978[2], ret_V_24_reg_978[2], ret_V_24_reg_978[2], ret_V_24_reg_978[2], ret_V_24_reg_978[2], ret_V_24_reg_978[2], ret_V_24_reg_978[2], ret_V_24_reg_978[2], ret_V_24_reg_978[2], ret_V_24_reg_978[2], ret_V_24_reg_978[2], ret_V_24_reg_978[2], ret_V_24_reg_978[2], ret_V_24_reg_978[2], ret_V_24_reg_978[2], ret_V_24_reg_978[2], ret_V_24_reg_978[2], ret_V_24_reg_978[2], ret_V_24_reg_978[2], ret_V_24_reg_978[2], ret_V_24_reg_978[2], ret_V_24_reg_978 };
assign \ashr_32s_16ns_32_7_1_U18.din1  = { 16'h0000, sh_V_1_reg_1005[3], sh_V_1_reg_1005[3], sh_V_1_reg_1005[3], sh_V_1_reg_1005[3], sh_V_1_reg_1005[3], sh_V_1_reg_1005[3], sh_V_1_reg_1005[3], sh_V_1_reg_1005[3], sh_V_1_reg_1005[3], sh_V_1_reg_1005[3], sh_V_1_reg_1005[3], sh_V_1_reg_1005[3], sh_V_1_reg_1005 };
assign grp_fu_582_p2 = \ashr_32s_16ns_32_7_1_U18.dout ;
assign \ashr_32s_16ns_32_7_1_U18.reset  = ap_rst;
assign \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_8_U.ain_s0  = \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_8_U.a ;
assign \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_8_U.bin_s0  = \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_8_U.b ;
assign \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_8_U.s  = { \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_8_U.fas_s2 , \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_8_U.sum_s1  };
assign \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_8_U.u2.a  = \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_8_U.ain_s1 ;
assign \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_8_U.u2.b  = \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_8_U.bin_s1 ;
assign \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_8_U.u2.cin  = \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_8_U.carry_s1 ;
assign \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_8_U.facout_s2  = \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_8_U.u2.cout ;
assign \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_8_U.fas_s2  = \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_8_U.u2.s ;
assign \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_8_U.u1.a  = \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_8_U.a [2:0];
assign \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_8_U.u1.b  = \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_8_U.b [2:0];
assign \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_8_U.u1.cin  = 1'h0;
assign \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_8_U.facout_s1  = \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_8_U.u1.cout ;
assign \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_8_U.fas_s1  = \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_8_U.u1.s ;
assign \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_8_U.a  = \add_6s_6ns_6_2_1_U12.din0 ;
assign \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_8_U.b  = \add_6s_6ns_6_2_1_U12.din1 ;
assign \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_8_U.ce  = \add_6s_6ns_6_2_1_U12.ce ;
assign \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_8_U.clk  = \add_6s_6ns_6_2_1_U12.clk ;
assign \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_8_U.reset  = \add_6s_6ns_6_2_1_U12.reset ;
assign \add_6s_6ns_6_2_1_U12.dout  = \add_6s_6ns_6_2_1_U12.top_add_6s_6ns_6_2_1_Adder_8_U.s ;
assign \add_6s_6ns_6_2_1_U12.ce  = 1'h1;
assign \add_6s_6ns_6_2_1_U12.clk  = ap_clk;
assign \add_6s_6ns_6_2_1_U12.din0  = { add_ln69_1_reg_897[2], add_ln69_1_reg_897[2], add_ln69_1_reg_897[2], add_ln69_1_reg_897 };
assign \add_6s_6ns_6_2_1_U12.din1  = { 2'h0, op_8 };
assign grp_fu_462_p2 = \add_6s_6ns_6_2_1_U12.dout ;
assign \add_6s_6ns_6_2_1_U12.reset  = ap_rst;
assign \add_3s_3s_3_2_1_U9.top_add_3s_3s_3_2_1_Adder_5_U.ain_s0  = \add_3s_3s_3_2_1_U9.top_add_3s_3s_3_2_1_Adder_5_U.a ;
assign \add_3s_3s_3_2_1_U9.top_add_3s_3s_3_2_1_Adder_5_U.bin_s0  = \add_3s_3s_3_2_1_U9.top_add_3s_3s_3_2_1_Adder_5_U.b ;
assign \add_3s_3s_3_2_1_U9.top_add_3s_3s_3_2_1_Adder_5_U.s  = { \add_3s_3s_3_2_1_U9.top_add_3s_3s_3_2_1_Adder_5_U.fas_s2 , \add_3s_3s_3_2_1_U9.top_add_3s_3s_3_2_1_Adder_5_U.sum_s1  };
assign \add_3s_3s_3_2_1_U9.top_add_3s_3s_3_2_1_Adder_5_U.u2.a  = \add_3s_3s_3_2_1_U9.top_add_3s_3s_3_2_1_Adder_5_U.ain_s1 ;
assign \add_3s_3s_3_2_1_U9.top_add_3s_3s_3_2_1_Adder_5_U.u2.b  = \add_3s_3s_3_2_1_U9.top_add_3s_3s_3_2_1_Adder_5_U.bin_s1 ;
assign \add_3s_3s_3_2_1_U9.top_add_3s_3s_3_2_1_Adder_5_U.u2.cin  = \add_3s_3s_3_2_1_U9.top_add_3s_3s_3_2_1_Adder_5_U.carry_s1 ;
assign \add_3s_3s_3_2_1_U9.top_add_3s_3s_3_2_1_Adder_5_U.facout_s2  = \add_3s_3s_3_2_1_U9.top_add_3s_3s_3_2_1_Adder_5_U.u2.cout ;
assign \add_3s_3s_3_2_1_U9.top_add_3s_3s_3_2_1_Adder_5_U.fas_s2  = \add_3s_3s_3_2_1_U9.top_add_3s_3s_3_2_1_Adder_5_U.u2.s ;
assign \add_3s_3s_3_2_1_U9.top_add_3s_3s_3_2_1_Adder_5_U.u1.a  = \add_3s_3s_3_2_1_U9.top_add_3s_3s_3_2_1_Adder_5_U.a [0];
assign \add_3s_3s_3_2_1_U9.top_add_3s_3s_3_2_1_Adder_5_U.u1.b  = \add_3s_3s_3_2_1_U9.top_add_3s_3s_3_2_1_Adder_5_U.b [0];
assign \add_3s_3s_3_2_1_U9.top_add_3s_3s_3_2_1_Adder_5_U.u1.cin  = 1'h0;
assign \add_3s_3s_3_2_1_U9.top_add_3s_3s_3_2_1_Adder_5_U.facout_s1  = \add_3s_3s_3_2_1_U9.top_add_3s_3s_3_2_1_Adder_5_U.u1.cout ;
assign \add_3s_3s_3_2_1_U9.top_add_3s_3s_3_2_1_Adder_5_U.fas_s1  = \add_3s_3s_3_2_1_U9.top_add_3s_3s_3_2_1_Adder_5_U.u1.s ;
assign \add_3s_3s_3_2_1_U9.top_add_3s_3s_3_2_1_Adder_5_U.a  = \add_3s_3s_3_2_1_U9.din0 ;
assign \add_3s_3s_3_2_1_U9.top_add_3s_3s_3_2_1_Adder_5_U.b  = \add_3s_3s_3_2_1_U9.din1 ;
assign \add_3s_3s_3_2_1_U9.top_add_3s_3s_3_2_1_Adder_5_U.ce  = \add_3s_3s_3_2_1_U9.ce ;
assign \add_3s_3s_3_2_1_U9.top_add_3s_3s_3_2_1_Adder_5_U.clk  = \add_3s_3s_3_2_1_U9.clk ;
assign \add_3s_3s_3_2_1_U9.top_add_3s_3s_3_2_1_Adder_5_U.reset  = \add_3s_3s_3_2_1_U9.reset ;
assign \add_3s_3s_3_2_1_U9.dout  = \add_3s_3s_3_2_1_U9.top_add_3s_3s_3_2_1_Adder_5_U.s ;
assign \add_3s_3s_3_2_1_U9.ce  = 1'h1;
assign \add_3s_3s_3_2_1_U9.clk  = ap_clk;
assign \add_3s_3s_3_2_1_U9.din0  = { ret_V_21_reg_828[1], ret_V_21_reg_828 };
assign \add_3s_3s_3_2_1_U9.din1  = { op_0[1], op_0 };
assign grp_fu_409_p2 = \add_3s_3s_3_2_1_U9.dout ;
assign \add_3s_3s_3_2_1_U9.reset  = ap_rst;
assign \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.ain_s0  = \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.a ;
assign \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.bin_s0  = \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.b ;
assign \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.s  = { \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.fas_s2 , \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.sum_s1  };
assign \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.u2.a  = \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.ain_s1 ;
assign \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.u2.b  = \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.bin_s1 ;
assign \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.u2.cin  = \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.carry_s1 ;
assign \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.facout_s2  = \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.u2.cout ;
assign \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.fas_s2  = \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.u2.s ;
assign \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.u1.a  = \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.a [0];
assign \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.u1.b  = \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.b [0];
assign \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.u1.cin  = 1'h0;
assign \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.facout_s1  = \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.u1.cout ;
assign \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.fas_s1  = \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.u1.s ;
assign \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.a  = \add_3s_3ns_3_2_1_U10.din0 ;
assign \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.b  = \add_3s_3ns_3_2_1_U10.din1 ;
assign \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.ce  = \add_3s_3ns_3_2_1_U10.ce ;
assign \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.clk  = \add_3s_3ns_3_2_1_U10.clk ;
assign \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.reset  = \add_3s_3ns_3_2_1_U10.reset ;
assign \add_3s_3ns_3_2_1_U10.dout  = \add_3s_3ns_3_2_1_U10.top_add_3s_3ns_3_2_1_Adder_6_U.s ;
assign \add_3s_3ns_3_2_1_U10.ce  = 1'h1;
assign \add_3s_3ns_3_2_1_U10.clk  = ap_clk;
assign \add_3s_3ns_3_2_1_U10.din0  = { op_12[1], op_12 };
assign \add_3s_3ns_3_2_1_U10.din1  = { 2'h0, icmp_ln1499_reg_726 };
assign grp_fu_422_p2 = \add_3s_3ns_3_2_1_U10.dout ;
assign \add_3s_3ns_3_2_1_U10.reset  = ap_rst;
assign \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_10_U.ain_s0  = \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_10_U.a ;
assign \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_10_U.bin_s0  = \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_10_U.b ;
assign \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_10_U.s  = { \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_10_U.fas_s2 , \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_10_U.sum_s1  };
assign \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_10_U.u2.a  = \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_10_U.ain_s1 ;
assign \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_10_U.u2.b  = \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_10_U.bin_s1 ;
assign \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_10_U.u2.cin  = \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_10_U.carry_s1 ;
assign \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_10_U.facout_s2  = \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_10_U.u2.cout ;
assign \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_10_U.fas_s2  = \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_10_U.u2.s ;
assign \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_10_U.u1.a  = \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_10_U.a [0];
assign \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_10_U.u1.b  = \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_10_U.b [0];
assign \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_10_U.u1.cin  = 1'h0;
assign \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_10_U.facout_s1  = \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_10_U.u1.cout ;
assign \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_10_U.fas_s1  = \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_10_U.u1.s ;
assign \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_10_U.a  = \add_3ns_3ns_3_2_1_U15.din0 ;
assign \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_10_U.b  = \add_3ns_3ns_3_2_1_U15.din1 ;
assign \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_10_U.ce  = \add_3ns_3ns_3_2_1_U15.ce ;
assign \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_10_U.clk  = \add_3ns_3ns_3_2_1_U15.clk ;
assign \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_10_U.reset  = \add_3ns_3ns_3_2_1_U15.reset ;
assign \add_3ns_3ns_3_2_1_U15.dout  = \add_3ns_3ns_3_2_1_U15.top_add_3ns_3ns_3_2_1_Adder_10_U.s ;
assign \add_3ns_3ns_3_2_1_U15.ce  = 1'h1;
assign \add_3ns_3ns_3_2_1_U15.clk  = ap_clk;
assign \add_3ns_3ns_3_2_1_U15.din0  = ret_V_11_reg_958;
assign \add_3ns_3ns_3_2_1_U15.din1  = 3'h1;
assign grp_fu_503_p2 = \add_3ns_3ns_3_2_1_U15.dout ;
assign \add_3ns_3ns_3_2_1_U15.reset  = ap_rst;
assign \add_35s_35s_35_2_1_U22.top_add_35s_35s_35_2_1_Adder_12_U.ain_s0  = \add_35s_35s_35_2_1_U22.top_add_35s_35s_35_2_1_Adder_12_U.a ;
assign \add_35s_35s_35_2_1_U22.top_add_35s_35s_35_2_1_Adder_12_U.bin_s0  = \add_35s_35s_35_2_1_U22.top_add_35s_35s_35_2_1_Adder_12_U.b ;
assign \add_35s_35s_35_2_1_U22.top_add_35s_35s_35_2_1_Adder_12_U.s  = { \add_35s_35s_35_2_1_U22.top_add_35s_35s_35_2_1_Adder_12_U.fas_s2 , \add_35s_35s_35_2_1_U22.top_add_35s_35s_35_2_1_Adder_12_U.sum_s1  };
assign \add_35s_35s_35_2_1_U22.top_add_35s_35s_35_2_1_Adder_12_U.u2.a  = \add_35s_35s_35_2_1_U22.top_add_35s_35s_35_2_1_Adder_12_U.ain_s1 ;
assign \add_35s_35s_35_2_1_U22.top_add_35s_35s_35_2_1_Adder_12_U.u2.b  = \add_35s_35s_35_2_1_U22.top_add_35s_35s_35_2_1_Adder_12_U.bin_s1 ;
assign \add_35s_35s_35_2_1_U22.top_add_35s_35s_35_2_1_Adder_12_U.u2.cin  = \add_35s_35s_35_2_1_U22.top_add_35s_35s_35_2_1_Adder_12_U.carry_s1 ;
assign \add_35s_35s_35_2_1_U22.top_add_35s_35s_35_2_1_Adder_12_U.facout_s2  = \add_35s_35s_35_2_1_U22.top_add_35s_35s_35_2_1_Adder_12_U.u2.cout ;
assign \add_35s_35s_35_2_1_U22.top_add_35s_35s_35_2_1_Adder_12_U.fas_s2  = \add_35s_35s_35_2_1_U22.top_add_35s_35s_35_2_1_Adder_12_U.u2.s ;
assign \add_35s_35s_35_2_1_U22.top_add_35s_35s_35_2_1_Adder_12_U.u1.a  = \add_35s_35s_35_2_1_U22.top_add_35s_35s_35_2_1_Adder_12_U.a [16:0];
assign \add_35s_35s_35_2_1_U22.top_add_35s_35s_35_2_1_Adder_12_U.u1.b  = \add_35s_35s_35_2_1_U22.top_add_35s_35s_35_2_1_Adder_12_U.b [16:0];
assign \add_35s_35s_35_2_1_U22.top_add_35s_35s_35_2_1_Adder_12_U.u1.cin  = 1'h0;
assign \add_35s_35s_35_2_1_U22.top_add_35s_35s_35_2_1_Adder_12_U.facout_s1  = \add_35s_35s_35_2_1_U22.top_add_35s_35s_35_2_1_Adder_12_U.u1.cout ;
assign \add_35s_35s_35_2_1_U22.top_add_35s_35s_35_2_1_Adder_12_U.fas_s1  = \add_35s_35s_35_2_1_U22.top_add_35s_35s_35_2_1_Adder_12_U.u1.s ;
assign \add_35s_35s_35_2_1_U22.top_add_35s_35s_35_2_1_Adder_12_U.a  = \add_35s_35s_35_2_1_U22.din0 ;
assign \add_35s_35s_35_2_1_U22.top_add_35s_35s_35_2_1_Adder_12_U.b  = \add_35s_35s_35_2_1_U22.din1 ;
assign \add_35s_35s_35_2_1_U22.top_add_35s_35s_35_2_1_Adder_12_U.ce  = \add_35s_35s_35_2_1_U22.ce ;
assign \add_35s_35s_35_2_1_U22.top_add_35s_35s_35_2_1_Adder_12_U.clk  = \add_35s_35s_35_2_1_U22.clk ;
assign \add_35s_35s_35_2_1_U22.top_add_35s_35s_35_2_1_Adder_12_U.reset  = \add_35s_35s_35_2_1_U22.reset ;
assign \add_35s_35s_35_2_1_U22.dout  = \add_35s_35s_35_2_1_U22.top_add_35s_35s_35_2_1_Adder_12_U.s ;
assign \add_35s_35s_35_2_1_U22.ce  = 1'h1;
assign \add_35s_35s_35_2_1_U22.clk  = ap_clk;
assign \add_35s_35s_35_2_1_U22.din0  = { ret_V_27_reg_1056[10], ret_V_27_reg_1056[10], ret_V_27_reg_1056[10], ret_V_27_reg_1056[10], ret_V_27_reg_1056[10], ret_V_27_reg_1056[10], ret_V_27_reg_1056[10], ret_V_27_reg_1056[10], ret_V_27_reg_1056[10], ret_V_27_reg_1056[10], ret_V_27_reg_1056[10], ret_V_27_reg_1056[10], ret_V_27_reg_1056[10], ret_V_27_reg_1056[10], ret_V_27_reg_1056[10], ret_V_27_reg_1056[10], ret_V_27_reg_1056[10], ret_V_27_reg_1056[10], ret_V_27_reg_1056[10], ret_V_27_reg_1056[10], ret_V_27_reg_1056[10], ret_V_27_reg_1056[10], ret_V_27_reg_1056, 2'h0 };
assign \add_35s_35s_35_2_1_U22.din1  = { op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18[3], op_18 };
assign grp_fu_650_p2 = \add_35s_35s_35_2_1_U22.dout ;
assign \add_35s_35s_35_2_1_U22.reset  = ap_rst;
assign \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_13_U.ain_s0  = \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_13_U.a ;
assign \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_13_U.bin_s0  = \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_13_U.b ;
assign \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_13_U.s  = { \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_13_U.fas_s2 , \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_13_U.sum_s1  };
assign \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_13_U.u2.a  = \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_13_U.ain_s1 ;
assign \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_13_U.u2.b  = \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_13_U.bin_s1 ;
assign \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_13_U.u2.cin  = \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_13_U.carry_s1 ;
assign \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_13_U.facout_s2  = \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_13_U.u2.cout ;
assign \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_13_U.fas_s2  = \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_13_U.u2.s ;
assign \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_13_U.u1.a  = \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_13_U.a [15:0];
assign \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_13_U.u1.b  = \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_13_U.b [15:0];
assign \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_13_U.u1.cin  = 1'h0;
assign \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_13_U.facout_s1  = \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_13_U.u1.cout ;
assign \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_13_U.fas_s1  = \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_13_U.u1.s ;
assign \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_13_U.a  = \add_32ns_32ns_32_2_1_U23.din0 ;
assign \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_13_U.b  = \add_32ns_32ns_32_2_1_U23.din1 ;
assign \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_13_U.ce  = \add_32ns_32ns_32_2_1_U23.ce ;
assign \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_13_U.clk  = \add_32ns_32ns_32_2_1_U23.clk ;
assign \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_13_U.reset  = \add_32ns_32ns_32_2_1_U23.reset ;
assign \add_32ns_32ns_32_2_1_U23.dout  = \add_32ns_32ns_32_2_1_U23.top_add_32ns_32ns_32_2_1_Adder_13_U.s ;
assign \add_32ns_32ns_32_2_1_U23.ce  = 1'h1;
assign \add_32ns_32ns_32_2_1_U23.clk  = ap_clk;
assign \add_32ns_32ns_32_2_1_U23.din0  = ret_V_30_cast_reg_1081;
assign \add_32ns_32ns_32_2_1_U23.din1  = 32'd1;
assign grp_fu_676_p2 = \add_32ns_32ns_32_2_1_U23.dout ;
assign \add_32ns_32ns_32_2_1_U23.reset  = ap_rst;
assign \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_3_U.ain_s0  = \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_3_U.a ;
assign \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_3_U.bin_s0  = \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_3_U.b ;
assign \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_3_U.s  = { \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_3_U.fas_s2 , \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_3_U.sum_s1  };
assign \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_3_U.u2.a  = \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_3_U.ain_s1 ;
assign \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_3_U.u2.b  = \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_3_U.bin_s1 ;
assign \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_3_U.u2.cin  = \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_3_U.carry_s1 ;
assign \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_3_U.facout_s2  = \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_3_U.u2.cout ;
assign \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_3_U.fas_s2  = \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_3_U.u2.s ;
assign \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_3_U.u1.a  = \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_3_U.a [0];
assign \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_3_U.u1.b  = \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_3_U.b [0];
assign \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_3_U.u1.cin  = 1'h0;
assign \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_3_U.facout_s1  = \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_3_U.u1.cout ;
assign \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_3_U.fas_s1  = \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_3_U.u1.s ;
assign \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_3_U.a  = \add_2ns_2ns_2_2_1_U5.din0 ;
assign \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_3_U.b  = \add_2ns_2ns_2_2_1_U5.din1 ;
assign \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_3_U.ce  = \add_2ns_2ns_2_2_1_U5.ce ;
assign \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_3_U.clk  = \add_2ns_2ns_2_2_1_U5.clk ;
assign \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_3_U.reset  = \add_2ns_2ns_2_2_1_U5.reset ;
assign \add_2ns_2ns_2_2_1_U5.dout  = \add_2ns_2ns_2_2_1_U5.top_add_2ns_2ns_2_2_1_Adder_3_U.s ;
assign \add_2ns_2ns_2_2_1_U5.ce  = 1'h1;
assign \add_2ns_2ns_2_2_1_U5.clk  = ap_clk;
assign \add_2ns_2ns_2_2_1_U5.din0  = ret_V_3_reg_780;
assign \add_2ns_2ns_2_2_1_U5.din1  = 2'h1;
assign grp_fu_307_p2 = \add_2ns_2ns_2_2_1_U5.dout ;
assign \add_2ns_2ns_2_2_1_U5.reset  = ap_rst;
assign \add_12ns_12s_12_2_1_U1.top_add_12ns_12s_12_2_1_Adder_0_U.ain_s0  = \add_12ns_12s_12_2_1_U1.top_add_12ns_12s_12_2_1_Adder_0_U.a ;
assign \add_12ns_12s_12_2_1_U1.top_add_12ns_12s_12_2_1_Adder_0_U.bin_s0  = \add_12ns_12s_12_2_1_U1.top_add_12ns_12s_12_2_1_Adder_0_U.b ;
assign \add_12ns_12s_12_2_1_U1.top_add_12ns_12s_12_2_1_Adder_0_U.s  = { \add_12ns_12s_12_2_1_U1.top_add_12ns_12s_12_2_1_Adder_0_U.fas_s2 , \add_12ns_12s_12_2_1_U1.top_add_12ns_12s_12_2_1_Adder_0_U.sum_s1  };
assign \add_12ns_12s_12_2_1_U1.top_add_12ns_12s_12_2_1_Adder_0_U.u2.a  = \add_12ns_12s_12_2_1_U1.top_add_12ns_12s_12_2_1_Adder_0_U.ain_s1 ;
assign \add_12ns_12s_12_2_1_U1.top_add_12ns_12s_12_2_1_Adder_0_U.u2.b  = \add_12ns_12s_12_2_1_U1.top_add_12ns_12s_12_2_1_Adder_0_U.bin_s1 ;
assign \add_12ns_12s_12_2_1_U1.top_add_12ns_12s_12_2_1_Adder_0_U.u2.cin  = \add_12ns_12s_12_2_1_U1.top_add_12ns_12s_12_2_1_Adder_0_U.carry_s1 ;
assign \add_12ns_12s_12_2_1_U1.top_add_12ns_12s_12_2_1_Adder_0_U.facout_s2  = \add_12ns_12s_12_2_1_U1.top_add_12ns_12s_12_2_1_Adder_0_U.u2.cout ;
assign \add_12ns_12s_12_2_1_U1.top_add_12ns_12s_12_2_1_Adder_0_U.fas_s2  = \add_12ns_12s_12_2_1_U1.top_add_12ns_12s_12_2_1_Adder_0_U.u2.s ;
assign \add_12ns_12s_12_2_1_U1.top_add_12ns_12s_12_2_1_Adder_0_U.u1.a  = \add_12ns_12s_12_2_1_U1.top_add_12ns_12s_12_2_1_Adder_0_U.a [5:0];
assign \add_12ns_12s_12_2_1_U1.top_add_12ns_12s_12_2_1_Adder_0_U.u1.b  = \add_12ns_12s_12_2_1_U1.top_add_12ns_12s_12_2_1_Adder_0_U.b [5:0];
assign \add_12ns_12s_12_2_1_U1.top_add_12ns_12s_12_2_1_Adder_0_U.u1.cin  = 1'h0;
assign \add_12ns_12s_12_2_1_U1.top_add_12ns_12s_12_2_1_Adder_0_U.facout_s1  = \add_12ns_12s_12_2_1_U1.top_add_12ns_12s_12_2_1_Adder_0_U.u1.cout ;
assign \add_12ns_12s_12_2_1_U1.top_add_12ns_12s_12_2_1_Adder_0_U.fas_s1  = \add_12ns_12s_12_2_1_U1.top_add_12ns_12s_12_2_1_Adder_0_U.u1.s ;
assign \add_12ns_12s_12_2_1_U1.top_add_12ns_12s_12_2_1_Adder_0_U.a  = \add_12ns_12s_12_2_1_U1.din0 ;
assign \add_12ns_12s_12_2_1_U1.top_add_12ns_12s_12_2_1_Adder_0_U.b  = \add_12ns_12s_12_2_1_U1.din1 ;
assign \add_12ns_12s_12_2_1_U1.top_add_12ns_12s_12_2_1_Adder_0_U.ce  = \add_12ns_12s_12_2_1_U1.ce ;
assign \add_12ns_12s_12_2_1_U1.top_add_12ns_12s_12_2_1_Adder_0_U.clk  = \add_12ns_12s_12_2_1_U1.clk ;
assign \add_12ns_12s_12_2_1_U1.top_add_12ns_12s_12_2_1_Adder_0_U.reset  = \add_12ns_12s_12_2_1_U1.reset ;
assign \add_12ns_12s_12_2_1_U1.dout  = \add_12ns_12s_12_2_1_U1.top_add_12ns_12s_12_2_1_Adder_0_U.s ;
assign \add_12ns_12s_12_2_1_U1.ce  = 1'h1;
assign \add_12ns_12s_12_2_1_U1.clk  = ap_clk;
assign \add_12ns_12s_12_2_1_U1.din0  = { 2'h0, op_2, 2'h0 };
assign \add_12ns_12s_12_2_1_U1.din1  = { op_1[3], op_1[3], op_1[3], op_1[3], op_1[3], op_1[3], op_1[3], op_1[3], op_1 };
assign grp_fu_189_p2 = \add_12ns_12s_12_2_1_U1.dout ;
assign \add_12ns_12s_12_2_1_U1.reset  = ap_rst;
assign \add_11s_11ns_11_2_1_U6.top_add_11s_11ns_11_2_1_Adder_4_U.ain_s0  = \add_11s_11ns_11_2_1_U6.top_add_11s_11ns_11_2_1_Adder_4_U.a ;
assign \add_11s_11ns_11_2_1_U6.top_add_11s_11ns_11_2_1_Adder_4_U.bin_s0  = \add_11s_11ns_11_2_1_U6.top_add_11s_11ns_11_2_1_Adder_4_U.b ;
assign \add_11s_11ns_11_2_1_U6.top_add_11s_11ns_11_2_1_Adder_4_U.s  = { \add_11s_11ns_11_2_1_U6.top_add_11s_11ns_11_2_1_Adder_4_U.fas_s2 , \add_11s_11ns_11_2_1_U6.top_add_11s_11ns_11_2_1_Adder_4_U.sum_s1  };
assign \add_11s_11ns_11_2_1_U6.top_add_11s_11ns_11_2_1_Adder_4_U.u2.a  = \add_11s_11ns_11_2_1_U6.top_add_11s_11ns_11_2_1_Adder_4_U.ain_s1 ;
assign \add_11s_11ns_11_2_1_U6.top_add_11s_11ns_11_2_1_Adder_4_U.u2.b  = \add_11s_11ns_11_2_1_U6.top_add_11s_11ns_11_2_1_Adder_4_U.bin_s1 ;
assign \add_11s_11ns_11_2_1_U6.top_add_11s_11ns_11_2_1_Adder_4_U.u2.cin  = \add_11s_11ns_11_2_1_U6.top_add_11s_11ns_11_2_1_Adder_4_U.carry_s1 ;
assign \add_11s_11ns_11_2_1_U6.top_add_11s_11ns_11_2_1_Adder_4_U.facout_s2  = \add_11s_11ns_11_2_1_U6.top_add_11s_11ns_11_2_1_Adder_4_U.u2.cout ;
assign \add_11s_11ns_11_2_1_U6.top_add_11s_11ns_11_2_1_Adder_4_U.fas_s2  = \add_11s_11ns_11_2_1_U6.top_add_11s_11ns_11_2_1_Adder_4_U.u2.s ;
assign \add_11s_11ns_11_2_1_U6.top_add_11s_11ns_11_2_1_Adder_4_U.u1.a  = \add_11s_11ns_11_2_1_U6.top_add_11s_11ns_11_2_1_Adder_4_U.a [4:0];
assign \add_11s_11ns_11_2_1_U6.top_add_11s_11ns_11_2_1_Adder_4_U.u1.b  = \add_11s_11ns_11_2_1_U6.top_add_11s_11ns_11_2_1_Adder_4_U.b [4:0];
assign \add_11s_11ns_11_2_1_U6.top_add_11s_11ns_11_2_1_Adder_4_U.u1.cin  = 1'h0;
assign \add_11s_11ns_11_2_1_U6.top_add_11s_11ns_11_2_1_Adder_4_U.facout_s1  = \add_11s_11ns_11_2_1_U6.top_add_11s_11ns_11_2_1_Adder_4_U.u1.cout ;
assign \add_11s_11ns_11_2_1_U6.top_add_11s_11ns_11_2_1_Adder_4_U.fas_s1  = \add_11s_11ns_11_2_1_U6.top_add_11s_11ns_11_2_1_Adder_4_U.u1.s ;
assign \add_11s_11ns_11_2_1_U6.top_add_11s_11ns_11_2_1_Adder_4_U.a  = \add_11s_11ns_11_2_1_U6.din0 ;
assign \add_11s_11ns_11_2_1_U6.top_add_11s_11ns_11_2_1_Adder_4_U.b  = \add_11s_11ns_11_2_1_U6.din1 ;
assign \add_11s_11ns_11_2_1_U6.top_add_11s_11ns_11_2_1_Adder_4_U.ce  = \add_11s_11ns_11_2_1_U6.ce ;
assign \add_11s_11ns_11_2_1_U6.top_add_11s_11ns_11_2_1_Adder_4_U.clk  = \add_11s_11ns_11_2_1_U6.clk ;
assign \add_11s_11ns_11_2_1_U6.top_add_11s_11ns_11_2_1_Adder_4_U.reset  = \add_11s_11ns_11_2_1_U6.reset ;
assign \add_11s_11ns_11_2_1_U6.dout  = \add_11s_11ns_11_2_1_U6.top_add_11s_11ns_11_2_1_Adder_4_U.s ;
assign \add_11s_11ns_11_2_1_U6.ce  = 1'h1;
assign \add_11s_11ns_11_2_1_U6.clk  = ap_clk;
assign \add_11s_11ns_11_2_1_U6.din0  = { ret_V_8_reg_813[9], ret_V_8_reg_813 };
assign \add_11s_11ns_11_2_1_U6.din1  = 11'h001;
assign grp_fu_377_p2 = \add_11s_11ns_11_2_1_U6.dout ;
assign \add_11s_11ns_11_2_1_U6.reset  = ap_rst;
assign \add_11s_11ns_11_2_1_U13.top_add_11s_11ns_11_2_1_Adder_4_U.ain_s0  = \add_11s_11ns_11_2_1_U13.top_add_11s_11ns_11_2_1_Adder_4_U.a ;
assign \add_11s_11ns_11_2_1_U13.top_add_11s_11ns_11_2_1_Adder_4_U.bin_s0  = \add_11s_11ns_11_2_1_U13.top_add_11s_11ns_11_2_1_Adder_4_U.b ;
assign \add_11s_11ns_11_2_1_U13.top_add_11s_11ns_11_2_1_Adder_4_U.s  = { \add_11s_11ns_11_2_1_U13.top_add_11s_11ns_11_2_1_Adder_4_U.fas_s2 , \add_11s_11ns_11_2_1_U13.top_add_11s_11ns_11_2_1_Adder_4_U.sum_s1  };
assign \add_11s_11ns_11_2_1_U13.top_add_11s_11ns_11_2_1_Adder_4_U.u2.a  = \add_11s_11ns_11_2_1_U13.top_add_11s_11ns_11_2_1_Adder_4_U.ain_s1 ;
assign \add_11s_11ns_11_2_1_U13.top_add_11s_11ns_11_2_1_Adder_4_U.u2.b  = \add_11s_11ns_11_2_1_U13.top_add_11s_11ns_11_2_1_Adder_4_U.bin_s1 ;
assign \add_11s_11ns_11_2_1_U13.top_add_11s_11ns_11_2_1_Adder_4_U.u2.cin  = \add_11s_11ns_11_2_1_U13.top_add_11s_11ns_11_2_1_Adder_4_U.carry_s1 ;
assign \add_11s_11ns_11_2_1_U13.top_add_11s_11ns_11_2_1_Adder_4_U.facout_s2  = \add_11s_11ns_11_2_1_U13.top_add_11s_11ns_11_2_1_Adder_4_U.u2.cout ;
assign \add_11s_11ns_11_2_1_U13.top_add_11s_11ns_11_2_1_Adder_4_U.fas_s2  = \add_11s_11ns_11_2_1_U13.top_add_11s_11ns_11_2_1_Adder_4_U.u2.s ;
assign \add_11s_11ns_11_2_1_U13.top_add_11s_11ns_11_2_1_Adder_4_U.u1.a  = \add_11s_11ns_11_2_1_U13.top_add_11s_11ns_11_2_1_Adder_4_U.a [4:0];
assign \add_11s_11ns_11_2_1_U13.top_add_11s_11ns_11_2_1_Adder_4_U.u1.b  = \add_11s_11ns_11_2_1_U13.top_add_11s_11ns_11_2_1_Adder_4_U.b [4:0];
assign \add_11s_11ns_11_2_1_U13.top_add_11s_11ns_11_2_1_Adder_4_U.u1.cin  = 1'h0;
assign \add_11s_11ns_11_2_1_U13.top_add_11s_11ns_11_2_1_Adder_4_U.facout_s1  = \add_11s_11ns_11_2_1_U13.top_add_11s_11ns_11_2_1_Adder_4_U.u1.cout ;
assign \add_11s_11ns_11_2_1_U13.top_add_11s_11ns_11_2_1_Adder_4_U.fas_s1  = \add_11s_11ns_11_2_1_U13.top_add_11s_11ns_11_2_1_Adder_4_U.u1.s ;
assign \add_11s_11ns_11_2_1_U13.top_add_11s_11ns_11_2_1_Adder_4_U.a  = \add_11s_11ns_11_2_1_U13.din0 ;
assign \add_11s_11ns_11_2_1_U13.top_add_11s_11ns_11_2_1_Adder_4_U.b  = \add_11s_11ns_11_2_1_U13.din1 ;
assign \add_11s_11ns_11_2_1_U13.top_add_11s_11ns_11_2_1_Adder_4_U.ce  = \add_11s_11ns_11_2_1_U13.ce ;
assign \add_11s_11ns_11_2_1_U13.top_add_11s_11ns_11_2_1_Adder_4_U.clk  = \add_11s_11ns_11_2_1_U13.clk ;
assign \add_11s_11ns_11_2_1_U13.top_add_11s_11ns_11_2_1_Adder_4_U.reset  = \add_11s_11ns_11_2_1_U13.reset ;
assign \add_11s_11ns_11_2_1_U13.dout  = \add_11s_11ns_11_2_1_U13.top_add_11s_11ns_11_2_1_Adder_4_U.s ;
assign \add_11s_11ns_11_2_1_U13.ce  = 1'h1;
assign \add_11s_11ns_11_2_1_U13.clk  = ap_clk;
assign \add_11s_11ns_11_2_1_U13.din0  = { add_ln69_2_reg_922[5], add_ln69_2_reg_922[5], add_ln69_2_reg_922[5], add_ln69_2_reg_922[5], add_ln69_2_reg_922[5], add_ln69_2_reg_922 };
assign \add_11s_11ns_11_2_1_U13.din1  = add_ln69_reg_917;
assign grp_fu_471_p2 = \add_11s_11ns_11_2_1_U13.dout ;
assign \add_11s_11ns_11_2_1_U13.reset  = ap_rst;
assign \add_11ns_11s_11_2_1_U21.top_add_11ns_11s_11_2_1_Adder_7_U.ain_s0  = \add_11ns_11s_11_2_1_U21.top_add_11ns_11s_11_2_1_Adder_7_U.a ;
assign \add_11ns_11s_11_2_1_U21.top_add_11ns_11s_11_2_1_Adder_7_U.bin_s0  = \add_11ns_11s_11_2_1_U21.top_add_11ns_11s_11_2_1_Adder_7_U.b ;
assign \add_11ns_11s_11_2_1_U21.top_add_11ns_11s_11_2_1_Adder_7_U.s  = { \add_11ns_11s_11_2_1_U21.top_add_11ns_11s_11_2_1_Adder_7_U.fas_s2 , \add_11ns_11s_11_2_1_U21.top_add_11ns_11s_11_2_1_Adder_7_U.sum_s1  };
assign \add_11ns_11s_11_2_1_U21.top_add_11ns_11s_11_2_1_Adder_7_U.u2.a  = \add_11ns_11s_11_2_1_U21.top_add_11ns_11s_11_2_1_Adder_7_U.ain_s1 ;
assign \add_11ns_11s_11_2_1_U21.top_add_11ns_11s_11_2_1_Adder_7_U.u2.b  = \add_11ns_11s_11_2_1_U21.top_add_11ns_11s_11_2_1_Adder_7_U.bin_s1 ;
assign \add_11ns_11s_11_2_1_U21.top_add_11ns_11s_11_2_1_Adder_7_U.u2.cin  = \add_11ns_11s_11_2_1_U21.top_add_11ns_11s_11_2_1_Adder_7_U.carry_s1 ;
assign \add_11ns_11s_11_2_1_U21.top_add_11ns_11s_11_2_1_Adder_7_U.facout_s2  = \add_11ns_11s_11_2_1_U21.top_add_11ns_11s_11_2_1_Adder_7_U.u2.cout ;
assign \add_11ns_11s_11_2_1_U21.top_add_11ns_11s_11_2_1_Adder_7_U.fas_s2  = \add_11ns_11s_11_2_1_U21.top_add_11ns_11s_11_2_1_Adder_7_U.u2.s ;
assign \add_11ns_11s_11_2_1_U21.top_add_11ns_11s_11_2_1_Adder_7_U.u1.a  = \add_11ns_11s_11_2_1_U21.top_add_11ns_11s_11_2_1_Adder_7_U.a [4:0];
assign \add_11ns_11s_11_2_1_U21.top_add_11ns_11s_11_2_1_Adder_7_U.u1.b  = \add_11ns_11s_11_2_1_U21.top_add_11ns_11s_11_2_1_Adder_7_U.b [4:0];
assign \add_11ns_11s_11_2_1_U21.top_add_11ns_11s_11_2_1_Adder_7_U.u1.cin  = 1'h0;
assign \add_11ns_11s_11_2_1_U21.top_add_11ns_11s_11_2_1_Adder_7_U.facout_s1  = \add_11ns_11s_11_2_1_U21.top_add_11ns_11s_11_2_1_Adder_7_U.u1.cout ;
assign \add_11ns_11s_11_2_1_U21.top_add_11ns_11s_11_2_1_Adder_7_U.fas_s1  = \add_11ns_11s_11_2_1_U21.top_add_11ns_11s_11_2_1_Adder_7_U.u1.s ;
assign \add_11ns_11s_11_2_1_U21.top_add_11ns_11s_11_2_1_Adder_7_U.a  = \add_11ns_11s_11_2_1_U21.din0 ;
assign \add_11ns_11s_11_2_1_U21.top_add_11ns_11s_11_2_1_Adder_7_U.b  = \add_11ns_11s_11_2_1_U21.din1 ;
assign \add_11ns_11s_11_2_1_U21.top_add_11ns_11s_11_2_1_Adder_7_U.ce  = \add_11ns_11s_11_2_1_U21.ce ;
assign \add_11ns_11s_11_2_1_U21.top_add_11ns_11s_11_2_1_Adder_7_U.clk  = \add_11ns_11s_11_2_1_U21.clk ;
assign \add_11ns_11s_11_2_1_U21.top_add_11ns_11s_11_2_1_Adder_7_U.reset  = \add_11ns_11s_11_2_1_U21.reset ;
assign \add_11ns_11s_11_2_1_U21.dout  = \add_11ns_11s_11_2_1_U21.top_add_11ns_11s_11_2_1_Adder_7_U.s ;
assign \add_11ns_11s_11_2_1_U21.ce  = 1'h1;
assign \add_11ns_11s_11_2_1_U21.clk  = ap_clk;
assign \add_11ns_11s_11_2_1_U21.din0  = op_27_V_reg_1046;
assign \add_11ns_11s_11_2_1_U21.din1  = { r_reg_1041[5], r_reg_1041[5], r_reg_1041[5], r_reg_1041[5], r_reg_1041[5], r_reg_1041 };
assign grp_fu_630_p2 = \add_11ns_11s_11_2_1_U21.dout ;
assign \add_11ns_11s_11_2_1_U21.reset  = ap_rst;
assign \add_11ns_11s_11_2_1_U20.top_add_11ns_11s_11_2_1_Adder_7_U.ain_s0  = \add_11ns_11s_11_2_1_U20.top_add_11ns_11s_11_2_1_Adder_7_U.a ;
assign \add_11ns_11s_11_2_1_U20.top_add_11ns_11s_11_2_1_Adder_7_U.bin_s0  = \add_11ns_11s_11_2_1_U20.top_add_11ns_11s_11_2_1_Adder_7_U.b ;
assign \add_11ns_11s_11_2_1_U20.top_add_11ns_11s_11_2_1_Adder_7_U.s  = { \add_11ns_11s_11_2_1_U20.top_add_11ns_11s_11_2_1_Adder_7_U.fas_s2 , \add_11ns_11s_11_2_1_U20.top_add_11ns_11s_11_2_1_Adder_7_U.sum_s1  };
assign \add_11ns_11s_11_2_1_U20.top_add_11ns_11s_11_2_1_Adder_7_U.u2.a  = \add_11ns_11s_11_2_1_U20.top_add_11ns_11s_11_2_1_Adder_7_U.ain_s1 ;
assign \add_11ns_11s_11_2_1_U20.top_add_11ns_11s_11_2_1_Adder_7_U.u2.b  = \add_11ns_11s_11_2_1_U20.top_add_11ns_11s_11_2_1_Adder_7_U.bin_s1 ;
assign \add_11ns_11s_11_2_1_U20.top_add_11ns_11s_11_2_1_Adder_7_U.u2.cin  = \add_11ns_11s_11_2_1_U20.top_add_11ns_11s_11_2_1_Adder_7_U.carry_s1 ;
assign \add_11ns_11s_11_2_1_U20.top_add_11ns_11s_11_2_1_Adder_7_U.facout_s2  = \add_11ns_11s_11_2_1_U20.top_add_11ns_11s_11_2_1_Adder_7_U.u2.cout ;
assign \add_11ns_11s_11_2_1_U20.top_add_11ns_11s_11_2_1_Adder_7_U.fas_s2  = \add_11ns_11s_11_2_1_U20.top_add_11ns_11s_11_2_1_Adder_7_U.u2.s ;
assign \add_11ns_11s_11_2_1_U20.top_add_11ns_11s_11_2_1_Adder_7_U.u1.a  = \add_11ns_11s_11_2_1_U20.top_add_11ns_11s_11_2_1_Adder_7_U.a [4:0];
assign \add_11ns_11s_11_2_1_U20.top_add_11ns_11s_11_2_1_Adder_7_U.u1.b  = \add_11ns_11s_11_2_1_U20.top_add_11ns_11s_11_2_1_Adder_7_U.b [4:0];
assign \add_11ns_11s_11_2_1_U20.top_add_11ns_11s_11_2_1_Adder_7_U.u1.cin  = 1'h0;
assign \add_11ns_11s_11_2_1_U20.top_add_11ns_11s_11_2_1_Adder_7_U.facout_s1  = \add_11ns_11s_11_2_1_U20.top_add_11ns_11s_11_2_1_Adder_7_U.u1.cout ;
assign \add_11ns_11s_11_2_1_U20.top_add_11ns_11s_11_2_1_Adder_7_U.fas_s1  = \add_11ns_11s_11_2_1_U20.top_add_11ns_11s_11_2_1_Adder_7_U.u1.s ;
assign \add_11ns_11s_11_2_1_U20.top_add_11ns_11s_11_2_1_Adder_7_U.a  = \add_11ns_11s_11_2_1_U20.din0 ;
assign \add_11ns_11s_11_2_1_U20.top_add_11ns_11s_11_2_1_Adder_7_U.b  = \add_11ns_11s_11_2_1_U20.din1 ;
assign \add_11ns_11s_11_2_1_U20.top_add_11ns_11s_11_2_1_Adder_7_U.ce  = \add_11ns_11s_11_2_1_U20.ce ;
assign \add_11ns_11s_11_2_1_U20.top_add_11ns_11s_11_2_1_Adder_7_U.clk  = \add_11ns_11s_11_2_1_U20.clk ;
assign \add_11ns_11s_11_2_1_U20.top_add_11ns_11s_11_2_1_Adder_7_U.reset  = \add_11ns_11s_11_2_1_U20.reset ;
assign \add_11ns_11s_11_2_1_U20.dout  = \add_11ns_11s_11_2_1_U20.top_add_11ns_11s_11_2_1_Adder_7_U.s ;
assign \add_11ns_11s_11_2_1_U20.ce  = 1'h1;
assign \add_11ns_11s_11_2_1_U20.clk  = ap_clk;
assign \add_11ns_11s_11_2_1_U20.din0  = ret_V_26_reg_1000;
assign \add_11ns_11s_11_2_1_U20.din1  = { op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16[3], op_16 };
assign grp_fu_613_p2 = \add_11ns_11s_11_2_1_U20.dout ;
assign \add_11ns_11s_11_2_1_U20.reset  = ap_rst;
assign \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_7_U.ain_s0  = \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_7_U.a ;
assign \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_7_U.bin_s0  = \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_7_U.b ;
assign \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_7_U.s  = { \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_7_U.fas_s2 , \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_7_U.sum_s1  };
assign \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_7_U.u2.a  = \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_7_U.ain_s1 ;
assign \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_7_U.u2.b  = \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_7_U.bin_s1 ;
assign \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_7_U.u2.cin  = \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_7_U.carry_s1 ;
assign \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_7_U.facout_s2  = \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_7_U.u2.cout ;
assign \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_7_U.fas_s2  = \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_7_U.u2.s ;
assign \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_7_U.u1.a  = \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_7_U.a [4:0];
assign \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_7_U.u1.b  = \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_7_U.b [4:0];
assign \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_7_U.u1.cin  = 1'h0;
assign \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_7_U.facout_s1  = \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_7_U.u1.cout ;
assign \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_7_U.fas_s1  = \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_7_U.u1.s ;
assign \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_7_U.a  = \add_11ns_11s_11_2_1_U11.din0 ;
assign \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_7_U.b  = \add_11ns_11s_11_2_1_U11.din1 ;
assign \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_7_U.ce  = \add_11ns_11s_11_2_1_U11.ce ;
assign \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_7_U.clk  = \add_11ns_11s_11_2_1_U11.clk ;
assign \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_7_U.reset  = \add_11ns_11s_11_2_1_U11.reset ;
assign \add_11ns_11s_11_2_1_U11.dout  = \add_11ns_11s_11_2_1_U11.top_add_11ns_11s_11_2_1_Adder_7_U.s ;
assign \add_11ns_11s_11_2_1_U11.ce  = 1'h1;
assign \add_11ns_11s_11_2_1_U11.clk  = ap_clk;
assign \add_11ns_11s_11_2_1_U11.din0  = ret_V_23_reg_887;
assign \add_11ns_11s_11_2_1_U11.din1  = { ret_reg_892[2], ret_reg_892[2], ret_reg_892[2], ret_reg_892[2], ret_reg_892[2], ret_reg_892[2], ret_reg_892[2], ret_reg_892[2], ret_reg_892 };
assign grp_fu_454_p2 = \add_11ns_11s_11_2_1_U11.dout ;
assign \add_11ns_11s_11_2_1_U11.reset  = ap_rst;
assign \add_11ns_11ns_11_2_1_U16.top_add_11ns_11ns_11_2_1_Adder_9_U.ain_s0  = \add_11ns_11ns_11_2_1_U16.top_add_11ns_11ns_11_2_1_Adder_9_U.a ;
assign \add_11ns_11ns_11_2_1_U16.top_add_11ns_11ns_11_2_1_Adder_9_U.bin_s0  = \add_11ns_11ns_11_2_1_U16.top_add_11ns_11ns_11_2_1_Adder_9_U.b ;
assign \add_11ns_11ns_11_2_1_U16.top_add_11ns_11ns_11_2_1_Adder_9_U.s  = { \add_11ns_11ns_11_2_1_U16.top_add_11ns_11ns_11_2_1_Adder_9_U.fas_s2 , \add_11ns_11ns_11_2_1_U16.top_add_11ns_11ns_11_2_1_Adder_9_U.sum_s1  };
assign \add_11ns_11ns_11_2_1_U16.top_add_11ns_11ns_11_2_1_Adder_9_U.u2.a  = \add_11ns_11ns_11_2_1_U16.top_add_11ns_11ns_11_2_1_Adder_9_U.ain_s1 ;
assign \add_11ns_11ns_11_2_1_U16.top_add_11ns_11ns_11_2_1_Adder_9_U.u2.b  = \add_11ns_11ns_11_2_1_U16.top_add_11ns_11ns_11_2_1_Adder_9_U.bin_s1 ;
assign \add_11ns_11ns_11_2_1_U16.top_add_11ns_11ns_11_2_1_Adder_9_U.u2.cin  = \add_11ns_11ns_11_2_1_U16.top_add_11ns_11ns_11_2_1_Adder_9_U.carry_s1 ;
assign \add_11ns_11ns_11_2_1_U16.top_add_11ns_11ns_11_2_1_Adder_9_U.facout_s2  = \add_11ns_11ns_11_2_1_U16.top_add_11ns_11ns_11_2_1_Adder_9_U.u2.cout ;
assign \add_11ns_11ns_11_2_1_U16.top_add_11ns_11ns_11_2_1_Adder_9_U.fas_s2  = \add_11ns_11ns_11_2_1_U16.top_add_11ns_11ns_11_2_1_Adder_9_U.u2.s ;
assign \add_11ns_11ns_11_2_1_U16.top_add_11ns_11ns_11_2_1_Adder_9_U.u1.a  = \add_11ns_11ns_11_2_1_U16.top_add_11ns_11ns_11_2_1_Adder_9_U.a [4:0];
assign \add_11ns_11ns_11_2_1_U16.top_add_11ns_11ns_11_2_1_Adder_9_U.u1.b  = \add_11ns_11ns_11_2_1_U16.top_add_11ns_11ns_11_2_1_Adder_9_U.b [4:0];
assign \add_11ns_11ns_11_2_1_U16.top_add_11ns_11ns_11_2_1_Adder_9_U.u1.cin  = 1'h0;
assign \add_11ns_11ns_11_2_1_U16.top_add_11ns_11ns_11_2_1_Adder_9_U.facout_s1  = \add_11ns_11ns_11_2_1_U16.top_add_11ns_11ns_11_2_1_Adder_9_U.u1.cout ;
assign \add_11ns_11ns_11_2_1_U16.top_add_11ns_11ns_11_2_1_Adder_9_U.fas_s1  = \add_11ns_11ns_11_2_1_U16.top_add_11ns_11ns_11_2_1_Adder_9_U.u1.s ;
assign \add_11ns_11ns_11_2_1_U16.top_add_11ns_11ns_11_2_1_Adder_9_U.a  = \add_11ns_11ns_11_2_1_U16.din0 ;
assign \add_11ns_11ns_11_2_1_U16.top_add_11ns_11ns_11_2_1_Adder_9_U.b  = \add_11ns_11ns_11_2_1_U16.din1 ;
assign \add_11ns_11ns_11_2_1_U16.top_add_11ns_11ns_11_2_1_Adder_9_U.ce  = \add_11ns_11ns_11_2_1_U16.ce ;
assign \add_11ns_11ns_11_2_1_U16.top_add_11ns_11ns_11_2_1_Adder_9_U.clk  = \add_11ns_11ns_11_2_1_U16.clk ;
assign \add_11ns_11ns_11_2_1_U16.top_add_11ns_11ns_11_2_1_Adder_9_U.reset  = \add_11ns_11ns_11_2_1_U16.reset ;
assign \add_11ns_11ns_11_2_1_U16.dout  = \add_11ns_11ns_11_2_1_U16.top_add_11ns_11ns_11_2_1_Adder_9_U.s ;
assign \add_11ns_11ns_11_2_1_U16.ce  = 1'h1;
assign \add_11ns_11ns_11_2_1_U16.clk  = ap_clk;
assign \add_11ns_11ns_11_2_1_U16.din0  = ret_V_25_reg_965;
assign \add_11ns_11ns_11_2_1_U16.din1  = 11'h001;
assign grp_fu_508_p2 = \add_11ns_11ns_11_2_1_U16.dout ;
assign \add_11ns_11ns_11_2_1_U16.reset  = ap_rst;
assign \add_11ns_11ns_11_2_1_U14.top_add_11ns_11ns_11_2_1_Adder_9_U.ain_s0  = \add_11ns_11ns_11_2_1_U14.top_add_11ns_11ns_11_2_1_Adder_9_U.a ;
assign \add_11ns_11ns_11_2_1_U14.top_add_11ns_11ns_11_2_1_Adder_9_U.bin_s0  = \add_11ns_11ns_11_2_1_U14.top_add_11ns_11ns_11_2_1_Adder_9_U.b ;
assign \add_11ns_11ns_11_2_1_U14.top_add_11ns_11ns_11_2_1_Adder_9_U.s  = { \add_11ns_11ns_11_2_1_U14.top_add_11ns_11ns_11_2_1_Adder_9_U.fas_s2 , \add_11ns_11ns_11_2_1_U14.top_add_11ns_11ns_11_2_1_Adder_9_U.sum_s1  };
assign \add_11ns_11ns_11_2_1_U14.top_add_11ns_11ns_11_2_1_Adder_9_U.u2.a  = \add_11ns_11ns_11_2_1_U14.top_add_11ns_11ns_11_2_1_Adder_9_U.ain_s1 ;
assign \add_11ns_11ns_11_2_1_U14.top_add_11ns_11ns_11_2_1_Adder_9_U.u2.b  = \add_11ns_11ns_11_2_1_U14.top_add_11ns_11ns_11_2_1_Adder_9_U.bin_s1 ;
assign \add_11ns_11ns_11_2_1_U14.top_add_11ns_11ns_11_2_1_Adder_9_U.u2.cin  = \add_11ns_11ns_11_2_1_U14.top_add_11ns_11ns_11_2_1_Adder_9_U.carry_s1 ;
assign \add_11ns_11ns_11_2_1_U14.top_add_11ns_11ns_11_2_1_Adder_9_U.facout_s2  = \add_11ns_11ns_11_2_1_U14.top_add_11ns_11ns_11_2_1_Adder_9_U.u2.cout ;
assign \add_11ns_11ns_11_2_1_U14.top_add_11ns_11ns_11_2_1_Adder_9_U.fas_s2  = \add_11ns_11ns_11_2_1_U14.top_add_11ns_11ns_11_2_1_Adder_9_U.u2.s ;
assign \add_11ns_11ns_11_2_1_U14.top_add_11ns_11ns_11_2_1_Adder_9_U.u1.a  = \add_11ns_11ns_11_2_1_U14.top_add_11ns_11ns_11_2_1_Adder_9_U.a [4:0];
assign \add_11ns_11ns_11_2_1_U14.top_add_11ns_11ns_11_2_1_Adder_9_U.u1.b  = \add_11ns_11ns_11_2_1_U14.top_add_11ns_11ns_11_2_1_Adder_9_U.b [4:0];
assign \add_11ns_11ns_11_2_1_U14.top_add_11ns_11ns_11_2_1_Adder_9_U.u1.cin  = 1'h0;
assign \add_11ns_11ns_11_2_1_U14.top_add_11ns_11ns_11_2_1_Adder_9_U.facout_s1  = \add_11ns_11ns_11_2_1_U14.top_add_11ns_11ns_11_2_1_Adder_9_U.u1.cout ;
assign \add_11ns_11ns_11_2_1_U14.top_add_11ns_11ns_11_2_1_Adder_9_U.fas_s1  = \add_11ns_11ns_11_2_1_U14.top_add_11ns_11ns_11_2_1_Adder_9_U.u1.s ;
assign \add_11ns_11ns_11_2_1_U14.top_add_11ns_11ns_11_2_1_Adder_9_U.a  = \add_11ns_11ns_11_2_1_U14.din0 ;
assign \add_11ns_11ns_11_2_1_U14.top_add_11ns_11ns_11_2_1_Adder_9_U.b  = \add_11ns_11ns_11_2_1_U14.din1 ;
assign \add_11ns_11ns_11_2_1_U14.top_add_11ns_11ns_11_2_1_Adder_9_U.ce  = \add_11ns_11ns_11_2_1_U14.ce ;
assign \add_11ns_11ns_11_2_1_U14.top_add_11ns_11ns_11_2_1_Adder_9_U.clk  = \add_11ns_11ns_11_2_1_U14.clk ;
assign \add_11ns_11ns_11_2_1_U14.top_add_11ns_11ns_11_2_1_Adder_9_U.reset  = \add_11ns_11ns_11_2_1_U14.reset ;
assign \add_11ns_11ns_11_2_1_U14.dout  = \add_11ns_11ns_11_2_1_U14.top_add_11ns_11ns_11_2_1_Adder_9_U.s ;
assign \add_11ns_11ns_11_2_1_U14.ce  = 1'h1;
assign \add_11ns_11ns_11_2_1_U14.clk  = ap_clk;
assign \add_11ns_11ns_11_2_1_U14.din0  = op_24_V_reg_942;
assign \add_11ns_11ns_11_2_1_U14.din1  = select_ln1192_reg_947;
assign grp_fu_499_p2 = \add_11ns_11ns_11_2_1_U14.dout ;
assign \add_11ns_11ns_11_2_1_U14.reset  = ap_rst;
assign \add_10ns_10ns_10_2_1_U3.top_add_10ns_10ns_10_2_1_Adder_1_U.ain_s0  = \add_10ns_10ns_10_2_1_U3.top_add_10ns_10ns_10_2_1_Adder_1_U.a ;
assign \add_10ns_10ns_10_2_1_U3.top_add_10ns_10ns_10_2_1_Adder_1_U.bin_s0  = \add_10ns_10ns_10_2_1_U3.top_add_10ns_10ns_10_2_1_Adder_1_U.b ;
assign \add_10ns_10ns_10_2_1_U3.top_add_10ns_10ns_10_2_1_Adder_1_U.s  = { \add_10ns_10ns_10_2_1_U3.top_add_10ns_10ns_10_2_1_Adder_1_U.fas_s2 , \add_10ns_10ns_10_2_1_U3.top_add_10ns_10ns_10_2_1_Adder_1_U.sum_s1  };
assign \add_10ns_10ns_10_2_1_U3.top_add_10ns_10ns_10_2_1_Adder_1_U.u2.a  = \add_10ns_10ns_10_2_1_U3.top_add_10ns_10ns_10_2_1_Adder_1_U.ain_s1 ;
assign \add_10ns_10ns_10_2_1_U3.top_add_10ns_10ns_10_2_1_Adder_1_U.u2.b  = \add_10ns_10ns_10_2_1_U3.top_add_10ns_10ns_10_2_1_Adder_1_U.bin_s1 ;
assign \add_10ns_10ns_10_2_1_U3.top_add_10ns_10ns_10_2_1_Adder_1_U.u2.cin  = \add_10ns_10ns_10_2_1_U3.top_add_10ns_10ns_10_2_1_Adder_1_U.carry_s1 ;
assign \add_10ns_10ns_10_2_1_U3.top_add_10ns_10ns_10_2_1_Adder_1_U.facout_s2  = \add_10ns_10ns_10_2_1_U3.top_add_10ns_10ns_10_2_1_Adder_1_U.u2.cout ;
assign \add_10ns_10ns_10_2_1_U3.top_add_10ns_10ns_10_2_1_Adder_1_U.fas_s2  = \add_10ns_10ns_10_2_1_U3.top_add_10ns_10ns_10_2_1_Adder_1_U.u2.s ;
assign \add_10ns_10ns_10_2_1_U3.top_add_10ns_10ns_10_2_1_Adder_1_U.u1.a  = \add_10ns_10ns_10_2_1_U3.top_add_10ns_10ns_10_2_1_Adder_1_U.a [4:0];
assign \add_10ns_10ns_10_2_1_U3.top_add_10ns_10ns_10_2_1_Adder_1_U.u1.b  = \add_10ns_10ns_10_2_1_U3.top_add_10ns_10ns_10_2_1_Adder_1_U.b [4:0];
assign \add_10ns_10ns_10_2_1_U3.top_add_10ns_10ns_10_2_1_Adder_1_U.u1.cin  = 1'h0;
assign \add_10ns_10ns_10_2_1_U3.top_add_10ns_10ns_10_2_1_Adder_1_U.facout_s1  = \add_10ns_10ns_10_2_1_U3.top_add_10ns_10ns_10_2_1_Adder_1_U.u1.cout ;
assign \add_10ns_10ns_10_2_1_U3.top_add_10ns_10ns_10_2_1_Adder_1_U.fas_s1  = \add_10ns_10ns_10_2_1_U3.top_add_10ns_10ns_10_2_1_Adder_1_U.u1.s ;
assign \add_10ns_10ns_10_2_1_U3.top_add_10ns_10ns_10_2_1_Adder_1_U.a  = \add_10ns_10ns_10_2_1_U3.din0 ;
assign \add_10ns_10ns_10_2_1_U3.top_add_10ns_10ns_10_2_1_Adder_1_U.b  = \add_10ns_10ns_10_2_1_U3.din1 ;
assign \add_10ns_10ns_10_2_1_U3.top_add_10ns_10ns_10_2_1_Adder_1_U.ce  = \add_10ns_10ns_10_2_1_U3.ce ;
assign \add_10ns_10ns_10_2_1_U3.top_add_10ns_10ns_10_2_1_Adder_1_U.clk  = \add_10ns_10ns_10_2_1_U3.clk ;
assign \add_10ns_10ns_10_2_1_U3.top_add_10ns_10ns_10_2_1_Adder_1_U.reset  = \add_10ns_10ns_10_2_1_U3.reset ;
assign \add_10ns_10ns_10_2_1_U3.dout  = \add_10ns_10ns_10_2_1_U3.top_add_10ns_10ns_10_2_1_Adder_1_U.s ;
assign \add_10ns_10ns_10_2_1_U3.ce  = 1'h1;
assign \add_10ns_10ns_10_2_1_U3.clk  = ap_clk;
assign \add_10ns_10ns_10_2_1_U3.din0  = ret_V_reg_741;
assign \add_10ns_10ns_10_2_1_U3.din1  = 10'h001;
assign grp_fu_239_p2 = \add_10ns_10ns_10_2_1_U3.dout ;
assign \add_10ns_10ns_10_2_1_U3.reset  = ap_rst;
endmodule


// Product machine:
module top_A_times_top_B (ap_start, op_0, op_1, op_12, op_14, op_16, op_18, op_2, op_5, op_8, ap_clk, unsafe_signal);
input ap_start;
input [1:0] op_0;
input [3:0] op_1;
input [1:0] op_12;
input op_14;
input [3:0] op_16;
input [3:0] op_18;
input [7:0] op_2;
input [3:0] op_5;
input [3:0] op_8;
input ap_clk;
output unsafe_signal;
reg _setup;
initial _setup = 1'b0;
always @ (posedge ap_clk) _setup <= 1'b1;
reg ap_start_internal;
always @ (posedge ap_clk) if (!_setup) ap_start_internal <= ap_start;
reg [1:0] op_0_internal;
always @ (posedge ap_clk) if (!_setup) op_0_internal <= op_0;
reg [3:0] op_1_internal;
always @ (posedge ap_clk) if (!_setup) op_1_internal <= op_1;
reg [1:0] op_12_internal;
always @ (posedge ap_clk) if (!_setup) op_12_internal <= op_12;
reg op_14_internal;
always @ (posedge ap_clk) if (!_setup) op_14_internal <= op_14;
reg [3:0] op_16_internal;
always @ (posedge ap_clk) if (!_setup) op_16_internal <= op_16;
reg [3:0] op_18_internal;
always @ (posedge ap_clk) if (!_setup) op_18_internal <= op_18;
reg [7:0] op_2_internal;
always @ (posedge ap_clk) if (!_setup) op_2_internal <= op_2;
reg [3:0] op_5_internal;
always @ (posedge ap_clk) if (!_setup) op_5_internal <= op_5;
reg [3:0] op_8_internal;
always @ (posedge ap_clk) if (!_setup) op_8_internal <= op_8;
wire ap_done_A;
wire ap_done_B;
wire ap_done_eq;
assign ap_done_eq = ap_done_A == ap_done_B;
wire ap_idle_A;
wire ap_idle_B;
wire ap_idle_eq;
assign ap_idle_eq = ap_idle_A == ap_idle_B;
wire ap_ready_A;
wire ap_ready_B;
wire ap_ready_eq;
assign ap_ready_eq = ap_ready_A == ap_ready_B;
wire [31:0] op_30_A;
wire [31:0] op_30_B;
wire op_30_eq;
assign op_30_eq = op_30_A == op_30_B;
wire op_30_ap_vld_A;
wire op_30_ap_vld_B;
wire clk_enable_A;
wire clk_enable_B;
assign clk_enable_A = _setup & (~op_30_ap_vld_A | op_30_ap_vld_B);
assign clk_enable_B = _setup;
wire divergent;
assign divergent = ~(ap_done_eq & ap_idle_eq & ap_ready_eq & op_30_eq);
assign unsafe_signal = op_30_ap_vld_A & op_30_ap_vld_B & divergent;
top_A instance_A (
    .ap_clk(ap_clk),
    .clk_enable(clk_enable_A),
    .ap_start(ap_start_internal),
    .op_0(op_0_internal),
    .op_1(op_1_internal),
    .op_12(op_12_internal),
    .op_14(op_14_internal),
    .op_16(op_16_internal),
    .op_18(op_18_internal),
    .op_2(op_2_internal),
    .op_5(op_5_internal),
    .op_8(op_8_internal),
    .ap_done(ap_done_A),
    .ap_idle(ap_idle_A),
    .ap_ready(ap_ready_A),
    .op_30(op_30_A),
    .op_30_ap_vld(op_30_ap_vld_A)
);
top_B instance_B (
    .ap_clk(ap_clk),
    .clk_enable(clk_enable_B),
    .ap_start(ap_start_internal),
    .op_0(op_0_internal),
    .op_1(op_1_internal),
    .op_12(op_12_internal),
    .op_14(op_14_internal),
    .op_16(op_16_internal),
    .op_18(op_18_internal),
    .op_2(op_2_internal),
    .op_5(op_5_internal),
    .op_8(op_8_internal),
    .ap_done(ap_done_B),
    .ap_idle(ap_idle_B),
    .ap_ready(ap_ready_B),
    .op_30(op_30_B),
    .op_30_ap_vld(op_30_ap_vld_B)
);
endmodule
