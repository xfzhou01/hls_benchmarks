// Processed by function `construct_kairos` in `verilog_tricks.py`.
// Machine A:
// Processed by function `add_clk_enable_signal` in `verilog_tricks.py`.
// Processed by function `remove_reset_signal` in `verilog_tricks.py`.
module top_A (
  ap_clk,
  ap_start,
  ap_done,
  ap_idle,
  ap_ready,
  op_0,
  op_5,
  op_7,
  op_9,
  op_10,
  op_11,
  op_12,
  op_13,
  op_14,
  op_18,
  op_30,
  op_30_ap_vld,
clk_enable
);
input clk_enable;


input ap_clk;
wire ap_rst;
assign ap_rst = op_30_ap_vld;
input ap_start;
input [1:0] op_0;
input [15:0] op_10;
input [1:0] op_11;
input [7:0] op_12;
input [3:0] op_13;
input [1:0] op_14;
input [3:0] op_18;
input [1:0] op_5;
input [7:0] op_7;
input [15:0] op_9;
output ap_done;
output ap_idle;
output ap_ready;
output [31:0] op_30;
output op_30_ap_vld;


reg [8:0] \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.ain_s1 ;
reg [8:0] \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.bin_s1 ;
reg \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.carry_s1 ;
reg [7:0] \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.sum_s1 ;
reg [8:0] \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.ain_s1 ;
reg [8:0] \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.bin_s1 ;
reg \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.carry_s1 ;
reg [8:0] \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.sum_s1 ;
reg [9:0] \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.ain_s1 ;
reg [9:0] \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.bin_s1 ;
reg \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.carry_s1 ;
reg [8:0] \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.sum_s1 ;
reg [9:0] \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.ain_s1 ;
reg [9:0] \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.bin_s1 ;
reg \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.carry_s1 ;
reg [8:0] \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.sum_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.ain_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.bin_s1 ;
reg \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.carry_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.sum_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.ain_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.bin_s1 ;
reg \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.carry_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.sum_s1 ;
reg [16:0] \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.ain_s1 ;
reg [16:0] \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.bin_s1 ;
reg \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.carry_s1 ;
reg [16:0] \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.sum_s1 ;
reg [2:0] \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.ain_s1 ;
reg [2:0] \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.bin_s1 ;
reg \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.carry_s1 ;
reg [1:0] \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.sum_s1 ;
reg [2:0] \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.ain_s1 ;
reg [2:0] \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.bin_s1 ;
reg \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.carry_s1 ;
reg [1:0] \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.sum_s1 ;
reg [2:0] \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.ain_s1 ;
reg [2:0] \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.bin_s1 ;
reg \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.carry_s1 ;
reg [1:0] \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.sum_s1 ;
reg [2:0] \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.ain_s1 ;
reg [2:0] \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.bin_s1 ;
reg \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.carry_s1 ;
reg [2:0] \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.sum_s1 ;
reg [4:0] \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.ain_s1 ;
reg [4:0] \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.bin_s1 ;
reg \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.carry_s1 ;
reg [3:0] \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.sum_s1 ;
reg [18:0] add_ln691_reg_533;
reg [4:0] add_ln69_1_reg_451;
reg [5:0] add_ln69_2_reg_481;
reg [31:0] add_ln69_4_reg_573;
reg [4:0] add_ln69_6_reg_578;
reg [16:0] add_ln69_reg_476;
reg [19:0] ap_CS_fsm = 20'h00001;
reg icmp_ln1495_reg_548;
reg icmp_ln851_reg_431;
reg [17:0] op_24_V_reg_496;
reg [31:0] op_26_V_reg_553;
reg [4:0] ret_V_2_reg_436;
reg [8:0] ret_V_6_reg_414;
reg [4:0] ret_V_7_reg_446;
reg [18:0] ret_V_8_reg_516;
reg [4:0] ret_V_reg_419;
reg [18:0] select_ln353_reg_538;
reg [31:0] select_ln69_reg_558;
reg [18:0] sext_ln850_reg_526;
reg [17:0] tmp_reg_521;
reg [3:0] trunc_ln851_reg_426;
wire [18:0] _000_;
wire [4:0] _001_;
wire [5:0] _002_;
wire [31:0] _003_;
wire [4:0] _004_;
wire [16:0] _005_;
wire [19:0] _006_;
wire _007_;
wire _008_;
wire [17:0] _009_;
wire [31:0] _010_;
wire [4:0] _011_;
wire [8:0] _012_;
wire [4:0] _013_;
wire [18:0] _014_;
wire [4:0] _015_;
wire [18:0] _016_;
wire [31:0] _017_;
wire [18:0] _018_;
wire [17:0] _019_;
wire [3:0] _020_;
wire [1:0] _021_;
wire _022_;
wire _023_;
wire _024_;
wire _025_;
wire [8:0] _026_;
wire [8:0] _027_;
wire _028_;
wire [7:0] _029_;
wire [8:0] _030_;
wire [9:0] _031_;
wire [8:0] _032_;
wire [8:0] _033_;
wire _034_;
wire [8:0] _035_;
wire [9:0] _036_;
wire [9:0] _037_;
wire [9:0] _038_;
wire [9:0] _039_;
wire _040_;
wire [8:0] _041_;
wire [9:0] _042_;
wire [10:0] _043_;
wire [9:0] _044_;
wire [9:0] _045_;
wire _046_;
wire [8:0] _047_;
wire [9:0] _048_;
wire [10:0] _049_;
wire [15:0] _050_;
wire [15:0] _051_;
wire _052_;
wire [15:0] _053_;
wire [16:0] _054_;
wire [16:0] _055_;
wire [15:0] _056_;
wire [15:0] _057_;
wire _058_;
wire [15:0] _059_;
wire [16:0] _060_;
wire [16:0] _061_;
wire [16:0] _062_;
wire [16:0] _063_;
wire _064_;
wire [16:0] _065_;
wire [17:0] _066_;
wire [17:0] _067_;
wire [2:0] _068_;
wire [2:0] _069_;
wire _070_;
wire [1:0] _071_;
wire [2:0] _072_;
wire [3:0] _073_;
wire [2:0] _074_;
wire [2:0] _075_;
wire _076_;
wire [1:0] _077_;
wire [2:0] _078_;
wire [3:0] _079_;
wire [2:0] _080_;
wire [2:0] _081_;
wire _082_;
wire [1:0] _083_;
wire [2:0] _084_;
wire [3:0] _085_;
wire [2:0] _086_;
wire [2:0] _087_;
wire _088_;
wire [2:0] _089_;
wire [3:0] _090_;
wire [3:0] _091_;
wire [4:0] _092_;
wire [4:0] _093_;
wire _094_;
wire [3:0] _095_;
wire [4:0] _096_;
wire [5:0] _097_;
wire _098_;
wire _099_;
wire _100_;
wire _101_;
wire _102_;
wire _103_;
wire _104_;
wire _105_;
wire _106_;
wire _107_;
wire _108_;
wire _109_;
wire _110_;
wire _111_;
wire _112_;
wire _113_;
wire _114_;
wire _115_;
wire _116_;
wire _117_;
wire _118_;
wire \add_17s_17s_17_2_1_U4.ce ;
wire \add_17s_17s_17_2_1_U4.clk ;
wire [16:0] \add_17s_17s_17_2_1_U4.din0 ;
wire [16:0] \add_17s_17s_17_2_1_U4.din1 ;
wire [16:0] \add_17s_17s_17_2_1_U4.dout ;
wire \add_17s_17s_17_2_1_U4.reset ;
wire [16:0] \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.a ;
wire [16:0] \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.ain_s0 ;
wire [16:0] \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.b ;
wire [16:0] \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.bin_s0 ;
wire \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.ce ;
wire \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.clk ;
wire \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.facout_s1 ;
wire \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.facout_s2 ;
wire [7:0] \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.fas_s1 ;
wire [8:0] \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.fas_s2 ;
wire \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.reset ;
wire [16:0] \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.s ;
wire [7:0] \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.u1.a ;
wire [7:0] \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.u1.b ;
wire \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.u1.cin ;
wire \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.u1.cout ;
wire [7:0] \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.u1.s ;
wire [8:0] \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.u2.a ;
wire [8:0] \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.u2.b ;
wire \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.u2.cin ;
wire \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.u2.cout ;
wire [8:0] \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.u2.s ;
wire \add_18s_18s_18_2_1_U6.ce ;
wire \add_18s_18s_18_2_1_U6.clk ;
wire [17:0] \add_18s_18s_18_2_1_U6.din0 ;
wire [17:0] \add_18s_18s_18_2_1_U6.din1 ;
wire [17:0] \add_18s_18s_18_2_1_U6.dout ;
wire \add_18s_18s_18_2_1_U6.reset ;
wire [17:0] \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.a ;
wire [17:0] \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.ain_s0 ;
wire [17:0] \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.b ;
wire [17:0] \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.bin_s0 ;
wire \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.ce ;
wire \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.clk ;
wire \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.facout_s1 ;
wire \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.facout_s2 ;
wire [8:0] \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.fas_s1 ;
wire [8:0] \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.fas_s2 ;
wire \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.reset ;
wire [17:0] \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.s ;
wire [8:0] \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.u1.a ;
wire [8:0] \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.u1.b ;
wire \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.u1.cin ;
wire \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.u1.cout ;
wire [8:0] \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.u1.s ;
wire [8:0] \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.u2.a ;
wire [8:0] \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.u2.b ;
wire \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.u2.cin ;
wire \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.u2.cout ;
wire [8:0] \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.u2.s ;
wire \add_19ns_19s_19_2_1_U7.ce ;
wire \add_19ns_19s_19_2_1_U7.clk ;
wire [18:0] \add_19ns_19s_19_2_1_U7.din0 ;
wire [18:0] \add_19ns_19s_19_2_1_U7.din1 ;
wire [18:0] \add_19ns_19s_19_2_1_U7.dout ;
wire \add_19ns_19s_19_2_1_U7.reset ;
wire [18:0] \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.a ;
wire [18:0] \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.ain_s0 ;
wire [18:0] \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.b ;
wire [18:0] \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.bin_s0 ;
wire \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.ce ;
wire \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.clk ;
wire \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.facout_s1 ;
wire \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.facout_s2 ;
wire [8:0] \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.fas_s1 ;
wire [9:0] \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.fas_s2 ;
wire \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.reset ;
wire [18:0] \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.s ;
wire [8:0] \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.u1.a ;
wire [8:0] \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.u1.b ;
wire \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.u1.cin ;
wire \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.u1.cout ;
wire [8:0] \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.u1.s ;
wire [9:0] \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.u2.a ;
wire [9:0] \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.u2.b ;
wire \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.u2.cin ;
wire \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.u2.cout ;
wire [9:0] \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.u2.s ;
wire \add_19s_19ns_19_2_1_U8.ce ;
wire \add_19s_19ns_19_2_1_U8.clk ;
wire [18:0] \add_19s_19ns_19_2_1_U8.din0 ;
wire [18:0] \add_19s_19ns_19_2_1_U8.din1 ;
wire [18:0] \add_19s_19ns_19_2_1_U8.dout ;
wire \add_19s_19ns_19_2_1_U8.reset ;
wire [18:0] \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.a ;
wire [18:0] \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.ain_s0 ;
wire [18:0] \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.b ;
wire [18:0] \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.bin_s0 ;
wire \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.ce ;
wire \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.clk ;
wire \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.facout_s1 ;
wire \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.facout_s2 ;
wire [8:0] \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.fas_s1 ;
wire [9:0] \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.fas_s2 ;
wire \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.reset ;
wire [18:0] \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.s ;
wire [8:0] \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.u1.a ;
wire [8:0] \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.u1.b ;
wire \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.u1.cin ;
wire \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.u1.cout ;
wire [8:0] \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.u1.s ;
wire [9:0] \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.u2.a ;
wire [9:0] \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.u2.b ;
wire \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.u2.cin ;
wire \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.u2.cout ;
wire [9:0] \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.u2.s ;
wire \add_32ns_32ns_32_2_1_U10.ce ;
wire \add_32ns_32ns_32_2_1_U10.clk ;
wire [31:0] \add_32ns_32ns_32_2_1_U10.din0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U10.din1 ;
wire [31:0] \add_32ns_32ns_32_2_1_U10.dout ;
wire \add_32ns_32ns_32_2_1_U10.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.a ;
wire [31:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.ain_s0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.b ;
wire [31:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.bin_s0 ;
wire \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.ce ;
wire \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.clk ;
wire \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.facout_s1 ;
wire \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.facout_s2 ;
wire [15:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.fas_s1 ;
wire [15:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.fas_s2 ;
wire \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.u1.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.u1.b ;
wire \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.u1.cin ;
wire \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.u1.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.u1.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.u2.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.u2.b ;
wire \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.u2.cin ;
wire \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.u2.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.u2.s ;
wire \add_32ns_32ns_32_2_1_U12.ce ;
wire \add_32ns_32ns_32_2_1_U12.clk ;
wire [31:0] \add_32ns_32ns_32_2_1_U12.din0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U12.din1 ;
wire [31:0] \add_32ns_32ns_32_2_1_U12.dout ;
wire \add_32ns_32ns_32_2_1_U12.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.a ;
wire [31:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.ain_s0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.b ;
wire [31:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.bin_s0 ;
wire \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.ce ;
wire \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.clk ;
wire \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.facout_s1 ;
wire \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.facout_s2 ;
wire [15:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.fas_s1 ;
wire [15:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.fas_s2 ;
wire \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.u1.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.u1.b ;
wire \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.u1.cin ;
wire \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.u1.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.u1.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.u2.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.u2.b ;
wire \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.u2.cin ;
wire \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.u2.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.u2.s ;
wire \add_34s_34ns_34_2_1_U9.ce ;
wire \add_34s_34ns_34_2_1_U9.clk ;
wire [33:0] \add_34s_34ns_34_2_1_U9.din0 ;
wire [33:0] \add_34s_34ns_34_2_1_U9.din1 ;
wire [33:0] \add_34s_34ns_34_2_1_U9.dout ;
wire \add_34s_34ns_34_2_1_U9.reset ;
wire [33:0] \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.a ;
wire [33:0] \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.ain_s0 ;
wire [33:0] \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.b ;
wire [33:0] \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.bin_s0 ;
wire \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.ce ;
wire \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.clk ;
wire \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.facout_s1 ;
wire \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.facout_s2 ;
wire [16:0] \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.fas_s1 ;
wire [16:0] \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.fas_s2 ;
wire \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.reset ;
wire [33:0] \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.s ;
wire [16:0] \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.u1.a ;
wire [16:0] \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.u1.b ;
wire \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.u1.cin ;
wire \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.u1.cout ;
wire [16:0] \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.u1.s ;
wire [16:0] \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.u2.a ;
wire [16:0] \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.u2.b ;
wire \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.u2.cin ;
wire \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.u2.cout ;
wire [16:0] \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.u2.s ;
wire \add_5ns_5ns_5_2_1_U11.ce ;
wire \add_5ns_5ns_5_2_1_U11.clk ;
wire [4:0] \add_5ns_5ns_5_2_1_U11.din0 ;
wire [4:0] \add_5ns_5ns_5_2_1_U11.din1 ;
wire [4:0] \add_5ns_5ns_5_2_1_U11.dout ;
wire \add_5ns_5ns_5_2_1_U11.reset ;
wire [4:0] \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.a ;
wire [4:0] \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.ain_s0 ;
wire [4:0] \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.b ;
wire [4:0] \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.bin_s0 ;
wire \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.ce ;
wire \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.clk ;
wire \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.facout_s1 ;
wire \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.facout_s2 ;
wire [1:0] \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.fas_s1 ;
wire [2:0] \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.fas_s2 ;
wire \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.reset ;
wire [4:0] \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.s ;
wire [1:0] \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.u1.a ;
wire [1:0] \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.u1.b ;
wire \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.u1.cin ;
wire \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.u1.cout ;
wire [1:0] \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.u1.s ;
wire [2:0] \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.u2.a ;
wire [2:0] \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.u2.b ;
wire \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.u2.cin ;
wire \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.u2.cout ;
wire [2:0] \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.u2.s ;
wire \add_5ns_5ns_5_2_1_U2.ce ;
wire \add_5ns_5ns_5_2_1_U2.clk ;
wire [4:0] \add_5ns_5ns_5_2_1_U2.din0 ;
wire [4:0] \add_5ns_5ns_5_2_1_U2.din1 ;
wire [4:0] \add_5ns_5ns_5_2_1_U2.dout ;
wire \add_5ns_5ns_5_2_1_U2.reset ;
wire [4:0] \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.a ;
wire [4:0] \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.ain_s0 ;
wire [4:0] \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.b ;
wire [4:0] \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.bin_s0 ;
wire \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.ce ;
wire \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.clk ;
wire \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.facout_s1 ;
wire \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.facout_s2 ;
wire [1:0] \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.fas_s1 ;
wire [2:0] \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.fas_s2 ;
wire \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.reset ;
wire [4:0] \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.s ;
wire [1:0] \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.u1.a ;
wire [1:0] \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.u1.b ;
wire \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.u1.cin ;
wire \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.u1.cout ;
wire [1:0] \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.u1.s ;
wire [2:0] \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.u2.a ;
wire [2:0] \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.u2.b ;
wire \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.u2.cin ;
wire \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.u2.cout ;
wire [2:0] \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.u2.s ;
wire \add_5s_5ns_5_2_1_U3.ce ;
wire \add_5s_5ns_5_2_1_U3.clk ;
wire [4:0] \add_5s_5ns_5_2_1_U3.din0 ;
wire [4:0] \add_5s_5ns_5_2_1_U3.din1 ;
wire [4:0] \add_5s_5ns_5_2_1_U3.dout ;
wire \add_5s_5ns_5_2_1_U3.reset ;
wire [4:0] \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.a ;
wire [4:0] \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.ain_s0 ;
wire [4:0] \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.b ;
wire [4:0] \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.bin_s0 ;
wire \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.ce ;
wire \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.clk ;
wire \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.facout_s1 ;
wire \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.facout_s2 ;
wire [1:0] \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.fas_s1 ;
wire [2:0] \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.fas_s2 ;
wire \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.reset ;
wire [4:0] \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.s ;
wire [1:0] \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.u1.a ;
wire [1:0] \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.u1.b ;
wire \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.u1.cin ;
wire \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.u1.cout ;
wire [1:0] \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.u1.s ;
wire [2:0] \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.u2.a ;
wire [2:0] \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.u2.b ;
wire \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.u2.cin ;
wire \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.u2.cout ;
wire [2:0] \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.u2.s ;
wire \add_6s_6s_6_2_1_U5.ce ;
wire \add_6s_6s_6_2_1_U5.clk ;
wire [5:0] \add_6s_6s_6_2_1_U5.din0 ;
wire [5:0] \add_6s_6s_6_2_1_U5.din1 ;
wire [5:0] \add_6s_6s_6_2_1_U5.dout ;
wire \add_6s_6s_6_2_1_U5.reset ;
wire [5:0] \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.a ;
wire [5:0] \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.ain_s0 ;
wire [5:0] \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.b ;
wire [5:0] \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.bin_s0 ;
wire \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.ce ;
wire \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.clk ;
wire \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.facout_s1 ;
wire \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.facout_s2 ;
wire [2:0] \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.fas_s1 ;
wire [2:0] \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.fas_s2 ;
wire \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.reset ;
wire [5:0] \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.s ;
wire [2:0] \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.u1.a ;
wire [2:0] \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.u1.b ;
wire \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.u1.cin ;
wire \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.u1.cout ;
wire [2:0] \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.u1.s ;
wire [2:0] \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.u2.a ;
wire [2:0] \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.u2.b ;
wire \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.u2.cin ;
wire \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.u2.cout ;
wire [2:0] \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.u2.s ;
wire \add_9s_9s_9_2_1_U1.ce ;
wire \add_9s_9s_9_2_1_U1.clk ;
wire [8:0] \add_9s_9s_9_2_1_U1.din0 ;
wire [8:0] \add_9s_9s_9_2_1_U1.din1 ;
wire [8:0] \add_9s_9s_9_2_1_U1.dout ;
wire \add_9s_9s_9_2_1_U1.reset ;
wire [8:0] \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.a ;
wire [8:0] \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.ain_s0 ;
wire [8:0] \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.b ;
wire [8:0] \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.bin_s0 ;
wire \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.ce ;
wire \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.clk ;
wire \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.facout_s1 ;
wire \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.facout_s2 ;
wire [3:0] \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.fas_s1 ;
wire [4:0] \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.fas_s2 ;
wire \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.reset ;
wire [8:0] \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.s ;
wire [3:0] \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.u1.a ;
wire [3:0] \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.u1.b ;
wire \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.u1.cin ;
wire \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.u1.cout ;
wire [3:0] \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.u1.s ;
wire [4:0] \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.u2.a ;
wire [4:0] \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.u2.b ;
wire \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.u2.cin ;
wire \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.u2.cout ;
wire [4:0] \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.u2.s ;
wire ap_CS_fsm_state1;
wire ap_CS_fsm_state10;
wire ap_CS_fsm_state11;
wire ap_CS_fsm_state12;
wire ap_CS_fsm_state13;
wire ap_CS_fsm_state14;
wire ap_CS_fsm_state15;
wire ap_CS_fsm_state16;
wire ap_CS_fsm_state17;
wire ap_CS_fsm_state18;
wire ap_CS_fsm_state19;
wire ap_CS_fsm_state2;
wire ap_CS_fsm_state20;
wire ap_CS_fsm_state3;
wire ap_CS_fsm_state4;
wire ap_CS_fsm_state5;
wire ap_CS_fsm_state6;
wire ap_CS_fsm_state7;
wire ap_CS_fsm_state8;
wire ap_CS_fsm_state9;
wire [19:0] ap_NS_fsm;
wire ap_clk;
wire ap_done;
wire ap_idle;
wire ap_ready;
wire ap_rst;
wire ap_start;
wire [8:0] grp_fu_171_p0;
wire [8:0] grp_fu_171_p1;
wire [8:0] grp_fu_171_p2;
wire [4:0] grp_fu_196_p2;
wire [4:0] grp_fu_205_p0;
wire [4:0] grp_fu_205_p2;
wire [16:0] grp_fu_241_p0;
wire [16:0] grp_fu_241_p1;
wire [16:0] grp_fu_241_p2;
wire [5:0] grp_fu_250_p0;
wire [5:0] grp_fu_250_p1;
wire [5:0] grp_fu_250_p2;
wire [17:0] grp_fu_262_p0;
wire [17:0] grp_fu_262_p1;
wire [17:0] grp_fu_262_p2;
wire [18:0] grp_fu_279_p0;
wire [18:0] grp_fu_279_p1;
wire [18:0] grp_fu_279_p2;
wire [18:0] grp_fu_298_p0;
wire [18:0] grp_fu_298_p2;
wire [33:0] grp_fu_338_p0;
wire [33:0] grp_fu_338_p2;
wire [31:0] grp_fu_385_p2;
wire [4:0] grp_fu_389_p0;
wire [4:0] grp_fu_389_p1;
wire [4:0] grp_fu_389_p2;
wire [31:0] grp_fu_398_p0;
wire [31:0] grp_fu_398_p2;
wire icmp_ln1495_fu_348_p2;
wire icmp_ln851_fu_191_p2;
wire [4:0] lhs_fu_155_p3;
wire [1:0] op_0;
wire [15:0] op_10;
wire [1:0] op_11;
wire [7:0] op_12;
wire [3:0] op_13;
wire [1:0] op_14;
wire op_17_V_fu_344_p1;
wire [3:0] op_18;
wire [31:0] op_30;
wire op_30_ap_vld;
wire [1:0] op_5;
wire [7:0] op_7;
wire [15:0] op_9;
wire p_Result_1_fu_304_p3;
wire p_Result_s_fu_211_p3;
wire [4:0] ret_V_7_fu_223_p3;
wire [18:0] select_ln353_fu_320_p3;
wire [31:0] select_ln69_fu_370_p3;
wire [18:0] select_ln850_2_fu_314_p3;
wire [4:0] select_ln850_fu_218_p3;
wire [1:0] sext_ln1192_1_fu_268_p0;
wire [18:0] sext_ln850_fu_295_p1;
wire [20:0] tmp_3_fu_327_p3;
wire [1:0] trunc_ln851_1_fu_311_p0;
wire trunc_ln851_1_fu_311_p1;
wire [3:0] trunc_ln851_fu_187_p1;


assign _022_ = _024_ & ap_CS_fsm[0];
assign _023_ = ap_start & ap_CS_fsm[0];
assign _024_ = ~ ap_start;
assign _025_ = ! trunc_ln851_reg_426;
always @(posedge \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.clk )
\add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.bin_s1  <= _027_;
always @(posedge \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.clk )
\add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.ain_s1  <= _026_;
always @(posedge \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.clk )
\add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.sum_s1  <= _029_;
always @(posedge \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.clk )
\add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.carry_s1  <= _028_;
assign _027_ = \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.ce  ? \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.b [16:8] : \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.bin_s1 ;
assign _026_ = \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.ce  ? \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.a [16:8] : \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.ain_s1 ;
assign _028_ = \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.ce  ? \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.facout_s1  : \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.carry_s1 ;
assign _029_ = \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.ce  ? \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.fas_s1  : \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.sum_s1 ;
assign _030_ = \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.u1.a  + \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.u1.b ;
assign { \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.u1.cout , \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.u1.s  } = _030_ + \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.u1.cin ;
assign _031_ = \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.u2.a  + \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.u2.b ;
assign { \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.u2.cout , \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.u2.s  } = _031_ + \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.u2.cin ;
always @(posedge \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.clk )
\add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.bin_s1  <= _033_;
always @(posedge \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.clk )
\add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.ain_s1  <= _032_;
always @(posedge \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.clk )
\add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.sum_s1  <= _035_;
always @(posedge \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.clk )
\add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.carry_s1  <= _034_;
assign _033_ = \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.ce  ? \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.b [17:9] : \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.bin_s1 ;
assign _032_ = \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.ce  ? \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.a [17:9] : \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.ain_s1 ;
assign _034_ = \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.ce  ? \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.facout_s1  : \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.carry_s1 ;
assign _035_ = \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.ce  ? \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.fas_s1  : \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.sum_s1 ;
assign _036_ = \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.u1.a  + \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.u1.b ;
assign { \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.u1.cout , \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.u1.s  } = _036_ + \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.u1.cin ;
assign _037_ = \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.u2.a  + \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.u2.b ;
assign { \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.u2.cout , \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.u2.s  } = _037_ + \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.u2.cin ;
always @(posedge \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.clk )
\add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.bin_s1  <= _039_;
always @(posedge \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.clk )
\add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.ain_s1  <= _038_;
always @(posedge \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.clk )
\add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.sum_s1  <= _041_;
always @(posedge \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.clk )
\add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.carry_s1  <= _040_;
assign _039_ = \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.ce  ? \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.b [18:9] : \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.bin_s1 ;
assign _038_ = \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.ce  ? \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.a [18:9] : \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.ain_s1 ;
assign _040_ = \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.ce  ? \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.facout_s1  : \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.carry_s1 ;
assign _041_ = \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.ce  ? \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.fas_s1  : \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.sum_s1 ;
assign _042_ = \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.u1.a  + \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.u1.b ;
assign { \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.u1.cout , \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.u1.s  } = _042_ + \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.u1.cin ;
assign { \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.u2.cout , \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.u2.s  } = _043_ + \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.u2.cin ;
assign _043_ = \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.u2.a  + \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.u2.b ;
always @(posedge \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.clk )
\add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.bin_s1  <= _045_;
always @(posedge \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.clk )
\add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.ain_s1  <= _044_;
always @(posedge \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.clk )
\add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.sum_s1  <= _047_;
always @(posedge \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.clk )
\add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.carry_s1  <= _046_;
assign _045_ = \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.ce  ? \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.b [18:9] : \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.bin_s1 ;
assign _044_ = \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.ce  ? \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.a [18:9] : \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.ain_s1 ;
assign _046_ = \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.ce  ? \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.facout_s1  : \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.carry_s1 ;
assign _047_ = \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.ce  ? \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.fas_s1  : \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.sum_s1 ;
assign _048_ = \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.u1.a  + \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.u1.b ;
assign { \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.u1.cout , \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.u1.s  } = _048_ + \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.u1.cin ;
assign _049_ = \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.u2.a  + \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.u2.b ;
assign { \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.u2.cout , \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.u2.s  } = _049_ + \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.u2.cin ;
always @(posedge \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.clk )
\add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.bin_s1  <= _051_;
always @(posedge \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.clk )
\add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.ain_s1  <= _050_;
always @(posedge \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.clk )
\add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.sum_s1  <= _053_;
always @(posedge \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.clk )
\add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.carry_s1  <= _052_;
assign _051_ = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.ce  ? \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.b [31:16] : \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.bin_s1 ;
assign _050_ = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.ce  ? \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.a [31:16] : \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.ain_s1 ;
assign _052_ = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.ce  ? \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.facout_s1  : \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.carry_s1 ;
assign _053_ = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.ce  ? \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.fas_s1  : \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.sum_s1 ;
assign _054_ = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.u1.a  + \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.u1.b ;
assign { \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.u1.cout , \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.u1.s  } = _054_ + \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.u1.cin ;
assign _055_ = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.u2.a  + \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.u2.b ;
assign { \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.u2.cout , \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.u2.s  } = _055_ + \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.u2.cin ;
always @(posedge \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.clk )
\add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.bin_s1  <= _057_;
always @(posedge \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.clk )
\add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.ain_s1  <= _056_;
always @(posedge \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.clk )
\add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.sum_s1  <= _059_;
always @(posedge \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.clk )
\add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.carry_s1  <= _058_;
assign _057_ = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.ce  ? \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.b [31:16] : \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.bin_s1 ;
assign _056_ = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.ce  ? \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.a [31:16] : \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.ain_s1 ;
assign _058_ = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.ce  ? \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.facout_s1  : \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.carry_s1 ;
assign _059_ = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.ce  ? \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.fas_s1  : \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.sum_s1 ;
assign _060_ = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.u1.a  + \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.u1.b ;
assign { \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.u1.cout , \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.u1.s  } = _060_ + \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.u1.cin ;
assign _061_ = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.u2.a  + \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.u2.b ;
assign { \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.u2.cout , \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.u2.s  } = _061_ + \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.u2.cin ;
always @(posedge \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.clk )
\add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.bin_s1  <= _063_;
always @(posedge \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.clk )
\add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.ain_s1  <= _062_;
always @(posedge \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.clk )
\add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.sum_s1  <= _065_;
always @(posedge \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.clk )
\add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.carry_s1  <= _064_;
assign _063_ = \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.ce  ? \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.b [33:17] : \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.bin_s1 ;
assign _062_ = \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.ce  ? \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.a [33:17] : \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.ain_s1 ;
assign _064_ = \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.ce  ? \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.facout_s1  : \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.carry_s1 ;
assign _065_ = \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.ce  ? \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.fas_s1  : \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.sum_s1 ;
assign _066_ = \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.u1.a  + \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.u1.b ;
assign { \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.u1.cout , \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.u1.s  } = _066_ + \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.u1.cin ;
assign _067_ = \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.u2.a  + \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.u2.b ;
assign { \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.u2.cout , \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.u2.s  } = _067_ + \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.u2.cin ;
always @(posedge \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.clk )
\add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.bin_s1  <= _069_;
always @(posedge \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.clk )
\add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.ain_s1  <= _068_;
always @(posedge \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.clk )
\add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.sum_s1  <= _071_;
always @(posedge \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.clk )
\add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.carry_s1  <= _070_;
assign _069_ = \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.ce  ? \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.b [4:2] : \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.bin_s1 ;
assign _068_ = \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.ce  ? \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.a [4:2] : \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.ain_s1 ;
assign _070_ = \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.ce  ? \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.facout_s1  : \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.carry_s1 ;
assign _071_ = \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.ce  ? \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.fas_s1  : \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.sum_s1 ;
assign _072_ = \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.u1.a  + \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.u1.b ;
assign { \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.u1.cout , \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.u1.s  } = _072_ + \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.u1.cin ;
assign _073_ = \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.u2.a  + \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.u2.b ;
assign { \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.u2.cout , \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.u2.s  } = _073_ + \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.u2.cin ;
always @(posedge \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.clk )
\add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.bin_s1  <= _075_;
always @(posedge \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.clk )
\add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.ain_s1  <= _074_;
always @(posedge \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.clk )
\add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.sum_s1  <= _077_;
always @(posedge \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.clk )
\add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.carry_s1  <= _076_;
assign _075_ = \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.ce  ? \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.b [4:2] : \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.bin_s1 ;
assign _074_ = \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.ce  ? \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.a [4:2] : \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.ain_s1 ;
assign _076_ = \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.ce  ? \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.facout_s1  : \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.carry_s1 ;
assign _077_ = \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.ce  ? \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.fas_s1  : \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.sum_s1 ;
assign _078_ = \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.u1.a  + \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.u1.b ;
assign { \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.u1.cout , \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.u1.s  } = _078_ + \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.u1.cin ;
assign _079_ = \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.u2.a  + \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.u2.b ;
assign { \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.u2.cout , \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.u2.s  } = _079_ + \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.u2.cin ;
always @(posedge \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.clk )
\add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.bin_s1  <= _081_;
always @(posedge \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.clk )
\add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.ain_s1  <= _080_;
always @(posedge \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.clk )
\add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.sum_s1  <= _083_;
always @(posedge \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.clk )
\add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.carry_s1  <= _082_;
assign _081_ = \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.ce  ? \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.b [4:2] : \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.bin_s1 ;
assign _080_ = \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.ce  ? \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.a [4:2] : \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.ain_s1 ;
assign _082_ = \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.ce  ? \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.facout_s1  : \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.carry_s1 ;
assign _083_ = \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.ce  ? \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.fas_s1  : \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.sum_s1 ;
assign _084_ = \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.u1.a  + \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.u1.b ;
assign { \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.u1.cout , \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.u1.s  } = _084_ + \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.u1.cin ;
assign _085_ = \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.u2.a  + \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.u2.b ;
assign { \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.u2.cout , \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.u2.s  } = _085_ + \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.u2.cin ;
always @(posedge \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.clk )
\add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.bin_s1  <= _087_;
always @(posedge \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.clk )
\add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.ain_s1  <= _086_;
always @(posedge \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.clk )
\add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.sum_s1  <= _089_;
always @(posedge \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.clk )
\add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.carry_s1  <= _088_;
assign _087_ = \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.ce  ? \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.b [5:3] : \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.bin_s1 ;
assign _086_ = \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.ce  ? \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.a [5:3] : \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.ain_s1 ;
assign _088_ = \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.ce  ? \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.facout_s1  : \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.carry_s1 ;
assign _089_ = \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.ce  ? \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.fas_s1  : \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.sum_s1 ;
assign _090_ = \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.u1.a  + \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.u1.b ;
assign { \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.u1.cout , \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.u1.s  } = _090_ + \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.u1.cin ;
assign _091_ = \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.u2.a  + \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.u2.b ;
assign { \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.u2.cout , \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.u2.s  } = _091_ + \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.u2.cin ;
always @(posedge \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.clk )
\add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.bin_s1  <= _093_;
always @(posedge \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.clk )
\add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.ain_s1  <= _092_;
always @(posedge \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.clk )
\add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.sum_s1  <= _095_;
always @(posedge \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.clk )
\add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.carry_s1  <= _094_;
assign _093_ = \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.ce  ? \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.b [8:4] : \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.bin_s1 ;
assign _092_ = \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.ce  ? \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.a [8:4] : \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.ain_s1 ;
assign _094_ = \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.ce  ? \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.facout_s1  : \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.carry_s1 ;
assign _095_ = \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.ce  ? \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.fas_s1  : \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.sum_s1 ;
assign _096_ = \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.u1.a  + \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.u1.b ;
assign { \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.u1.cout , \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.u1.s  } = _096_ + \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.u1.cin ;
assign _097_ = \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.u2.a  + \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.u2.b ;
assign { \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.u2.cout , \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.u2.s  } = _097_ + \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.u2.cin ;
assign _098_ = $signed(op_12) > $signed(1'h0);
always @(posedge ap_clk)
sext_ln850_reg_526 <= _018_;
always @(posedge ap_clk)
select_ln353_reg_538 <= _016_;
always @(posedge ap_clk)
ret_V_8_reg_516 <= _014_;
always @(posedge ap_clk)
tmp_reg_521 <= _019_;
always @(posedge ap_clk)
ret_V_6_reg_414 <= _012_;
always @(posedge ap_clk)
ret_V_reg_419 <= _015_;
always @(posedge ap_clk)
trunc_ln851_reg_426 <= _020_;
always @(posedge ap_clk)
ret_V_2_reg_436 <= _011_;
always @(posedge ap_clk)
op_24_V_reg_496 <= _009_;
always @(posedge ap_clk)
icmp_ln851_reg_431 <= _008_;
always @(posedge ap_clk)
icmp_ln1495_reg_548 <= _007_;
always @(posedge ap_clk)
op_26_V_reg_553 <= _010_;
always @(posedge ap_clk)
select_ln69_reg_558 <= _017_;
always @(posedge ap_clk)
add_ln69_4_reg_573 <= _003_;
always @(posedge ap_clk)
add_ln69_6_reg_578 <= _004_;
always @(posedge ap_clk)
add_ln69_reg_476 <= _005_;
always @(posedge ap_clk)
add_ln69_2_reg_481 <= _002_;
always @(posedge ap_clk)
ret_V_7_reg_446 <= _013_;
always @(posedge ap_clk)
add_ln69_1_reg_451 <= _001_;
always @(posedge ap_clk)
add_ln691_reg_533 <= _000_;
always @(posedge ap_clk)
ap_CS_fsm <= _006_;
assign _021_ = _023_ ? 2'h2 : 2'h1;
assign _099_ = ap_CS_fsm == 1'h1;
function [19:0] _291_;
input [19:0] a;
input [399:0] b;
input [19:0] s;
case (s)
20'b00000000000000000001:
_291_ = b[19:0];
20'b00000000000000000010:
_291_ = b[39:20];
20'b00000000000000000100:
_291_ = b[59:40];
20'b00000000000000001000:
_291_ = b[79:60];
20'b00000000000000010000:
_291_ = b[99:80];
20'b00000000000000100000:
_291_ = b[119:100];
20'b00000000000001000000:
_291_ = b[139:120];
20'b00000000000010000000:
_291_ = b[159:140];
20'b00000000000100000000:
_291_ = b[179:160];
20'b00000000001000000000:
_291_ = b[199:180];
20'b00000000010000000000:
_291_ = b[219:200];
20'b00000000100000000000:
_291_ = b[239:220];
20'b00000001000000000000:
_291_ = b[259:240];
20'b00000010000000000000:
_291_ = b[279:260];
20'b00000100000000000000:
_291_ = b[299:280];
20'b00001000000000000000:
_291_ = b[319:300];
20'b00010000000000000000:
_291_ = b[339:320];
20'b00100000000000000000:
_291_ = b[359:340];
20'b01000000000000000000:
_291_ = b[379:360];
20'b10000000000000000000:
_291_ = b[399:380];
20'b00000000000000000000:
_291_ = a;
default:
_291_ = 20'bx;
endcase
endfunction
assign ap_NS_fsm = _291_(20'hxxxxx, { 18'h00000, _021_, 380'h00004000080001000020000400008000100002000040000800010000200004000080001000020000400008000000001 }, { _099_, _118_, _117_, _116_, _115_, _114_, _113_, _112_, _111_, _110_, _109_, _108_, _107_, _106_, _105_, _104_, _103_, _102_, _101_, _100_ });
assign _100_ = ap_CS_fsm == 20'h80000;
assign _101_ = ap_CS_fsm == 19'h40000;
assign _102_ = ap_CS_fsm == 18'h20000;
assign _103_ = ap_CS_fsm == 17'h10000;
assign _104_ = ap_CS_fsm == 16'h8000;
assign _105_ = ap_CS_fsm == 15'h4000;
assign _106_ = ap_CS_fsm == 14'h2000;
assign _107_ = ap_CS_fsm == 13'h1000;
assign _108_ = ap_CS_fsm == 12'h800;
assign _109_ = ap_CS_fsm == 11'h400;
assign _110_ = ap_CS_fsm == 10'h200;
assign _111_ = ap_CS_fsm == 9'h100;
assign _112_ = ap_CS_fsm == 8'h80;
assign _113_ = ap_CS_fsm == 7'h40;
assign _114_ = ap_CS_fsm == 6'h20;
assign _115_ = ap_CS_fsm == 5'h10;
assign _116_ = ap_CS_fsm == 4'h8;
assign _117_ = ap_CS_fsm == 3'h4;
assign _118_ = ap_CS_fsm == 2'h2;
assign op_30_ap_vld = ap_CS_fsm[19] ? 1'h1 : 1'h0;
assign ap_idle = _022_ ? 1'h1 : 1'h0;
assign _018_ = ap_CS_fsm[11] ? { tmp_reg_521[17], tmp_reg_521 } : sext_ln850_reg_526;
assign _016_ = ap_CS_fsm[13] ? select_ln353_fu_320_p3 : select_ln353_reg_538;
assign _019_ = ap_CS_fsm[10] ? grp_fu_279_p2[18:1] : tmp_reg_521;
assign _014_ = ap_CS_fsm[10] ? grp_fu_279_p2 : ret_V_8_reg_516;
assign _020_ = ap_CS_fsm[1] ? grp_fu_171_p2[3:0] : trunc_ln851_reg_426;
assign _015_ = ap_CS_fsm[1] ? grp_fu_171_p2[8:4] : ret_V_reg_419;
assign _012_ = ap_CS_fsm[1] ? grp_fu_171_p2 : ret_V_6_reg_414;
assign _011_ = ap_CS_fsm[3] ? grp_fu_196_p2 : ret_V_2_reg_436;
assign _009_ = ap_CS_fsm[8] ? grp_fu_262_p2 : op_24_V_reg_496;
assign _008_ = ap_CS_fsm[2] ? icmp_ln851_fu_191_p2 : icmp_ln851_reg_431;
assign _017_ = ap_CS_fsm[15] ? select_ln69_fu_370_p3 : select_ln69_reg_558;
assign _010_ = ap_CS_fsm[15] ? grp_fu_338_p2[33:2] : op_26_V_reg_553;
assign _007_ = ap_CS_fsm[15] ? icmp_ln1495_fu_348_p2 : icmp_ln1495_reg_548;
assign _004_ = ap_CS_fsm[17] ? grp_fu_389_p2 : add_ln69_6_reg_578;
assign _003_ = ap_CS_fsm[17] ? grp_fu_385_p2 : add_ln69_4_reg_573;
assign _002_ = ap_CS_fsm[6] ? grp_fu_250_p2 : add_ln69_2_reg_481;
assign _005_ = ap_CS_fsm[6] ? grp_fu_241_p2 : add_ln69_reg_476;
assign _001_ = ap_CS_fsm[4] ? grp_fu_205_p2 : add_ln69_1_reg_451;
assign _013_ = ap_CS_fsm[4] ? ret_V_7_fu_223_p3 : ret_V_7_reg_446;
assign _000_ = ap_CS_fsm[12] ? grp_fu_298_p2 : add_ln691_reg_533;
assign _006_ = ap_rst ? 20'h00001 : ap_NS_fsm;
assign icmp_ln1495_fu_348_p2 = _098_ ? 1'h1 : 1'h0;
assign icmp_ln851_fu_191_p2 = _025_ ? 1'h1 : 1'h0;
assign ret_V_7_fu_223_p3 = ret_V_6_reg_414[8] ? select_ln850_fu_218_p3 : ret_V_reg_419;
assign select_ln353_fu_320_p3 = ret_V_8_reg_516[18] ? select_ln850_2_fu_314_p3 : sext_ln850_reg_526;
assign select_ln69_fu_370_p3 = op_11[0] ? 32'd0 : 32'd4294967295;
assign select_ln850_2_fu_314_p3 = op_14[0] ? add_ln691_reg_533 : sext_ln850_reg_526;
assign select_ln850_fu_218_p3 = icmp_ln851_reg_431 ? ret_V_reg_419 : ret_V_2_reg_436;
assign ap_CS_fsm_state1 = ap_CS_fsm[0];
assign ap_CS_fsm_state10 = ap_CS_fsm[9];
assign ap_CS_fsm_state11 = ap_CS_fsm[10];
assign ap_CS_fsm_state12 = ap_CS_fsm[11];
assign ap_CS_fsm_state13 = ap_CS_fsm[12];
assign ap_CS_fsm_state14 = ap_CS_fsm[13];
assign ap_CS_fsm_state15 = ap_CS_fsm[14];
assign ap_CS_fsm_state16 = ap_CS_fsm[15];
assign ap_CS_fsm_state17 = ap_CS_fsm[16];
assign ap_CS_fsm_state18 = ap_CS_fsm[17];
assign ap_CS_fsm_state19 = ap_CS_fsm[18];
assign ap_CS_fsm_state2 = ap_CS_fsm[1];
assign ap_CS_fsm_state20 = ap_CS_fsm[19];
assign ap_CS_fsm_state3 = ap_CS_fsm[2];
assign ap_CS_fsm_state4 = ap_CS_fsm[3];
assign ap_CS_fsm_state5 = ap_CS_fsm[4];
assign ap_CS_fsm_state6 = ap_CS_fsm[5];
assign ap_CS_fsm_state7 = ap_CS_fsm[6];
assign ap_CS_fsm_state8 = ap_CS_fsm[7];
assign ap_CS_fsm_state9 = ap_CS_fsm[8];
assign ap_done = op_30_ap_vld;
assign ap_ready = op_30_ap_vld;
assign grp_fu_171_p0 = { op_5[1], op_5[1], op_5[1], op_5[1], op_5, 3'h0 };
assign grp_fu_171_p1 = { op_7[7], op_7 };
assign grp_fu_205_p0 = { op_13[3], op_13 };
assign grp_fu_241_p0 = { op_9[15], op_9 };
assign grp_fu_241_p1 = { op_10[15], op_10 };
assign grp_fu_250_p0 = { add_ln69_1_reg_451[4], add_ln69_1_reg_451 };
assign grp_fu_250_p1 = { ret_V_7_reg_446[4], ret_V_7_reg_446 };
assign grp_fu_262_p0 = { add_ln69_2_reg_481[5], add_ln69_2_reg_481[5], add_ln69_2_reg_481[5], add_ln69_2_reg_481[5], add_ln69_2_reg_481[5], add_ln69_2_reg_481[5], add_ln69_2_reg_481[5], add_ln69_2_reg_481[5], add_ln69_2_reg_481[5], add_ln69_2_reg_481[5], add_ln69_2_reg_481[5], add_ln69_2_reg_481[5], add_ln69_2_reg_481 };
assign grp_fu_262_p1 = { add_ln69_reg_476[16], add_ln69_reg_476 };
assign grp_fu_279_p0 = { op_24_V_reg_496, 1'h0 };
assign grp_fu_279_p1 = { op_14[1], op_14[1], op_14[1], op_14[1], op_14[1], op_14[1], op_14[1], op_14[1], op_14[1], op_14[1], op_14[1], op_14[1], op_14[1], op_14[1], op_14[1], op_14[1], op_14[1], op_14 };
assign grp_fu_298_p0 = { tmp_reg_521[17], tmp_reg_521 };
assign grp_fu_338_p0 = { select_ln353_reg_538[18], select_ln353_reg_538[18], select_ln353_reg_538[18], select_ln353_reg_538[18], select_ln353_reg_538[18], select_ln353_reg_538[18], select_ln353_reg_538[18], select_ln353_reg_538[18], select_ln353_reg_538[18], select_ln353_reg_538[18], select_ln353_reg_538[18], select_ln353_reg_538[18], select_ln353_reg_538[18], select_ln353_reg_538, 2'h0 };
assign grp_fu_389_p0 = { 1'h0, op_18 };
assign grp_fu_389_p1 = { 4'h0, icmp_ln1495_reg_548 };
assign grp_fu_398_p0 = { 27'h0000000, add_ln69_6_reg_578 };
assign lhs_fu_155_p3 = { op_5, 3'h0 };
assign op_17_V_fu_344_p1 = op_11[0];
assign op_30 = grp_fu_398_p2;
assign p_Result_1_fu_304_p3 = ret_V_8_reg_516[18];
assign p_Result_s_fu_211_p3 = ret_V_6_reg_414[8];
assign sext_ln1192_1_fu_268_p0 = op_14;
assign sext_ln850_fu_295_p1 = { tmp_reg_521[17], tmp_reg_521 };
assign tmp_3_fu_327_p3 = { select_ln353_reg_538, 2'h0 };
assign trunc_ln851_1_fu_311_p0 = op_14;
assign trunc_ln851_1_fu_311_p1 = op_14[0];
assign trunc_ln851_fu_187_p1 = grp_fu_171_p2[3:0];
assign \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.ain_s0  = \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.a ;
assign \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.bin_s0  = \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.b ;
assign \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.s  = { \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.fas_s2 , \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.sum_s1  };
assign \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.u2.a  = \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.ain_s1 ;
assign \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.u2.b  = \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.bin_s1 ;
assign \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.u2.cin  = \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.carry_s1 ;
assign \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.facout_s2  = \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.u2.cout ;
assign \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.fas_s2  = \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.u2.s ;
assign \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.u1.a  = \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.a [3:0];
assign \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.u1.b  = \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.b [3:0];
assign \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.u1.cin  = 1'h0;
assign \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.facout_s1  = \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.u1.cout ;
assign \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.fas_s1  = \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.u1.s ;
assign \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.a  = \add_9s_9s_9_2_1_U1.din0 ;
assign \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.b  = \add_9s_9s_9_2_1_U1.din1 ;
assign \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.ce  = \add_9s_9s_9_2_1_U1.ce ;
assign \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.clk  = \add_9s_9s_9_2_1_U1.clk ;
assign \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.reset  = \add_9s_9s_9_2_1_U1.reset ;
assign \add_9s_9s_9_2_1_U1.dout  = \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.s ;
assign \add_9s_9s_9_2_1_U1.ce  = 1'h1;
assign \add_9s_9s_9_2_1_U1.clk  = ap_clk;
assign \add_9s_9s_9_2_1_U1.din0  = { op_5[1], op_5[1], op_5[1], op_5[1], op_5, 3'h0 };
assign \add_9s_9s_9_2_1_U1.din1  = { op_7[7], op_7 };
assign grp_fu_171_p2 = \add_9s_9s_9_2_1_U1.dout ;
assign \add_9s_9s_9_2_1_U1.reset  = ap_rst;
assign \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.ain_s0  = \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.a ;
assign \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.bin_s0  = \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.b ;
assign \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.s  = { \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.fas_s2 , \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.sum_s1  };
assign \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.u2.a  = \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.ain_s1 ;
assign \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.u2.b  = \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.bin_s1 ;
assign \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.u2.cin  = \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.carry_s1 ;
assign \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.facout_s2  = \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.u2.cout ;
assign \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.fas_s2  = \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.u2.s ;
assign \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.u1.a  = \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.a [2:0];
assign \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.u1.b  = \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.b [2:0];
assign \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.u1.cin  = 1'h0;
assign \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.facout_s1  = \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.u1.cout ;
assign \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.fas_s1  = \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.u1.s ;
assign \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.a  = \add_6s_6s_6_2_1_U5.din0 ;
assign \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.b  = \add_6s_6s_6_2_1_U5.din1 ;
assign \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.ce  = \add_6s_6s_6_2_1_U5.ce ;
assign \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.clk  = \add_6s_6s_6_2_1_U5.clk ;
assign \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.reset  = \add_6s_6s_6_2_1_U5.reset ;
assign \add_6s_6s_6_2_1_U5.dout  = \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.s ;
assign \add_6s_6s_6_2_1_U5.ce  = 1'h1;
assign \add_6s_6s_6_2_1_U5.clk  = ap_clk;
assign \add_6s_6s_6_2_1_U5.din0  = { add_ln69_1_reg_451[4], add_ln69_1_reg_451 };
assign \add_6s_6s_6_2_1_U5.din1  = { ret_V_7_reg_446[4], ret_V_7_reg_446 };
assign grp_fu_250_p2 = \add_6s_6s_6_2_1_U5.dout ;
assign \add_6s_6s_6_2_1_U5.reset  = ap_rst;
assign \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.ain_s0  = \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.a ;
assign \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.bin_s0  = \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.b ;
assign \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.s  = { \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.fas_s2 , \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.sum_s1  };
assign \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.u2.a  = \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.ain_s1 ;
assign \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.u2.b  = \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.bin_s1 ;
assign \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.u2.cin  = \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.carry_s1 ;
assign \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.facout_s2  = \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.u2.cout ;
assign \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.fas_s2  = \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.u2.s ;
assign \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.u1.a  = \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.a [1:0];
assign \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.u1.b  = \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.b [1:0];
assign \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.u1.cin  = 1'h0;
assign \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.facout_s1  = \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.u1.cout ;
assign \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.fas_s1  = \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.u1.s ;
assign \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.a  = \add_5s_5ns_5_2_1_U3.din0 ;
assign \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.b  = \add_5s_5ns_5_2_1_U3.din1 ;
assign \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.ce  = \add_5s_5ns_5_2_1_U3.ce ;
assign \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.clk  = \add_5s_5ns_5_2_1_U3.clk ;
assign \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.reset  = \add_5s_5ns_5_2_1_U3.reset ;
assign \add_5s_5ns_5_2_1_U3.dout  = \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.s ;
assign \add_5s_5ns_5_2_1_U3.ce  = 1'h1;
assign \add_5s_5ns_5_2_1_U3.clk  = ap_clk;
assign \add_5s_5ns_5_2_1_U3.din0  = { op_13[3], op_13 };
assign \add_5s_5ns_5_2_1_U3.din1  = 5'h01;
assign grp_fu_205_p2 = \add_5s_5ns_5_2_1_U3.dout ;
assign \add_5s_5ns_5_2_1_U3.reset  = ap_rst;
assign \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.ain_s0  = \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.a ;
assign \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.bin_s0  = \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.b ;
assign \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.s  = { \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.fas_s2 , \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.sum_s1  };
assign \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.u2.a  = \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.ain_s1 ;
assign \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.u2.b  = \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.bin_s1 ;
assign \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.u2.cin  = \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.carry_s1 ;
assign \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.facout_s2  = \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.u2.cout ;
assign \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.fas_s2  = \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.u2.s ;
assign \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.u1.a  = \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.a [1:0];
assign \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.u1.b  = \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.b [1:0];
assign \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.u1.cin  = 1'h0;
assign \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.facout_s1  = \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.u1.cout ;
assign \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.fas_s1  = \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.u1.s ;
assign \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.a  = \add_5ns_5ns_5_2_1_U2.din0 ;
assign \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.b  = \add_5ns_5ns_5_2_1_U2.din1 ;
assign \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.ce  = \add_5ns_5ns_5_2_1_U2.ce ;
assign \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.clk  = \add_5ns_5ns_5_2_1_U2.clk ;
assign \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.reset  = \add_5ns_5ns_5_2_1_U2.reset ;
assign \add_5ns_5ns_5_2_1_U2.dout  = \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.s ;
assign \add_5ns_5ns_5_2_1_U2.ce  = 1'h1;
assign \add_5ns_5ns_5_2_1_U2.clk  = ap_clk;
assign \add_5ns_5ns_5_2_1_U2.din0  = ret_V_reg_419;
assign \add_5ns_5ns_5_2_1_U2.din1  = 5'h01;
assign grp_fu_196_p2 = \add_5ns_5ns_5_2_1_U2.dout ;
assign \add_5ns_5ns_5_2_1_U2.reset  = ap_rst;
assign \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.ain_s0  = \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.a ;
assign \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.bin_s0  = \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.b ;
assign \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.s  = { \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.fas_s2 , \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.sum_s1  };
assign \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.u2.a  = \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.ain_s1 ;
assign \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.u2.b  = \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.bin_s1 ;
assign \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.u2.cin  = \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.carry_s1 ;
assign \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.facout_s2  = \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.u2.cout ;
assign \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.fas_s2  = \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.u2.s ;
assign \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.u1.a  = \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.a [1:0];
assign \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.u1.b  = \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.b [1:0];
assign \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.u1.cin  = 1'h0;
assign \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.facout_s1  = \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.u1.cout ;
assign \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.fas_s1  = \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.u1.s ;
assign \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.a  = \add_5ns_5ns_5_2_1_U11.din0 ;
assign \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.b  = \add_5ns_5ns_5_2_1_U11.din1 ;
assign \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.ce  = \add_5ns_5ns_5_2_1_U11.ce ;
assign \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.clk  = \add_5ns_5ns_5_2_1_U11.clk ;
assign \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.reset  = \add_5ns_5ns_5_2_1_U11.reset ;
assign \add_5ns_5ns_5_2_1_U11.dout  = \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.s ;
assign \add_5ns_5ns_5_2_1_U11.ce  = 1'h1;
assign \add_5ns_5ns_5_2_1_U11.clk  = ap_clk;
assign \add_5ns_5ns_5_2_1_U11.din0  = { 1'h0, op_18 };
assign \add_5ns_5ns_5_2_1_U11.din1  = { 4'h0, icmp_ln1495_reg_548 };
assign grp_fu_389_p2 = \add_5ns_5ns_5_2_1_U11.dout ;
assign \add_5ns_5ns_5_2_1_U11.reset  = ap_rst;
assign \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.ain_s0  = \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.a ;
assign \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.bin_s0  = \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.b ;
assign \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.s  = { \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.fas_s2 , \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.sum_s1  };
assign \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.u2.a  = \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.ain_s1 ;
assign \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.u2.b  = \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.bin_s1 ;
assign \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.u2.cin  = \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.carry_s1 ;
assign \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.facout_s2  = \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.u2.cout ;
assign \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.fas_s2  = \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.u2.s ;
assign \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.u1.a  = \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.a [16:0];
assign \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.u1.b  = \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.b [16:0];
assign \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.u1.cin  = 1'h0;
assign \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.facout_s1  = \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.u1.cout ;
assign \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.fas_s1  = \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.u1.s ;
assign \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.a  = \add_34s_34ns_34_2_1_U9.din0 ;
assign \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.b  = \add_34s_34ns_34_2_1_U9.din1 ;
assign \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.ce  = \add_34s_34ns_34_2_1_U9.ce ;
assign \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.clk  = \add_34s_34ns_34_2_1_U9.clk ;
assign \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.reset  = \add_34s_34ns_34_2_1_U9.reset ;
assign \add_34s_34ns_34_2_1_U9.dout  = \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.s ;
assign \add_34s_34ns_34_2_1_U9.ce  = 1'h1;
assign \add_34s_34ns_34_2_1_U9.clk  = ap_clk;
assign \add_34s_34ns_34_2_1_U9.din0  = { select_ln353_reg_538[18], select_ln353_reg_538[18], select_ln353_reg_538[18], select_ln353_reg_538[18], select_ln353_reg_538[18], select_ln353_reg_538[18], select_ln353_reg_538[18], select_ln353_reg_538[18], select_ln353_reg_538[18], select_ln353_reg_538[18], select_ln353_reg_538[18], select_ln353_reg_538[18], select_ln353_reg_538[18], select_ln353_reg_538, 2'h0 };
assign \add_34s_34ns_34_2_1_U9.din1  = 34'h000000004;
assign grp_fu_338_p2 = \add_34s_34ns_34_2_1_U9.dout ;
assign \add_34s_34ns_34_2_1_U9.reset  = ap_rst;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.ain_s0  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.a ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.bin_s0  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.b ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.s  = { \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.fas_s2 , \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.sum_s1  };
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.u2.a  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.ain_s1 ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.u2.b  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.bin_s1 ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.u2.cin  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.carry_s1 ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.facout_s2  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.u2.cout ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.fas_s2  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.u2.s ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.u1.a  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.a [15:0];
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.u1.b  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.b [15:0];
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.u1.cin  = 1'h0;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.facout_s1  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.u1.cout ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.fas_s1  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.u1.s ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.a  = \add_32ns_32ns_32_2_1_U12.din0 ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.b  = \add_32ns_32ns_32_2_1_U12.din1 ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.ce  = \add_32ns_32ns_32_2_1_U12.ce ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.clk  = \add_32ns_32ns_32_2_1_U12.clk ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.reset  = \add_32ns_32ns_32_2_1_U12.reset ;
assign \add_32ns_32ns_32_2_1_U12.dout  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.s ;
assign \add_32ns_32ns_32_2_1_U12.ce  = 1'h1;
assign \add_32ns_32ns_32_2_1_U12.clk  = ap_clk;
assign \add_32ns_32ns_32_2_1_U12.din0  = { 27'h0000000, add_ln69_6_reg_578 };
assign \add_32ns_32ns_32_2_1_U12.din1  = add_ln69_4_reg_573;
assign grp_fu_398_p2 = \add_32ns_32ns_32_2_1_U12.dout ;
assign \add_32ns_32ns_32_2_1_U12.reset  = ap_rst;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.ain_s0  = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.a ;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.bin_s0  = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.b ;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.s  = { \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.fas_s2 , \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.sum_s1  };
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.u2.a  = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.ain_s1 ;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.u2.b  = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.bin_s1 ;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.u2.cin  = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.carry_s1 ;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.facout_s2  = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.u2.cout ;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.fas_s2  = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.u2.s ;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.u1.a  = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.a [15:0];
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.u1.b  = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.b [15:0];
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.u1.cin  = 1'h0;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.facout_s1  = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.u1.cout ;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.fas_s1  = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.u1.s ;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.a  = \add_32ns_32ns_32_2_1_U10.din0 ;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.b  = \add_32ns_32ns_32_2_1_U10.din1 ;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.ce  = \add_32ns_32ns_32_2_1_U10.ce ;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.clk  = \add_32ns_32ns_32_2_1_U10.clk ;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.reset  = \add_32ns_32ns_32_2_1_U10.reset ;
assign \add_32ns_32ns_32_2_1_U10.dout  = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.s ;
assign \add_32ns_32ns_32_2_1_U10.ce  = 1'h1;
assign \add_32ns_32ns_32_2_1_U10.clk  = ap_clk;
assign \add_32ns_32ns_32_2_1_U10.din0  = op_26_V_reg_553;
assign \add_32ns_32ns_32_2_1_U10.din1  = select_ln69_reg_558;
assign grp_fu_385_p2 = \add_32ns_32ns_32_2_1_U10.dout ;
assign \add_32ns_32ns_32_2_1_U10.reset  = ap_rst;
assign \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.ain_s0  = \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.a ;
assign \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.bin_s0  = \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.b ;
assign \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.s  = { \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.fas_s2 , \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.sum_s1  };
assign \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.u2.a  = \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.ain_s1 ;
assign \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.u2.b  = \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.bin_s1 ;
assign \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.u2.cin  = \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.carry_s1 ;
assign \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.facout_s2  = \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.u2.cout ;
assign \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.fas_s2  = \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.u2.s ;
assign \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.u1.a  = \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.a [8:0];
assign \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.u1.b  = \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.b [8:0];
assign \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.u1.cin  = 1'h0;
assign \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.facout_s1  = \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.u1.cout ;
assign \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.fas_s1  = \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.u1.s ;
assign \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.a  = \add_19s_19ns_19_2_1_U8.din0 ;
assign \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.b  = \add_19s_19ns_19_2_1_U8.din1 ;
assign \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.ce  = \add_19s_19ns_19_2_1_U8.ce ;
assign \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.clk  = \add_19s_19ns_19_2_1_U8.clk ;
assign \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.reset  = \add_19s_19ns_19_2_1_U8.reset ;
assign \add_19s_19ns_19_2_1_U8.dout  = \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.s ;
assign \add_19s_19ns_19_2_1_U8.ce  = 1'h1;
assign \add_19s_19ns_19_2_1_U8.clk  = ap_clk;
assign \add_19s_19ns_19_2_1_U8.din0  = { tmp_reg_521[17], tmp_reg_521 };
assign \add_19s_19ns_19_2_1_U8.din1  = 19'h00001;
assign grp_fu_298_p2 = \add_19s_19ns_19_2_1_U8.dout ;
assign \add_19s_19ns_19_2_1_U8.reset  = ap_rst;
assign \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.ain_s0  = \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.a ;
assign \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.bin_s0  = \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.b ;
assign \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.s  = { \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.fas_s2 , \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.sum_s1  };
assign \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.u2.a  = \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.ain_s1 ;
assign \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.u2.b  = \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.bin_s1 ;
assign \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.u2.cin  = \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.carry_s1 ;
assign \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.facout_s2  = \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.u2.cout ;
assign \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.fas_s2  = \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.u2.s ;
assign \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.u1.a  = \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.a [8:0];
assign \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.u1.b  = \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.b [8:0];
assign \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.u1.cin  = 1'h0;
assign \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.facout_s1  = \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.u1.cout ;
assign \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.fas_s1  = \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.u1.s ;
assign \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.a  = \add_19ns_19s_19_2_1_U7.din0 ;
assign \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.b  = \add_19ns_19s_19_2_1_U7.din1 ;
assign \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.ce  = \add_19ns_19s_19_2_1_U7.ce ;
assign \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.clk  = \add_19ns_19s_19_2_1_U7.clk ;
assign \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.reset  = \add_19ns_19s_19_2_1_U7.reset ;
assign \add_19ns_19s_19_2_1_U7.dout  = \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.s ;
assign \add_19ns_19s_19_2_1_U7.ce  = 1'h1;
assign \add_19ns_19s_19_2_1_U7.clk  = ap_clk;
assign \add_19ns_19s_19_2_1_U7.din0  = { op_24_V_reg_496, 1'h0 };
assign \add_19ns_19s_19_2_1_U7.din1  = { op_14[1], op_14[1], op_14[1], op_14[1], op_14[1], op_14[1], op_14[1], op_14[1], op_14[1], op_14[1], op_14[1], op_14[1], op_14[1], op_14[1], op_14[1], op_14[1], op_14[1], op_14 };
assign grp_fu_279_p2 = \add_19ns_19s_19_2_1_U7.dout ;
assign \add_19ns_19s_19_2_1_U7.reset  = ap_rst;
assign \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.ain_s0  = \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.a ;
assign \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.bin_s0  = \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.b ;
assign \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.s  = { \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.fas_s2 , \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.sum_s1  };
assign \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.u2.a  = \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.ain_s1 ;
assign \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.u2.b  = \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.bin_s1 ;
assign \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.u2.cin  = \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.carry_s1 ;
assign \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.facout_s2  = \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.u2.cout ;
assign \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.fas_s2  = \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.u2.s ;
assign \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.u1.a  = \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.a [8:0];
assign \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.u1.b  = \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.b [8:0];
assign \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.u1.cin  = 1'h0;
assign \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.facout_s1  = \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.u1.cout ;
assign \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.fas_s1  = \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.u1.s ;
assign \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.a  = \add_18s_18s_18_2_1_U6.din0 ;
assign \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.b  = \add_18s_18s_18_2_1_U6.din1 ;
assign \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.ce  = \add_18s_18s_18_2_1_U6.ce ;
assign \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.clk  = \add_18s_18s_18_2_1_U6.clk ;
assign \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.reset  = \add_18s_18s_18_2_1_U6.reset ;
assign \add_18s_18s_18_2_1_U6.dout  = \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.s ;
assign \add_18s_18s_18_2_1_U6.ce  = 1'h1;
assign \add_18s_18s_18_2_1_U6.clk  = ap_clk;
assign \add_18s_18s_18_2_1_U6.din0  = { add_ln69_2_reg_481[5], add_ln69_2_reg_481[5], add_ln69_2_reg_481[5], add_ln69_2_reg_481[5], add_ln69_2_reg_481[5], add_ln69_2_reg_481[5], add_ln69_2_reg_481[5], add_ln69_2_reg_481[5], add_ln69_2_reg_481[5], add_ln69_2_reg_481[5], add_ln69_2_reg_481[5], add_ln69_2_reg_481[5], add_ln69_2_reg_481 };
assign \add_18s_18s_18_2_1_U6.din1  = { add_ln69_reg_476[16], add_ln69_reg_476 };
assign grp_fu_262_p2 = \add_18s_18s_18_2_1_U6.dout ;
assign \add_18s_18s_18_2_1_U6.reset  = ap_rst;
assign \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.ain_s0  = \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.a ;
assign \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.bin_s0  = \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.b ;
assign \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.s  = { \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.fas_s2 , \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.sum_s1  };
assign \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.u2.a  = \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.ain_s1 ;
assign \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.u2.b  = \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.bin_s1 ;
assign \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.u2.cin  = \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.carry_s1 ;
assign \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.facout_s2  = \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.u2.cout ;
assign \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.fas_s2  = \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.u2.s ;
assign \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.u1.a  = \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.a [7:0];
assign \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.u1.b  = \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.b [7:0];
assign \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.u1.cin  = 1'h0;
assign \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.facout_s1  = \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.u1.cout ;
assign \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.fas_s1  = \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.u1.s ;
assign \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.a  = \add_17s_17s_17_2_1_U4.din0 ;
assign \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.b  = \add_17s_17s_17_2_1_U4.din1 ;
assign \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.ce  = \add_17s_17s_17_2_1_U4.ce ;
assign \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.clk  = \add_17s_17s_17_2_1_U4.clk ;
assign \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.reset  = \add_17s_17s_17_2_1_U4.reset ;
assign \add_17s_17s_17_2_1_U4.dout  = \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.s ;
assign \add_17s_17s_17_2_1_U4.ce  = 1'h1;
assign \add_17s_17s_17_2_1_U4.clk  = ap_clk;
assign \add_17s_17s_17_2_1_U4.din0  = { op_9[15], op_9 };
assign \add_17s_17s_17_2_1_U4.din1  = { op_10[15], op_10 };
assign grp_fu_241_p2 = \add_17s_17s_17_2_1_U4.dout ;
assign \add_17s_17s_17_2_1_U4.reset  = ap_rst;
endmodule


// Machine B:
// Processed by function `add_clk_enable_signal` in `verilog_tricks.py`.
// Processed by function `remove_reset_signal` in `verilog_tricks.py`.
module top_B (
  ap_clk,
  ap_start,
  ap_done,
  ap_idle,
  ap_ready,
  op_0,
  op_5,
  op_7,
  op_9,
  op_10,
  op_11,
  op_12,
  op_13,
  op_14,
  op_18,
  op_30,
  op_30_ap_vld,
clk_enable
);
input clk_enable;


input ap_clk;
wire ap_rst;
assign ap_rst = op_30_ap_vld;
input ap_start;
input [1:0] op_0;
input [15:0] op_10;
input [1:0] op_11;
input [7:0] op_12;
input [3:0] op_13;
input [1:0] op_14;
input [3:0] op_18;
input [1:0] op_5;
input [7:0] op_7;
input [15:0] op_9;
output ap_done;
output ap_idle;
output ap_ready;
output [31:0] op_30;
output op_30_ap_vld;


reg [8:0] \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.ain_s1 ;
reg [8:0] \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.bin_s1 ;
reg \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.carry_s1 ;
reg [7:0] \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.sum_s1 ;
reg [8:0] \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.ain_s1 ;
reg [8:0] \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.bin_s1 ;
reg \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.carry_s1 ;
reg [8:0] \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.sum_s1 ;
reg [9:0] \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.ain_s1 ;
reg [9:0] \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.bin_s1 ;
reg \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.carry_s1 ;
reg [8:0] \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.sum_s1 ;
reg [9:0] \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.ain_s1 ;
reg [9:0] \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.bin_s1 ;
reg \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.carry_s1 ;
reg [8:0] \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.sum_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.ain_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.bin_s1 ;
reg \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.carry_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.sum_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.ain_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.bin_s1 ;
reg \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.carry_s1 ;
reg [15:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.sum_s1 ;
reg [16:0] \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.ain_s1 ;
reg [16:0] \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.bin_s1 ;
reg \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.carry_s1 ;
reg [16:0] \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.sum_s1 ;
reg [2:0] \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.ain_s1 ;
reg [2:0] \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.bin_s1 ;
reg \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.carry_s1 ;
reg [1:0] \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.sum_s1 ;
reg [2:0] \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.ain_s1 ;
reg [2:0] \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.bin_s1 ;
reg \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.carry_s1 ;
reg [1:0] \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.sum_s1 ;
reg [2:0] \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.ain_s1 ;
reg [2:0] \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.bin_s1 ;
reg \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.carry_s1 ;
reg [1:0] \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.sum_s1 ;
reg [2:0] \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.ain_s1 ;
reg [2:0] \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.bin_s1 ;
reg \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.carry_s1 ;
reg [2:0] \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.sum_s1 ;
reg [4:0] \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.ain_s1 ;
reg [4:0] \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.bin_s1 ;
reg \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.carry_s1 ;
reg [3:0] \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.sum_s1 ;
reg [18:0] add_ln691_reg_533;
reg [4:0] add_ln69_1_reg_451;
reg [5:0] add_ln69_2_reg_481;
reg [31:0] add_ln69_4_reg_573;
reg [4:0] add_ln69_6_reg_578;
reg [16:0] add_ln69_reg_476;
reg [19:0] ap_CS_fsm = 20'h00001;
reg icmp_ln1495_reg_548;
reg icmp_ln851_reg_431;
reg [17:0] op_24_V_reg_496;
reg [31:0] op_26_V_reg_553;
reg [4:0] ret_V_2_reg_436;
reg [8:0] ret_V_6_reg_414;
reg [4:0] ret_V_7_reg_446;
reg [18:0] ret_V_8_reg_516;
reg [4:0] ret_V_reg_419;
reg [18:0] select_ln353_reg_538;
reg [31:0] select_ln69_reg_558;
reg [18:0] sext_ln850_reg_526;
reg [17:0] tmp_reg_521;
reg [3:0] trunc_ln851_reg_426;
wire [18:0] _000_;
wire [4:0] _001_;
wire [5:0] _002_;
wire [31:0] _003_;
wire [4:0] _004_;
wire [16:0] _005_;
wire [19:0] _006_;
wire _007_;
wire _008_;
wire [17:0] _009_;
wire [31:0] _010_;
wire [4:0] _011_;
wire [8:0] _012_;
wire [4:0] _013_;
wire [18:0] _014_;
wire [4:0] _015_;
wire [18:0] _016_;
wire [31:0] _017_;
wire [18:0] _018_;
wire [17:0] _019_;
wire [3:0] _020_;
wire [1:0] _021_;
wire _022_;
wire _023_;
wire _024_;
wire _025_;
wire [8:0] _026_;
wire [8:0] _027_;
wire _028_;
wire [7:0] _029_;
wire [8:0] _030_;
wire [9:0] _031_;
wire [8:0] _032_;
wire [8:0] _033_;
wire _034_;
wire [8:0] _035_;
wire [9:0] _036_;
wire [9:0] _037_;
wire [9:0] _038_;
wire [9:0] _039_;
wire _040_;
wire [8:0] _041_;
wire [9:0] _042_;
wire [10:0] _043_;
wire [9:0] _044_;
wire [9:0] _045_;
wire _046_;
wire [8:0] _047_;
wire [9:0] _048_;
wire [10:0] _049_;
wire [15:0] _050_;
wire [15:0] _051_;
wire _052_;
wire [15:0] _053_;
wire [16:0] _054_;
wire [16:0] _055_;
wire [15:0] _056_;
wire [15:0] _057_;
wire _058_;
wire [15:0] _059_;
wire [16:0] _060_;
wire [16:0] _061_;
wire [16:0] _062_;
wire [16:0] _063_;
wire _064_;
wire [16:0] _065_;
wire [17:0] _066_;
wire [17:0] _067_;
wire [2:0] _068_;
wire [2:0] _069_;
wire _070_;
wire [1:0] _071_;
wire [2:0] _072_;
wire [3:0] _073_;
wire [2:0] _074_;
wire [2:0] _075_;
wire _076_;
wire [1:0] _077_;
wire [2:0] _078_;
wire [3:0] _079_;
wire [2:0] _080_;
wire [2:0] _081_;
wire _082_;
wire [1:0] _083_;
wire [2:0] _084_;
wire [3:0] _085_;
wire [2:0] _086_;
wire [2:0] _087_;
wire _088_;
wire [2:0] _089_;
wire [3:0] _090_;
wire [3:0] _091_;
wire [4:0] _092_;
wire [4:0] _093_;
wire _094_;
wire [3:0] _095_;
wire [4:0] _096_;
wire [5:0] _097_;
wire _098_;
wire _099_;
wire _100_;
wire _101_;
wire _102_;
wire _103_;
wire _104_;
wire _105_;
wire _106_;
wire _107_;
wire _108_;
wire _109_;
wire _110_;
wire _111_;
wire _112_;
wire _113_;
wire _114_;
wire _115_;
wire _116_;
wire _117_;
wire _118_;
wire \add_17s_17s_17_2_1_U4.ce ;
wire \add_17s_17s_17_2_1_U4.clk ;
wire [16:0] \add_17s_17s_17_2_1_U4.din0 ;
wire [16:0] \add_17s_17s_17_2_1_U4.din1 ;
wire [16:0] \add_17s_17s_17_2_1_U4.dout ;
wire \add_17s_17s_17_2_1_U4.reset ;
wire [16:0] \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.a ;
wire [16:0] \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.ain_s0 ;
wire [16:0] \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.b ;
wire [16:0] \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.bin_s0 ;
wire \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.ce ;
wire \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.clk ;
wire \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.facout_s1 ;
wire \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.facout_s2 ;
wire [7:0] \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.fas_s1 ;
wire [8:0] \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.fas_s2 ;
wire \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.reset ;
wire [16:0] \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.s ;
wire [7:0] \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.u1.a ;
wire [7:0] \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.u1.b ;
wire \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.u1.cin ;
wire \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.u1.cout ;
wire [7:0] \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.u1.s ;
wire [8:0] \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.u2.a ;
wire [8:0] \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.u2.b ;
wire \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.u2.cin ;
wire \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.u2.cout ;
wire [8:0] \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.u2.s ;
wire \add_18s_18s_18_2_1_U6.ce ;
wire \add_18s_18s_18_2_1_U6.clk ;
wire [17:0] \add_18s_18s_18_2_1_U6.din0 ;
wire [17:0] \add_18s_18s_18_2_1_U6.din1 ;
wire [17:0] \add_18s_18s_18_2_1_U6.dout ;
wire \add_18s_18s_18_2_1_U6.reset ;
wire [17:0] \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.a ;
wire [17:0] \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.ain_s0 ;
wire [17:0] \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.b ;
wire [17:0] \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.bin_s0 ;
wire \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.ce ;
wire \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.clk ;
wire \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.facout_s1 ;
wire \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.facout_s2 ;
wire [8:0] \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.fas_s1 ;
wire [8:0] \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.fas_s2 ;
wire \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.reset ;
wire [17:0] \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.s ;
wire [8:0] \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.u1.a ;
wire [8:0] \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.u1.b ;
wire \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.u1.cin ;
wire \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.u1.cout ;
wire [8:0] \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.u1.s ;
wire [8:0] \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.u2.a ;
wire [8:0] \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.u2.b ;
wire \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.u2.cin ;
wire \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.u2.cout ;
wire [8:0] \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.u2.s ;
wire \add_19ns_19s_19_2_1_U7.ce ;
wire \add_19ns_19s_19_2_1_U7.clk ;
wire [18:0] \add_19ns_19s_19_2_1_U7.din0 ;
wire [18:0] \add_19ns_19s_19_2_1_U7.din1 ;
wire [18:0] \add_19ns_19s_19_2_1_U7.dout ;
wire \add_19ns_19s_19_2_1_U7.reset ;
wire [18:0] \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.a ;
wire [18:0] \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.ain_s0 ;
wire [18:0] \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.b ;
wire [18:0] \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.bin_s0 ;
wire \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.ce ;
wire \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.clk ;
wire \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.facout_s1 ;
wire \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.facout_s2 ;
wire [8:0] \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.fas_s1 ;
wire [9:0] \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.fas_s2 ;
wire \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.reset ;
wire [18:0] \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.s ;
wire [8:0] \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.u1.a ;
wire [8:0] \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.u1.b ;
wire \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.u1.cin ;
wire \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.u1.cout ;
wire [8:0] \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.u1.s ;
wire [9:0] \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.u2.a ;
wire [9:0] \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.u2.b ;
wire \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.u2.cin ;
wire \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.u2.cout ;
wire [9:0] \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.u2.s ;
wire \add_19s_19ns_19_2_1_U8.ce ;
wire \add_19s_19ns_19_2_1_U8.clk ;
wire [18:0] \add_19s_19ns_19_2_1_U8.din0 ;
wire [18:0] \add_19s_19ns_19_2_1_U8.din1 ;
wire [18:0] \add_19s_19ns_19_2_1_U8.dout ;
wire \add_19s_19ns_19_2_1_U8.reset ;
wire [18:0] \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.a ;
wire [18:0] \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.ain_s0 ;
wire [18:0] \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.b ;
wire [18:0] \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.bin_s0 ;
wire \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.ce ;
wire \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.clk ;
wire \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.facout_s1 ;
wire \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.facout_s2 ;
wire [8:0] \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.fas_s1 ;
wire [9:0] \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.fas_s2 ;
wire \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.reset ;
wire [18:0] \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.s ;
wire [8:0] \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.u1.a ;
wire [8:0] \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.u1.b ;
wire \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.u1.cin ;
wire \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.u1.cout ;
wire [8:0] \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.u1.s ;
wire [9:0] \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.u2.a ;
wire [9:0] \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.u2.b ;
wire \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.u2.cin ;
wire \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.u2.cout ;
wire [9:0] \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.u2.s ;
wire \add_32ns_32ns_32_2_1_U10.ce ;
wire \add_32ns_32ns_32_2_1_U10.clk ;
wire [31:0] \add_32ns_32ns_32_2_1_U10.din0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U10.din1 ;
wire [31:0] \add_32ns_32ns_32_2_1_U10.dout ;
wire \add_32ns_32ns_32_2_1_U10.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.a ;
wire [31:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.ain_s0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.b ;
wire [31:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.bin_s0 ;
wire \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.ce ;
wire \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.clk ;
wire \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.facout_s1 ;
wire \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.facout_s2 ;
wire [15:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.fas_s1 ;
wire [15:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.fas_s2 ;
wire \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.u1.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.u1.b ;
wire \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.u1.cin ;
wire \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.u1.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.u1.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.u2.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.u2.b ;
wire \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.u2.cin ;
wire \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.u2.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.u2.s ;
wire \add_32ns_32ns_32_2_1_U12.ce ;
wire \add_32ns_32ns_32_2_1_U12.clk ;
wire [31:0] \add_32ns_32ns_32_2_1_U12.din0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U12.din1 ;
wire [31:0] \add_32ns_32ns_32_2_1_U12.dout ;
wire \add_32ns_32ns_32_2_1_U12.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.a ;
wire [31:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.ain_s0 ;
wire [31:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.b ;
wire [31:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.bin_s0 ;
wire \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.ce ;
wire \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.clk ;
wire \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.facout_s1 ;
wire \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.facout_s2 ;
wire [15:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.fas_s1 ;
wire [15:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.fas_s2 ;
wire \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.reset ;
wire [31:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.u1.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.u1.b ;
wire \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.u1.cin ;
wire \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.u1.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.u1.s ;
wire [15:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.u2.a ;
wire [15:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.u2.b ;
wire \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.u2.cin ;
wire \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.u2.cout ;
wire [15:0] \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.u2.s ;
wire \add_34s_34ns_34_2_1_U9.ce ;
wire \add_34s_34ns_34_2_1_U9.clk ;
wire [33:0] \add_34s_34ns_34_2_1_U9.din0 ;
wire [33:0] \add_34s_34ns_34_2_1_U9.din1 ;
wire [33:0] \add_34s_34ns_34_2_1_U9.dout ;
wire \add_34s_34ns_34_2_1_U9.reset ;
wire [33:0] \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.a ;
wire [33:0] \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.ain_s0 ;
wire [33:0] \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.b ;
wire [33:0] \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.bin_s0 ;
wire \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.ce ;
wire \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.clk ;
wire \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.facout_s1 ;
wire \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.facout_s2 ;
wire [16:0] \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.fas_s1 ;
wire [16:0] \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.fas_s2 ;
wire \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.reset ;
wire [33:0] \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.s ;
wire [16:0] \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.u1.a ;
wire [16:0] \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.u1.b ;
wire \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.u1.cin ;
wire \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.u1.cout ;
wire [16:0] \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.u1.s ;
wire [16:0] \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.u2.a ;
wire [16:0] \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.u2.b ;
wire \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.u2.cin ;
wire \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.u2.cout ;
wire [16:0] \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.u2.s ;
wire \add_5ns_5ns_5_2_1_U11.ce ;
wire \add_5ns_5ns_5_2_1_U11.clk ;
wire [4:0] \add_5ns_5ns_5_2_1_U11.din0 ;
wire [4:0] \add_5ns_5ns_5_2_1_U11.din1 ;
wire [4:0] \add_5ns_5ns_5_2_1_U11.dout ;
wire \add_5ns_5ns_5_2_1_U11.reset ;
wire [4:0] \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.a ;
wire [4:0] \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.ain_s0 ;
wire [4:0] \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.b ;
wire [4:0] \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.bin_s0 ;
wire \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.ce ;
wire \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.clk ;
wire \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.facout_s1 ;
wire \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.facout_s2 ;
wire [1:0] \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.fas_s1 ;
wire [2:0] \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.fas_s2 ;
wire \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.reset ;
wire [4:0] \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.s ;
wire [1:0] \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.u1.a ;
wire [1:0] \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.u1.b ;
wire \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.u1.cin ;
wire \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.u1.cout ;
wire [1:0] \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.u1.s ;
wire [2:0] \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.u2.a ;
wire [2:0] \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.u2.b ;
wire \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.u2.cin ;
wire \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.u2.cout ;
wire [2:0] \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.u2.s ;
wire \add_5ns_5ns_5_2_1_U2.ce ;
wire \add_5ns_5ns_5_2_1_U2.clk ;
wire [4:0] \add_5ns_5ns_5_2_1_U2.din0 ;
wire [4:0] \add_5ns_5ns_5_2_1_U2.din1 ;
wire [4:0] \add_5ns_5ns_5_2_1_U2.dout ;
wire \add_5ns_5ns_5_2_1_U2.reset ;
wire [4:0] \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.a ;
wire [4:0] \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.ain_s0 ;
wire [4:0] \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.b ;
wire [4:0] \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.bin_s0 ;
wire \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.ce ;
wire \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.clk ;
wire \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.facout_s1 ;
wire \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.facout_s2 ;
wire [1:0] \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.fas_s1 ;
wire [2:0] \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.fas_s2 ;
wire \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.reset ;
wire [4:0] \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.s ;
wire [1:0] \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.u1.a ;
wire [1:0] \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.u1.b ;
wire \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.u1.cin ;
wire \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.u1.cout ;
wire [1:0] \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.u1.s ;
wire [2:0] \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.u2.a ;
wire [2:0] \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.u2.b ;
wire \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.u2.cin ;
wire \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.u2.cout ;
wire [2:0] \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.u2.s ;
wire \add_5s_5ns_5_2_1_U3.ce ;
wire \add_5s_5ns_5_2_1_U3.clk ;
wire [4:0] \add_5s_5ns_5_2_1_U3.din0 ;
wire [4:0] \add_5s_5ns_5_2_1_U3.din1 ;
wire [4:0] \add_5s_5ns_5_2_1_U3.dout ;
wire \add_5s_5ns_5_2_1_U3.reset ;
wire [4:0] \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.a ;
wire [4:0] \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.ain_s0 ;
wire [4:0] \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.b ;
wire [4:0] \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.bin_s0 ;
wire \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.ce ;
wire \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.clk ;
wire \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.facout_s1 ;
wire \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.facout_s2 ;
wire [1:0] \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.fas_s1 ;
wire [2:0] \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.fas_s2 ;
wire \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.reset ;
wire [4:0] \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.s ;
wire [1:0] \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.u1.a ;
wire [1:0] \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.u1.b ;
wire \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.u1.cin ;
wire \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.u1.cout ;
wire [1:0] \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.u1.s ;
wire [2:0] \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.u2.a ;
wire [2:0] \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.u2.b ;
wire \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.u2.cin ;
wire \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.u2.cout ;
wire [2:0] \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.u2.s ;
wire \add_6s_6s_6_2_1_U5.ce ;
wire \add_6s_6s_6_2_1_U5.clk ;
wire [5:0] \add_6s_6s_6_2_1_U5.din0 ;
wire [5:0] \add_6s_6s_6_2_1_U5.din1 ;
wire [5:0] \add_6s_6s_6_2_1_U5.dout ;
wire \add_6s_6s_6_2_1_U5.reset ;
wire [5:0] \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.a ;
wire [5:0] \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.ain_s0 ;
wire [5:0] \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.b ;
wire [5:0] \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.bin_s0 ;
wire \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.ce ;
wire \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.clk ;
wire \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.facout_s1 ;
wire \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.facout_s2 ;
wire [2:0] \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.fas_s1 ;
wire [2:0] \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.fas_s2 ;
wire \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.reset ;
wire [5:0] \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.s ;
wire [2:0] \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.u1.a ;
wire [2:0] \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.u1.b ;
wire \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.u1.cin ;
wire \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.u1.cout ;
wire [2:0] \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.u1.s ;
wire [2:0] \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.u2.a ;
wire [2:0] \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.u2.b ;
wire \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.u2.cin ;
wire \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.u2.cout ;
wire [2:0] \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.u2.s ;
wire \add_9s_9s_9_2_1_U1.ce ;
wire \add_9s_9s_9_2_1_U1.clk ;
wire [8:0] \add_9s_9s_9_2_1_U1.din0 ;
wire [8:0] \add_9s_9s_9_2_1_U1.din1 ;
wire [8:0] \add_9s_9s_9_2_1_U1.dout ;
wire \add_9s_9s_9_2_1_U1.reset ;
wire [8:0] \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.a ;
wire [8:0] \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.ain_s0 ;
wire [8:0] \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.b ;
wire [8:0] \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.bin_s0 ;
wire \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.ce ;
wire \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.clk ;
wire \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.facout_s1 ;
wire \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.facout_s2 ;
wire [3:0] \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.fas_s1 ;
wire [4:0] \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.fas_s2 ;
wire \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.reset ;
wire [8:0] \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.s ;
wire [3:0] \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.u1.a ;
wire [3:0] \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.u1.b ;
wire \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.u1.cin ;
wire \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.u1.cout ;
wire [3:0] \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.u1.s ;
wire [4:0] \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.u2.a ;
wire [4:0] \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.u2.b ;
wire \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.u2.cin ;
wire \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.u2.cout ;
wire [4:0] \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.u2.s ;
wire ap_CS_fsm_state1;
wire ap_CS_fsm_state10;
wire ap_CS_fsm_state11;
wire ap_CS_fsm_state12;
wire ap_CS_fsm_state13;
wire ap_CS_fsm_state14;
wire ap_CS_fsm_state15;
wire ap_CS_fsm_state16;
wire ap_CS_fsm_state17;
wire ap_CS_fsm_state18;
wire ap_CS_fsm_state19;
wire ap_CS_fsm_state2;
wire ap_CS_fsm_state20;
wire ap_CS_fsm_state3;
wire ap_CS_fsm_state4;
wire ap_CS_fsm_state5;
wire ap_CS_fsm_state6;
wire ap_CS_fsm_state7;
wire ap_CS_fsm_state8;
wire ap_CS_fsm_state9;
wire [19:0] ap_NS_fsm;
wire ap_clk;
wire ap_done;
wire ap_idle;
wire ap_ready;
wire ap_rst;
wire ap_start;
wire [8:0] grp_fu_171_p0;
wire [8:0] grp_fu_171_p1;
wire [8:0] grp_fu_171_p2;
wire [4:0] grp_fu_196_p2;
wire [4:0] grp_fu_205_p0;
wire [4:0] grp_fu_205_p2;
wire [16:0] grp_fu_241_p0;
wire [16:0] grp_fu_241_p1;
wire [16:0] grp_fu_241_p2;
wire [5:0] grp_fu_250_p0;
wire [5:0] grp_fu_250_p1;
wire [5:0] grp_fu_250_p2;
wire [17:0] grp_fu_262_p0;
wire [17:0] grp_fu_262_p1;
wire [17:0] grp_fu_262_p2;
wire [18:0] grp_fu_279_p0;
wire [18:0] grp_fu_279_p1;
wire [18:0] grp_fu_279_p2;
wire [18:0] grp_fu_298_p0;
wire [18:0] grp_fu_298_p2;
wire [33:0] grp_fu_338_p0;
wire [33:0] grp_fu_338_p2;
wire [31:0] grp_fu_385_p2;
wire [4:0] grp_fu_389_p0;
wire [4:0] grp_fu_389_p1;
wire [4:0] grp_fu_389_p2;
wire [31:0] grp_fu_398_p0;
wire [31:0] grp_fu_398_p2;
wire icmp_ln1495_fu_348_p2;
wire icmp_ln851_fu_191_p2;
wire [4:0] lhs_fu_155_p3;
wire [1:0] op_0;
wire [15:0] op_10;
wire [1:0] op_11;
wire [7:0] op_12;
wire [3:0] op_13;
wire [1:0] op_14;
wire op_17_V_fu_344_p1;
wire [3:0] op_18;
wire [31:0] op_30;
wire op_30_ap_vld;
wire [1:0] op_5;
wire [7:0] op_7;
wire [15:0] op_9;
wire p_Result_1_fu_304_p3;
wire p_Result_s_fu_211_p3;
wire [4:0] ret_V_7_fu_223_p3;
wire [18:0] select_ln353_fu_320_p3;
wire [31:0] select_ln69_fu_370_p3;
wire [18:0] select_ln850_2_fu_314_p3;
wire [4:0] select_ln850_fu_218_p3;
wire [1:0] sext_ln1192_1_fu_268_p0;
wire [18:0] sext_ln850_fu_295_p1;
wire [20:0] tmp_3_fu_327_p3;
wire [1:0] trunc_ln851_1_fu_311_p0;
wire trunc_ln851_1_fu_311_p1;
wire [3:0] trunc_ln851_fu_187_p1;


assign _022_ = _024_ & ap_CS_fsm[0];
assign _023_ = ap_start & ap_CS_fsm[0];
assign _024_ = ~ ap_start;
assign _025_ = ! trunc_ln851_reg_426;
always @(posedge \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.clk )
\add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.bin_s1  <= _027_;
always @(posedge \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.clk )
\add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.ain_s1  <= _026_;
always @(posedge \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.clk )
\add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.sum_s1  <= _029_;
always @(posedge \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.clk )
\add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.carry_s1  <= _028_;
assign _027_ = \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.ce  ? \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.b [16:8] : \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.bin_s1 ;
assign _026_ = \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.ce  ? \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.a [16:8] : \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.ain_s1 ;
assign _028_ = \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.ce  ? \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.facout_s1  : \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.carry_s1 ;
assign _029_ = \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.ce  ? \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.fas_s1  : \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.sum_s1 ;
assign _030_ = \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.u1.a  + \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.u1.b ;
assign { \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.u1.cout , \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.u1.s  } = _030_ + \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.u1.cin ;
assign _031_ = \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.u2.a  + \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.u2.b ;
assign { \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.u2.cout , \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.u2.s  } = _031_ + \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.u2.cin ;
always @(posedge \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.clk )
\add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.bin_s1  <= _033_;
always @(posedge \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.clk )
\add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.ain_s1  <= _032_;
always @(posedge \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.clk )
\add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.sum_s1  <= _035_;
always @(posedge \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.clk )
\add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.carry_s1  <= _034_;
assign _033_ = \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.ce  ? \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.b [17:9] : \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.bin_s1 ;
assign _032_ = \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.ce  ? \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.a [17:9] : \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.ain_s1 ;
assign _034_ = \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.ce  ? \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.facout_s1  : \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.carry_s1 ;
assign _035_ = \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.ce  ? \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.fas_s1  : \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.sum_s1 ;
assign _036_ = \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.u1.a  + \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.u1.b ;
assign { \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.u1.cout , \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.u1.s  } = _036_ + \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.u1.cin ;
assign _037_ = \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.u2.a  + \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.u2.b ;
assign { \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.u2.cout , \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.u2.s  } = _037_ + \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.u2.cin ;
always @(posedge \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.clk )
\add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.bin_s1  <= _039_;
always @(posedge \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.clk )
\add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.ain_s1  <= _038_;
always @(posedge \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.clk )
\add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.sum_s1  <= _041_;
always @(posedge \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.clk )
\add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.carry_s1  <= _040_;
assign _039_ = \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.ce  ? \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.b [18:9] : \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.bin_s1 ;
assign _038_ = \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.ce  ? \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.a [18:9] : \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.ain_s1 ;
assign _040_ = \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.ce  ? \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.facout_s1  : \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.carry_s1 ;
assign _041_ = \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.ce  ? \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.fas_s1  : \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.sum_s1 ;
assign _042_ = \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.u1.a  + \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.u1.b ;
assign { \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.u1.cout , \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.u1.s  } = _042_ + \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.u1.cin ;
assign { \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.u2.cout , \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.u2.s  } = _043_ + \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.u2.cin ;
assign _043_ = \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.u2.a  + \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.u2.b ;
always @(posedge \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.clk )
\add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.bin_s1  <= _045_;
always @(posedge \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.clk )
\add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.ain_s1  <= _044_;
always @(posedge \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.clk )
\add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.sum_s1  <= _047_;
always @(posedge \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.clk )
\add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.carry_s1  <= _046_;
assign _045_ = \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.ce  ? \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.b [18:9] : \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.bin_s1 ;
assign _044_ = \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.ce  ? \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.a [18:9] : \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.ain_s1 ;
assign _046_ = \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.ce  ? \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.facout_s1  : \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.carry_s1 ;
assign _047_ = \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.ce  ? \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.fas_s1  : \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.sum_s1 ;
assign _048_ = \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.u1.a  + \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.u1.b ;
assign { \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.u1.cout , \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.u1.s  } = _048_ + \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.u1.cin ;
assign _049_ = \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.u2.a  + \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.u2.b ;
assign { \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.u2.cout , \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.u2.s  } = _049_ + \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.u2.cin ;
always @(posedge \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.clk )
\add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.bin_s1  <= _051_;
always @(posedge \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.clk )
\add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.ain_s1  <= _050_;
always @(posedge \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.clk )
\add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.sum_s1  <= _053_;
always @(posedge \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.clk )
\add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.carry_s1  <= _052_;
assign _051_ = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.ce  ? \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.b [31:16] : \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.bin_s1 ;
assign _050_ = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.ce  ? \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.a [31:16] : \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.ain_s1 ;
assign _052_ = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.ce  ? \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.facout_s1  : \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.carry_s1 ;
assign _053_ = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.ce  ? \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.fas_s1  : \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.sum_s1 ;
assign _054_ = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.u1.a  + \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.u1.b ;
assign { \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.u1.cout , \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.u1.s  } = _054_ + \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.u1.cin ;
assign _055_ = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.u2.a  + \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.u2.b ;
assign { \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.u2.cout , \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.u2.s  } = _055_ + \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.u2.cin ;
always @(posedge \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.clk )
\add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.bin_s1  <= _057_;
always @(posedge \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.clk )
\add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.ain_s1  <= _056_;
always @(posedge \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.clk )
\add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.sum_s1  <= _059_;
always @(posedge \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.clk )
\add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.carry_s1  <= _058_;
assign _057_ = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.ce  ? \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.b [31:16] : \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.bin_s1 ;
assign _056_ = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.ce  ? \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.a [31:16] : \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.ain_s1 ;
assign _058_ = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.ce  ? \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.facout_s1  : \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.carry_s1 ;
assign _059_ = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.ce  ? \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.fas_s1  : \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.sum_s1 ;
assign _060_ = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.u1.a  + \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.u1.b ;
assign { \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.u1.cout , \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.u1.s  } = _060_ + \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.u1.cin ;
assign _061_ = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.u2.a  + \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.u2.b ;
assign { \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.u2.cout , \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.u2.s  } = _061_ + \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.u2.cin ;
always @(posedge \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.clk )
\add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.bin_s1  <= _063_;
always @(posedge \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.clk )
\add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.ain_s1  <= _062_;
always @(posedge \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.clk )
\add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.sum_s1  <= _065_;
always @(posedge \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.clk )
\add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.carry_s1  <= _064_;
assign _063_ = \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.ce  ? \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.b [33:17] : \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.bin_s1 ;
assign _062_ = \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.ce  ? \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.a [33:17] : \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.ain_s1 ;
assign _064_ = \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.ce  ? \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.facout_s1  : \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.carry_s1 ;
assign _065_ = \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.ce  ? \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.fas_s1  : \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.sum_s1 ;
assign _066_ = \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.u1.a  + \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.u1.b ;
assign { \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.u1.cout , \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.u1.s  } = _066_ + \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.u1.cin ;
assign _067_ = \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.u2.a  + \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.u2.b ;
assign { \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.u2.cout , \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.u2.s  } = _067_ + \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.u2.cin ;
always @(posedge \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.clk )
\add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.bin_s1  <= _069_;
always @(posedge \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.clk )
\add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.ain_s1  <= _068_;
always @(posedge \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.clk )
\add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.sum_s1  <= _071_;
always @(posedge \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.clk )
\add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.carry_s1  <= _070_;
assign _069_ = \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.ce  ? \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.b [4:2] : \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.bin_s1 ;
assign _068_ = \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.ce  ? \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.a [4:2] : \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.ain_s1 ;
assign _070_ = \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.ce  ? \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.facout_s1  : \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.carry_s1 ;
assign _071_ = \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.ce  ? \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.fas_s1  : \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.sum_s1 ;
assign _072_ = \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.u1.a  + \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.u1.b ;
assign { \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.u1.cout , \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.u1.s  } = _072_ + \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.u1.cin ;
assign _073_ = \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.u2.a  + \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.u2.b ;
assign { \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.u2.cout , \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.u2.s  } = _073_ + \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.u2.cin ;
always @(posedge \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.clk )
\add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.bin_s1  <= _075_;
always @(posedge \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.clk )
\add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.ain_s1  <= _074_;
always @(posedge \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.clk )
\add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.sum_s1  <= _077_;
always @(posedge \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.clk )
\add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.carry_s1  <= _076_;
assign _075_ = \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.ce  ? \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.b [4:2] : \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.bin_s1 ;
assign _074_ = \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.ce  ? \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.a [4:2] : \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.ain_s1 ;
assign _076_ = \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.ce  ? \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.facout_s1  : \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.carry_s1 ;
assign _077_ = \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.ce  ? \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.fas_s1  : \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.sum_s1 ;
assign _078_ = \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.u1.a  + \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.u1.b ;
assign { \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.u1.cout , \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.u1.s  } = _078_ + \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.u1.cin ;
assign _079_ = \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.u2.a  + \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.u2.b ;
assign { \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.u2.cout , \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.u2.s  } = _079_ + \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.u2.cin ;
always @(posedge \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.clk )
\add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.bin_s1  <= _081_;
always @(posedge \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.clk )
\add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.ain_s1  <= _080_;
always @(posedge \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.clk )
\add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.sum_s1  <= _083_;
always @(posedge \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.clk )
\add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.carry_s1  <= _082_;
assign _081_ = \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.ce  ? \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.b [4:2] : \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.bin_s1 ;
assign _080_ = \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.ce  ? \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.a [4:2] : \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.ain_s1 ;
assign _082_ = \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.ce  ? \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.facout_s1  : \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.carry_s1 ;
assign _083_ = \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.ce  ? \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.fas_s1  : \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.sum_s1 ;
assign _084_ = \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.u1.a  + \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.u1.b ;
assign { \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.u1.cout , \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.u1.s  } = _084_ + \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.u1.cin ;
assign _085_ = \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.u2.a  + \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.u2.b ;
assign { \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.u2.cout , \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.u2.s  } = _085_ + \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.u2.cin ;
always @(posedge \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.clk )
\add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.bin_s1  <= _087_;
always @(posedge \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.clk )
\add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.ain_s1  <= _086_;
always @(posedge \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.clk )
\add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.sum_s1  <= _089_;
always @(posedge \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.clk )
\add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.carry_s1  <= _088_;
assign _087_ = \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.ce  ? \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.b [5:3] : \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.bin_s1 ;
assign _086_ = \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.ce  ? \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.a [5:3] : \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.ain_s1 ;
assign _088_ = \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.ce  ? \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.facout_s1  : \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.carry_s1 ;
assign _089_ = \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.ce  ? \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.fas_s1  : \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.sum_s1 ;
assign _090_ = \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.u1.a  + \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.u1.b ;
assign { \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.u1.cout , \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.u1.s  } = _090_ + \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.u1.cin ;
assign _091_ = \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.u2.a  + \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.u2.b ;
assign { \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.u2.cout , \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.u2.s  } = _091_ + \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.u2.cin ;
always @(posedge \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.clk )
\add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.bin_s1  <= _093_;
always @(posedge \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.clk )
\add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.ain_s1  <= _092_;
always @(posedge \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.clk )
\add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.sum_s1  <= _095_;
always @(posedge \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.clk )
\add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.carry_s1  <= _094_;
assign _093_ = \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.ce  ? \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.b [8:4] : \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.bin_s1 ;
assign _092_ = \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.ce  ? \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.a [8:4] : \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.ain_s1 ;
assign _094_ = \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.ce  ? \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.facout_s1  : \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.carry_s1 ;
assign _095_ = \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.ce  ? \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.fas_s1  : \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.sum_s1 ;
assign _096_ = \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.u1.a  + \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.u1.b ;
assign { \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.u1.cout , \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.u1.s  } = _096_ + \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.u1.cin ;
assign _097_ = \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.u2.a  + \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.u2.b ;
assign { \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.u2.cout , \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.u2.s  } = _097_ + \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.u2.cin ;
assign _098_ = $signed(op_12) > $signed(1'h0);
always @(posedge ap_clk)
sext_ln850_reg_526 <= _018_;
always @(posedge ap_clk)
select_ln353_reg_538 <= _016_;
always @(posedge ap_clk)
ret_V_8_reg_516 <= _014_;
always @(posedge ap_clk)
tmp_reg_521 <= _019_;
always @(posedge ap_clk)
ret_V_6_reg_414 <= _012_;
always @(posedge ap_clk)
ret_V_reg_419 <= _015_;
always @(posedge ap_clk)
trunc_ln851_reg_426 <= _020_;
always @(posedge ap_clk)
ret_V_2_reg_436 <= _011_;
always @(posedge ap_clk)
op_24_V_reg_496 <= _009_;
always @(posedge ap_clk)
icmp_ln851_reg_431 <= _008_;
always @(posedge ap_clk)
icmp_ln1495_reg_548 <= _007_;
always @(posedge ap_clk)
op_26_V_reg_553 <= _010_;
always @(posedge ap_clk)
select_ln69_reg_558 <= _017_;
always @(posedge ap_clk)
add_ln69_4_reg_573 <= _003_;
always @(posedge ap_clk)
add_ln69_6_reg_578 <= _004_;
always @(posedge ap_clk)
add_ln69_reg_476 <= _005_;
always @(posedge ap_clk)
add_ln69_2_reg_481 <= _002_;
always @(posedge ap_clk)
ret_V_7_reg_446 <= _013_;
always @(posedge ap_clk)
add_ln69_1_reg_451 <= _001_;
always @(posedge ap_clk)
add_ln691_reg_533 <= _000_;
always @(posedge ap_clk)
ap_CS_fsm <= _006_;
assign _021_ = _023_ ? 2'h2 : 2'h1;
assign _099_ = ap_CS_fsm == 1'h1;
function [19:0] _291_;
input [19:0] a;
input [399:0] b;
input [19:0] s;
case (s)
20'b00000000000000000001:
_291_ = b[19:0];
20'b00000000000000000010:
_291_ = b[39:20];
20'b00000000000000000100:
_291_ = b[59:40];
20'b00000000000000001000:
_291_ = b[79:60];
20'b00000000000000010000:
_291_ = b[99:80];
20'b00000000000000100000:
_291_ = b[119:100];
20'b00000000000001000000:
_291_ = b[139:120];
20'b00000000000010000000:
_291_ = b[159:140];
20'b00000000000100000000:
_291_ = b[179:160];
20'b00000000001000000000:
_291_ = b[199:180];
20'b00000000010000000000:
_291_ = b[219:200];
20'b00000000100000000000:
_291_ = b[239:220];
20'b00000001000000000000:
_291_ = b[259:240];
20'b00000010000000000000:
_291_ = b[279:260];
20'b00000100000000000000:
_291_ = b[299:280];
20'b00001000000000000000:
_291_ = b[319:300];
20'b00010000000000000000:
_291_ = b[339:320];
20'b00100000000000000000:
_291_ = b[359:340];
20'b01000000000000000000:
_291_ = b[379:360];
20'b10000000000000000000:
_291_ = b[399:380];
20'b00000000000000000000:
_291_ = a;
default:
_291_ = 20'bx;
endcase
endfunction
assign ap_NS_fsm = _291_(20'hxxxxx, { 18'h00000, _021_, 380'h00004000080001000020000400008000100002000040000800010000200004000080001000020000400008000000001 }, { _099_, _118_, _117_, _116_, _115_, _114_, _113_, _112_, _111_, _110_, _109_, _108_, _107_, _106_, _105_, _104_, _103_, _102_, _101_, _100_ });
assign _100_ = ap_CS_fsm == 20'h80000;
assign _101_ = ap_CS_fsm == 19'h40000;
assign _102_ = ap_CS_fsm == 18'h20000;
assign _103_ = ap_CS_fsm == 17'h10000;
assign _104_ = ap_CS_fsm == 16'h8000;
assign _105_ = ap_CS_fsm == 15'h4000;
assign _106_ = ap_CS_fsm == 14'h2000;
assign _107_ = ap_CS_fsm == 13'h1000;
assign _108_ = ap_CS_fsm == 12'h800;
assign _109_ = ap_CS_fsm == 11'h400;
assign _110_ = ap_CS_fsm == 10'h200;
assign _111_ = ap_CS_fsm == 9'h100;
assign _112_ = ap_CS_fsm == 8'h80;
assign _113_ = ap_CS_fsm == 7'h40;
assign _114_ = ap_CS_fsm == 6'h20;
assign _115_ = ap_CS_fsm == 5'h10;
assign _116_ = ap_CS_fsm == 4'h8;
assign _117_ = ap_CS_fsm == 3'h4;
assign _118_ = ap_CS_fsm == 2'h2;
assign op_30_ap_vld = ap_CS_fsm[19] ? 1'h1 : 1'h0;
assign ap_idle = _022_ ? 1'h1 : 1'h0;
assign _018_ = ap_CS_fsm[11] ? { tmp_reg_521[17], tmp_reg_521 } : sext_ln850_reg_526;
assign _016_ = ap_CS_fsm[13] ? select_ln353_fu_320_p3 : select_ln353_reg_538;
assign _019_ = ap_CS_fsm[10] ? grp_fu_279_p2[18:1] : tmp_reg_521;
assign _014_ = ap_CS_fsm[10] ? grp_fu_279_p2 : ret_V_8_reg_516;
assign _020_ = ap_CS_fsm[1] ? grp_fu_171_p2[3:0] : trunc_ln851_reg_426;
assign _015_ = ap_CS_fsm[1] ? grp_fu_171_p2[8:4] : ret_V_reg_419;
assign _012_ = ap_CS_fsm[1] ? grp_fu_171_p2 : ret_V_6_reg_414;
assign _011_ = ap_CS_fsm[3] ? grp_fu_196_p2 : ret_V_2_reg_436;
assign _009_ = ap_CS_fsm[8] ? grp_fu_262_p2 : op_24_V_reg_496;
assign _008_ = ap_CS_fsm[2] ? icmp_ln851_fu_191_p2 : icmp_ln851_reg_431;
assign _017_ = ap_CS_fsm[15] ? select_ln69_fu_370_p3 : select_ln69_reg_558;
assign _010_ = ap_CS_fsm[15] ? grp_fu_338_p2[33:2] : op_26_V_reg_553;
assign _007_ = ap_CS_fsm[15] ? icmp_ln1495_fu_348_p2 : icmp_ln1495_reg_548;
assign _004_ = ap_CS_fsm[17] ? grp_fu_389_p2 : add_ln69_6_reg_578;
assign _003_ = ap_CS_fsm[17] ? grp_fu_385_p2 : add_ln69_4_reg_573;
assign _002_ = ap_CS_fsm[6] ? grp_fu_250_p2 : add_ln69_2_reg_481;
assign _005_ = ap_CS_fsm[6] ? grp_fu_241_p2 : add_ln69_reg_476;
assign _001_ = ap_CS_fsm[4] ? grp_fu_205_p2 : add_ln69_1_reg_451;
assign _013_ = ap_CS_fsm[4] ? ret_V_7_fu_223_p3 : ret_V_7_reg_446;
assign _000_ = ap_CS_fsm[12] ? grp_fu_298_p2 : add_ln691_reg_533;
assign _006_ = ap_rst ? 20'h00001 : ap_NS_fsm;
assign icmp_ln1495_fu_348_p2 = _098_ ? 1'h1 : 1'h0;
assign icmp_ln851_fu_191_p2 = _025_ ? 1'h1 : 1'h0;
assign ret_V_7_fu_223_p3 = ret_V_6_reg_414[8] ? select_ln850_fu_218_p3 : ret_V_reg_419;
assign select_ln353_fu_320_p3 = ret_V_8_reg_516[18] ? select_ln850_2_fu_314_p3 : sext_ln850_reg_526;
assign select_ln69_fu_370_p3 = op_11[0] ? 32'd0 : 32'd4294967295;
assign select_ln850_2_fu_314_p3 = op_14[0] ? add_ln691_reg_533 : sext_ln850_reg_526;
assign select_ln850_fu_218_p3 = icmp_ln851_reg_431 ? ret_V_reg_419 : ret_V_2_reg_436;
assign ap_CS_fsm_state1 = ap_CS_fsm[0];
assign ap_CS_fsm_state10 = ap_CS_fsm[9];
assign ap_CS_fsm_state11 = ap_CS_fsm[10];
assign ap_CS_fsm_state12 = ap_CS_fsm[11];
assign ap_CS_fsm_state13 = ap_CS_fsm[12];
assign ap_CS_fsm_state14 = ap_CS_fsm[13];
assign ap_CS_fsm_state15 = ap_CS_fsm[14];
assign ap_CS_fsm_state16 = ap_CS_fsm[15];
assign ap_CS_fsm_state17 = ap_CS_fsm[16];
assign ap_CS_fsm_state18 = ap_CS_fsm[17];
assign ap_CS_fsm_state19 = ap_CS_fsm[18];
assign ap_CS_fsm_state2 = ap_CS_fsm[1];
assign ap_CS_fsm_state20 = ap_CS_fsm[19];
assign ap_CS_fsm_state3 = ap_CS_fsm[2];
assign ap_CS_fsm_state4 = ap_CS_fsm[3];
assign ap_CS_fsm_state5 = ap_CS_fsm[4];
assign ap_CS_fsm_state6 = ap_CS_fsm[5];
assign ap_CS_fsm_state7 = ap_CS_fsm[6];
assign ap_CS_fsm_state8 = ap_CS_fsm[7];
assign ap_CS_fsm_state9 = ap_CS_fsm[8];
assign ap_done = op_30_ap_vld;
assign ap_ready = op_30_ap_vld;
assign grp_fu_171_p0 = { op_5[1], op_5[1], op_5[1], op_5[1], op_5, 3'h0 };
assign grp_fu_171_p1 = { op_7[7], op_7 };
assign grp_fu_205_p0 = { op_13[3], op_13 };
assign grp_fu_241_p0 = { op_9[15], op_9 };
assign grp_fu_241_p1 = { op_10[15], op_10 };
assign grp_fu_250_p0 = { add_ln69_1_reg_451[4], add_ln69_1_reg_451 };
assign grp_fu_250_p1 = { ret_V_7_reg_446[4], ret_V_7_reg_446 };
assign grp_fu_262_p0 = { add_ln69_2_reg_481[5], add_ln69_2_reg_481[5], add_ln69_2_reg_481[5], add_ln69_2_reg_481[5], add_ln69_2_reg_481[5], add_ln69_2_reg_481[5], add_ln69_2_reg_481[5], add_ln69_2_reg_481[5], add_ln69_2_reg_481[5], add_ln69_2_reg_481[5], add_ln69_2_reg_481[5], add_ln69_2_reg_481[5], add_ln69_2_reg_481 };
assign grp_fu_262_p1 = { add_ln69_reg_476[16], add_ln69_reg_476 };
assign grp_fu_279_p0 = { op_24_V_reg_496, 1'h0 };
assign grp_fu_279_p1 = { op_14[1], op_14[1], op_14[1], op_14[1], op_14[1], op_14[1], op_14[1], op_14[1], op_14[1], op_14[1], op_14[1], op_14[1], op_14[1], op_14[1], op_14[1], op_14[1], op_14[1], op_14 };
assign grp_fu_298_p0 = { tmp_reg_521[17], tmp_reg_521 };
assign grp_fu_338_p0 = { select_ln353_reg_538[18], select_ln353_reg_538[18], select_ln353_reg_538[18], select_ln353_reg_538[18], select_ln353_reg_538[18], select_ln353_reg_538[18], select_ln353_reg_538[18], select_ln353_reg_538[18], select_ln353_reg_538[18], select_ln353_reg_538[18], select_ln353_reg_538[18], select_ln353_reg_538[18], select_ln353_reg_538[18], select_ln353_reg_538, 2'h0 };
assign grp_fu_389_p0 = { 1'h0, op_18 };
assign grp_fu_389_p1 = { 4'h0, icmp_ln1495_reg_548 };
assign grp_fu_398_p0 = { 27'h0000000, add_ln69_6_reg_578 };
assign lhs_fu_155_p3 = { op_5, 3'h0 };
assign op_17_V_fu_344_p1 = op_11[0];
assign op_30 = grp_fu_398_p2;
assign p_Result_1_fu_304_p3 = ret_V_8_reg_516[18];
assign p_Result_s_fu_211_p3 = ret_V_6_reg_414[8];
assign sext_ln1192_1_fu_268_p0 = op_14;
assign sext_ln850_fu_295_p1 = { tmp_reg_521[17], tmp_reg_521 };
assign tmp_3_fu_327_p3 = { select_ln353_reg_538, 2'h0 };
assign trunc_ln851_1_fu_311_p0 = op_14;
assign trunc_ln851_1_fu_311_p1 = op_14[0];
assign trunc_ln851_fu_187_p1 = grp_fu_171_p2[3:0];
assign \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.ain_s0  = \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.a ;
assign \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.bin_s0  = \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.b ;
assign \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.s  = { \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.fas_s2 , \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.sum_s1  };
assign \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.u2.a  = \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.ain_s1 ;
assign \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.u2.b  = \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.bin_s1 ;
assign \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.u2.cin  = \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.carry_s1 ;
assign \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.facout_s2  = \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.u2.cout ;
assign \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.fas_s2  = \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.u2.s ;
assign \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.u1.a  = \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.a [3:0];
assign \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.u1.b  = \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.b [3:0];
assign \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.u1.cin  = 1'h0;
assign \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.facout_s1  = \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.u1.cout ;
assign \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.fas_s1  = \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.u1.s ;
assign \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.a  = \add_9s_9s_9_2_1_U1.din0 ;
assign \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.b  = \add_9s_9s_9_2_1_U1.din1 ;
assign \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.ce  = \add_9s_9s_9_2_1_U1.ce ;
assign \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.clk  = \add_9s_9s_9_2_1_U1.clk ;
assign \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.reset  = \add_9s_9s_9_2_1_U1.reset ;
assign \add_9s_9s_9_2_1_U1.dout  = \add_9s_9s_9_2_1_U1.top_add_9s_9s_9_2_1_Adder_0_U.s ;
assign \add_9s_9s_9_2_1_U1.ce  = 1'h1;
assign \add_9s_9s_9_2_1_U1.clk  = ap_clk;
assign \add_9s_9s_9_2_1_U1.din0  = { op_5[1], op_5[1], op_5[1], op_5[1], op_5, 3'h0 };
assign \add_9s_9s_9_2_1_U1.din1  = { op_7[7], op_7 };
assign grp_fu_171_p2 = \add_9s_9s_9_2_1_U1.dout ;
assign \add_9s_9s_9_2_1_U1.reset  = ap_rst;
assign \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.ain_s0  = \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.a ;
assign \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.bin_s0  = \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.b ;
assign \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.s  = { \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.fas_s2 , \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.sum_s1  };
assign \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.u2.a  = \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.ain_s1 ;
assign \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.u2.b  = \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.bin_s1 ;
assign \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.u2.cin  = \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.carry_s1 ;
assign \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.facout_s2  = \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.u2.cout ;
assign \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.fas_s2  = \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.u2.s ;
assign \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.u1.a  = \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.a [2:0];
assign \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.u1.b  = \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.b [2:0];
assign \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.u1.cin  = 1'h0;
assign \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.facout_s1  = \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.u1.cout ;
assign \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.fas_s1  = \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.u1.s ;
assign \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.a  = \add_6s_6s_6_2_1_U5.din0 ;
assign \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.b  = \add_6s_6s_6_2_1_U5.din1 ;
assign \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.ce  = \add_6s_6s_6_2_1_U5.ce ;
assign \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.clk  = \add_6s_6s_6_2_1_U5.clk ;
assign \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.reset  = \add_6s_6s_6_2_1_U5.reset ;
assign \add_6s_6s_6_2_1_U5.dout  = \add_6s_6s_6_2_1_U5.top_add_6s_6s_6_2_1_Adder_4_U.s ;
assign \add_6s_6s_6_2_1_U5.ce  = 1'h1;
assign \add_6s_6s_6_2_1_U5.clk  = ap_clk;
assign \add_6s_6s_6_2_1_U5.din0  = { add_ln69_1_reg_451[4], add_ln69_1_reg_451 };
assign \add_6s_6s_6_2_1_U5.din1  = { ret_V_7_reg_446[4], ret_V_7_reg_446 };
assign grp_fu_250_p2 = \add_6s_6s_6_2_1_U5.dout ;
assign \add_6s_6s_6_2_1_U5.reset  = ap_rst;
assign \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.ain_s0  = \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.a ;
assign \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.bin_s0  = \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.b ;
assign \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.s  = { \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.fas_s2 , \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.sum_s1  };
assign \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.u2.a  = \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.ain_s1 ;
assign \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.u2.b  = \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.bin_s1 ;
assign \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.u2.cin  = \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.carry_s1 ;
assign \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.facout_s2  = \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.u2.cout ;
assign \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.fas_s2  = \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.u2.s ;
assign \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.u1.a  = \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.a [1:0];
assign \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.u1.b  = \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.b [1:0];
assign \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.u1.cin  = 1'h0;
assign \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.facout_s1  = \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.u1.cout ;
assign \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.fas_s1  = \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.u1.s ;
assign \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.a  = \add_5s_5ns_5_2_1_U3.din0 ;
assign \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.b  = \add_5s_5ns_5_2_1_U3.din1 ;
assign \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.ce  = \add_5s_5ns_5_2_1_U3.ce ;
assign \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.clk  = \add_5s_5ns_5_2_1_U3.clk ;
assign \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.reset  = \add_5s_5ns_5_2_1_U3.reset ;
assign \add_5s_5ns_5_2_1_U3.dout  = \add_5s_5ns_5_2_1_U3.top_add_5s_5ns_5_2_1_Adder_2_U.s ;
assign \add_5s_5ns_5_2_1_U3.ce  = 1'h1;
assign \add_5s_5ns_5_2_1_U3.clk  = ap_clk;
assign \add_5s_5ns_5_2_1_U3.din0  = { op_13[3], op_13 };
assign \add_5s_5ns_5_2_1_U3.din1  = 5'h01;
assign grp_fu_205_p2 = \add_5s_5ns_5_2_1_U3.dout ;
assign \add_5s_5ns_5_2_1_U3.reset  = ap_rst;
assign \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.ain_s0  = \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.a ;
assign \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.bin_s0  = \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.b ;
assign \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.s  = { \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.fas_s2 , \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.sum_s1  };
assign \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.u2.a  = \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.ain_s1 ;
assign \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.u2.b  = \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.bin_s1 ;
assign \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.u2.cin  = \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.carry_s1 ;
assign \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.facout_s2  = \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.u2.cout ;
assign \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.fas_s2  = \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.u2.s ;
assign \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.u1.a  = \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.a [1:0];
assign \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.u1.b  = \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.b [1:0];
assign \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.u1.cin  = 1'h0;
assign \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.facout_s1  = \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.u1.cout ;
assign \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.fas_s1  = \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.u1.s ;
assign \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.a  = \add_5ns_5ns_5_2_1_U2.din0 ;
assign \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.b  = \add_5ns_5ns_5_2_1_U2.din1 ;
assign \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.ce  = \add_5ns_5ns_5_2_1_U2.ce ;
assign \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.clk  = \add_5ns_5ns_5_2_1_U2.clk ;
assign \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.reset  = \add_5ns_5ns_5_2_1_U2.reset ;
assign \add_5ns_5ns_5_2_1_U2.dout  = \add_5ns_5ns_5_2_1_U2.top_add_5ns_5ns_5_2_1_Adder_1_U.s ;
assign \add_5ns_5ns_5_2_1_U2.ce  = 1'h1;
assign \add_5ns_5ns_5_2_1_U2.clk  = ap_clk;
assign \add_5ns_5ns_5_2_1_U2.din0  = ret_V_reg_419;
assign \add_5ns_5ns_5_2_1_U2.din1  = 5'h01;
assign grp_fu_196_p2 = \add_5ns_5ns_5_2_1_U2.dout ;
assign \add_5ns_5ns_5_2_1_U2.reset  = ap_rst;
assign \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.ain_s0  = \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.a ;
assign \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.bin_s0  = \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.b ;
assign \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.s  = { \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.fas_s2 , \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.sum_s1  };
assign \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.u2.a  = \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.ain_s1 ;
assign \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.u2.b  = \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.bin_s1 ;
assign \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.u2.cin  = \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.carry_s1 ;
assign \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.facout_s2  = \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.u2.cout ;
assign \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.fas_s2  = \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.u2.s ;
assign \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.u1.a  = \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.a [1:0];
assign \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.u1.b  = \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.b [1:0];
assign \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.u1.cin  = 1'h0;
assign \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.facout_s1  = \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.u1.cout ;
assign \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.fas_s1  = \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.u1.s ;
assign \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.a  = \add_5ns_5ns_5_2_1_U11.din0 ;
assign \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.b  = \add_5ns_5ns_5_2_1_U11.din1 ;
assign \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.ce  = \add_5ns_5ns_5_2_1_U11.ce ;
assign \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.clk  = \add_5ns_5ns_5_2_1_U11.clk ;
assign \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.reset  = \add_5ns_5ns_5_2_1_U11.reset ;
assign \add_5ns_5ns_5_2_1_U11.dout  = \add_5ns_5ns_5_2_1_U11.top_add_5ns_5ns_5_2_1_Adder_1_U.s ;
assign \add_5ns_5ns_5_2_1_U11.ce  = 1'h1;
assign \add_5ns_5ns_5_2_1_U11.clk  = ap_clk;
assign \add_5ns_5ns_5_2_1_U11.din0  = { 1'h0, op_18 };
assign \add_5ns_5ns_5_2_1_U11.din1  = { 4'h0, icmp_ln1495_reg_548 };
assign grp_fu_389_p2 = \add_5ns_5ns_5_2_1_U11.dout ;
assign \add_5ns_5ns_5_2_1_U11.reset  = ap_rst;
assign \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.ain_s0  = \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.a ;
assign \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.bin_s0  = \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.b ;
assign \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.s  = { \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.fas_s2 , \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.sum_s1  };
assign \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.u2.a  = \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.ain_s1 ;
assign \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.u2.b  = \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.bin_s1 ;
assign \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.u2.cin  = \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.carry_s1 ;
assign \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.facout_s2  = \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.u2.cout ;
assign \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.fas_s2  = \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.u2.s ;
assign \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.u1.a  = \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.a [16:0];
assign \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.u1.b  = \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.b [16:0];
assign \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.u1.cin  = 1'h0;
assign \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.facout_s1  = \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.u1.cout ;
assign \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.fas_s1  = \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.u1.s ;
assign \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.a  = \add_34s_34ns_34_2_1_U9.din0 ;
assign \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.b  = \add_34s_34ns_34_2_1_U9.din1 ;
assign \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.ce  = \add_34s_34ns_34_2_1_U9.ce ;
assign \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.clk  = \add_34s_34ns_34_2_1_U9.clk ;
assign \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.reset  = \add_34s_34ns_34_2_1_U9.reset ;
assign \add_34s_34ns_34_2_1_U9.dout  = \add_34s_34ns_34_2_1_U9.top_add_34s_34ns_34_2_1_Adder_8_U.s ;
assign \add_34s_34ns_34_2_1_U9.ce  = 1'h1;
assign \add_34s_34ns_34_2_1_U9.clk  = ap_clk;
assign \add_34s_34ns_34_2_1_U9.din0  = { select_ln353_reg_538[18], select_ln353_reg_538[18], select_ln353_reg_538[18], select_ln353_reg_538[18], select_ln353_reg_538[18], select_ln353_reg_538[18], select_ln353_reg_538[18], select_ln353_reg_538[18], select_ln353_reg_538[18], select_ln353_reg_538[18], select_ln353_reg_538[18], select_ln353_reg_538[18], select_ln353_reg_538[18], select_ln353_reg_538, 2'h0 };
assign \add_34s_34ns_34_2_1_U9.din1  = 34'h000000004;
assign grp_fu_338_p2 = \add_34s_34ns_34_2_1_U9.dout ;
assign \add_34s_34ns_34_2_1_U9.reset  = ap_rst;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.ain_s0  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.a ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.bin_s0  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.b ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.s  = { \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.fas_s2 , \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.sum_s1  };
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.u2.a  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.ain_s1 ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.u2.b  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.bin_s1 ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.u2.cin  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.carry_s1 ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.facout_s2  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.u2.cout ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.fas_s2  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.u2.s ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.u1.a  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.a [15:0];
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.u1.b  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.b [15:0];
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.u1.cin  = 1'h0;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.facout_s1  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.u1.cout ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.fas_s1  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.u1.s ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.a  = \add_32ns_32ns_32_2_1_U12.din0 ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.b  = \add_32ns_32ns_32_2_1_U12.din1 ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.ce  = \add_32ns_32ns_32_2_1_U12.ce ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.clk  = \add_32ns_32ns_32_2_1_U12.clk ;
assign \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.reset  = \add_32ns_32ns_32_2_1_U12.reset ;
assign \add_32ns_32ns_32_2_1_U12.dout  = \add_32ns_32ns_32_2_1_U12.top_add_32ns_32ns_32_2_1_Adder_9_U.s ;
assign \add_32ns_32ns_32_2_1_U12.ce  = 1'h1;
assign \add_32ns_32ns_32_2_1_U12.clk  = ap_clk;
assign \add_32ns_32ns_32_2_1_U12.din0  = { 27'h0000000, add_ln69_6_reg_578 };
assign \add_32ns_32ns_32_2_1_U12.din1  = add_ln69_4_reg_573;
assign grp_fu_398_p2 = \add_32ns_32ns_32_2_1_U12.dout ;
assign \add_32ns_32ns_32_2_1_U12.reset  = ap_rst;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.ain_s0  = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.a ;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.bin_s0  = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.b ;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.s  = { \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.fas_s2 , \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.sum_s1  };
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.u2.a  = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.ain_s1 ;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.u2.b  = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.bin_s1 ;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.u2.cin  = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.carry_s1 ;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.facout_s2  = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.u2.cout ;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.fas_s2  = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.u2.s ;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.u1.a  = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.a [15:0];
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.u1.b  = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.b [15:0];
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.u1.cin  = 1'h0;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.facout_s1  = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.u1.cout ;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.fas_s1  = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.u1.s ;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.a  = \add_32ns_32ns_32_2_1_U10.din0 ;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.b  = \add_32ns_32ns_32_2_1_U10.din1 ;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.ce  = \add_32ns_32ns_32_2_1_U10.ce ;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.clk  = \add_32ns_32ns_32_2_1_U10.clk ;
assign \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.reset  = \add_32ns_32ns_32_2_1_U10.reset ;
assign \add_32ns_32ns_32_2_1_U10.dout  = \add_32ns_32ns_32_2_1_U10.top_add_32ns_32ns_32_2_1_Adder_9_U.s ;
assign \add_32ns_32ns_32_2_1_U10.ce  = 1'h1;
assign \add_32ns_32ns_32_2_1_U10.clk  = ap_clk;
assign \add_32ns_32ns_32_2_1_U10.din0  = op_26_V_reg_553;
assign \add_32ns_32ns_32_2_1_U10.din1  = select_ln69_reg_558;
assign grp_fu_385_p2 = \add_32ns_32ns_32_2_1_U10.dout ;
assign \add_32ns_32ns_32_2_1_U10.reset  = ap_rst;
assign \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.ain_s0  = \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.a ;
assign \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.bin_s0  = \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.b ;
assign \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.s  = { \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.fas_s2 , \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.sum_s1  };
assign \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.u2.a  = \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.ain_s1 ;
assign \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.u2.b  = \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.bin_s1 ;
assign \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.u2.cin  = \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.carry_s1 ;
assign \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.facout_s2  = \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.u2.cout ;
assign \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.fas_s2  = \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.u2.s ;
assign \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.u1.a  = \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.a [8:0];
assign \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.u1.b  = \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.b [8:0];
assign \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.u1.cin  = 1'h0;
assign \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.facout_s1  = \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.u1.cout ;
assign \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.fas_s1  = \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.u1.s ;
assign \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.a  = \add_19s_19ns_19_2_1_U8.din0 ;
assign \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.b  = \add_19s_19ns_19_2_1_U8.din1 ;
assign \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.ce  = \add_19s_19ns_19_2_1_U8.ce ;
assign \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.clk  = \add_19s_19ns_19_2_1_U8.clk ;
assign \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.reset  = \add_19s_19ns_19_2_1_U8.reset ;
assign \add_19s_19ns_19_2_1_U8.dout  = \add_19s_19ns_19_2_1_U8.top_add_19s_19ns_19_2_1_Adder_7_U.s ;
assign \add_19s_19ns_19_2_1_U8.ce  = 1'h1;
assign \add_19s_19ns_19_2_1_U8.clk  = ap_clk;
assign \add_19s_19ns_19_2_1_U8.din0  = { tmp_reg_521[17], tmp_reg_521 };
assign \add_19s_19ns_19_2_1_U8.din1  = 19'h00001;
assign grp_fu_298_p2 = \add_19s_19ns_19_2_1_U8.dout ;
assign \add_19s_19ns_19_2_1_U8.reset  = ap_rst;
assign \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.ain_s0  = \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.a ;
assign \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.bin_s0  = \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.b ;
assign \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.s  = { \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.fas_s2 , \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.sum_s1  };
assign \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.u2.a  = \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.ain_s1 ;
assign \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.u2.b  = \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.bin_s1 ;
assign \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.u2.cin  = \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.carry_s1 ;
assign \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.facout_s2  = \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.u2.cout ;
assign \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.fas_s2  = \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.u2.s ;
assign \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.u1.a  = \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.a [8:0];
assign \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.u1.b  = \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.b [8:0];
assign \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.u1.cin  = 1'h0;
assign \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.facout_s1  = \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.u1.cout ;
assign \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.fas_s1  = \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.u1.s ;
assign \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.a  = \add_19ns_19s_19_2_1_U7.din0 ;
assign \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.b  = \add_19ns_19s_19_2_1_U7.din1 ;
assign \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.ce  = \add_19ns_19s_19_2_1_U7.ce ;
assign \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.clk  = \add_19ns_19s_19_2_1_U7.clk ;
assign \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.reset  = \add_19ns_19s_19_2_1_U7.reset ;
assign \add_19ns_19s_19_2_1_U7.dout  = \add_19ns_19s_19_2_1_U7.top_add_19ns_19s_19_2_1_Adder_6_U.s ;
assign \add_19ns_19s_19_2_1_U7.ce  = 1'h1;
assign \add_19ns_19s_19_2_1_U7.clk  = ap_clk;
assign \add_19ns_19s_19_2_1_U7.din0  = { op_24_V_reg_496, 1'h0 };
assign \add_19ns_19s_19_2_1_U7.din1  = { op_14[1], op_14[1], op_14[1], op_14[1], op_14[1], op_14[1], op_14[1], op_14[1], op_14[1], op_14[1], op_14[1], op_14[1], op_14[1], op_14[1], op_14[1], op_14[1], op_14[1], op_14 };
assign grp_fu_279_p2 = \add_19ns_19s_19_2_1_U7.dout ;
assign \add_19ns_19s_19_2_1_U7.reset  = ap_rst;
assign \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.ain_s0  = \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.a ;
assign \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.bin_s0  = \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.b ;
assign \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.s  = { \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.fas_s2 , \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.sum_s1  };
assign \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.u2.a  = \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.ain_s1 ;
assign \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.u2.b  = \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.bin_s1 ;
assign \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.u2.cin  = \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.carry_s1 ;
assign \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.facout_s2  = \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.u2.cout ;
assign \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.fas_s2  = \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.u2.s ;
assign \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.u1.a  = \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.a [8:0];
assign \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.u1.b  = \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.b [8:0];
assign \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.u1.cin  = 1'h0;
assign \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.facout_s1  = \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.u1.cout ;
assign \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.fas_s1  = \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.u1.s ;
assign \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.a  = \add_18s_18s_18_2_1_U6.din0 ;
assign \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.b  = \add_18s_18s_18_2_1_U6.din1 ;
assign \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.ce  = \add_18s_18s_18_2_1_U6.ce ;
assign \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.clk  = \add_18s_18s_18_2_1_U6.clk ;
assign \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.reset  = \add_18s_18s_18_2_1_U6.reset ;
assign \add_18s_18s_18_2_1_U6.dout  = \add_18s_18s_18_2_1_U6.top_add_18s_18s_18_2_1_Adder_5_U.s ;
assign \add_18s_18s_18_2_1_U6.ce  = 1'h1;
assign \add_18s_18s_18_2_1_U6.clk  = ap_clk;
assign \add_18s_18s_18_2_1_U6.din0  = { add_ln69_2_reg_481[5], add_ln69_2_reg_481[5], add_ln69_2_reg_481[5], add_ln69_2_reg_481[5], add_ln69_2_reg_481[5], add_ln69_2_reg_481[5], add_ln69_2_reg_481[5], add_ln69_2_reg_481[5], add_ln69_2_reg_481[5], add_ln69_2_reg_481[5], add_ln69_2_reg_481[5], add_ln69_2_reg_481[5], add_ln69_2_reg_481 };
assign \add_18s_18s_18_2_1_U6.din1  = { add_ln69_reg_476[16], add_ln69_reg_476 };
assign grp_fu_262_p2 = \add_18s_18s_18_2_1_U6.dout ;
assign \add_18s_18s_18_2_1_U6.reset  = ap_rst;
assign \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.ain_s0  = \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.a ;
assign \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.bin_s0  = \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.b ;
assign \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.s  = { \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.fas_s2 , \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.sum_s1  };
assign \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.u2.a  = \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.ain_s1 ;
assign \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.u2.b  = \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.bin_s1 ;
assign \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.u2.cin  = \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.carry_s1 ;
assign \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.facout_s2  = \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.u2.cout ;
assign \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.fas_s2  = \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.u2.s ;
assign \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.u1.a  = \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.a [7:0];
assign \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.u1.b  = \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.b [7:0];
assign \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.u1.cin  = 1'h0;
assign \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.facout_s1  = \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.u1.cout ;
assign \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.fas_s1  = \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.u1.s ;
assign \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.a  = \add_17s_17s_17_2_1_U4.din0 ;
assign \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.b  = \add_17s_17s_17_2_1_U4.din1 ;
assign \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.ce  = \add_17s_17s_17_2_1_U4.ce ;
assign \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.clk  = \add_17s_17s_17_2_1_U4.clk ;
assign \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.reset  = \add_17s_17s_17_2_1_U4.reset ;
assign \add_17s_17s_17_2_1_U4.dout  = \add_17s_17s_17_2_1_U4.top_add_17s_17s_17_2_1_Adder_3_U.s ;
assign \add_17s_17s_17_2_1_U4.ce  = 1'h1;
assign \add_17s_17s_17_2_1_U4.clk  = ap_clk;
assign \add_17s_17s_17_2_1_U4.din0  = { op_9[15], op_9 };
assign \add_17s_17s_17_2_1_U4.din1  = { op_10[15], op_10 };
assign grp_fu_241_p2 = \add_17s_17s_17_2_1_U4.dout ;
assign \add_17s_17s_17_2_1_U4.reset  = ap_rst;
endmodule


// Product machine:
module top_A_times_top_B (ap_start, op_0, op_10, op_11, op_12, op_13, op_14, op_18, op_5, op_7, op_9, ap_clk, unsafe_signal);
input ap_start;
input [1:0] op_0;
input [15:0] op_10;
input [1:0] op_11;
input [7:0] op_12;
input [3:0] op_13;
input [1:0] op_14;
input [3:0] op_18;
input [1:0] op_5;
input [7:0] op_7;
input [15:0] op_9;
input ap_clk;
output unsafe_signal;
reg _setup;
initial _setup = 1'b0;
always @ (posedge ap_clk) _setup <= 1'b1;
reg ap_start_internal;
always @ (posedge ap_clk) if (!_setup) ap_start_internal <= ap_start;
reg [1:0] op_0_internal;
always @ (posedge ap_clk) if (!_setup) op_0_internal <= op_0;
reg [15:0] op_10_internal;
always @ (posedge ap_clk) if (!_setup) op_10_internal <= op_10;
reg [1:0] op_11_internal;
always @ (posedge ap_clk) if (!_setup) op_11_internal <= op_11;
reg [7:0] op_12_internal;
always @ (posedge ap_clk) if (!_setup) op_12_internal <= op_12;
reg [3:0] op_13_internal;
always @ (posedge ap_clk) if (!_setup) op_13_internal <= op_13;
reg [1:0] op_14_internal;
always @ (posedge ap_clk) if (!_setup) op_14_internal <= op_14;
reg [3:0] op_18_internal;
always @ (posedge ap_clk) if (!_setup) op_18_internal <= op_18;
reg [1:0] op_5_internal;
always @ (posedge ap_clk) if (!_setup) op_5_internal <= op_5;
reg [7:0] op_7_internal;
always @ (posedge ap_clk) if (!_setup) op_7_internal <= op_7;
reg [15:0] op_9_internal;
always @ (posedge ap_clk) if (!_setup) op_9_internal <= op_9;
wire ap_done_A;
wire ap_done_B;
wire ap_done_eq;
assign ap_done_eq = ap_done_A == ap_done_B;
wire ap_idle_A;
wire ap_idle_B;
wire ap_idle_eq;
assign ap_idle_eq = ap_idle_A == ap_idle_B;
wire ap_ready_A;
wire ap_ready_B;
wire ap_ready_eq;
assign ap_ready_eq = ap_ready_A == ap_ready_B;
wire [31:0] op_30_A;
wire [31:0] op_30_B;
wire op_30_eq;
assign op_30_eq = op_30_A == op_30_B;
wire op_30_ap_vld_A;
wire op_30_ap_vld_B;
wire clk_enable_A;
wire clk_enable_B;
assign clk_enable_A = _setup & (~op_30_ap_vld_A | op_30_ap_vld_B);
assign clk_enable_B = _setup;
wire divergent;
assign divergent = ~(ap_done_eq & ap_idle_eq & ap_ready_eq & op_30_eq);
assign unsafe_signal = op_30_ap_vld_A & op_30_ap_vld_B & divergent;
top_A instance_A (
    .ap_clk(ap_clk),
    .clk_enable(clk_enable_A),
    .ap_start(ap_start_internal),
    .op_0(op_0_internal),
    .op_10(op_10_internal),
    .op_11(op_11_internal),
    .op_12(op_12_internal),
    .op_13(op_13_internal),
    .op_14(op_14_internal),
    .op_18(op_18_internal),
    .op_5(op_5_internal),
    .op_7(op_7_internal),
    .op_9(op_9_internal),
    .ap_done(ap_done_A),
    .ap_idle(ap_idle_A),
    .ap_ready(ap_ready_A),
    .op_30(op_30_A),
    .op_30_ap_vld(op_30_ap_vld_A)
);
top_B instance_B (
    .ap_clk(ap_clk),
    .clk_enable(clk_enable_B),
    .ap_start(ap_start_internal),
    .op_0(op_0_internal),
    .op_10(op_10_internal),
    .op_11(op_11_internal),
    .op_12(op_12_internal),
    .op_13(op_13_internal),
    .op_14(op_14_internal),
    .op_18(op_18_internal),
    .op_5(op_5_internal),
    .op_7(op_7_internal),
    .op_9(op_9_internal),
    .ap_done(ap_done_B),
    .ap_idle(ap_idle_B),
    .ap_ready(ap_ready_B),
    .op_30(op_30_B),
    .op_30_ap_vld(op_30_ap_vld_B)
);
endmodule
